`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  reg [0:0] PI_wbs_cyc_i;
  reg [0:0] PI_wb_rst_i;
  reg [0:0] PI_rst_i;
  reg [7:0] PI_hb_dq_i;
  reg [31:0] PI_wbs_dat_i;
  reg [0:0] PI_wbs_we_i;
  reg [0:0] PI_wb_clk_i;
  reg [0:0] PI_hb_rwds_i;
  reg [0:0] PI_wbs_stb_i;
  reg [3:0] PI_wbs_sel_i;
  reg [31:0] PI_wbs_addr_i;
  wb_hyperram UUT (
    .wbs_cyc_i(PI_wbs_cyc_i),
    .wb_rst_i(PI_wb_rst_i),
    .rst_i(PI_rst_i),
    .hb_dq_i(PI_hb_dq_i),
    .wbs_dat_i(PI_wbs_dat_i),
    .wbs_we_i(PI_wbs_we_i),
    .wb_clk_i(PI_wb_clk_i),
    .hb_rwds_i(PI_hb_rwds_i),
    .wbs_stb_i(PI_wbs_stb_i),
    .wbs_sel_i(PI_wbs_sel_i),
    .wbs_addr_i(PI_wbs_addr_i)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    // UUT.$and$wb_hyperram.\v:0$463_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$472_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$476_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$494_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$507_Y  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:156:execute$6225  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:156:execute$6235  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:156:execute$6245  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:168:execute$6227  = 1'b1;
    // UUT.$auto$clk2fflogic.\cc:192:execute$6231  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:192:execute$6241  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:192:execute$6251  = 1'b0;
    // UUT.$eq$wb_hyperram.\v:435$654_Y  = 1'b0;
    // UUT.$eq$wb_hyperram.\v:544$796_Y  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:270$128_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:270$128_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:272$129_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:272$129_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:276$130_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:276$130_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:281$131_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:281$131_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:283$132_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:283$132_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:288$133_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:288$133_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:290$134_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:290$134_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:322$135_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:322$135_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:323$136_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:327$137_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:327$137_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:328$138_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:329$139_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:330$140_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:331$141_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:332$142_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:336$143_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:336$143_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:337$144_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:338$145_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:339$146_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:340$147_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:349$148_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:350$149_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:351$150_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:352$151_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:356$152_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:359$153_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:362$154_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:365$155_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:370$156_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:386$157_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:400$158_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:415$159_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:429$160_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:445$161_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:461$162_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:474$163_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:490$164_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:510$165_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:524$166_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:524$166_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:531$167_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:531$167_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:533$168_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:533$168_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:535$169_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:535$169_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:537$170_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:537$170_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:539$171_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:539$171_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:546$172_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:546$172_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:548$173_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:548$173_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:550$174_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:550$174_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:552$175_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:552$175_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:559$176_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:559$176_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:561$177_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:561$177_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:567$178_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:567$178_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:569$179_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:569$179_EN  = 1'b0;
    // UUT.$past$wb_hyperram.\v:330$17$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:331$18$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:332$19$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:333$20$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:349$25$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:350$26$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:351$28$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:374$30$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:375$31$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:381$36$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:381$37$0  = 6'b000000;
    // UUT.$past$wb_hyperram.\v:390$40$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:393$42$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:404$48$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:407$50$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:408$51$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:419$58$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:422$60$0  = 5'b00000;
    // UUT.$past$wb_hyperram.\v:447$72$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:448$73$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:454$77$0  = 3'b000;
    // UUT.$past$wb_hyperram.\v:492$91$0  = 1'b0;
    UUT.f_past_valid = 1'b0;
    // UUT.hram.$and$hyperram.\v:0$1779_Y  = 1'b0;
    // UUT.hram.$and$hyperram.\v:0$1788_Y  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6025  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6035  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6045  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6055  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6065  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6075  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6085  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6095  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6105  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6115  = 5'b00000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6125  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6135  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6145  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6155  = 48'b000000000000000000000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6165  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6175  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6185  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6195  = 3'b010;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6205  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$6215  = 6'b100000;
    // UUT.hram.$auto$clk2fflogic.\cc:168:execute$6027  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:168:execute$6077  = 1'b1;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6031  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6041  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6051  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6061  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6071  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6081  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6091  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6101  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6111  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6121  = 5'b00000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6131  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6141  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6151  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6161  = 48'b000000000000000000000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6171  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6181  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6191  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6201  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6211  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$6221  = 6'b000000;
    // UUT.hram.$formal$hyperram.\v:1000$1262_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1000$1262_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1003$1263_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1003$1263_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1006$1264_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1006$1264_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1010$1265_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1010$1265_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1012$1266_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1012$1266_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1016$1267_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1016$1267_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1018$1268_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1018$1268_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1020$1269_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1020$1269_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1024$1270_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1024$1270_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1027$1271_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1027$1271_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1030$1272_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1030$1272_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1036$1273_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1039$1274_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1039$1274_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1042$1275_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1042$1275_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1045$1276_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1045$1276_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1048$1277_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1048$1277_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1053$1278_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1057$1279_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1057$1279_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1059$1280_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1059$1280_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1072$1282_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1072$1282_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1084$1283_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1084$1283_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1085$1284_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1085$1284_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1086$1285_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1086$1285_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1087$1286_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1087$1286_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1095$1287_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1095$1287_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1096$1288_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1097$1289_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1098$1290_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:402$1192_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:402$1192_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:405$1193_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:405$1193_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:412$1194_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:415$1195_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:418$1196_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:421$1197_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:424$1198_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:430$1199_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:445$1200_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:462$1201_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:482$1202_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:502$1203_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:524$1204_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:540$1205_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:559$1206_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:580$1207_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:600$1208_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:622$1209_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:638$1210_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:655$1211_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:675$1212_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:695$1213_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:716$1214_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:733$1215_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:752$1216_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:768$1217_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:784$1218_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:803$1219_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:820$1220_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:838$1221_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:854$1222_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:854$1222_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:860$1223_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:861$1224_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:867$1225_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:867$1225_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:868$1226_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:869$1227_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:872$1228_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:872$1228_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:874$1229_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:874$1229_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:877$1230_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:877$1230_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:879$1231_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:879$1231_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:879$1232_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:881$1233_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:889$1234_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:889$1234_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:891$1235_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:891$1235_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:893$1236_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:893$1236_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:907$1237_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:907$1237_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:923$1238_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:923$1238_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:925$1239_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:925$1239_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:929$1240_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:929$1240_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:931$1241_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:931$1241_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:937$1242_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:937$1242_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:939$1243_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:939$1243_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:944$1244_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:944$1244_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:945$1245_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:946$1246_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:947$1247_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:949$1248_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:949$1248_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:955$1249_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:955$1249_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:959$1250_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:959$1250_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:962$1251_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:962$1251_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:965$1252_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:965$1252_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:968$1253_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:968$1253_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:972$1254_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:972$1254_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:974$1255_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:974$1255_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:978$1256_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:978$1256_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:981$1257_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:981$1257_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:984$1258_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:984$1258_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:987$1259_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:987$1259_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:990$1260_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:990$1260_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:997$1261_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:997$1261_EN  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1038$1163$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1038$1164$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1071$1173$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1078$1174$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1084$1176$0  = 8'b00000000;
    // UUT.hram.$past$hyperram.\v:1095$1184$0  = 32'b00000000000000000000000000000000;
    // UUT.hram.$past$hyperram.\v:1096$1185$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:1097$1186$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1098$1187$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:436$999$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:867$1112$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:868$1113$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:869$1114$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:871$1115$0  = 5'b00000;
    // UUT.hram.$past$hyperram.\v:876$1117$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:881$1119$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:882$1120$0  = 1'b0;
    UUT.hram.f_past_valid = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5635  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5645  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5655  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5665  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5675  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5685  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5695  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5705  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5715  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5725  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5735  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5745  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5755  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:168:execute$5637  = 1'b1;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5641  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5661  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5671  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5681  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5691  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5701  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5711  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5721  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5731  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5741  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5751  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5761  = 6'b000000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5505  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5515  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5525  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5535  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5545  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5555  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5565  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5575  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5585  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5595  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5605  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5615  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5625  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:168:execute$5507  = 1'b1;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5511  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5531  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5541  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5551  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5561  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5571  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5581  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5591  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5601  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5611  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5621  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5631  = 4'b0000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5765  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5775  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5785  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5795  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5805  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5815  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5825  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5835  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5845  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5855  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5865  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5875  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5885  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:168:execute$5767  = 1'b1;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5771  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5791  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5801  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5811  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5821  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5831  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5841  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5851  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5861  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5871  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5881  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5891  = 8'b00000000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5895  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5905  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5915  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5925  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5935  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5945  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5955  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5965  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5975  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5985  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$5995  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$6005  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$6015  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:168:execute$5897  = 1'b1;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5901  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5921  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5931  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5941  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5951  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5961  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5971  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5981  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$5991  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$6001  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$6011  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$6021  = 5'b00000;
    UUT.wb_state = 2'b00;

    // state 0
    PI_wbs_cyc_i = 1'b0;
    PI_wb_rst_i = 1'b1;
    PI_rst_i = 1'b1;
    PI_hb_dq_i = 8'b00000000;
    PI_wbs_dat_i = 32'b10000000000000000000000000000000;
    PI_wbs_we_i = 1'b0;
    PI_wb_clk_i = 1'b0;
    PI_hb_rwds_i = 1'b0;
    PI_wbs_stb_i = 1'b0;
    PI_wbs_sel_i = 4'b1000;
    PI_wbs_addr_i = 32'b00000000001000000000000000000000;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      PI_wbs_cyc_i <= 1'b0;
      PI_wb_rst_i <= 1'b1;
      PI_rst_i <= 1'b1;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
      PI_wbs_we_i <= 1'b0;
      PI_wb_clk_i <= 1'b1;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b0;
      PI_wbs_sel_i <= 4'b0000;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
    end

    // state 2
    if (cycle == 1) begin
      PI_wbs_cyc_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b10000000000000000000000000000000;
      PI_wbs_we_i <= 1'b0;
      PI_wb_clk_i <= 1'b0;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b0;
      PI_wbs_sel_i <= 4'b1000;
      PI_wbs_addr_i <= 32'b00000000001000000000000000000000;
    end

    // state 3
    if (cycle == 2) begin
      PI_wbs_cyc_i <= 1'b1;
      PI_wb_rst_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
      PI_wbs_we_i <= 1'b0;
      PI_wb_clk_i <= 1'b1;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_sel_i <= 4'b0000;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
    end

    // state 4
    if (cycle == 3) begin
      PI_wbs_cyc_i <= 1'b1;
      PI_wb_rst_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000011111100;
      PI_wbs_we_i <= 1'b1;
      PI_wb_clk_i <= 1'b0;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_sel_i <= 4'b0001;
      PI_wbs_addr_i <= 32'b00110000110000000000000000000100;
    end

    // state 5
    if (cycle == 4) begin
      PI_wbs_cyc_i <= 1'b1;
      PI_wb_rst_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000011111100;
      PI_wbs_we_i <= 1'b1;
      PI_wb_clk_i <= 1'b1;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_sel_i <= 4'b0001;
      PI_wbs_addr_i <= 32'b00110000110000000000000000000100;
    end

    // state 6
    if (cycle == 5) begin
      PI_wbs_cyc_i <= 1'b1;
      PI_wb_rst_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000011111100;
      PI_wbs_we_i <= 1'b1;
      PI_wb_clk_i <= 1'b0;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_sel_i <= 4'b0001;
      PI_wbs_addr_i <= 32'b00110000110000000000000000000100;
    end

    // state 7
    if (cycle == 6) begin
      PI_wbs_cyc_i <= 1'b1;
      PI_wb_rst_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000011111100;
      PI_wbs_we_i <= 1'b1;
      PI_wb_clk_i <= 1'b1;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b0;
      PI_wbs_sel_i <= 4'b0001;
      PI_wbs_addr_i <= 32'b00110000110000000000000000000100;
    end

    // state 8
    if (cycle == 7) begin
      PI_wbs_cyc_i <= 1'b1;
      PI_wb_rst_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000011111100;
      PI_wbs_we_i <= 1'b1;
      PI_wb_clk_i <= 1'b0;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b0;
      PI_wbs_sel_i <= 4'b0001;
      PI_wbs_addr_i <= 32'b00110000110000000000000000000100;
    end

    // state 9
    if (cycle == 8) begin
      PI_wbs_cyc_i <= 1'b1;
      PI_wb_rst_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000011111100;
      PI_wbs_we_i <= 1'b0;
      PI_wb_clk_i <= 1'b1;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_sel_i <= 4'b0001;
      PI_wbs_addr_i <= 32'b00110000100000000000000000000000;
    end

    // state 10
    if (cycle == 9) begin
      PI_wbs_cyc_i <= 1'b1;
      PI_wb_rst_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000011111100;
      PI_wbs_we_i <= 1'b0;
      PI_wb_clk_i <= 1'b0;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_sel_i <= 4'b0000;
      PI_wbs_addr_i <= 32'b00110000100000000000000000000000;
    end

    // state 11
    if (cycle == 10) begin
      PI_wbs_cyc_i <= 1'b1;
      PI_wb_rst_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000011111100;
      PI_wbs_we_i <= 1'b0;
      PI_wb_clk_i <= 1'b1;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_sel_i <= 4'b0000;
      PI_wbs_addr_i <= 32'b00110000100000000000000000000000;
    end

    // state 12
    if (cycle == 11) begin
      PI_wbs_cyc_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
      PI_wbs_we_i <= 1'b0;
      PI_wb_clk_i <= 1'b0;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_stb_i <= 1'b0;
      PI_wbs_sel_i <= 4'b0000;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
    end

    genclock <= cycle < 12;
    cycle <= cycle + 1;
  end
endmodule
