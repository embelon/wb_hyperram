`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  reg [0:0] PI_hb_rwds_i;
  reg [0:0] PI_wb_rst_i;
  reg [31:0] PI_wbs_addr_i;
  reg [0:0] PI_wbs_stb_i;
  reg [3:0] PI_wbs_sel_i;
  reg [0:0] PI_wb_clk_i;
  reg [7:0] PI_hb_dq_i;
  reg [0:0] PI_rst_i;
  reg [0:0] PI_wbs_cyc_i;
  reg [0:0] PI_wbs_we_i;
  reg [31:0] PI_wbs_dat_i;
  wb_hyperram UUT (
    .hb_rwds_i(PI_hb_rwds_i),
    .wb_rst_i(PI_wb_rst_i),
    .wbs_addr_i(PI_wbs_addr_i),
    .wbs_stb_i(PI_wbs_stb_i),
    .wbs_sel_i(PI_wbs_sel_i),
    .wb_clk_i(PI_wb_clk_i),
    .hb_dq_i(PI_hb_dq_i),
    .rst_i(PI_rst_i),
    .wbs_cyc_i(PI_wbs_cyc_i),
    .wbs_we_i(PI_wbs_we_i),
    .wbs_dat_i(PI_wbs_dat_i)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    // UUT.$and$wb_hyperram.\v:0$463_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$472_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$476_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$494_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$507_Y  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:156:execute$4812  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:156:execute$4822  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:156:execute$4832  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:168:execute$4814  = 1'b1;
    // UUT.$auto$clk2fflogic.\cc:192:execute$4818  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:192:execute$4828  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:192:execute$4838  = 1'b0;
    // UUT.$eq$wb_hyperram.\v:434$654_Y  = 1'b0;
    // UUT.$eq$wb_hyperram.\v:543$796_Y  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:269$128_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:269$128_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:271$129_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:271$129_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:275$130_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:275$130_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:280$131_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:280$131_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:282$132_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:282$132_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:287$133_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:287$133_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:289$134_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:289$134_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:321$135_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:321$135_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:322$136_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:326$137_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:326$137_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:327$138_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:328$139_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:329$140_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:330$141_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:331$142_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:335$143_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:335$143_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:336$144_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:337$145_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:338$146_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:339$147_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:348$148_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:349$149_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:350$150_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:351$151_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:355$152_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:358$153_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:361$154_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:364$155_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:369$156_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:385$157_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:399$158_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:414$159_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:428$160_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:444$161_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:460$162_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:473$163_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:489$164_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:509$165_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:523$166_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:523$166_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:530$167_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:530$167_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:532$168_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:532$168_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:534$169_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:534$169_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:536$170_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:536$170_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:538$171_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:538$171_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:545$172_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:545$172_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:547$173_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:547$173_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:549$174_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:549$174_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:551$175_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:551$175_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:558$176_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:558$176_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:560$177_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:560$177_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:566$178_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:566$178_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:568$179_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:568$179_EN  = 1'b0;
    // UUT.$past$wb_hyperram.\v:329$17$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:330$18$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:331$19$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:332$20$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:348$25$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:349$26$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:350$28$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:373$30$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:374$31$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:380$36$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:380$37$0  = 6'b000000;
    // UUT.$past$wb_hyperram.\v:389$40$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:392$42$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:403$48$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:406$50$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:407$51$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:418$58$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:421$60$0  = 5'b00000;
    // UUT.$past$wb_hyperram.\v:446$72$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:447$73$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:453$77$0  = 3'b000;
    // UUT.$past$wb_hyperram.\v:491$91$0  = 1'b0;
    UUT.f_past_valid = 1'b0;
    // UUT.hram.$and$hyperram.\v:0$1487_Y  = 1'b0;
    // UUT.hram.$and$hyperram.\v:0$1496_Y  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4612  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4622  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4632  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4642  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4652  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4662  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4672  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4682  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4692  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4702  = 5'b00000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4712  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4722  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4732  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4742  = 48'b000000000000000000000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4752  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4762  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4772  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4782  = 3'b010;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4792  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4802  = 6'b100000;
    // UUT.hram.$auto$clk2fflogic.\cc:168:execute$4614  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:168:execute$4664  = 1'b1;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4618  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4628  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4638  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4648  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4658  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4668  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4678  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4688  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4698  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4708  = 5'b00000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4718  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4728  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4738  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4748  = 48'b000000000000000000000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4758  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4768  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4778  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4788  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4798  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4808  = 6'b000000;
    // UUT.hram.$formal$hyperram.\v:1001$1129_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1001$1129_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1005$1130_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1005$1130_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1007$1131_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1007$1131_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1011$1132_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1011$1132_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1013$1133_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1013$1133_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1015$1134_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1015$1134_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1019$1135_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1019$1135_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1022$1136_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1022$1136_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1025$1137_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1025$1137_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1030$1138_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1033$1139_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1033$1139_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1036$1140_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1036$1140_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1039$1141_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1039$1141_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1042$1142_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1042$1142_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1047$1143_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1051$1144_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1051$1144_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1053$1145_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1053$1145_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1057$1146_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1057$1146_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1065$1148_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1065$1148_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1070$1149_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1070$1149_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1073$1150_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1073$1150_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1074$1151_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1074$1151_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1075$1152_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1075$1152_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1076$1153_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1076$1153_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1084$1154_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1084$1154_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1085$1155_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1086$1156_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1087$1157_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:402$1086_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:402$1086_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:405$1087_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:405$1087_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:854$1088_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:854$1088_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:860$1089_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:861$1090_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:867$1091_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:867$1091_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:868$1092_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:869$1093_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:872$1094_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:872$1094_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:874$1095_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:874$1095_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:877$1096_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:877$1096_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:879$1097_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:879$1097_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:879$1098_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:881$1099_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:889$1100_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:889$1100_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:891$1101_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:891$1101_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:893$1102_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:893$1102_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:907$1103_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:907$1103_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:923$1104_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:923$1104_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:925$1105_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:925$1105_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:929$1106_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:929$1106_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:931$1107_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:931$1107_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:937$1108_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:937$1108_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:939$1109_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:939$1109_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:944$1110_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:944$1110_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:945$1111_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:946$1112_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:947$1113_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:949$1114_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:949$1114_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:955$1115_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:955$1115_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:959$1116_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:959$1116_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:962$1117_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:962$1117_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:965$1118_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:965$1118_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:968$1119_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:968$1119_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:971$1120_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:971$1120_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:974$1121_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:974$1121_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:977$1122_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:977$1122_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:980$1123_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:980$1123_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:983$1124_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:983$1124_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:986$1125_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:986$1125_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:992$1126_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:992$1126_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:995$1127_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:995$1127_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:998$1128_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:998$1128_EN  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1032$1051$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1032$1052$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1064$1063$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1064$1064$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1069$1068$0  = 8'b00000000;
    // UUT.hram.$past$hyperram.\v:1084$1078$0  = 32'b00000000000000000000000000000000;
    // UUT.hram.$past$hyperram.\v:1085$1079$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:1086$1080$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1087$1081$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:867$1000$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:868$1001$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:869$1002$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:871$1003$0  = 5'b00000;
    // UUT.hram.$past$hyperram.\v:876$1005$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:881$1007$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:882$1008$0  = 1'b0;
    UUT.hram.f_past_valid = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4312  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4322  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4332  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4342  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4352  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4362  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4372  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4382  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4392  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4402  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4314  = 1'b1;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4318  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4328  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4338  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4348  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4368  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4378  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4388  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4398  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4408  = 6'b000000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4212  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4222  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4232  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4242  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4252  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4262  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4272  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4282  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4292  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4302  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4214  = 1'b1;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4218  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4228  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4238  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4248  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4268  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4278  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4288  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4298  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4308  = 4'b0000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4412  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4422  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4432  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4442  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4452  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4462  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4472  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4482  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4492  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4502  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4414  = 1'b1;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4418  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4428  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4438  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4448  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4468  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4478  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4488  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4498  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4508  = 8'b00000000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4512  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4522  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4532  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4542  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4552  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4562  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4572  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4582  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4592  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4602  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4514  = 1'b1;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4518  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4528  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4538  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4548  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4568  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4578  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4588  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4598  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4608  = 5'b00000;
    UUT.wb_state = 2'b00;

    // state 0
    PI_hb_rwds_i = 1'b0;
    PI_wb_rst_i = 1'b1;
    PI_wbs_addr_i = 32'b00000000000000000000000010000000;
    PI_wbs_stb_i = 1'b0;
    PI_wbs_sel_i = 4'b1000;
    PI_wb_clk_i = 1'b0;
    PI_hb_dq_i = 8'b00000000;
    PI_rst_i = 1'b1;
    PI_wbs_cyc_i = 1'b0;
    PI_wbs_we_i = 1'b0;
    PI_wbs_dat_i = 32'b10000000000000000000000000000000;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      PI_hb_rwds_i <= 1'b0;
      PI_wb_rst_i <= 1'b1;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
      PI_wbs_stb_i <= 1'b0;
      PI_wbs_sel_i <= 4'b0000;
      PI_wb_clk_i <= 1'b1;
      PI_hb_dq_i <= 8'b00000000;
      PI_rst_i <= 1'b1;
      PI_wbs_cyc_i <= 1'b0;
      PI_wbs_we_i <= 1'b0;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
    end

    // state 2
    if (cycle == 1) begin
      PI_hb_rwds_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_addr_i <= 32'b00000000000000000000000010000000;
      PI_wbs_stb_i <= 1'b0;
      PI_wbs_sel_i <= 4'b1000;
      PI_wb_clk_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_rst_i <= 1'b0;
      PI_wbs_cyc_i <= 1'b0;
      PI_wbs_we_i <= 1'b0;
      PI_wbs_dat_i <= 32'b10000000000000000000000000000000;
    end

    // state 3
    if (cycle == 2) begin
      PI_hb_rwds_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_sel_i <= 4'b0000;
      PI_wb_clk_i <= 1'b1;
      PI_hb_dq_i <= 8'b00000000;
      PI_rst_i <= 1'b0;
      PI_wbs_cyc_i <= 1'b1;
      PI_wbs_we_i <= 1'b0;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
    end

    // state 4
    if (cycle == 3) begin
      PI_hb_rwds_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_addr_i <= 32'b00110100000000100000000000000100;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_sel_i <= 4'b1001;
      PI_wb_clk_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_rst_i <= 1'b0;
      PI_wbs_cyc_i <= 1'b1;
      PI_wbs_we_i <= 1'b1;
      PI_wbs_dat_i <= 32'b00000000000000000000000000101101;
    end

    // state 5
    if (cycle == 4) begin
      PI_hb_rwds_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_addr_i <= 32'b00110100000000100000000000000100;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_sel_i <= 4'b1001;
      PI_wb_clk_i <= 1'b1;
      PI_hb_dq_i <= 8'b00000000;
      PI_rst_i <= 1'b0;
      PI_wbs_cyc_i <= 1'b1;
      PI_wbs_we_i <= 1'b1;
      PI_wbs_dat_i <= 32'b00000000000000000000000000101101;
    end

    // state 6
    if (cycle == 5) begin
      PI_hb_rwds_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
      PI_wbs_stb_i <= 1'b0;
      PI_wbs_sel_i <= 4'b0000;
      PI_wb_clk_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_rst_i <= 1'b0;
      PI_wbs_cyc_i <= 1'b0;
      PI_wbs_we_i <= 1'b0;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
    end

    genclock <= cycle < 6;
    cycle <= cycle + 1;
  end
endmodule
