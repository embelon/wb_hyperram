magic
tech sky130A
magscale 1 2
timestamp 1636528672
<< locali >>
rect 24225 40579 24259 40681
rect 21649 40375 21683 40477
rect 30941 39491 30975 43945
rect 31585 40987 31619 44081
rect 15393 35071 15427 35241
rect 19199 33949 19291 33983
rect 19257 33847 19291 33949
rect 11345 33371 11379 33473
rect 21005 31875 21039 31977
rect 17417 27319 17451 27421
rect 13829 26843 13863 27081
rect 18797 23511 18831 23681
rect 16313 20927 16347 21097
rect 12541 20315 12575 20485
rect 11713 19703 11747 20009
rect 21925 18275 21959 18377
rect 12633 17663 12667 17765
rect 12725 15351 12759 15521
rect 14749 11543 14783 11713
rect 27077 6103 27111 6273
<< viali >>
rect 6377 45577 6411 45611
rect 8033 45577 8067 45611
rect 16773 45577 16807 45611
rect 21097 45577 21131 45611
rect 30021 45577 30055 45611
rect 1593 45441 1627 45475
rect 2421 45441 2455 45475
rect 3801 45441 3835 45475
rect 5089 45441 5123 45475
rect 6561 45441 6595 45475
rect 7205 45441 7239 45475
rect 8217 45441 8251 45475
rect 8953 45441 8987 45475
rect 9229 45441 9263 45475
rect 10241 45441 10275 45475
rect 11529 45441 11563 45475
rect 12633 45441 12667 45475
rect 12909 45441 12943 45475
rect 13553 45441 13587 45475
rect 14657 45441 14691 45475
rect 15301 45441 15335 45475
rect 16957 45441 16991 45475
rect 17785 45441 17819 45475
rect 18429 45441 18463 45475
rect 19257 45441 19291 45475
rect 20637 45441 20671 45475
rect 21281 45441 21315 45475
rect 21833 45441 21867 45475
rect 23857 45441 23891 45475
rect 26157 45441 26191 45475
rect 27445 45441 27479 45475
rect 27721 45441 27755 45475
rect 28365 45441 28399 45475
rect 28549 45441 28583 45475
rect 29837 45441 29871 45475
rect 2697 45373 2731 45407
rect 4077 45373 4111 45407
rect 5365 45373 5399 45407
rect 15577 45373 15611 45407
rect 17233 45373 17267 45407
rect 18705 45373 18739 45407
rect 19349 45373 19383 45407
rect 22109 45373 22143 45407
rect 24409 45373 24443 45407
rect 24685 45373 24719 45407
rect 27537 45373 27571 45407
rect 12725 45305 12759 45339
rect 17877 45305 17911 45339
rect 18521 45305 18555 45339
rect 26341 45305 26375 45339
rect 27905 45305 27939 45339
rect 1409 45237 1443 45271
rect 7021 45237 7055 45271
rect 10425 45237 10459 45271
rect 11713 45237 11747 45271
rect 13369 45237 13403 45271
rect 14473 45237 14507 45271
rect 15117 45237 15151 45271
rect 15485 45237 15519 45271
rect 17141 45237 17175 45271
rect 18429 45237 18463 45271
rect 19257 45237 19291 45271
rect 19625 45237 19659 45271
rect 20453 45237 20487 45271
rect 23673 45237 23707 45271
rect 27445 45237 27479 45271
rect 28733 45237 28767 45271
rect 11897 45033 11931 45067
rect 15485 45033 15519 45067
rect 16589 45033 16623 45067
rect 17601 45033 17635 45067
rect 20729 45033 20763 45067
rect 28273 45033 28307 45067
rect 10517 44965 10551 44999
rect 12633 44965 12667 44999
rect 15945 44965 15979 44999
rect 18061 44965 18095 44999
rect 28457 44965 28491 44999
rect 15577 44897 15611 44931
rect 16681 44897 16715 44931
rect 17693 44897 17727 44931
rect 19717 44897 19751 44931
rect 22569 44897 22603 44931
rect 24409 44897 24443 44931
rect 2053 44829 2087 44863
rect 5089 44829 5123 44863
rect 7481 44829 7515 44863
rect 10333 44829 10367 44863
rect 12081 44829 12115 44863
rect 12817 44829 12851 44863
rect 13553 44829 13587 44863
rect 14749 44829 14783 44863
rect 14933 44829 14967 44863
rect 15025 44829 15059 44863
rect 15761 44829 15795 44863
rect 16589 44829 16623 44863
rect 16865 44829 16899 44863
rect 17877 44829 17911 44863
rect 18521 44829 18555 44863
rect 19901 44829 19935 44863
rect 20637 44829 20671 44863
rect 21005 44829 21039 44863
rect 21097 44829 21131 44863
rect 21917 44829 21951 44863
rect 22845 44829 22879 44863
rect 24685 44829 24719 44863
rect 25881 44829 25915 44863
rect 27905 44829 27939 44863
rect 29837 44829 29871 44863
rect 2421 44761 2455 44795
rect 15485 44761 15519 44795
rect 17601 44761 17635 44795
rect 26148 44761 26182 44795
rect 28273 44761 28307 44795
rect 5181 44693 5215 44727
rect 7297 44693 7331 44727
rect 13369 44693 13403 44727
rect 14565 44693 14599 44727
rect 17049 44693 17083 44727
rect 18613 44693 18647 44727
rect 20085 44693 20119 44727
rect 21281 44693 21315 44727
rect 21741 44693 21775 44727
rect 27261 44693 27295 44727
rect 30021 44693 30055 44727
rect 15945 44489 15979 44523
rect 17049 44489 17083 44523
rect 27353 44489 27387 44523
rect 28273 44489 28307 44523
rect 28457 44489 28491 44523
rect 30113 44489 30147 44523
rect 14933 44421 14967 44455
rect 17877 44421 17911 44455
rect 18061 44421 18095 44455
rect 22201 44421 22235 44455
rect 1593 44353 1627 44387
rect 2053 44353 2087 44387
rect 2237 44353 2271 44387
rect 13185 44353 13219 44387
rect 13461 44353 13495 44387
rect 14105 44353 14139 44387
rect 16129 44353 16163 44387
rect 18981 44353 19015 44387
rect 19533 44353 19567 44387
rect 20269 44353 20303 44387
rect 20729 44353 20763 44387
rect 21833 44353 21867 44387
rect 22017 44353 22051 44387
rect 22937 44353 22971 44387
rect 23848 44353 23882 44387
rect 25421 44353 25455 44387
rect 25697 44353 25731 44387
rect 27169 44353 27203 44387
rect 29561 44353 29595 44387
rect 29929 44353 29963 44387
rect 2605 44285 2639 44319
rect 15025 44285 15059 44319
rect 15209 44285 15243 44319
rect 17141 44285 17175 44319
rect 17325 44285 17359 44319
rect 19441 44285 19475 44319
rect 20545 44285 20579 44319
rect 23581 44285 23615 44319
rect 29469 44285 29503 44319
rect 1409 44217 1443 44251
rect 13277 44217 13311 44251
rect 19533 44217 19567 44251
rect 27905 44217 27939 44251
rect 13921 44149 13955 44183
rect 14565 44149 14599 44183
rect 16681 44149 16715 44183
rect 18153 44149 18187 44183
rect 20453 44149 20487 44183
rect 20913 44149 20947 44183
rect 23121 44149 23155 44183
rect 24961 44149 24995 44183
rect 28273 44149 28307 44183
rect 29837 44149 29871 44183
rect 31585 44081 31619 44115
rect 1409 43945 1443 43979
rect 19441 43945 19475 43979
rect 20453 43945 20487 43979
rect 20637 43945 20671 43979
rect 21097 43945 21131 43979
rect 22661 43945 22695 43979
rect 28273 43945 28307 43979
rect 30941 43945 30975 43979
rect 25145 43877 25179 43911
rect 30021 43877 30055 43911
rect 10885 43809 10919 43843
rect 11805 43809 11839 43843
rect 12173 43809 12207 43843
rect 15301 43809 15335 43843
rect 16313 43809 16347 43843
rect 16405 43809 16439 43843
rect 17417 43809 17451 43843
rect 19349 43809 19383 43843
rect 23489 43809 23523 43843
rect 24777 43809 24811 43843
rect 1593 43741 1627 43775
rect 11069 43741 11103 43775
rect 11989 43741 12023 43775
rect 13461 43741 13495 43775
rect 15117 43741 15151 43775
rect 17141 43741 17175 43775
rect 18429 43741 18463 43775
rect 19257 43741 19291 43775
rect 20361 43741 20395 43775
rect 20453 43741 20487 43775
rect 21097 43741 21131 43775
rect 21281 43741 21315 43775
rect 22477 43741 22511 43775
rect 23121 43741 23155 43775
rect 23305 43741 23339 43775
rect 23397 43741 23431 43775
rect 23673 43741 23707 43775
rect 24409 43741 24443 43775
rect 24581 43739 24615 43773
rect 24685 43741 24719 43775
rect 24961 43741 24995 43775
rect 25973 43741 26007 43775
rect 27905 43741 27939 43775
rect 29837 43741 29871 43775
rect 15025 43673 15059 43707
rect 20177 43673 20211 43707
rect 26240 43673 26274 43707
rect 11253 43605 11287 43639
rect 13277 43605 13311 43639
rect 14657 43605 14691 43639
rect 15853 43605 15887 43639
rect 16221 43605 16255 43639
rect 18613 43605 18647 43639
rect 19625 43605 19659 43639
rect 21465 43605 21499 43639
rect 23857 43605 23891 43639
rect 27353 43605 27387 43639
rect 28273 43605 28307 43639
rect 28457 43605 28491 43639
rect 13369 43401 13403 43435
rect 14197 43401 14231 43435
rect 15209 43401 15243 43435
rect 15301 43401 15335 43435
rect 16773 43401 16807 43435
rect 22937 43401 22971 43435
rect 24777 43401 24811 43435
rect 26249 43401 26283 43435
rect 29285 43401 29319 43435
rect 23664 43333 23698 43367
rect 28273 43333 28307 43367
rect 1593 43265 1627 43299
rect 13553 43265 13587 43299
rect 14381 43265 14415 43299
rect 16957 43265 16991 43299
rect 17693 43265 17727 43299
rect 18889 43265 18923 43299
rect 19625 43265 19659 43299
rect 20269 43265 20303 43299
rect 20453 43265 20487 43299
rect 21281 43265 21315 43299
rect 22293 43265 22327 43299
rect 22753 43265 22787 43299
rect 23397 43265 23431 43299
rect 25513 43265 25547 43299
rect 25697 43265 25731 43299
rect 25881 43265 25915 43299
rect 26065 43265 26099 43299
rect 26985 43265 27019 43299
rect 29101 43265 29135 43299
rect 29837 43265 29871 43299
rect 15393 43197 15427 43231
rect 17417 43197 17451 43231
rect 19165 43197 19199 43231
rect 25789 43197 25823 43231
rect 21097 43129 21131 43163
rect 27905 43129 27939 43163
rect 28457 43129 28491 43163
rect 1409 43061 1443 43095
rect 14841 43061 14875 43095
rect 18705 43061 18739 43095
rect 19073 43061 19107 43095
rect 19717 43061 19751 43095
rect 20453 43061 20487 43095
rect 20637 43061 20671 43095
rect 22109 43061 22143 43095
rect 27169 43061 27203 43095
rect 28273 43061 28307 43095
rect 30021 43061 30055 43095
rect 16405 42857 16439 42891
rect 16773 42857 16807 42891
rect 25053 42857 25087 42891
rect 10885 42721 10919 42755
rect 15485 42721 15519 42755
rect 15945 42721 15979 42755
rect 16865 42721 16899 42755
rect 17785 42721 17819 42755
rect 17969 42721 18003 42755
rect 11069 42653 11103 42687
rect 14749 42653 14783 42687
rect 14933 42653 14967 42687
rect 15025 42653 15059 42687
rect 15669 42653 15703 42687
rect 15853 42653 15887 42687
rect 16589 42653 16623 42687
rect 18705 42653 18739 42687
rect 19533 42653 19567 42687
rect 19625 42653 19659 42687
rect 20545 42653 20579 42687
rect 22753 42653 22787 42687
rect 23581 42653 23615 42687
rect 24869 42653 24903 42687
rect 25513 42653 25547 42687
rect 25697 42653 25731 42687
rect 25789 42653 25823 42687
rect 25881 42653 25915 42687
rect 26065 42653 26099 42687
rect 26249 42653 26283 42687
rect 26709 42653 26743 42687
rect 27353 42653 27387 42687
rect 28181 42653 28215 42687
rect 28825 42653 28859 42687
rect 29837 42653 29871 42687
rect 20812 42585 20846 42619
rect 11253 42517 11287 42551
rect 14565 42517 14599 42551
rect 17325 42517 17359 42551
rect 17693 42517 17727 42551
rect 18521 42517 18555 42551
rect 19809 42517 19843 42551
rect 21925 42517 21959 42551
rect 22937 42517 22971 42551
rect 23397 42517 23431 42551
rect 26893 42517 26927 42551
rect 27537 42517 27571 42551
rect 27997 42517 28031 42551
rect 28641 42517 28675 42551
rect 30021 42517 30055 42551
rect 18245 42313 18279 42347
rect 19165 42313 19199 42347
rect 21189 42313 21223 42347
rect 23857 42313 23891 42347
rect 25973 42313 26007 42347
rect 29101 42313 29135 42347
rect 15945 42245 15979 42279
rect 19625 42245 19659 42279
rect 27905 42245 27939 42279
rect 28917 42245 28951 42279
rect 15025 42177 15059 42211
rect 15209 42177 15243 42211
rect 15301 42177 15335 42211
rect 18429 42177 18463 42211
rect 19533 42177 19567 42211
rect 20453 42177 20487 42211
rect 20637 42177 20671 42211
rect 21097 42177 21131 42211
rect 21281 42177 21315 42211
rect 22017 42177 22051 42211
rect 23029 42177 23063 42211
rect 24041 42177 24075 42211
rect 25789 42177 25823 42211
rect 27537 42177 27571 42211
rect 28549 42177 28583 42211
rect 29837 42177 29871 42211
rect 16957 42109 16991 42143
rect 17233 42109 17267 42143
rect 18705 42109 18739 42143
rect 19809 42109 19843 42143
rect 24501 42109 24535 42143
rect 24777 42109 24811 42143
rect 21833 42041 21867 42075
rect 22845 42041 22879 42075
rect 28089 42041 28123 42075
rect 14841 41973 14875 42007
rect 16037 41973 16071 42007
rect 18613 41973 18647 42007
rect 27905 41973 27939 42007
rect 28917 41973 28951 42007
rect 30021 41973 30055 42007
rect 19073 41769 19107 41803
rect 23857 41769 23891 41803
rect 28825 41769 28859 41803
rect 29009 41769 29043 41803
rect 28457 41701 28491 41735
rect 14749 41633 14783 41667
rect 14933 41633 14967 41667
rect 16589 41633 16623 41667
rect 19717 41633 19751 41667
rect 20085 41633 20119 41667
rect 24961 41633 24995 41667
rect 14657 41565 14691 41599
rect 17233 41565 17267 41599
rect 17509 41565 17543 41599
rect 18889 41565 18923 41599
rect 19441 41565 19475 41599
rect 21925 41565 21959 41599
rect 23029 41565 23063 41599
rect 23673 41565 23707 41599
rect 24685 41565 24719 41599
rect 25973 41565 26007 41599
rect 27997 41565 28031 41599
rect 29837 41565 29871 41599
rect 16405 41497 16439 41531
rect 18705 41497 18739 41531
rect 20352 41497 20386 41531
rect 22201 41497 22235 41531
rect 26240 41497 26274 41531
rect 28825 41497 28859 41531
rect 14289 41429 14323 41463
rect 16037 41429 16071 41463
rect 16497 41429 16531 41463
rect 19257 41429 19291 41463
rect 21465 41429 21499 41463
rect 23213 41429 23247 41463
rect 27353 41429 27387 41463
rect 27813 41429 27847 41463
rect 30021 41429 30055 41463
rect 14841 41225 14875 41259
rect 16681 41225 16715 41259
rect 18153 41225 18187 41259
rect 26249 41225 26283 41259
rect 29377 41225 29411 41259
rect 18061 41157 18095 41191
rect 29193 41157 29227 41191
rect 1593 41089 1627 41123
rect 14749 41089 14783 41123
rect 15577 41089 15611 41123
rect 15669 41089 15703 41123
rect 16865 41089 16899 41123
rect 19257 41089 19291 41123
rect 22293 41089 22327 41123
rect 23756 41089 23790 41123
rect 25513 41089 25547 41123
rect 25685 41089 25719 41123
rect 25789 41089 25823 41123
rect 26065 41089 26099 41123
rect 27241 41089 27275 41123
rect 28825 41089 28859 41123
rect 29837 41089 29871 41123
rect 14933 41021 14967 41055
rect 17141 41021 17175 41055
rect 18337 41021 18371 41055
rect 19349 41021 19383 41055
rect 19441 41021 19475 41055
rect 20913 41021 20947 41055
rect 23489 41021 23523 41055
rect 25881 41021 25915 41055
rect 26985 41021 27019 41055
rect 20361 40953 20395 40987
rect 20821 40953 20855 40987
rect 22477 40953 22511 40987
rect 1409 40885 1443 40919
rect 14381 40885 14415 40919
rect 15577 40885 15611 40919
rect 15945 40885 15979 40919
rect 17049 40885 17083 40919
rect 17693 40885 17727 40919
rect 18889 40885 18923 40919
rect 20729 40885 20763 40919
rect 21189 40885 21223 40919
rect 24869 40885 24903 40919
rect 28365 40885 28399 40919
rect 29193 40885 29227 40919
rect 30021 40885 30055 40919
rect 18245 40681 18279 40715
rect 20269 40681 20303 40715
rect 21833 40681 21867 40715
rect 23765 40681 23799 40715
rect 24225 40681 24259 40715
rect 28825 40681 28859 40715
rect 16221 40613 16255 40647
rect 21005 40613 21039 40647
rect 23121 40613 23155 40647
rect 25789 40613 25823 40647
rect 28457 40613 28491 40647
rect 29009 40613 29043 40647
rect 15117 40545 15151 40579
rect 15301 40545 15335 40579
rect 16773 40545 16807 40579
rect 18613 40545 18647 40579
rect 24225 40545 24259 40579
rect 24409 40545 24443 40579
rect 18429 40477 18463 40511
rect 18705 40477 18739 40511
rect 19533 40477 19567 40511
rect 19809 40477 19843 40511
rect 20453 40477 20487 40511
rect 21189 40477 21223 40511
rect 21649 40477 21683 40511
rect 21741 40477 21775 40511
rect 22937 40477 22971 40511
rect 23581 40477 23615 40511
rect 26249 40477 26283 40511
rect 26893 40477 26927 40511
rect 27997 40477 28031 40511
rect 29837 40477 29871 40511
rect 15025 40409 15059 40443
rect 24676 40409 24710 40443
rect 28825 40409 28859 40443
rect 14657 40341 14691 40375
rect 16589 40341 16623 40375
rect 16681 40341 16715 40375
rect 19625 40341 19659 40375
rect 21649 40341 21683 40375
rect 26433 40341 26467 40375
rect 27077 40341 27111 40375
rect 27813 40341 27847 40375
rect 30021 40341 30055 40375
rect 14657 40137 14691 40171
rect 16681 40137 16715 40171
rect 21097 40137 21131 40171
rect 21925 40137 21959 40171
rect 22569 40137 22603 40171
rect 25237 40137 25271 40171
rect 25881 40137 25915 40171
rect 27169 40137 27203 40171
rect 12081 40001 12115 40035
rect 12265 40001 12299 40035
rect 14841 40001 14875 40035
rect 15117 40001 15151 40035
rect 16865 40001 16899 40035
rect 17141 40001 17175 40035
rect 19441 40001 19475 40035
rect 19625 40001 19659 40035
rect 19993 40001 20027 40035
rect 21281 40001 21315 40035
rect 22109 40001 22143 40035
rect 22753 40001 22787 40035
rect 23213 40001 23247 40035
rect 23857 40001 23891 40035
rect 24041 40001 24075 40035
rect 24409 40001 24443 40035
rect 24593 40001 24627 40035
rect 25053 40001 25087 40035
rect 25697 40001 25731 40035
rect 26985 40001 27019 40035
rect 28365 40001 28399 40035
rect 29009 40001 29043 40035
rect 29837 40001 29871 40035
rect 15025 39933 15059 39967
rect 17049 39933 17083 39967
rect 19717 39933 19751 39967
rect 19809 39933 19843 39967
rect 24133 39933 24167 39967
rect 24225 39933 24259 39967
rect 12449 39865 12483 39899
rect 23397 39865 23431 39899
rect 20177 39797 20211 39831
rect 28181 39797 28215 39831
rect 28825 39797 28859 39831
rect 30021 39797 30055 39831
rect 19625 39593 19659 39627
rect 22937 39593 22971 39627
rect 25145 39593 25179 39627
rect 29929 39593 29963 39627
rect 22109 39525 22143 39559
rect 30113 39525 30147 39559
rect 31585 40953 31619 40987
rect 17969 39457 18003 39491
rect 20269 39457 20303 39491
rect 23765 39457 23799 39491
rect 24777 39457 24811 39491
rect 26249 39457 26283 39491
rect 27445 39457 27479 39491
rect 30941 39457 30975 39491
rect 1593 39389 1627 39423
rect 15209 39389 15243 39423
rect 15393 39389 15427 39423
rect 15485 39389 15519 39423
rect 15623 39389 15657 39423
rect 15772 39389 15806 39423
rect 17693 39389 17727 39423
rect 17877 39389 17911 39423
rect 18061 39389 18095 39423
rect 18245 39389 18279 39423
rect 19809 39389 19843 39423
rect 22293 39389 22327 39423
rect 22753 39389 22787 39423
rect 23673 39389 23707 39423
rect 24409 39389 24443 39423
rect 24593 39389 24627 39423
rect 24685 39389 24719 39423
rect 24961 39389 24995 39423
rect 25881 39389 25915 39423
rect 26065 39389 26099 39423
rect 26157 39389 26191 39423
rect 26433 39389 26467 39423
rect 26617 39389 26651 39423
rect 27077 39389 27111 39423
rect 27261 39389 27295 39423
rect 27353 39389 27387 39423
rect 27629 39389 27663 39423
rect 28733 39389 28767 39423
rect 29561 39389 29595 39423
rect 20536 39321 20570 39355
rect 29929 39321 29963 39355
rect 1409 39253 1443 39287
rect 15945 39253 15979 39287
rect 18429 39253 18463 39287
rect 21649 39253 21683 39287
rect 27813 39253 27847 39287
rect 28917 39253 28951 39287
rect 16037 39049 16071 39083
rect 21097 39049 21131 39083
rect 22109 39049 22143 39083
rect 23029 39049 23063 39083
rect 23673 39049 23707 39083
rect 28549 39049 28583 39083
rect 29377 39049 29411 39083
rect 29561 39049 29595 39083
rect 18766 38981 18800 39015
rect 27436 38981 27470 39015
rect 12081 38913 12115 38947
rect 12265 38913 12299 38947
rect 14924 38913 14958 38947
rect 16681 38913 16715 38947
rect 16948 38913 16982 38947
rect 18521 38913 18555 38947
rect 20361 38913 20395 38947
rect 20545 38913 20579 38947
rect 20913 38913 20947 38947
rect 22293 38913 22327 38947
rect 23213 38913 23247 38947
rect 23857 38913 23891 38947
rect 24317 38913 24351 38947
rect 24501 38913 24535 38947
rect 24685 38913 24719 38947
rect 24869 38913 24903 38947
rect 25697 38913 25731 38947
rect 25881 38913 25915 38947
rect 25973 38913 26007 38947
rect 26249 38913 26283 38947
rect 27169 38913 27203 38947
rect 14657 38845 14691 38879
rect 20637 38845 20671 38879
rect 20729 38845 20763 38879
rect 24593 38845 24627 38879
rect 26065 38845 26099 38879
rect 29009 38777 29043 38811
rect 12449 38709 12483 38743
rect 18061 38709 18095 38743
rect 19901 38709 19935 38743
rect 25053 38709 25087 38743
rect 26433 38709 26467 38743
rect 29377 38709 29411 38743
rect 16865 38505 16899 38539
rect 26065 38505 26099 38539
rect 26709 38505 26743 38539
rect 28549 38505 28583 38539
rect 16405 38369 16439 38403
rect 16497 38369 16531 38403
rect 19809 38369 19843 38403
rect 27169 38369 27203 38403
rect 10149 38301 10183 38335
rect 14105 38301 14139 38335
rect 16129 38301 16163 38335
rect 16313 38301 16347 38335
rect 16681 38301 16715 38335
rect 17325 38301 17359 38335
rect 17969 38301 18003 38335
rect 18153 38301 18187 38335
rect 18245 38301 18279 38335
rect 18337 38301 18371 38335
rect 18521 38301 18555 38335
rect 21649 38301 21683 38335
rect 22661 38301 22695 38335
rect 23305 38301 23339 38335
rect 24685 38301 24719 38335
rect 24952 38301 24986 38335
rect 26525 38301 26559 38335
rect 27425 38301 27459 38335
rect 29837 38301 29871 38335
rect 10416 38233 10450 38267
rect 14372 38233 14406 38267
rect 20076 38233 20110 38267
rect 11529 38165 11563 38199
rect 15485 38165 15519 38199
rect 17417 38165 17451 38199
rect 18705 38165 18739 38199
rect 21189 38165 21223 38199
rect 21741 38165 21775 38199
rect 22845 38165 22879 38199
rect 23489 38165 23523 38199
rect 30021 38165 30055 38199
rect 22109 37961 22143 37995
rect 27169 37961 27203 37995
rect 29561 37961 29595 37995
rect 29377 37893 29411 37927
rect 10057 37825 10091 37859
rect 10241 37825 10275 37859
rect 10609 37825 10643 37859
rect 12265 37825 12299 37859
rect 12532 37825 12566 37859
rect 14749 37825 14783 37859
rect 14933 37825 14967 37859
rect 15301 37825 15335 37859
rect 15945 37825 15979 37859
rect 16681 37825 16715 37859
rect 17601 37825 17635 37859
rect 18245 37825 18279 37859
rect 18512 37825 18546 37859
rect 20085 37825 20119 37859
rect 20269 37825 20303 37859
rect 20637 37825 20671 37859
rect 21925 37825 21959 37859
rect 22569 37825 22603 37859
rect 22836 37825 22870 37859
rect 24777 37825 24811 37859
rect 25513 37825 25547 37859
rect 26985 37825 27019 37859
rect 27905 37825 27939 37859
rect 28549 37825 28583 37859
rect 10333 37757 10367 37791
rect 10425 37757 10459 37791
rect 15025 37757 15059 37791
rect 15117 37757 15151 37791
rect 15485 37757 15519 37791
rect 20361 37757 20395 37791
rect 20453 37757 20487 37791
rect 25237 37757 25271 37791
rect 29009 37757 29043 37791
rect 27721 37689 27755 37723
rect 10793 37621 10827 37655
rect 13645 37621 13679 37655
rect 16037 37621 16071 37655
rect 16773 37621 16807 37655
rect 17693 37621 17727 37655
rect 19625 37621 19659 37655
rect 20821 37621 20855 37655
rect 23949 37621 23983 37655
rect 24593 37621 24627 37655
rect 28365 37621 28399 37655
rect 29377 37621 29411 37655
rect 13185 37417 13219 37451
rect 23765 37417 23799 37451
rect 24593 37417 24627 37451
rect 28825 37417 28859 37451
rect 29929 37417 29963 37451
rect 16681 37349 16715 37383
rect 18429 37349 18463 37383
rect 29009 37349 29043 37383
rect 12817 37281 12851 37315
rect 15209 37281 15243 37315
rect 15669 37281 15703 37315
rect 19533 37281 19567 37315
rect 20637 37281 20671 37315
rect 23305 37281 23339 37315
rect 26985 37281 27019 37315
rect 28457 37281 28491 37315
rect 29561 37281 29595 37315
rect 1593 37213 1627 37247
rect 10425 37213 10459 37247
rect 10692 37213 10726 37247
rect 12449 37213 12483 37247
rect 12633 37213 12667 37247
rect 12725 37213 12759 37247
rect 13001 37213 13035 37247
rect 14933 37213 14967 37247
rect 15117 37213 15151 37247
rect 15301 37213 15335 37247
rect 15485 37213 15519 37247
rect 16497 37213 16531 37247
rect 17141 37213 17175 37247
rect 19257 37213 19291 37247
rect 23029 37213 23063 37247
rect 23201 37213 23235 37247
rect 23397 37213 23431 37247
rect 23581 37213 23615 37247
rect 24409 37213 24443 37247
rect 25329 37213 25363 37247
rect 25605 37213 25639 37247
rect 26617 37213 26651 37247
rect 26801 37213 26835 37247
rect 26887 37213 26921 37247
rect 27169 37213 27203 37247
rect 27813 37213 27847 37247
rect 18245 37145 18279 37179
rect 20904 37145 20938 37179
rect 29929 37145 29963 37179
rect 1409 37077 1443 37111
rect 11805 37077 11839 37111
rect 17233 37077 17267 37111
rect 22017 37077 22051 37111
rect 27353 37077 27387 37111
rect 27997 37077 28031 37111
rect 28825 37077 28859 37111
rect 30113 37077 30147 37111
rect 10609 36873 10643 36907
rect 28365 36873 28399 36907
rect 29653 36873 29687 36907
rect 23397 36805 23431 36839
rect 24102 36805 24136 36839
rect 26433 36805 26467 36839
rect 27230 36805 27264 36839
rect 29469 36805 29503 36839
rect 8677 36737 8711 36771
rect 8861 36737 8895 36771
rect 8953 36737 8987 36771
rect 9229 36737 9263 36771
rect 9873 36737 9907 36771
rect 10057 36737 10091 36771
rect 10425 36737 10459 36771
rect 11713 36737 11747 36771
rect 13645 36737 13679 36771
rect 14933 36737 14967 36771
rect 15209 36737 15243 36771
rect 17049 36737 17083 36771
rect 17233 36737 17267 36771
rect 17325 36737 17359 36771
rect 17601 36737 17635 36771
rect 18797 36737 18831 36771
rect 20361 36737 20395 36771
rect 22017 36737 22051 36771
rect 22661 36737 22695 36771
rect 22845 36737 22879 36771
rect 22937 36737 22971 36771
rect 23213 36737 23247 36771
rect 23857 36737 23891 36771
rect 25697 36737 25731 36771
rect 25881 36737 25915 36771
rect 25973 36737 26007 36771
rect 26249 36737 26283 36771
rect 9045 36669 9079 36703
rect 10149 36669 10183 36703
rect 10241 36669 10275 36703
rect 12357 36669 12391 36703
rect 12633 36669 12667 36703
rect 13921 36669 13955 36703
rect 17417 36669 17451 36703
rect 19073 36669 19107 36703
rect 20085 36669 20119 36703
rect 23029 36669 23063 36703
rect 26065 36669 26099 36703
rect 26985 36669 27019 36703
rect 25237 36601 25271 36635
rect 29101 36601 29135 36635
rect 9413 36533 9447 36567
rect 11805 36533 11839 36567
rect 17785 36533 17819 36567
rect 22201 36533 22235 36567
rect 29469 36533 29503 36567
rect 19717 36329 19751 36363
rect 28273 36329 28307 36363
rect 28917 36329 28951 36363
rect 22293 36261 22327 36295
rect 16865 36193 16899 36227
rect 20269 36193 20303 36227
rect 24685 36193 24719 36227
rect 25697 36193 25731 36227
rect 11069 36125 11103 36159
rect 12817 36125 12851 36159
rect 13001 36125 13035 36159
rect 13093 36125 13127 36159
rect 13185 36125 13219 36159
rect 13369 36125 13403 36159
rect 14565 36125 14599 36159
rect 17132 36125 17166 36159
rect 22109 36125 22143 36159
rect 23581 36125 23615 36159
rect 24593 36125 24627 36159
rect 25421 36125 25455 36159
rect 26893 36125 26927 36159
rect 28733 36125 28767 36159
rect 29837 36125 29871 36159
rect 10793 36057 10827 36091
rect 11161 36057 11195 36091
rect 11529 36057 11563 36091
rect 11897 36057 11931 36091
rect 14832 36057 14866 36091
rect 19625 36057 19659 36091
rect 20536 36057 20570 36091
rect 22937 36057 22971 36091
rect 27160 36057 27194 36091
rect 12081 35989 12115 36023
rect 13553 35989 13587 36023
rect 15945 35989 15979 36023
rect 18245 35989 18279 36023
rect 21649 35989 21683 36023
rect 23029 35989 23063 36023
rect 23765 35989 23799 36023
rect 30021 35989 30055 36023
rect 12449 35785 12483 35819
rect 25973 35785 26007 35819
rect 27813 35785 27847 35819
rect 29653 35785 29687 35819
rect 20168 35717 20202 35751
rect 29469 35717 29503 35751
rect 9045 35649 9079 35683
rect 9312 35649 9346 35683
rect 12081 35649 12115 35683
rect 12265 35649 12299 35683
rect 13001 35649 13035 35683
rect 15117 35649 15151 35683
rect 15301 35649 15335 35683
rect 15393 35649 15427 35683
rect 15669 35649 15703 35683
rect 16957 35649 16991 35683
rect 17969 35649 18003 35683
rect 18153 35649 18187 35683
rect 18613 35649 18647 35683
rect 19901 35649 19935 35683
rect 22569 35649 22603 35683
rect 23213 35649 23247 35683
rect 23949 35649 23983 35683
rect 24216 35649 24250 35683
rect 25789 35649 25823 35683
rect 26985 35649 27019 35683
rect 27629 35649 27663 35683
rect 28641 35649 28675 35683
rect 29101 35649 29135 35683
rect 13277 35581 13311 35615
rect 15485 35581 15519 35615
rect 15853 35581 15887 35615
rect 16681 35581 16715 35615
rect 18889 35581 18923 35615
rect 22753 35581 22787 35615
rect 25329 35513 25363 35547
rect 10425 35445 10459 35479
rect 14381 35445 14415 35479
rect 17969 35445 18003 35479
rect 21281 35445 21315 35479
rect 23397 35445 23431 35479
rect 27169 35445 27203 35479
rect 28457 35445 28491 35479
rect 29469 35445 29503 35479
rect 12449 35241 12483 35275
rect 14657 35241 14691 35275
rect 15393 35241 15427 35275
rect 16865 35241 16899 35275
rect 18613 35241 18647 35275
rect 21925 35241 21959 35275
rect 23397 35241 23431 35275
rect 25145 35241 25179 35275
rect 26617 35241 26651 35275
rect 29929 35241 29963 35275
rect 30113 35241 30147 35275
rect 17877 35173 17911 35207
rect 21281 35173 21315 35207
rect 25789 35173 25823 35207
rect 28089 35173 28123 35207
rect 29561 35173 29595 35207
rect 20821 35105 20855 35139
rect 24685 35105 24719 35139
rect 1593 35037 1627 35071
rect 10885 35037 10919 35071
rect 12081 35037 12115 35071
rect 12265 35037 12299 35071
rect 13369 35037 13403 35071
rect 15393 35037 15427 35071
rect 15485 35037 15519 35071
rect 17450 35037 17484 35071
rect 17969 35037 18003 35071
rect 19257 35037 19291 35071
rect 19533 35037 19567 35071
rect 20545 35037 20579 35071
rect 20729 35037 20763 35071
rect 20913 35037 20947 35071
rect 21097 35037 21131 35071
rect 22661 35037 22695 35071
rect 23305 35037 23339 35071
rect 24409 35037 24443 35071
rect 24593 35037 24627 35071
rect 24777 35037 24811 35071
rect 24961 35037 24995 35071
rect 25973 35037 26007 35071
rect 26433 35037 26467 35071
rect 27629 35037 27663 35071
rect 28273 35037 28307 35071
rect 28733 35037 28767 35071
rect 14565 34969 14599 35003
rect 15730 34969 15764 35003
rect 18521 34969 18555 35003
rect 21833 34969 21867 35003
rect 1409 34901 1443 34935
rect 11069 34901 11103 34935
rect 13461 34901 13495 34935
rect 17325 34901 17359 34935
rect 17509 34901 17543 34935
rect 22753 34901 22787 34935
rect 27445 34901 27479 34935
rect 28917 34901 28951 34935
rect 29929 34901 29963 34935
rect 10701 34697 10735 34731
rect 14841 34697 14875 34731
rect 17233 34697 17267 34731
rect 17417 34697 17451 34731
rect 21005 34697 21039 34731
rect 22569 34697 22603 34731
rect 24685 34697 24719 34731
rect 25329 34697 25363 34731
rect 28457 34697 28491 34731
rect 29561 34697 29595 34731
rect 13728 34629 13762 34663
rect 16037 34629 16071 34663
rect 20269 34629 20303 34663
rect 29377 34629 29411 34663
rect 10517 34561 10551 34595
rect 11796 34561 11830 34595
rect 13461 34561 13495 34595
rect 15301 34561 15335 34595
rect 15485 34561 15519 34595
rect 15577 34561 15611 34595
rect 15853 34561 15887 34595
rect 17358 34561 17392 34595
rect 17877 34561 17911 34595
rect 18337 34561 18371 34595
rect 18521 34561 18555 34595
rect 18613 34561 18647 34595
rect 18889 34561 18923 34595
rect 19073 34561 19107 34595
rect 19533 34561 19567 34595
rect 19717 34561 19751 34595
rect 19809 34561 19843 34595
rect 20068 34561 20102 34595
rect 20913 34561 20947 34595
rect 22385 34561 22419 34595
rect 23029 34561 23063 34595
rect 23857 34561 23891 34595
rect 24501 34561 24535 34595
rect 25145 34561 25179 34595
rect 25789 34561 25823 34595
rect 26985 34561 27019 34595
rect 27813 34561 27847 34595
rect 28273 34561 28307 34595
rect 29009 34561 29043 34595
rect 11529 34493 11563 34527
rect 15669 34493 15703 34527
rect 18705 34493 18739 34527
rect 19901 34493 19935 34527
rect 23121 34493 23155 34527
rect 24041 34425 24075 34459
rect 27629 34425 27663 34459
rect 12909 34357 12943 34391
rect 17785 34357 17819 34391
rect 25973 34357 26007 34391
rect 27169 34357 27203 34391
rect 29377 34357 29411 34391
rect 10977 34153 11011 34187
rect 13185 34153 13219 34187
rect 14841 34153 14875 34187
rect 24777 34153 24811 34187
rect 26617 34153 26651 34187
rect 29929 34153 29963 34187
rect 30113 34153 30147 34187
rect 11437 34085 11471 34119
rect 20729 34085 20763 34119
rect 29561 34085 29595 34119
rect 12081 34017 12115 34051
rect 12449 34017 12483 34051
rect 15393 34017 15427 34051
rect 18245 34017 18279 34051
rect 19717 34017 19751 34051
rect 21189 34017 21223 34051
rect 25237 34017 25271 34051
rect 27445 34017 27479 34051
rect 10149 33949 10183 33983
rect 10333 33949 10367 33983
rect 10793 33949 10827 33983
rect 11621 33949 11655 33983
rect 12265 33949 12299 33983
rect 14749 33949 14783 33983
rect 17325 33949 17359 33983
rect 17969 33949 18003 33983
rect 18153 33949 18187 33983
rect 18383 33949 18417 33983
rect 18521 33949 18555 33983
rect 19165 33949 19199 33983
rect 19349 33949 19383 33983
rect 19533 33949 19567 33983
rect 19625 33949 19659 33983
rect 19901 33949 19935 33983
rect 20545 33949 20579 33983
rect 23029 33949 23063 33983
rect 24593 33949 24627 33983
rect 27077 33949 27111 33983
rect 27261 33949 27295 33983
rect 27353 33949 27387 33983
rect 27629 33949 27663 33983
rect 28733 33949 28767 33983
rect 13093 33881 13127 33915
rect 15660 33881 15694 33915
rect 21456 33881 21490 33915
rect 25504 33881 25538 33915
rect 29929 33881 29963 33915
rect 10241 33813 10275 33847
rect 16773 33813 16807 33847
rect 17417 33813 17451 33847
rect 18705 33813 18739 33847
rect 19257 33813 19291 33847
rect 20085 33813 20119 33847
rect 22569 33813 22603 33847
rect 23213 33813 23247 33847
rect 27813 33813 27847 33847
rect 28917 33813 28951 33847
rect 1409 33609 1443 33643
rect 11805 33609 11839 33643
rect 11897 33609 11931 33643
rect 12725 33609 12759 33643
rect 19349 33609 19383 33643
rect 21281 33609 21315 33643
rect 22293 33609 22327 33643
rect 26157 33609 26191 33643
rect 28641 33609 28675 33643
rect 11529 33541 11563 33575
rect 1593 33473 1627 33507
rect 10057 33473 10091 33507
rect 11345 33473 11379 33507
rect 11713 33473 11747 33507
rect 12081 33473 12115 33507
rect 12633 33473 12667 33507
rect 13277 33473 13311 33507
rect 13921 33473 13955 33507
rect 15025 33473 15059 33507
rect 15209 33473 15243 33507
rect 15393 33473 15427 33507
rect 15577 33473 15611 33507
rect 15761 33473 15795 33507
rect 16681 33473 16715 33507
rect 16865 33473 16899 33507
rect 17233 33473 17267 33507
rect 17969 33473 18003 33507
rect 18245 33473 18279 33507
rect 20545 33473 20579 33507
rect 20729 33473 20763 33507
rect 20821 33473 20855 33507
rect 21097 33473 21131 33507
rect 22109 33473 22143 33507
rect 22753 33473 22787 33507
rect 23009 33473 23043 33507
rect 24593 33473 24627 33507
rect 25421 33473 25455 33507
rect 25605 33473 25639 33507
rect 25697 33473 25731 33507
rect 25973 33473 26007 33507
rect 27261 33473 27295 33507
rect 27528 33473 27562 33507
rect 29101 33473 29135 33507
rect 29837 33473 29871 33507
rect 10149 33405 10183 33439
rect 10241 33405 10275 33439
rect 15301 33405 15335 33439
rect 16957 33405 16991 33439
rect 17049 33405 17083 33439
rect 20913 33405 20947 33439
rect 25789 33405 25823 33439
rect 11345 33337 11379 33371
rect 13461 33337 13495 33371
rect 9689 33269 9723 33303
rect 14105 33269 14139 33303
rect 17417 33269 17451 33303
rect 24133 33269 24167 33303
rect 24777 33269 24811 33303
rect 29285 33269 29319 33303
rect 30021 33269 30055 33303
rect 9965 33065 9999 33099
rect 17785 33065 17819 33099
rect 22017 33065 22051 33099
rect 26525 33065 26559 33099
rect 28641 33065 28675 33099
rect 9413 32997 9447 33031
rect 11161 32997 11195 33031
rect 19533 32929 19567 32963
rect 22477 32929 22511 32963
rect 25053 32929 25087 32963
rect 25329 32929 25363 32963
rect 27261 32929 27295 32963
rect 9321 32861 9355 32895
rect 9505 32861 9539 32895
rect 10149 32861 10183 32895
rect 10425 32861 10459 32895
rect 11713 32861 11747 32895
rect 12173 32861 12207 32895
rect 14197 32861 14231 32895
rect 16405 32861 16439 32895
rect 18245 32861 18279 32895
rect 19789 32861 19823 32895
rect 21833 32861 21867 32895
rect 24593 32861 24627 32895
rect 26341 32861 26375 32895
rect 29837 32861 29871 32895
rect 11345 32793 11379 32827
rect 12440 32793 12474 32827
rect 14464 32793 14498 32827
rect 16672 32793 16706 32827
rect 22744 32793 22778 32827
rect 27528 32793 27562 32827
rect 10333 32725 10367 32759
rect 11437 32725 11471 32759
rect 11529 32725 11563 32759
rect 13553 32725 13587 32759
rect 15577 32725 15611 32759
rect 18337 32725 18371 32759
rect 20913 32725 20947 32759
rect 23857 32725 23891 32759
rect 24409 32725 24443 32759
rect 30021 32725 30055 32759
rect 11713 32521 11747 32555
rect 13001 32521 13035 32555
rect 17233 32521 17267 32555
rect 21281 32521 21315 32555
rect 22845 32521 22879 32555
rect 23489 32521 23523 32555
rect 26433 32521 26467 32555
rect 29469 32521 29503 32555
rect 10241 32453 10275 32487
rect 27721 32453 27755 32487
rect 29285 32453 29319 32487
rect 11621 32385 11655 32419
rect 12265 32385 12299 32419
rect 12449 32385 12483 32419
rect 12633 32385 12667 32419
rect 12817 32385 12851 32419
rect 13553 32385 13587 32419
rect 14473 32385 14507 32419
rect 14657 32385 14691 32419
rect 15025 32385 15059 32419
rect 15209 32385 15243 32419
rect 15945 32385 15979 32419
rect 17141 32385 17175 32419
rect 17785 32385 17819 32419
rect 19257 32385 19291 32419
rect 19524 32385 19558 32419
rect 21097 32385 21131 32419
rect 22109 32385 22143 32419
rect 22293 32385 22327 32419
rect 22661 32385 22695 32419
rect 23305 32385 23339 32419
rect 24501 32385 24535 32419
rect 25605 32385 25639 32419
rect 26249 32385 26283 32419
rect 26985 32385 27019 32419
rect 27169 32385 27203 32419
rect 27353 32385 27387 32419
rect 27537 32385 27571 32419
rect 28457 32385 28491 32419
rect 30113 32385 30147 32419
rect 10333 32317 10367 32351
rect 10517 32317 10551 32351
rect 12541 32317 12575 32351
rect 14749 32317 14783 32351
rect 14841 32317 14875 32351
rect 16129 32317 16163 32351
rect 22385 32317 22419 32351
rect 22477 32317 22511 32351
rect 27261 32317 27295 32351
rect 20637 32249 20671 32283
rect 24961 32249 24995 32283
rect 28273 32249 28307 32283
rect 28917 32249 28951 32283
rect 9873 32181 9907 32215
rect 13553 32181 13587 32215
rect 17877 32181 17911 32215
rect 24777 32181 24811 32215
rect 25789 32181 25823 32215
rect 29285 32181 29319 32215
rect 29929 32181 29963 32215
rect 10149 31977 10183 32011
rect 11805 31977 11839 32011
rect 21005 31977 21039 32011
rect 23121 31977 23155 32011
rect 24685 31977 24719 32011
rect 24869 31977 24903 32011
rect 28181 31977 28215 32011
rect 10517 31909 10551 31943
rect 18613 31909 18647 31943
rect 23857 31909 23891 31943
rect 25973 31909 26007 31943
rect 28825 31909 28859 31943
rect 11161 31841 11195 31875
rect 12265 31841 12299 31875
rect 12449 31841 12483 31875
rect 16773 31841 16807 31875
rect 19993 31841 20027 31875
rect 21005 31841 21039 31875
rect 21097 31841 21131 31875
rect 21373 31841 21407 31875
rect 22661 31841 22695 31875
rect 26709 31841 26743 31875
rect 10333 31773 10367 31807
rect 10609 31773 10643 31807
rect 11069 31773 11103 31807
rect 15761 31773 15795 31807
rect 16405 31773 16439 31807
rect 16589 31773 16623 31807
rect 16681 31773 16715 31807
rect 16957 31773 16991 31807
rect 18429 31773 18463 31807
rect 19901 31773 19935 31807
rect 22385 31773 22419 31807
rect 22569 31773 22603 31807
rect 22753 31773 22787 31807
rect 22937 31773 22971 31807
rect 23673 31773 23707 31807
rect 24409 31773 24443 31807
rect 25789 31773 25823 31807
rect 26433 31773 26467 31807
rect 26617 31773 26651 31807
rect 26801 31773 26835 31807
rect 26985 31773 27019 31807
rect 28365 31773 28399 31807
rect 29009 31773 29043 31807
rect 29837 31773 29871 31807
rect 12173 31705 12207 31739
rect 15853 31637 15887 31671
rect 17141 31637 17175 31671
rect 27169 31637 27203 31671
rect 30021 31637 30055 31671
rect 10977 31433 11011 31467
rect 12817 31433 12851 31467
rect 15577 31433 15611 31467
rect 23213 31433 23247 31467
rect 28549 31433 28583 31467
rect 29561 31433 29595 31467
rect 15393 31365 15427 31399
rect 18981 31365 19015 31399
rect 19257 31365 19291 31399
rect 21097 31365 21131 31399
rect 27436 31365 27470 31399
rect 29377 31365 29411 31399
rect 1685 31297 1719 31331
rect 7941 31297 7975 31331
rect 8852 31297 8886 31331
rect 10609 31297 10643 31331
rect 11621 31297 11655 31331
rect 11805 31297 11839 31331
rect 12909 31297 12943 31331
rect 15209 31297 15243 31331
rect 17785 31297 17819 31331
rect 17969 31297 18003 31331
rect 18061 31297 18095 31331
rect 18337 31297 18371 31331
rect 19165 31297 19199 31331
rect 19354 31297 19388 31331
rect 20361 31297 20395 31331
rect 21833 31297 21867 31331
rect 22017 31297 22051 31331
rect 22109 31297 22143 31331
rect 22385 31297 22419 31331
rect 23029 31297 23063 31331
rect 27169 31297 27203 31331
rect 1409 31229 1443 31263
rect 8585 31229 8619 31263
rect 10701 31229 10735 31263
rect 12817 31229 12851 31263
rect 18153 31229 18187 31263
rect 22201 31229 22235 31263
rect 23949 31229 23983 31263
rect 24225 31229 24259 31263
rect 25421 31229 25455 31263
rect 25697 31229 25731 31263
rect 8125 31161 8159 31195
rect 9965 31161 9999 31195
rect 12357 31161 12391 31195
rect 18981 31161 19015 31195
rect 29009 31161 29043 31195
rect 10609 31093 10643 31127
rect 11621 31093 11655 31127
rect 18521 31093 18555 31127
rect 20545 31093 20579 31127
rect 21189 31093 21223 31127
rect 22569 31093 22603 31127
rect 29377 31093 29411 31127
rect 10701 30889 10735 30923
rect 18245 30889 18279 30923
rect 23765 30889 23799 30923
rect 25973 30889 26007 30923
rect 29929 30889 29963 30923
rect 30113 30889 30147 30923
rect 21741 30821 21775 30855
rect 11713 30753 11747 30787
rect 14105 30753 14139 30787
rect 17325 30753 17359 30787
rect 17417 30753 17451 30787
rect 19257 30753 19291 30787
rect 20361 30753 20395 30787
rect 22477 30753 22511 30787
rect 9873 30685 9907 30719
rect 11437 30685 11471 30719
rect 11529 30685 11563 30719
rect 12265 30685 12299 30719
rect 13093 30685 13127 30719
rect 14381 30685 14415 30719
rect 17049 30685 17083 30719
rect 17221 30679 17255 30713
rect 17601 30685 17635 30719
rect 18649 30685 18683 30719
rect 19630 30685 19664 30719
rect 20628 30685 20662 30719
rect 22201 30685 22235 30719
rect 22385 30685 22419 30719
rect 22569 30685 22603 30719
rect 22753 30685 22787 30719
rect 23581 30685 23615 30719
rect 24593 30685 24627 30719
rect 26433 30685 26467 30719
rect 27077 30685 27111 30719
rect 29561 30685 29595 30719
rect 10517 30617 10551 30651
rect 11713 30617 11747 30651
rect 12449 30617 12483 30651
rect 12909 30617 12943 30651
rect 18245 30617 18279 30651
rect 18429 30617 18463 30651
rect 18521 30617 18555 30651
rect 19257 30617 19291 30651
rect 19441 30617 19475 30651
rect 19533 30617 19567 30651
rect 24860 30617 24894 30651
rect 27344 30617 27378 30651
rect 9965 30549 9999 30583
rect 10717 30549 10751 30583
rect 10885 30549 10919 30583
rect 13277 30549 13311 30583
rect 15485 30549 15519 30583
rect 17785 30549 17819 30583
rect 22937 30549 22971 30583
rect 26617 30549 26651 30583
rect 28457 30549 28491 30583
rect 29929 30549 29963 30583
rect 8953 30345 8987 30379
rect 12725 30345 12759 30379
rect 25145 30345 25179 30379
rect 28365 30345 28399 30379
rect 9873 30277 9907 30311
rect 12265 30277 12299 30311
rect 13093 30277 13127 30311
rect 18981 30277 19015 30311
rect 22376 30277 22410 30311
rect 27721 30277 27755 30311
rect 8861 30209 8895 30243
rect 9045 30209 9079 30243
rect 10149 30209 10183 30243
rect 10333 30209 10367 30243
rect 10609 30209 10643 30243
rect 11529 30209 11563 30243
rect 11713 30209 11747 30243
rect 11897 30209 11931 30243
rect 12081 30209 12115 30243
rect 14473 30209 14507 30243
rect 14740 30209 14774 30243
rect 17049 30209 17083 30243
rect 17233 30209 17267 30243
rect 17325 30209 17359 30243
rect 17601 30209 17635 30243
rect 18245 30209 18279 30243
rect 18429 30209 18463 30243
rect 18797 30209 18831 30243
rect 19441 30209 19475 30243
rect 20729 30209 20763 30243
rect 24409 30209 24443 30243
rect 24593 30209 24627 30243
rect 24685 30209 24719 30243
rect 24961 30209 24995 30243
rect 26985 30209 27019 30243
rect 27169 30209 27203 30243
rect 27261 30209 27295 30243
rect 27537 30209 27571 30243
rect 28181 30209 28215 30243
rect 29377 30209 29411 30243
rect 29837 30209 29871 30243
rect 10425 30141 10459 30175
rect 11805 30141 11839 30175
rect 13185 30141 13219 30175
rect 13369 30141 13403 30175
rect 17417 30141 17451 30175
rect 18521 30141 18555 30175
rect 18613 30141 18647 30175
rect 22109 30141 22143 30175
rect 24777 30141 24811 30175
rect 25605 30141 25639 30175
rect 25881 30141 25915 30175
rect 27353 30141 27387 30175
rect 19625 30073 19659 30107
rect 29193 30073 29227 30107
rect 10241 30005 10275 30039
rect 15853 30005 15887 30039
rect 17785 30005 17819 30039
rect 20913 30005 20947 30039
rect 23489 30005 23523 30039
rect 30021 30005 30055 30039
rect 9413 29801 9447 29835
rect 13553 29801 13587 29835
rect 14933 29801 14967 29835
rect 15301 29801 15335 29835
rect 19717 29801 19751 29835
rect 21695 29801 21729 29835
rect 23121 29801 23155 29835
rect 28825 29801 28859 29835
rect 29009 29801 29043 29835
rect 30021 29801 30055 29835
rect 11897 29733 11931 29767
rect 9965 29665 9999 29699
rect 15393 29665 15427 29699
rect 16865 29665 16899 29699
rect 23857 29665 23891 29699
rect 25145 29665 25179 29699
rect 25237 29665 25271 29699
rect 8217 29597 8251 29631
rect 8401 29597 8435 29631
rect 9594 29597 9628 29631
rect 10057 29597 10091 29631
rect 10517 29597 10551 29631
rect 11161 29597 11195 29631
rect 11344 29597 11378 29631
rect 11434 29597 11468 29631
rect 11529 29597 11563 29631
rect 11713 29597 11747 29631
rect 12909 29597 12943 29631
rect 13002 29597 13036 29631
rect 13185 29597 13219 29631
rect 13415 29597 13449 29631
rect 14105 29597 14139 29631
rect 15117 29597 15151 29631
rect 15853 29597 15887 29631
rect 16037 29597 16071 29631
rect 16497 29597 16531 29631
rect 16653 29599 16687 29633
rect 16773 29597 16807 29631
rect 17049 29597 17083 29631
rect 17233 29597 17267 29631
rect 17969 29597 18003 29631
rect 19533 29597 19567 29631
rect 20177 29597 20211 29631
rect 20821 29597 20855 29631
rect 21465 29597 21499 29631
rect 22937 29597 22971 29631
rect 24869 29597 24903 29631
rect 25053 29597 25087 29631
rect 25421 29597 25455 29631
rect 26065 29597 26099 29631
rect 28457 29597 28491 29631
rect 29837 29597 29871 29631
rect 13277 29529 13311 29563
rect 14197 29529 14231 29563
rect 18061 29529 18095 29563
rect 23673 29529 23707 29563
rect 26310 29529 26344 29563
rect 28825 29529 28859 29563
rect 8309 29461 8343 29495
rect 9597 29461 9631 29495
rect 10609 29461 10643 29495
rect 15945 29461 15979 29495
rect 20361 29461 20395 29495
rect 20913 29461 20947 29495
rect 25605 29461 25639 29495
rect 27445 29461 27479 29495
rect 10333 29257 10367 29291
rect 12725 29257 12759 29291
rect 16129 29257 16163 29291
rect 16911 29257 16945 29291
rect 18981 29257 19015 29291
rect 20269 29257 20303 29291
rect 25513 29257 25547 29291
rect 26157 29257 26191 29291
rect 27169 29257 27203 29291
rect 29009 29257 29043 29291
rect 29193 29257 29227 29291
rect 14013 29189 14047 29223
rect 14197 29189 14231 29223
rect 15209 29189 15243 29223
rect 1409 29121 1443 29155
rect 7665 29121 7699 29155
rect 8565 29121 8599 29155
rect 10274 29121 10308 29155
rect 10701 29121 10735 29155
rect 10793 29121 10827 29155
rect 11529 29121 11563 29155
rect 11694 29121 11728 29155
rect 11805 29121 11839 29155
rect 12081 29121 12115 29155
rect 13093 29121 13127 29155
rect 14841 29121 14875 29155
rect 15025 29121 15059 29155
rect 15669 29121 15703 29155
rect 18153 29121 18187 29155
rect 18337 29121 18371 29155
rect 18797 29121 18831 29155
rect 19441 29121 19475 29155
rect 20085 29121 20119 29155
rect 20821 29121 20855 29155
rect 22017 29121 22051 29155
rect 22273 29121 22307 29155
rect 23857 29121 23891 29155
rect 24777 29121 24811 29155
rect 24961 29121 24995 29155
rect 25329 29121 25363 29155
rect 25973 29121 26007 29155
rect 26985 29121 27019 29155
rect 27629 29121 27663 29155
rect 28641 29121 28675 29155
rect 29837 29121 29871 29155
rect 8309 29053 8343 29087
rect 11897 29053 11931 29087
rect 13185 29053 13219 29087
rect 13369 29053 13403 29087
rect 16681 29053 16715 29087
rect 25053 29053 25087 29087
rect 25145 29053 25179 29087
rect 1593 28985 1627 29019
rect 10149 28985 10183 29019
rect 12265 28985 12299 29019
rect 18153 28985 18187 29019
rect 19625 28985 19659 29019
rect 21005 28985 21039 29019
rect 23397 28985 23431 29019
rect 24317 28985 24351 29019
rect 27813 28985 27847 29019
rect 30021 28985 30055 29019
rect 7849 28917 7883 28951
rect 9689 28917 9723 28951
rect 15761 28917 15795 28951
rect 23949 28917 23983 28951
rect 29009 28917 29043 28951
rect 8125 28713 8159 28747
rect 10701 28713 10735 28747
rect 10885 28713 10919 28747
rect 12909 28713 12943 28747
rect 22937 28713 22971 28747
rect 24869 28713 24903 28747
rect 27353 28713 27387 28747
rect 9965 28645 9999 28679
rect 15025 28645 15059 28679
rect 18245 28645 18279 28679
rect 23857 28645 23891 28679
rect 21741 28577 21775 28611
rect 7941 28509 7975 28543
rect 9873 28509 9907 28543
rect 12081 28509 12115 28543
rect 12817 28509 12851 28543
rect 14197 28509 14231 28543
rect 14841 28509 14875 28543
rect 15577 28509 15611 28543
rect 15853 28509 15887 28543
rect 16865 28509 16899 28543
rect 19257 28509 19291 28543
rect 21373 28509 21407 28543
rect 21557 28509 21591 28543
rect 21649 28509 21683 28543
rect 21925 28509 21959 28543
rect 22753 28509 22787 28543
rect 23673 28509 23707 28543
rect 24777 28509 24811 28543
rect 25973 28509 26007 28543
rect 29837 28509 29871 28543
rect 10517 28441 10551 28475
rect 11437 28441 11471 28475
rect 17132 28441 17166 28475
rect 19524 28441 19558 28475
rect 26240 28441 26274 28475
rect 10717 28373 10751 28407
rect 11529 28373 11563 28407
rect 12265 28373 12299 28407
rect 14289 28373 14323 28407
rect 20637 28373 20671 28407
rect 22109 28373 22143 28407
rect 23213 28373 23247 28407
rect 30021 28373 30055 28407
rect 17877 28169 17911 28203
rect 19441 28169 19475 28203
rect 25789 28169 25823 28203
rect 11805 28101 11839 28135
rect 14556 28101 14590 28135
rect 20269 28101 20303 28135
rect 7941 28033 7975 28067
rect 9505 28033 9539 28067
rect 12449 28033 12483 28067
rect 12716 28033 12750 28067
rect 14289 28033 14323 28067
rect 17141 28033 17175 28067
rect 17325 28033 17359 28067
rect 17417 28033 17451 28067
rect 17509 28033 17543 28067
rect 17693 28033 17727 28067
rect 18705 28033 18739 28067
rect 18877 28033 18911 28067
rect 19073 28033 19107 28067
rect 19257 28033 19291 28067
rect 21097 28033 21131 28067
rect 21833 28033 21867 28067
rect 22017 28033 22051 28067
rect 22103 28033 22137 28067
rect 22385 28033 22419 28067
rect 23121 28033 23155 28067
rect 24225 28033 24259 28067
rect 24685 28033 24719 28067
rect 24869 28033 24903 28067
rect 25605 28033 25639 28067
rect 29837 28033 29871 28067
rect 9597 27965 9631 27999
rect 10149 27965 10183 27999
rect 10425 27965 10459 27999
rect 18981 27965 19015 27999
rect 20361 27965 20395 27999
rect 20453 27965 20487 27999
rect 22201 27965 22235 27999
rect 24777 27965 24811 27999
rect 19901 27897 19935 27931
rect 22569 27897 22603 27931
rect 24041 27897 24075 27931
rect 8125 27829 8159 27863
rect 11897 27829 11931 27863
rect 13829 27829 13863 27863
rect 15669 27829 15703 27863
rect 21281 27829 21315 27863
rect 23213 27829 23247 27863
rect 23581 27829 23615 27863
rect 30021 27829 30055 27863
rect 16497 27625 16531 27659
rect 22569 27625 22603 27659
rect 11621 27557 11655 27591
rect 15071 27557 15105 27591
rect 15209 27557 15243 27591
rect 23213 27557 23247 27591
rect 26341 27557 26375 27591
rect 9781 27489 9815 27523
rect 10241 27489 10275 27523
rect 14473 27489 14507 27523
rect 15301 27489 15335 27523
rect 17785 27489 17819 27523
rect 17877 27489 17911 27523
rect 18245 27489 18279 27523
rect 20177 27489 20211 27523
rect 25789 27489 25823 27523
rect 1409 27421 1443 27455
rect 8033 27421 8067 27455
rect 10425 27421 10459 27455
rect 10793 27421 10827 27455
rect 12081 27421 12115 27455
rect 12449 27421 12483 27455
rect 12909 27421 12943 27455
rect 16129 27421 16163 27455
rect 16313 27421 16347 27455
rect 17417 27421 17451 27455
rect 17509 27421 17543 27455
rect 17693 27421 17727 27455
rect 18061 27421 18095 27455
rect 19257 27421 19291 27455
rect 19901 27421 19935 27455
rect 21189 27421 21223 27455
rect 23029 27421 23063 27455
rect 23857 27421 23891 27455
rect 24593 27421 24627 27455
rect 25053 27421 25087 27455
rect 25237 27421 25271 27455
rect 25697 27421 25731 27455
rect 25881 27421 25915 27455
rect 26341 27421 26375 27455
rect 26525 27421 26559 27455
rect 9597 27353 9631 27387
rect 11253 27353 11287 27387
rect 11437 27353 11471 27387
rect 12265 27353 12299 27387
rect 14289 27353 14323 27387
rect 14933 27353 14967 27387
rect 21456 27353 21490 27387
rect 1593 27285 1627 27319
rect 8217 27285 8251 27319
rect 10517 27285 10551 27319
rect 10609 27285 10643 27319
rect 13093 27285 13127 27319
rect 15577 27285 15611 27319
rect 17417 27285 17451 27319
rect 19441 27285 19475 27319
rect 23673 27285 23707 27319
rect 24409 27285 24443 27319
rect 25145 27285 25179 27319
rect 11805 27081 11839 27115
rect 11897 27081 11931 27115
rect 13277 27081 13311 27115
rect 13829 27081 13863 27115
rect 15025 27081 15059 27115
rect 18797 27081 18831 27115
rect 19165 27081 19199 27115
rect 22385 27081 22419 27115
rect 23581 27081 23615 27115
rect 23949 27081 23983 27115
rect 25329 27081 25363 27115
rect 26157 27081 26191 27115
rect 12081 27013 12115 27047
rect 9321 26945 9355 26979
rect 9413 26945 9447 26979
rect 10333 26945 10367 26979
rect 10425 26945 10459 26979
rect 11713 26945 11747 26979
rect 12541 26945 12575 26979
rect 13185 26945 13219 26979
rect 13369 26945 13403 26979
rect 9505 26877 9539 26911
rect 10517 26877 10551 26911
rect 10609 26877 10643 26911
rect 15761 27013 15795 27047
rect 17224 27013 17258 27047
rect 14105 26945 14139 26979
rect 14289 26945 14323 26979
rect 14381 26945 14415 26979
rect 14933 26945 14967 26979
rect 16957 26945 16991 26979
rect 20545 26945 20579 26979
rect 20729 26945 20763 26979
rect 20821 26945 20855 26979
rect 21097 26945 21131 26979
rect 22293 26945 22327 26979
rect 22937 26945 22971 26979
rect 24041 26945 24075 26979
rect 26341 26945 26375 26979
rect 29837 26945 29871 26979
rect 19257 26877 19291 26911
rect 19349 26877 19383 26911
rect 20913 26877 20947 26911
rect 24225 26877 24259 26911
rect 25421 26877 25455 26911
rect 25513 26877 25547 26911
rect 11529 26809 11563 26843
rect 12633 26809 12667 26843
rect 13829 26809 13863 26843
rect 14197 26809 14231 26843
rect 18337 26809 18371 26843
rect 23121 26809 23155 26843
rect 30021 26809 30055 26843
rect 8953 26741 8987 26775
rect 10149 26741 10183 26775
rect 13921 26741 13955 26775
rect 16037 26741 16071 26775
rect 21281 26741 21315 26775
rect 24961 26741 24995 26775
rect 10885 26537 10919 26571
rect 12817 26537 12851 26571
rect 14565 26537 14599 26571
rect 19993 26537 20027 26571
rect 21925 26537 21959 26571
rect 22661 26537 22695 26571
rect 24869 26537 24903 26571
rect 13093 26469 13127 26503
rect 15301 26469 15335 26503
rect 26249 26469 26283 26503
rect 10701 26401 10735 26435
rect 13277 26401 13311 26435
rect 14197 26401 14231 26435
rect 20545 26401 20579 26435
rect 22937 26401 22971 26435
rect 25513 26401 25547 26435
rect 9045 26333 9079 26367
rect 9321 26333 9355 26367
rect 10333 26333 10367 26367
rect 12173 26333 12207 26367
rect 13001 26333 13035 26367
rect 13185 26333 13219 26367
rect 13461 26333 13495 26367
rect 14381 26333 14415 26367
rect 14657 26333 14691 26367
rect 15485 26333 15519 26367
rect 15945 26333 15979 26367
rect 16773 26333 16807 26367
rect 18521 26333 18555 26367
rect 19901 26333 19935 26367
rect 22477 26333 22511 26367
rect 23581 26333 23615 26367
rect 25237 26333 25271 26367
rect 26065 26333 26099 26367
rect 29837 26333 29871 26367
rect 12265 26265 12299 26299
rect 16037 26265 16071 26299
rect 17509 26265 17543 26299
rect 18613 26265 18647 26299
rect 20812 26265 20846 26299
rect 25329 26265 25363 26299
rect 10517 26197 10551 26231
rect 23397 26197 23431 26231
rect 30021 26197 30055 26231
rect 1685 25993 1719 26027
rect 2329 25993 2363 26027
rect 11529 25993 11563 26027
rect 14197 25993 14231 26027
rect 17049 25993 17083 26027
rect 20453 25993 20487 26027
rect 21005 25993 21039 26027
rect 23397 25993 23431 26027
rect 24317 25993 24351 26027
rect 25237 25993 25271 26027
rect 9781 25925 9815 25959
rect 10793 25925 10827 25959
rect 14473 25925 14507 25959
rect 18889 25925 18923 25959
rect 20269 25925 20303 25959
rect 27445 25925 27479 25959
rect 1593 25857 1627 25891
rect 1777 25857 1811 25891
rect 2237 25857 2271 25891
rect 2421 25857 2455 25891
rect 9137 25857 9171 25891
rect 9321 25857 9355 25891
rect 10609 25857 10643 25891
rect 11897 25857 11931 25891
rect 13277 25857 13311 25891
rect 13461 25857 13495 25891
rect 13553 25857 13587 25891
rect 13737 25857 13771 25891
rect 14197 25857 14231 25891
rect 15761 25857 15795 25891
rect 17233 25857 17267 25891
rect 17325 25857 17359 25891
rect 17601 25857 17635 25891
rect 18061 25857 18095 25891
rect 19165 25857 19199 25891
rect 20085 25857 20119 25891
rect 20913 25857 20947 25891
rect 21097 25857 21131 25891
rect 22017 25857 22051 25891
rect 22937 25857 22971 25891
rect 25145 25857 25179 25891
rect 25329 25857 25363 25891
rect 29837 25857 29871 25891
rect 9045 25789 9079 25823
rect 11989 25789 12023 25823
rect 12081 25789 12115 25823
rect 15853 25789 15887 25823
rect 15945 25789 15979 25823
rect 18981 25789 19015 25823
rect 24409 25789 24443 25823
rect 24593 25789 24627 25823
rect 10977 25721 11011 25755
rect 13369 25721 13403 25755
rect 14289 25721 14323 25755
rect 18245 25721 18279 25755
rect 23949 25721 23983 25755
rect 27629 25721 27663 25755
rect 13093 25653 13127 25687
rect 15393 25653 15427 25687
rect 17509 25653 17543 25687
rect 18889 25653 18923 25687
rect 19349 25653 19383 25687
rect 22293 25653 22327 25687
rect 22477 25653 22511 25687
rect 23029 25653 23063 25687
rect 30021 25653 30055 25687
rect 9321 25449 9355 25483
rect 10793 25449 10827 25483
rect 13461 25449 13495 25483
rect 18705 25449 18739 25483
rect 19257 25449 19291 25483
rect 20453 25449 20487 25483
rect 23121 25449 23155 25483
rect 13231 25381 13265 25415
rect 29929 25381 29963 25415
rect 11345 25313 11379 25347
rect 13369 25313 13403 25347
rect 16405 25313 16439 25347
rect 16497 25313 16531 25347
rect 17601 25313 17635 25347
rect 19349 25313 19383 25347
rect 22109 25313 22143 25347
rect 23673 25313 23707 25347
rect 1409 25245 1443 25279
rect 11161 25245 11195 25279
rect 13093 25245 13127 25279
rect 13553 25245 13587 25279
rect 14105 25245 14139 25279
rect 17325 25245 17359 25279
rect 17417 25245 17451 25279
rect 17693 25245 17727 25279
rect 18337 25245 18371 25279
rect 19257 25245 19291 25279
rect 19533 25245 19567 25279
rect 22017 25245 22051 25279
rect 23489 25245 23523 25279
rect 24409 25245 24443 25279
rect 24593 25245 24627 25279
rect 29009 25245 29043 25279
rect 30113 25245 30147 25279
rect 8953 25177 8987 25211
rect 9137 25177 9171 25211
rect 10149 25177 10183 25211
rect 11989 25177 12023 25211
rect 12173 25177 12207 25211
rect 14350 25177 14384 25211
rect 17141 25177 17175 25211
rect 18521 25177 18555 25211
rect 20269 25177 20303 25211
rect 21189 25177 21223 25211
rect 21373 25177 21407 25211
rect 21557 25177 21591 25211
rect 26065 25177 26099 25211
rect 26249 25177 26283 25211
rect 26801 25177 26835 25211
rect 1593 25109 1627 25143
rect 10241 25109 10275 25143
rect 11253 25109 11287 25143
rect 12357 25109 12391 25143
rect 15485 25109 15519 25143
rect 15945 25109 15979 25143
rect 16313 25109 16347 25143
rect 19717 25109 19751 25143
rect 20453 25109 20487 25143
rect 20637 25109 20671 25143
rect 23581 25109 23615 25143
rect 24501 25109 24535 25143
rect 26893 25109 26927 25143
rect 28825 25109 28859 25143
rect 1685 24905 1719 24939
rect 12357 24905 12391 24939
rect 19441 24905 19475 24939
rect 8953 24837 8987 24871
rect 10793 24837 10827 24871
rect 11529 24837 11563 24871
rect 13737 24837 13771 24871
rect 14565 24837 14599 24871
rect 1593 24769 1627 24803
rect 1777 24769 1811 24803
rect 8309 24769 8343 24803
rect 9137 24769 9171 24803
rect 9781 24769 9815 24803
rect 9965 24769 9999 24803
rect 10609 24769 10643 24803
rect 11713 24769 11747 24803
rect 12541 24769 12575 24803
rect 13001 24769 13035 24803
rect 13645 24769 13679 24803
rect 14473 24769 14507 24803
rect 14657 24769 14691 24803
rect 15209 24769 15243 24803
rect 15853 24769 15887 24803
rect 16773 24769 16807 24803
rect 18245 24769 18279 24803
rect 19073 24769 19107 24803
rect 19165 24769 19199 24803
rect 20453 24769 20487 24803
rect 22661 24769 22695 24803
rect 23673 24769 23707 24803
rect 24685 24769 24719 24803
rect 25513 24769 25547 24803
rect 25697 24769 25731 24803
rect 28365 24769 28399 24803
rect 29009 24769 29043 24803
rect 29837 24769 29871 24803
rect 9321 24701 9355 24735
rect 17049 24701 17083 24735
rect 18521 24701 18555 24735
rect 20729 24701 20763 24735
rect 22753 24701 22787 24735
rect 22937 24701 22971 24735
rect 24777 24701 24811 24735
rect 24869 24701 24903 24735
rect 25605 24701 25639 24735
rect 8401 24633 8435 24667
rect 13093 24633 13127 24667
rect 15393 24633 15427 24667
rect 16037 24633 16071 24667
rect 24317 24633 24351 24667
rect 30021 24633 30055 24667
rect 10149 24565 10183 24599
rect 10885 24565 10919 24599
rect 11805 24565 11839 24599
rect 19073 24565 19107 24599
rect 22293 24565 22327 24599
rect 23489 24565 23523 24599
rect 28181 24565 28215 24599
rect 28825 24565 28859 24599
rect 10517 24361 10551 24395
rect 11529 24361 11563 24395
rect 12357 24361 12391 24395
rect 16037 24361 16071 24395
rect 22477 24361 22511 24395
rect 23121 24361 23155 24395
rect 24409 24361 24443 24395
rect 12541 24293 12575 24327
rect 19625 24293 19659 24327
rect 11713 24225 11747 24259
rect 15117 24225 15151 24259
rect 17509 24225 17543 24259
rect 23673 24225 23707 24259
rect 25329 24225 25363 24259
rect 25421 24225 25455 24259
rect 26985 24225 27019 24259
rect 8953 24157 8987 24191
rect 9137 24157 9171 24191
rect 9229 24157 9263 24191
rect 9367 24157 9401 24191
rect 9505 24157 9539 24191
rect 10517 24157 10551 24191
rect 10701 24157 10735 24191
rect 11437 24157 11471 24191
rect 12173 24157 12207 24191
rect 12357 24157 12391 24191
rect 13001 24157 13035 24191
rect 15025 24157 15059 24191
rect 16221 24157 16255 24191
rect 17233 24157 17267 24191
rect 17325 24157 17359 24191
rect 17601 24157 17635 24191
rect 19533 24157 19567 24191
rect 20821 24157 20855 24191
rect 21005 24157 21039 24191
rect 22661 24157 22695 24191
rect 23489 24157 23523 24191
rect 24593 24157 24627 24191
rect 25053 24157 25087 24191
rect 25237 24157 25271 24191
rect 25605 24157 25639 24191
rect 26617 24157 26651 24191
rect 26801 24157 26835 24191
rect 26893 24157 26927 24191
rect 27169 24157 27203 24191
rect 27813 24157 27847 24191
rect 29009 24157 29043 24191
rect 29837 24157 29871 24191
rect 17049 24089 17083 24123
rect 18337 24089 18371 24123
rect 21189 24089 21223 24123
rect 9689 24021 9723 24055
rect 10885 24021 10919 24055
rect 11713 24021 11747 24055
rect 13185 24021 13219 24055
rect 18429 24021 18463 24055
rect 23581 24021 23615 24055
rect 25789 24021 25823 24055
rect 27353 24021 27387 24055
rect 27905 24021 27939 24055
rect 28825 24021 28859 24055
rect 30021 24021 30055 24055
rect 8677 23817 8711 23851
rect 13001 23817 13035 23851
rect 24317 23817 24351 23851
rect 29285 23817 29319 23851
rect 11529 23749 11563 23783
rect 18153 23749 18187 23783
rect 22293 23749 22327 23783
rect 23029 23749 23063 23783
rect 7564 23681 7598 23715
rect 9137 23681 9171 23715
rect 9404 23681 9438 23715
rect 11989 23681 12023 23715
rect 12633 23681 12667 23715
rect 12909 23681 12943 23715
rect 13645 23681 13679 23715
rect 15025 23681 15059 23715
rect 16129 23681 16163 23715
rect 17141 23681 17175 23715
rect 17233 23681 17267 23715
rect 17509 23681 17543 23715
rect 17969 23681 18003 23715
rect 18797 23681 18831 23715
rect 18889 23681 18923 23715
rect 19901 23681 19935 23715
rect 20177 23681 20211 23715
rect 20269 23681 20303 23715
rect 22937 23681 22971 23715
rect 23121 23681 23155 23715
rect 24501 23681 24535 23715
rect 24961 23681 24995 23715
rect 25228 23681 25262 23715
rect 27445 23681 27479 23715
rect 27712 23681 27746 23715
rect 29469 23681 29503 23715
rect 30113 23681 30147 23715
rect 7297 23613 7331 23647
rect 11897 23613 11931 23647
rect 13001 23613 13035 23647
rect 15117 23613 15151 23647
rect 15209 23613 15243 23647
rect 12173 23545 12207 23579
rect 17417 23545 17451 23579
rect 19809 23613 19843 23647
rect 22477 23613 22511 23647
rect 10517 23477 10551 23511
rect 11989 23477 12023 23511
rect 12725 23477 12759 23511
rect 13645 23477 13679 23511
rect 14657 23477 14691 23511
rect 15945 23477 15979 23511
rect 16957 23477 16991 23511
rect 18337 23477 18371 23511
rect 18797 23477 18831 23511
rect 19073 23477 19107 23511
rect 19625 23477 19659 23511
rect 26341 23477 26375 23511
rect 28825 23477 28859 23511
rect 29929 23477 29963 23511
rect 8309 23273 8343 23307
rect 9689 23273 9723 23307
rect 11897 23273 11931 23307
rect 12357 23273 12391 23307
rect 20361 23273 20395 23307
rect 22017 23273 22051 23307
rect 24501 23273 24535 23307
rect 24869 23273 24903 23307
rect 25329 23273 25363 23307
rect 15945 23205 15979 23239
rect 19349 23205 19383 23239
rect 27537 23205 27571 23239
rect 9229 23137 9263 23171
rect 9321 23137 9355 23171
rect 10333 23137 10367 23171
rect 10609 23137 10643 23171
rect 12081 23137 12115 23171
rect 13369 23137 13403 23171
rect 14375 23137 14409 23171
rect 16497 23137 16531 23171
rect 17325 23137 17359 23171
rect 21557 23137 21591 23171
rect 21649 23137 21683 23171
rect 26157 23137 26191 23171
rect 28273 23137 28307 23171
rect 1409 23069 1443 23103
rect 2145 23069 2179 23103
rect 2329 23069 2363 23103
rect 8217 23069 8251 23103
rect 8953 23069 8987 23103
rect 9137 23069 9171 23103
rect 9505 23069 9539 23103
rect 11713 23069 11747 23103
rect 12173 23069 12207 23103
rect 13093 23069 13127 23103
rect 13466 23069 13500 23103
rect 14105 23069 14139 23103
rect 14289 23069 14323 23103
rect 14473 23069 14507 23103
rect 14657 23069 14691 23103
rect 16313 23069 16347 23103
rect 19257 23069 19291 23103
rect 20085 23069 20119 23103
rect 20177 23069 20211 23103
rect 20453 23069 20487 23103
rect 21281 23069 21315 23103
rect 21465 23069 21499 23103
rect 21833 23069 21867 23103
rect 22477 23069 22511 23103
rect 23673 23069 23707 23103
rect 24409 23069 24443 23103
rect 25513 23069 25547 23103
rect 26424 23069 26458 23103
rect 27997 23069 28031 23103
rect 29561 23069 29595 23103
rect 2237 23001 2271 23035
rect 13277 23001 13311 23035
rect 13369 23001 13403 23035
rect 16405 23001 16439 23035
rect 17592 23001 17626 23035
rect 19901 23001 19935 23035
rect 22569 23001 22603 23035
rect 1593 22933 1627 22967
rect 14841 22933 14875 22967
rect 18705 22933 18739 22967
rect 23765 22933 23799 22967
rect 29653 22933 29687 22967
rect 9689 22729 9723 22763
rect 11621 22729 11655 22763
rect 14013 22729 14047 22763
rect 14473 22729 14507 22763
rect 19717 22729 19751 22763
rect 24685 22729 24719 22763
rect 27997 22729 28031 22763
rect 8861 22661 8895 22695
rect 18429 22661 18463 22695
rect 21005 22661 21039 22695
rect 23765 22661 23799 22695
rect 8493 22593 8527 22627
rect 8585 22593 8619 22627
rect 8769 22593 8803 22627
rect 8953 22593 8987 22627
rect 9597 22593 9631 22627
rect 10517 22593 10551 22627
rect 10793 22593 10827 22627
rect 11529 22593 11563 22627
rect 12173 22593 12207 22627
rect 13369 22593 13403 22627
rect 14381 22593 14415 22627
rect 15209 22593 15243 22627
rect 15393 22593 15427 22627
rect 15485 22593 15519 22627
rect 15761 22593 15795 22627
rect 17049 22593 17083 22627
rect 17141 22593 17175 22627
rect 20821 22593 20855 22627
rect 21833 22593 21867 22627
rect 22100 22593 22134 22627
rect 24501 22593 24535 22627
rect 25329 22593 25363 22627
rect 26249 22593 26283 22627
rect 27261 22593 27295 22627
rect 27445 22593 27479 22627
rect 27813 22593 27847 22627
rect 28457 22593 28491 22627
rect 28724 22593 28758 22627
rect 14657 22525 14691 22559
rect 17233 22525 17267 22559
rect 25513 22525 25547 22559
rect 27537 22525 27571 22559
rect 27629 22525 27663 22559
rect 10701 22457 10735 22491
rect 15669 22457 15703 22491
rect 16681 22457 16715 22491
rect 23949 22457 23983 22491
rect 8493 22389 8527 22423
rect 10333 22389 10367 22423
rect 12265 22389 12299 22423
rect 13461 22389 13495 22423
rect 15577 22389 15611 22423
rect 21189 22389 21223 22423
rect 23213 22389 23247 22423
rect 26341 22389 26375 22423
rect 29837 22389 29871 22423
rect 8309 22185 8343 22219
rect 9505 22185 9539 22219
rect 23029 22185 23063 22219
rect 24501 22185 24535 22219
rect 24869 22185 24903 22219
rect 9873 22117 9907 22151
rect 21833 22117 21867 22151
rect 9781 22049 9815 22083
rect 15577 22049 15611 22083
rect 16681 22049 16715 22083
rect 16865 22049 16899 22083
rect 25697 22049 25731 22083
rect 25789 22049 25823 22083
rect 29009 22049 29043 22083
rect 29653 22049 29687 22083
rect 8217 21981 8251 22015
rect 9689 21981 9723 22015
rect 9965 21981 9999 22015
rect 10149 21981 10183 22015
rect 10885 21981 10919 22015
rect 10977 21981 11011 22015
rect 11069 21981 11103 22015
rect 11253 21981 11287 22015
rect 11897 21981 11931 22015
rect 12081 21981 12115 22015
rect 12173 21981 12207 22015
rect 12633 21981 12667 22015
rect 12725 21981 12759 22015
rect 15393 21981 15427 22015
rect 17969 21981 18003 22015
rect 18153 21981 18187 22015
rect 18245 21981 18279 22015
rect 18337 21981 18371 22015
rect 18521 21981 18555 22015
rect 19625 21981 19659 22015
rect 20453 21981 20487 22015
rect 22937 21981 22971 22015
rect 24409 21981 24443 22015
rect 25421 21981 25455 22015
rect 25605 21981 25639 22015
rect 25973 21981 26007 22015
rect 26709 21981 26743 22015
rect 26893 21981 26927 22015
rect 26979 21981 27013 22015
rect 27123 21981 27157 22015
rect 27261 21981 27295 22015
rect 28273 21981 28307 22015
rect 28457 21981 28491 22015
rect 28549 21981 28583 22015
rect 28641 21981 28675 22015
rect 28825 21981 28859 22015
rect 29561 21981 29595 22015
rect 10609 21913 10643 21947
rect 14105 21913 14139 21947
rect 14289 21913 14323 21947
rect 18705 21913 18739 21947
rect 20720 21913 20754 21947
rect 26157 21913 26191 21947
rect 11713 21845 11747 21879
rect 14473 21845 14507 21879
rect 15025 21845 15059 21879
rect 15485 21845 15519 21879
rect 16221 21845 16255 21879
rect 16589 21845 16623 21879
rect 19809 21845 19843 21879
rect 23397 21845 23431 21879
rect 27445 21845 27479 21879
rect 9137 21641 9171 21675
rect 13369 21641 13403 21675
rect 16865 21641 16899 21675
rect 21189 21641 21223 21675
rect 26249 21641 26283 21675
rect 2237 21573 2271 21607
rect 8024 21573 8058 21607
rect 14657 21573 14691 21607
rect 14841 21573 14875 21607
rect 19625 21573 19659 21607
rect 19809 21573 19843 21607
rect 20269 21573 20303 21607
rect 20453 21573 20487 21607
rect 20637 21573 20671 21607
rect 21833 21573 21867 21607
rect 26157 21573 26191 21607
rect 28273 21573 28307 21607
rect 28978 21573 29012 21607
rect 1409 21505 1443 21539
rect 2145 21505 2179 21539
rect 2329 21505 2363 21539
rect 7757 21505 7791 21539
rect 9965 21505 9999 21539
rect 10333 21505 10367 21539
rect 11794 21505 11828 21539
rect 14013 21505 14047 21539
rect 15485 21505 15519 21539
rect 16681 21505 16715 21539
rect 17693 21505 17727 21539
rect 17785 21505 17819 21539
rect 18061 21505 18095 21539
rect 18705 21505 18739 21539
rect 18797 21505 18831 21539
rect 19073 21505 19107 21539
rect 21097 21505 21131 21539
rect 22017 21505 22051 21539
rect 22661 21505 22695 21539
rect 22917 21505 22951 21539
rect 25053 21505 25087 21539
rect 27537 21505 27571 21539
rect 27721 21505 27755 21539
rect 27905 21505 27939 21539
rect 28089 21505 28123 21539
rect 28733 21505 28767 21539
rect 10057 21437 10091 21471
rect 12081 21437 12115 21471
rect 18521 21437 18555 21471
rect 18981 21437 19015 21471
rect 22201 21437 22235 21471
rect 24777 21437 24811 21471
rect 27813 21437 27847 21471
rect 9965 21369 9999 21403
rect 15577 21369 15611 21403
rect 1593 21301 1627 21335
rect 14105 21301 14139 21335
rect 14933 21301 14967 21335
rect 17509 21301 17543 21335
rect 17969 21301 18003 21335
rect 24041 21301 24075 21335
rect 30113 21301 30147 21335
rect 12173 21097 12207 21131
rect 14381 21097 14415 21131
rect 14749 21097 14783 21131
rect 16313 21097 16347 21131
rect 22661 21097 22695 21131
rect 23857 21097 23891 21131
rect 15669 21029 15703 21063
rect 11713 20961 11747 20995
rect 11805 20961 11839 20995
rect 25237 21029 25271 21063
rect 29929 21029 29963 21063
rect 23489 20961 23523 20995
rect 24869 20961 24903 20995
rect 25697 20961 25731 20995
rect 25973 20961 26007 20995
rect 27997 20961 28031 20995
rect 8953 20893 8987 20927
rect 9965 20893 9999 20927
rect 10609 20893 10643 20927
rect 10793 20893 10827 20927
rect 11437 20871 11471 20905
rect 11621 20893 11655 20927
rect 11989 20893 12023 20927
rect 12725 20893 12759 20927
rect 14381 20893 14415 20927
rect 14473 20893 14507 20927
rect 15485 20893 15519 20927
rect 16313 20893 16347 20927
rect 16497 20893 16531 20927
rect 17141 20893 17175 20927
rect 17417 20893 17451 20927
rect 18521 20893 18555 20927
rect 19441 20893 19475 20927
rect 20729 20893 20763 20927
rect 21373 20893 21407 20927
rect 22017 20893 22051 20927
rect 22165 20893 22199 20927
rect 22482 20893 22516 20927
rect 23121 20893 23155 20927
rect 23305 20893 23339 20927
rect 23397 20893 23431 20927
rect 23673 20893 23707 20927
rect 24501 20893 24535 20927
rect 24685 20893 24719 20927
rect 24777 20893 24811 20927
rect 25053 20893 25087 20927
rect 27353 20893 27387 20927
rect 28273 20893 28307 20927
rect 30113 20893 30147 20927
rect 10977 20825 11011 20859
rect 13001 20825 13035 20859
rect 15301 20825 15335 20859
rect 16681 20825 16715 20859
rect 18705 20825 18739 20859
rect 20545 20825 20579 20859
rect 20913 20825 20947 20859
rect 22293 20825 22327 20859
rect 22385 20825 22419 20859
rect 9137 20757 9171 20791
rect 10057 20757 10091 20791
rect 19625 20757 19659 20791
rect 21465 20757 21499 20791
rect 27445 20757 27479 20791
rect 8861 20553 8895 20587
rect 13001 20553 13035 20587
rect 19717 20553 19751 20587
rect 25237 20553 25271 20587
rect 26433 20553 26467 20587
rect 30113 20553 30147 20587
rect 9505 20485 9539 20519
rect 10241 20485 10275 20519
rect 10425 20485 10459 20519
rect 11713 20485 11747 20519
rect 11897 20485 11931 20519
rect 12081 20485 12115 20519
rect 12541 20485 12575 20519
rect 12817 20485 12851 20519
rect 15025 20485 15059 20519
rect 15669 20485 15703 20519
rect 17141 20485 17175 20519
rect 21281 20485 21315 20519
rect 23121 20485 23155 20519
rect 28273 20485 28307 20519
rect 28978 20485 29012 20519
rect 8677 20417 8711 20451
rect 12633 20417 12667 20451
rect 13829 20417 13863 20451
rect 14197 20417 14231 20451
rect 14381 20417 14415 20451
rect 14749 20417 14783 20451
rect 15485 20417 15519 20451
rect 17049 20417 17083 20451
rect 18337 20417 18371 20451
rect 18604 20417 18638 20451
rect 20545 20417 20579 20451
rect 20729 20417 20763 20451
rect 20821 20417 20855 20451
rect 20913 20417 20947 20451
rect 21080 20417 21114 20451
rect 21833 20417 21867 20451
rect 22017 20417 22051 20451
rect 22109 20417 22143 20451
rect 22385 20417 22419 20451
rect 23765 20417 23799 20451
rect 24501 20417 24535 20451
rect 24685 20417 24719 20451
rect 24777 20417 24811 20451
rect 25053 20417 25087 20451
rect 25697 20417 25731 20451
rect 25881 20417 25915 20451
rect 26249 20417 26283 20451
rect 27537 20417 27571 20451
rect 27725 20415 27759 20449
rect 27905 20417 27939 20451
rect 28089 20417 28123 20451
rect 28733 20417 28767 20451
rect 17233 20349 17267 20383
rect 22201 20349 22235 20383
rect 23857 20349 23891 20383
rect 24869 20349 24903 20383
rect 25973 20349 26007 20383
rect 26065 20349 26099 20383
rect 27813 20349 27847 20383
rect 12541 20281 12575 20315
rect 15853 20281 15887 20315
rect 22569 20281 22603 20315
rect 23305 20281 23339 20315
rect 9597 20213 9631 20247
rect 16681 20213 16715 20247
rect 11713 20009 11747 20043
rect 11805 20009 11839 20043
rect 12173 20009 12207 20043
rect 13369 20009 13403 20043
rect 14197 20009 14231 20043
rect 14565 20009 14599 20043
rect 19993 20009 20027 20043
rect 25789 20009 25823 20043
rect 28917 20009 28951 20043
rect 1593 19805 1627 19839
rect 1777 19805 1811 19839
rect 8953 19805 8987 19839
rect 9220 19737 9254 19771
rect 29653 19941 29687 19975
rect 11897 19873 11931 19907
rect 14197 19873 14231 19907
rect 15485 19873 15519 19907
rect 15577 19873 15611 19907
rect 16865 19873 16899 19907
rect 17877 19873 17911 19907
rect 23489 19873 23523 19907
rect 26801 19873 26835 19907
rect 11805 19805 11839 19839
rect 13185 19805 13219 19839
rect 13369 19805 13403 19839
rect 14381 19805 14415 19839
rect 16589 19805 16623 19839
rect 17601 19805 17635 19839
rect 17693 19805 17727 19839
rect 17969 19805 18003 19839
rect 19257 19805 19291 19839
rect 19441 19805 19475 19839
rect 19533 19805 19567 19839
rect 19625 19805 19659 19839
rect 19809 19805 19843 19839
rect 20545 19805 20579 19839
rect 21465 19805 21499 19839
rect 21613 19805 21647 19839
rect 21741 19805 21775 19839
rect 21971 19805 22005 19839
rect 23121 19805 23155 19839
rect 23305 19805 23339 19839
rect 23397 19805 23431 19839
rect 23673 19805 23707 19839
rect 24409 19805 24443 19839
rect 26433 19805 26467 19839
rect 26617 19805 26651 19839
rect 26709 19805 26743 19839
rect 26985 19805 27019 19839
rect 27629 19805 27663 19839
rect 27813 19805 27847 19839
rect 27905 19805 27939 19839
rect 27997 19805 28031 19839
rect 28181 19805 28215 19839
rect 28825 19805 28859 19839
rect 29561 19805 29595 19839
rect 14105 19737 14139 19771
rect 16681 19737 16715 19771
rect 20729 19737 20763 19771
rect 21833 19737 21867 19771
rect 23857 19737 23891 19771
rect 24654 19737 24688 19771
rect 27169 19737 27203 19771
rect 1685 19669 1719 19703
rect 10333 19669 10367 19703
rect 11713 19669 11747 19703
rect 13553 19669 13587 19703
rect 15025 19669 15059 19703
rect 15393 19669 15427 19703
rect 16221 19669 16255 19703
rect 17417 19669 17451 19703
rect 22109 19669 22143 19703
rect 28365 19669 28399 19703
rect 10333 19465 10367 19499
rect 13461 19465 13495 19499
rect 14841 19465 14875 19499
rect 25329 19465 25363 19499
rect 30113 19465 30147 19499
rect 9965 19397 9999 19431
rect 15577 19397 15611 19431
rect 16957 19397 16991 19431
rect 17969 19397 18003 19431
rect 1409 19329 1443 19363
rect 9689 19329 9723 19363
rect 9837 19329 9871 19363
rect 10057 19329 10091 19363
rect 10154 19329 10188 19363
rect 11989 19329 12023 19363
rect 12449 19329 12483 19363
rect 13093 19329 13127 19363
rect 13277 19329 13311 19363
rect 13921 19329 13955 19363
rect 14749 19329 14783 19363
rect 14933 19329 14967 19363
rect 15485 19329 15519 19363
rect 16681 19329 16715 19363
rect 17601 19329 17635 19363
rect 17749 19329 17783 19363
rect 17877 19329 17911 19363
rect 18066 19329 18100 19363
rect 19533 19329 19567 19363
rect 20821 19329 20855 19363
rect 21833 19329 21867 19363
rect 22100 19329 22134 19363
rect 24216 19329 24250 19363
rect 26249 19329 26283 19363
rect 27445 19329 27479 19363
rect 28733 19329 28767 19363
rect 29000 19329 29034 19363
rect 12357 19261 12391 19295
rect 21005 19261 21039 19295
rect 23949 19261 23983 19295
rect 27169 19261 27203 19295
rect 26433 19193 26467 19227
rect 1593 19125 1627 19159
rect 12633 19125 12667 19159
rect 18245 19125 18279 19159
rect 19717 19125 19751 19159
rect 23213 19125 23247 19159
rect 11253 18921 11287 18955
rect 15393 18921 15427 18955
rect 19993 18921 20027 18955
rect 23765 18921 23799 18955
rect 29929 18921 29963 18955
rect 21465 18853 21499 18887
rect 25881 18853 25915 18887
rect 12173 18785 12207 18819
rect 14381 18785 14415 18819
rect 16865 18785 16899 18819
rect 22385 18785 22419 18819
rect 22661 18785 22695 18819
rect 25513 18785 25547 18819
rect 9873 18717 9907 18751
rect 11805 18717 11839 18751
rect 11989 18717 12023 18751
rect 12081 18717 12115 18751
rect 12357 18717 12391 18751
rect 13369 18717 13403 18751
rect 13461 18717 13495 18751
rect 14105 18717 14139 18751
rect 14197 18717 14231 18751
rect 15209 18717 15243 18751
rect 15301 18717 15335 18751
rect 15485 18717 15519 18751
rect 15577 18717 15611 18751
rect 16589 18717 16623 18751
rect 17601 18717 17635 18751
rect 17749 18717 17783 18751
rect 18107 18717 18141 18751
rect 19533 18717 19567 18751
rect 20177 18717 20211 18751
rect 20729 18717 20763 18751
rect 21373 18717 21407 18751
rect 23673 18717 23707 18751
rect 25145 18717 25179 18751
rect 25329 18717 25363 18751
rect 25421 18717 25455 18751
rect 25697 18717 25731 18751
rect 26341 18717 26375 18751
rect 26617 18717 26651 18751
rect 27629 18717 27663 18751
rect 30113 18717 30147 18751
rect 10140 18649 10174 18683
rect 12541 18649 12575 18683
rect 17877 18649 17911 18683
rect 17969 18649 18003 18683
rect 24501 18649 24535 18683
rect 27896 18649 27930 18683
rect 14381 18581 14415 18615
rect 16221 18581 16255 18615
rect 16681 18581 16715 18615
rect 18245 18581 18279 18615
rect 19349 18581 19383 18615
rect 20821 18581 20855 18615
rect 24593 18581 24627 18615
rect 29009 18581 29043 18615
rect 13001 18377 13035 18411
rect 15485 18377 15519 18411
rect 16037 18377 16071 18411
rect 19073 18377 19107 18411
rect 21925 18377 21959 18411
rect 24133 18377 24167 18411
rect 29745 18377 29779 18411
rect 16681 18309 16715 18343
rect 7757 18241 7791 18275
rect 8024 18241 8058 18275
rect 11713 18241 11747 18275
rect 12265 18241 12299 18275
rect 13185 18241 13219 18275
rect 14749 18241 14783 18275
rect 14937 18239 14971 18273
rect 15025 18241 15059 18275
rect 15301 18241 15335 18275
rect 15945 18241 15979 18275
rect 16865 18241 16899 18275
rect 16957 18241 16991 18275
rect 17233 18241 17267 18275
rect 17693 18241 17727 18275
rect 17960 18241 17994 18275
rect 19800 18241 19834 18275
rect 21925 18241 21959 18275
rect 22017 18241 22051 18275
rect 22753 18241 22787 18275
rect 23397 18241 23431 18275
rect 23581 18241 23615 18275
rect 23949 18241 23983 18275
rect 25053 18241 25087 18275
rect 25320 18241 25354 18275
rect 27436 18241 27470 18275
rect 28997 18241 29031 18275
rect 29193 18241 29227 18275
rect 29561 18241 29595 18275
rect 15117 18173 15151 18207
rect 19533 18173 19567 18207
rect 23673 18173 23707 18207
rect 23765 18173 23799 18207
rect 27169 18173 27203 18207
rect 29285 18173 29319 18207
rect 29377 18173 29411 18207
rect 22937 18105 22971 18139
rect 26433 18105 26467 18139
rect 28549 18105 28583 18139
rect 9137 18037 9171 18071
rect 11529 18037 11563 18071
rect 12449 18037 12483 18071
rect 17141 18037 17175 18071
rect 20913 18037 20947 18071
rect 22109 18037 22143 18071
rect 8217 17833 8251 17867
rect 12725 17833 12759 17867
rect 15301 17833 15335 17867
rect 15853 17833 15887 17867
rect 20821 17833 20855 17867
rect 22385 17833 22419 17867
rect 23581 17833 23615 17867
rect 25605 17833 25639 17867
rect 26893 17833 26927 17867
rect 10057 17765 10091 17799
rect 12633 17765 12667 17799
rect 19533 17765 19567 17799
rect 11805 17697 11839 17731
rect 13369 17697 13403 17731
rect 14381 17697 14415 17731
rect 14473 17697 14507 17731
rect 16405 17697 16439 17731
rect 21925 17697 21959 17731
rect 23121 17697 23155 17731
rect 23213 17697 23247 17731
rect 26525 17697 26559 17731
rect 27537 17697 27571 17731
rect 27813 17697 27847 17731
rect 1593 17629 1627 17663
rect 1777 17629 1811 17663
rect 8401 17629 8435 17663
rect 9413 17629 9447 17663
rect 10701 17629 10735 17663
rect 10793 17629 10827 17663
rect 11621 17629 11655 17663
rect 11713 17629 11747 17663
rect 12633 17629 12667 17663
rect 14289 17629 14323 17663
rect 14565 17629 14599 17663
rect 15209 17629 15243 17663
rect 16221 17629 16255 17663
rect 17325 17629 17359 17663
rect 19717 17629 19751 17663
rect 20177 17629 20211 17663
rect 20270 17629 20304 17663
rect 20453 17629 20487 17663
rect 20661 17629 20695 17663
rect 21649 17629 21683 17663
rect 21833 17629 21867 17663
rect 22017 17629 22051 17663
rect 22201 17629 22235 17663
rect 22845 17629 22879 17663
rect 23033 17623 23067 17657
rect 23397 17629 23431 17663
rect 24409 17629 24443 17663
rect 25513 17629 25547 17663
rect 26157 17629 26191 17663
rect 26345 17629 26379 17663
rect 26433 17629 26467 17663
rect 26709 17629 26743 17663
rect 29009 17629 29043 17663
rect 30113 17629 30147 17663
rect 9689 17561 9723 17595
rect 9898 17561 9932 17595
rect 13093 17561 13127 17595
rect 17592 17561 17626 17595
rect 20553 17561 20587 17595
rect 1685 17493 1719 17527
rect 9781 17493 9815 17527
rect 11253 17493 11287 17527
rect 13185 17493 13219 17527
rect 14105 17493 14139 17527
rect 16313 17493 16347 17527
rect 18705 17493 18739 17527
rect 24501 17493 24535 17527
rect 28825 17493 28859 17527
rect 29929 17493 29963 17527
rect 11989 17289 12023 17323
rect 12449 17289 12483 17323
rect 13737 17289 13771 17323
rect 14197 17289 14231 17323
rect 15577 17289 15611 17323
rect 17141 17289 17175 17323
rect 17969 17289 18003 17323
rect 20729 17289 20763 17323
rect 25145 17289 25179 17323
rect 26341 17289 26375 17323
rect 28089 17289 28123 17323
rect 17049 17221 17083 17255
rect 21925 17221 21959 17255
rect 23305 17221 23339 17255
rect 24010 17221 24044 17255
rect 1409 17153 1443 17187
rect 2145 17153 2179 17187
rect 8769 17153 8803 17187
rect 12357 17153 12391 17187
rect 14105 17153 14139 17187
rect 14933 17153 14967 17187
rect 15761 17153 15795 17187
rect 15853 17153 15887 17187
rect 16129 17153 16163 17187
rect 17877 17153 17911 17187
rect 19441 17153 19475 17187
rect 20085 17153 20119 17187
rect 20913 17153 20947 17187
rect 21005 17153 21039 17187
rect 21281 17153 21315 17187
rect 21833 17153 21867 17187
rect 22569 17153 22603 17187
rect 22753 17153 22787 17187
rect 22845 17153 22879 17187
rect 23121 17153 23155 17187
rect 26249 17153 26283 17187
rect 27353 17153 27387 17187
rect 27537 17153 27571 17187
rect 27905 17153 27939 17187
rect 28641 17153 28675 17187
rect 28897 17153 28931 17187
rect 9045 17085 9079 17119
rect 12541 17085 12575 17119
rect 14289 17085 14323 17119
rect 17325 17085 17359 17119
rect 21189 17085 21223 17119
rect 22937 17085 22971 17119
rect 23765 17085 23799 17119
rect 27629 17085 27663 17119
rect 27721 17085 27755 17119
rect 16681 17017 16715 17051
rect 20177 17017 20211 17051
rect 1593 16949 1627 16983
rect 2237 16949 2271 16983
rect 10149 16949 10183 16983
rect 15025 16949 15059 16983
rect 16037 16949 16071 16983
rect 19533 16949 19567 16983
rect 30021 16949 30055 16983
rect 10425 16745 10459 16779
rect 13461 16745 13495 16779
rect 15669 16745 15703 16779
rect 23305 16745 23339 16779
rect 24409 16745 24443 16779
rect 26525 16745 26559 16779
rect 27813 16745 27847 16779
rect 29009 16745 29043 16779
rect 21097 16677 21131 16711
rect 9965 16609 9999 16643
rect 11345 16609 11379 16643
rect 11529 16609 11563 16643
rect 12081 16609 12115 16643
rect 12633 16609 12667 16643
rect 14565 16609 14599 16643
rect 14749 16609 14783 16643
rect 19257 16609 19291 16643
rect 21557 16609 21591 16643
rect 22845 16609 22879 16643
rect 22937 16609 22971 16643
rect 24869 16609 24903 16643
rect 27353 16609 27387 16643
rect 28641 16609 28675 16643
rect 9689 16541 9723 16575
rect 9873 16541 9907 16575
rect 10057 16541 10091 16575
rect 10241 16541 10275 16575
rect 11253 16541 11287 16575
rect 12265 16541 12299 16575
rect 13461 16541 13495 16575
rect 15301 16541 15335 16575
rect 21281 16541 21315 16575
rect 21373 16541 21407 16575
rect 21649 16541 21683 16575
rect 22569 16541 22603 16575
rect 22753 16541 22787 16575
rect 23121 16541 23155 16575
rect 24593 16541 24627 16575
rect 24685 16541 24719 16575
rect 24961 16541 24995 16575
rect 25697 16541 25731 16575
rect 26341 16541 26375 16575
rect 27077 16541 27111 16575
rect 27261 16541 27295 16575
rect 27445 16541 27479 16575
rect 27629 16541 27663 16575
rect 28273 16541 28307 16575
rect 28457 16541 28491 16575
rect 28549 16541 28583 16575
rect 28825 16541 28859 16575
rect 29561 16541 29595 16575
rect 15485 16473 15519 16507
rect 19524 16473 19558 16507
rect 25789 16473 25823 16507
rect 10885 16405 10919 16439
rect 12265 16405 12299 16439
rect 14105 16405 14139 16439
rect 14473 16405 14507 16439
rect 20637 16405 20671 16439
rect 29653 16405 29687 16439
rect 12081 16201 12115 16235
rect 15393 16201 15427 16235
rect 15761 16201 15795 16235
rect 17049 16201 17083 16235
rect 19533 16201 19567 16235
rect 21833 16201 21867 16235
rect 23121 16201 23155 16235
rect 24317 16201 24351 16235
rect 17969 16133 18003 16167
rect 21097 16133 21131 16167
rect 28978 16133 29012 16167
rect 10609 16065 10643 16099
rect 10701 16065 10735 16099
rect 10977 16065 11011 16099
rect 12449 16065 12483 16099
rect 12541 16065 12575 16099
rect 13645 16065 13679 16099
rect 13829 16065 13863 16099
rect 13921 16065 13955 16099
rect 14197 16065 14231 16099
rect 15853 16065 15887 16099
rect 17877 16065 17911 16099
rect 18797 16065 18831 16099
rect 18981 16065 19015 16099
rect 19073 16065 19107 16099
rect 19349 16065 19383 16099
rect 20361 16065 20395 16099
rect 22017 16065 22051 16099
rect 22109 16065 22143 16099
rect 22385 16065 22419 16099
rect 23029 16065 23063 16099
rect 24133 16065 24167 16099
rect 25136 16065 25170 16099
rect 27445 16065 27479 16099
rect 28733 16065 28767 16099
rect 12725 15997 12759 16031
rect 16037 15997 16071 16031
rect 17141 15997 17175 16031
rect 17325 15997 17359 16031
rect 19165 15997 19199 16031
rect 22293 15997 22327 16031
rect 24869 15997 24903 16031
rect 27721 15997 27755 16031
rect 10425 15929 10459 15963
rect 14013 15929 14047 15963
rect 16681 15929 16715 15963
rect 10885 15861 10919 15895
rect 14105 15861 14139 15895
rect 20453 15861 20487 15895
rect 21189 15861 21223 15895
rect 26249 15861 26283 15895
rect 30113 15861 30147 15895
rect 11253 15657 11287 15691
rect 13553 15657 13587 15691
rect 14197 15657 14231 15691
rect 18521 15657 18555 15691
rect 25329 15657 25363 15691
rect 28641 15657 28675 15691
rect 11621 15589 11655 15623
rect 28089 15589 28123 15623
rect 11529 15521 11563 15555
rect 12725 15521 12759 15555
rect 13093 15521 13127 15555
rect 14841 15521 14875 15555
rect 16037 15521 16071 15555
rect 19533 15521 19567 15555
rect 20913 15521 20947 15555
rect 23121 15521 23155 15555
rect 24961 15521 24995 15555
rect 1593 15453 1627 15487
rect 1777 15453 1811 15487
rect 10609 15453 10643 15487
rect 11437 15453 11471 15487
rect 11713 15453 11747 15487
rect 11897 15453 11931 15487
rect 10793 15385 10827 15419
rect 12817 15453 12851 15487
rect 13001 15453 13035 15487
rect 13185 15453 13219 15487
rect 13369 15453 13403 15487
rect 14565 15453 14599 15487
rect 17141 15453 17175 15487
rect 19257 15453 19291 15487
rect 19441 15453 19475 15487
rect 19625 15453 19659 15487
rect 19809 15453 19843 15487
rect 22753 15453 22787 15487
rect 22937 15453 22971 15487
rect 23029 15453 23063 15487
rect 23305 15453 23339 15487
rect 24593 15453 24627 15487
rect 24777 15453 24811 15487
rect 24869 15453 24903 15487
rect 25145 15453 25179 15487
rect 26065 15453 26099 15487
rect 26709 15453 26743 15487
rect 28549 15453 28583 15487
rect 30113 15453 30147 15487
rect 15761 15385 15795 15419
rect 17408 15385 17442 15419
rect 21180 15385 21214 15419
rect 26157 15385 26191 15419
rect 26976 15385 27010 15419
rect 1685 15317 1719 15351
rect 12725 15317 12759 15351
rect 14657 15317 14691 15351
rect 15393 15317 15427 15351
rect 15853 15317 15887 15351
rect 19993 15317 20027 15351
rect 22293 15317 22327 15351
rect 23489 15317 23523 15351
rect 29929 15317 29963 15351
rect 12265 15113 12299 15147
rect 12909 15113 12943 15147
rect 13369 15113 13403 15147
rect 19349 15113 19383 15147
rect 22569 15113 22603 15147
rect 24317 15113 24351 15147
rect 9680 15045 9714 15079
rect 15945 15045 15979 15079
rect 25329 15045 25363 15079
rect 25513 15045 25547 15079
rect 26157 15045 26191 15079
rect 1409 14977 1443 15011
rect 11529 14977 11563 15011
rect 11717 14977 11751 15011
rect 12081 14977 12115 15011
rect 13277 14977 13311 15011
rect 14657 14977 14691 15011
rect 14841 14977 14875 15011
rect 15209 14977 15243 15011
rect 17040 14977 17074 15011
rect 18613 14977 18647 15011
rect 18797 14977 18831 15011
rect 18889 14977 18923 15011
rect 19165 14977 19199 15011
rect 20168 14977 20202 15011
rect 21833 14977 21867 15011
rect 22017 14977 22051 15011
rect 22385 14977 22419 15011
rect 23029 14977 23063 15011
rect 23213 14977 23247 15011
rect 23397 14977 23431 15011
rect 23581 14977 23615 15011
rect 24225 14977 24259 15011
rect 25973 14977 26007 15011
rect 26249 14977 26283 15011
rect 26377 14977 26411 15011
rect 27721 14977 27755 15011
rect 28733 14977 28767 15011
rect 29000 14977 29034 15011
rect 9413 14909 9447 14943
rect 11805 14909 11839 14943
rect 11897 14909 11931 14943
rect 13461 14909 13495 14943
rect 14933 14909 14967 14943
rect 15025 14909 15059 14943
rect 15393 14909 15427 14943
rect 16773 14909 16807 14943
rect 18981 14909 19015 14943
rect 19901 14909 19935 14943
rect 22109 14909 22143 14943
rect 22201 14909 22235 14943
rect 23305 14909 23339 14943
rect 26157 14909 26191 14943
rect 27445 14909 27479 14943
rect 1593 14841 1627 14875
rect 10793 14841 10827 14875
rect 16037 14773 16071 14807
rect 18153 14773 18187 14807
rect 21281 14773 21315 14807
rect 23765 14773 23799 14807
rect 30113 14773 30147 14807
rect 12357 14569 12391 14603
rect 13277 14569 13311 14603
rect 15301 14569 15335 14603
rect 16681 14569 16715 14603
rect 18705 14569 18739 14603
rect 27445 14569 27479 14603
rect 29653 14501 29687 14535
rect 8953 14433 8987 14467
rect 11529 14433 11563 14467
rect 14749 14433 14783 14467
rect 15945 14433 15979 14467
rect 21373 14433 21407 14467
rect 21465 14433 21499 14467
rect 26985 14433 27019 14467
rect 27905 14433 27939 14467
rect 11437 14365 11471 14399
rect 12265 14365 12299 14399
rect 12909 14365 12943 14399
rect 14473 14365 14507 14399
rect 15761 14365 15795 14399
rect 16589 14365 16623 14399
rect 17233 14365 17267 14399
rect 17969 14365 18003 14399
rect 18153 14365 18187 14399
rect 18248 14365 18282 14399
rect 18337 14365 18371 14399
rect 18521 14365 18555 14399
rect 19257 14365 19291 14399
rect 19524 14365 19558 14399
rect 21097 14365 21131 14399
rect 21281 14365 21315 14399
rect 21649 14365 21683 14399
rect 22477 14365 22511 14399
rect 24501 14365 24535 14399
rect 26709 14365 26743 14399
rect 26893 14365 26927 14399
rect 27077 14365 27111 14399
rect 27261 14365 27295 14399
rect 28181 14365 28215 14399
rect 29561 14365 29595 14399
rect 9220 14297 9254 14331
rect 12081 14297 12115 14331
rect 13093 14297 13127 14331
rect 14565 14297 14599 14331
rect 17325 14297 17359 14331
rect 22744 14297 22778 14331
rect 24768 14297 24802 14331
rect 10333 14229 10367 14263
rect 14105 14229 14139 14263
rect 15669 14229 15703 14263
rect 20637 14229 20671 14263
rect 21833 14229 21867 14263
rect 23857 14229 23891 14263
rect 25881 14229 25915 14263
rect 10241 14025 10275 14059
rect 14749 14025 14783 14059
rect 15669 14025 15703 14059
rect 17325 14025 17359 14059
rect 21925 14025 21959 14059
rect 24317 14025 24351 14059
rect 28181 14025 28215 14059
rect 14381 13957 14415 13991
rect 18429 13957 18463 13991
rect 25973 13957 26007 13991
rect 9505 13889 9539 13923
rect 9689 13889 9723 13923
rect 10057 13889 10091 13923
rect 10701 13889 10735 13923
rect 11805 13889 11839 13923
rect 11897 13889 11931 13923
rect 14565 13889 14599 13923
rect 15577 13889 15611 13923
rect 16681 13889 16715 13923
rect 16865 13889 16899 13923
rect 17509 13889 17543 13923
rect 18245 13889 18279 13923
rect 21833 13889 21867 13923
rect 22937 13889 22971 13923
rect 23204 13889 23238 13923
rect 24961 13889 24995 13923
rect 25605 13889 25639 13923
rect 25789 13889 25823 13923
rect 26157 13889 26191 13923
rect 26341 13889 26375 13923
rect 27445 13889 27479 13923
rect 27629 13889 27663 13923
rect 27997 13889 28031 13923
rect 29000 13889 29034 13923
rect 9781 13821 9815 13855
rect 9873 13821 9907 13855
rect 10793 13821 10827 13855
rect 12081 13821 12115 13855
rect 16773 13821 16807 13855
rect 25145 13821 25179 13855
rect 27721 13821 27755 13855
rect 27813 13821 27847 13855
rect 28733 13821 28767 13855
rect 11989 13685 12023 13719
rect 30113 13685 30147 13719
rect 11437 13481 11471 13515
rect 12449 13481 12483 13515
rect 14749 13481 14783 13515
rect 16313 13481 16347 13515
rect 19901 13481 19935 13515
rect 22845 13481 22879 13515
rect 23489 13481 23523 13515
rect 25145 13481 25179 13515
rect 25881 13481 25915 13515
rect 29009 13481 29043 13515
rect 18245 13413 18279 13447
rect 29653 13413 29687 13447
rect 10425 13345 10459 13379
rect 10977 13345 11011 13379
rect 15209 13345 15243 13379
rect 15301 13345 15335 13379
rect 21097 13345 21131 13379
rect 24685 13345 24719 13379
rect 27353 13345 27387 13379
rect 1409 13277 1443 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 10517 13277 10551 13311
rect 11161 13277 11195 13311
rect 11253 13277 11287 13311
rect 11529 13277 11563 13311
rect 12173 13277 12207 13311
rect 12265 13277 12299 13311
rect 12541 13277 12575 13311
rect 14105 13277 14139 13311
rect 16129 13277 16163 13311
rect 20453 13277 20487 13311
rect 21373 13277 21407 13311
rect 22753 13277 22787 13311
rect 23397 13277 23431 13311
rect 24409 13277 24443 13311
rect 24593 13277 24627 13311
rect 24777 13277 24811 13311
rect 24961 13277 24995 13311
rect 26285 13277 26319 13311
rect 27077 13277 27111 13311
rect 27261 13277 27295 13311
rect 27445 13277 27479 13311
rect 27629 13277 27663 13311
rect 28273 13277 28307 13311
rect 28461 13277 28495 13311
rect 28552 13277 28586 13311
rect 28641 13277 28675 13311
rect 28825 13277 28859 13311
rect 29561 13277 29595 13311
rect 14197 13209 14231 13243
rect 15945 13209 15979 13243
rect 18061 13209 18095 13243
rect 19809 13209 19843 13243
rect 25881 13209 25915 13243
rect 26065 13209 26099 13243
rect 26157 13209 26191 13243
rect 1593 13141 1627 13175
rect 9965 13141 9999 13175
rect 11989 13141 12023 13175
rect 15117 13141 15151 13175
rect 20545 13141 20579 13175
rect 27813 13141 27847 13175
rect 10057 12937 10091 12971
rect 13829 12937 13863 12971
rect 14197 12937 14231 12971
rect 15577 12937 15611 12971
rect 16773 12937 16807 12971
rect 23581 12937 23615 12971
rect 28549 12937 28583 12971
rect 29745 12937 29779 12971
rect 23489 12869 23523 12903
rect 25973 12869 26007 12903
rect 9413 12801 9447 12835
rect 9597 12801 9631 12835
rect 10425 12801 10459 12835
rect 11713 12801 11747 12835
rect 12725 12801 12759 12835
rect 15761 12801 15795 12835
rect 15853 12801 15887 12835
rect 16129 12801 16163 12835
rect 16681 12801 16715 12835
rect 18153 12801 18187 12835
rect 18337 12801 18371 12835
rect 18705 12801 18739 12835
rect 19533 12801 19567 12835
rect 19809 12801 19843 12835
rect 20545 12801 20579 12835
rect 20821 12801 20855 12835
rect 21833 12801 21867 12835
rect 24133 12801 24167 12835
rect 24317 12801 24351 12835
rect 24501 12801 24535 12835
rect 24685 12801 24719 12835
rect 25605 12801 25639 12835
rect 25789 12801 25823 12835
rect 26157 12801 26191 12835
rect 26433 12801 26467 12835
rect 27169 12801 27203 12835
rect 27436 12801 27470 12835
rect 29009 12801 29043 12835
rect 29193 12801 29227 12835
rect 29377 12801 29411 12835
rect 29561 12801 29595 12835
rect 9505 12733 9539 12767
rect 10517 12733 10551 12767
rect 10701 12733 10735 12767
rect 11805 12733 11839 12767
rect 12817 12733 12851 12767
rect 13001 12733 13035 12767
rect 14289 12733 14323 12767
rect 14473 12733 14507 12767
rect 18429 12733 18463 12767
rect 18521 12733 18555 12767
rect 19625 12733 19659 12767
rect 20637 12733 20671 12767
rect 22109 12733 22143 12767
rect 24409 12733 24443 12767
rect 29285 12733 29319 12767
rect 19349 12665 19383 12699
rect 19717 12665 19751 12699
rect 20729 12665 20763 12699
rect 12357 12597 12391 12631
rect 16037 12597 16071 12631
rect 18889 12597 18923 12631
rect 20361 12597 20395 12631
rect 24869 12597 24903 12631
rect 10333 12393 10367 12427
rect 11529 12393 11563 12427
rect 18705 12393 18739 12427
rect 14105 12325 14139 12359
rect 21189 12325 21223 12359
rect 26525 12325 26559 12359
rect 10793 12257 10827 12291
rect 10885 12257 10919 12291
rect 12081 12257 12115 12291
rect 14749 12257 14783 12291
rect 17325 12257 17359 12291
rect 21373 12257 21407 12291
rect 24685 12257 24719 12291
rect 10701 12189 10735 12223
rect 12817 12189 12851 12223
rect 12909 12189 12943 12223
rect 15393 12189 15427 12223
rect 16221 12189 16255 12223
rect 16369 12189 16403 12223
rect 16727 12189 16761 12223
rect 17592 12189 17626 12223
rect 19257 12189 19291 12223
rect 21097 12189 21131 12223
rect 22006 12189 22040 12223
rect 24409 12189 24443 12223
rect 24593 12189 24627 12223
rect 24777 12189 24811 12223
rect 24961 12189 24995 12223
rect 26249 12189 26283 12223
rect 26341 12189 26375 12223
rect 26617 12189 26651 12223
rect 26801 12189 26835 12223
rect 27537 12189 27571 12223
rect 27813 12189 27847 12223
rect 29009 12189 29043 12223
rect 30113 12189 30147 12223
rect 16497 12121 16531 12155
rect 16589 12121 16623 12155
rect 19524 12121 19558 12155
rect 22284 12121 22318 12155
rect 11897 12053 11931 12087
rect 11989 12053 12023 12087
rect 13093 12053 13127 12087
rect 14473 12053 14507 12087
rect 14565 12053 14599 12087
rect 15669 12053 15703 12087
rect 16865 12053 16899 12087
rect 20637 12053 20671 12087
rect 21373 12053 21407 12087
rect 23397 12053 23431 12087
rect 25145 12053 25179 12087
rect 28825 12053 28859 12087
rect 29929 12053 29963 12087
rect 12081 11849 12115 11883
rect 12909 11849 12943 11883
rect 13553 11849 13587 11883
rect 13921 11849 13955 11883
rect 15117 11849 15151 11883
rect 18061 11849 18095 11883
rect 19533 11849 19567 11883
rect 21281 11849 21315 11883
rect 23489 11849 23523 11883
rect 25329 11849 25363 11883
rect 9873 11781 9907 11815
rect 10057 11781 10091 11815
rect 24216 11781 24250 11815
rect 25881 11781 25915 11815
rect 11989 11713 12023 11747
rect 12173 11713 12207 11747
rect 13093 11713 13127 11747
rect 14749 11713 14783 11747
rect 14841 11713 14875 11747
rect 15761 11713 15795 11747
rect 15945 11713 15979 11747
rect 16681 11713 16715 11747
rect 16948 11713 16982 11747
rect 18797 11713 18831 11747
rect 18981 11713 19015 11747
rect 19073 11713 19107 11747
rect 19349 11713 19383 11747
rect 20545 11713 20579 11747
rect 20729 11713 20763 11747
rect 20959 11713 20993 11747
rect 21097 11713 21131 11747
rect 22109 11713 22143 11747
rect 22376 11713 22410 11747
rect 23949 11713 23983 11747
rect 27537 11713 27571 11747
rect 27721 11713 27755 11747
rect 27813 11713 27847 11747
rect 28089 11713 28123 11747
rect 29000 11713 29034 11747
rect 14013 11645 14047 11679
rect 14197 11645 14231 11679
rect 15117 11645 15151 11679
rect 16037 11645 16071 11679
rect 19165 11645 19199 11679
rect 20821 11645 20855 11679
rect 27905 11645 27939 11679
rect 28733 11645 28767 11679
rect 14933 11577 14967 11611
rect 15577 11577 15611 11611
rect 26065 11577 26099 11611
rect 10241 11509 10275 11543
rect 14749 11509 14783 11543
rect 28273 11509 28307 11543
rect 30113 11509 30147 11543
rect 10517 11305 10551 11339
rect 11897 11305 11931 11339
rect 15301 11305 15335 11339
rect 16129 11305 16163 11339
rect 16865 11305 16899 11339
rect 20821 11305 20855 11339
rect 22109 11305 22143 11339
rect 23765 11305 23799 11339
rect 25789 11305 25823 11339
rect 29745 11305 29779 11339
rect 9413 11237 9447 11271
rect 10609 11237 10643 11271
rect 11989 11237 12023 11271
rect 26709 11237 26743 11271
rect 27629 11237 27663 11271
rect 29009 11237 29043 11271
rect 19625 11169 19659 11203
rect 21649 11169 21683 11203
rect 24409 11169 24443 11203
rect 28549 11169 28583 11203
rect 1409 11101 1443 11135
rect 2145 11101 2179 11135
rect 2329 11101 2363 11135
rect 9597 11101 9631 11135
rect 10149 11101 10183 11135
rect 10333 11101 10367 11135
rect 10425 11101 10459 11135
rect 10701 11101 10735 11135
rect 11529 11101 11563 11135
rect 11713 11101 11747 11135
rect 11805 11101 11839 11135
rect 12081 11101 12115 11135
rect 15209 11101 15243 11135
rect 15945 11101 15979 11135
rect 16129 11101 16163 11135
rect 16773 11101 16807 11135
rect 19257 11101 19291 11135
rect 19441 11101 19475 11135
rect 19533 11101 19567 11135
rect 19809 11101 19843 11135
rect 20729 11101 20763 11135
rect 21373 11101 21407 11135
rect 21557 11101 21591 11135
rect 21741 11101 21775 11135
rect 21925 11101 21959 11135
rect 23673 11101 23707 11135
rect 24676 11101 24710 11135
rect 26341 11101 26375 11135
rect 26617 11101 26651 11135
rect 26801 11101 26835 11135
rect 26985 11101 27019 11135
rect 27813 11101 27847 11135
rect 28273 11101 28307 11135
rect 28457 11101 28491 11135
rect 28641 11101 28675 11135
rect 28825 11101 28859 11135
rect 2237 11033 2271 11067
rect 29653 11033 29687 11067
rect 1593 10965 1627 10999
rect 16313 10965 16347 10999
rect 19993 10965 20027 10999
rect 10793 10761 10827 10795
rect 11897 10761 11931 10795
rect 12357 10761 12391 10795
rect 12725 10761 12759 10795
rect 21925 10761 21959 10795
rect 30113 10761 30147 10795
rect 10425 10693 10459 10727
rect 20913 10693 20947 10727
rect 29000 10693 29034 10727
rect 10609 10625 10643 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 14933 10625 14967 10659
rect 15577 10625 15611 10659
rect 15761 10625 15795 10659
rect 15945 10625 15979 10659
rect 16681 10625 16715 10659
rect 17601 10625 17635 10659
rect 18521 10625 18555 10659
rect 19809 10625 19843 10659
rect 21833 10625 21867 10659
rect 24041 10625 24075 10659
rect 25605 10625 25639 10659
rect 25789 10625 25823 10659
rect 26157 10625 26191 10659
rect 26433 10625 26467 10659
rect 26985 10625 27019 10659
rect 27169 10625 27203 10659
rect 27537 10625 27571 10659
rect 27629 10625 27663 10659
rect 12817 10557 12851 10591
rect 13001 10557 13035 10591
rect 18245 10557 18279 10591
rect 19533 10557 19567 10591
rect 21097 10557 21131 10591
rect 24317 10557 24351 10591
rect 27077 10557 27111 10591
rect 28733 10557 28767 10591
rect 17785 10489 17819 10523
rect 25605 10489 25639 10523
rect 15025 10421 15059 10455
rect 16773 10421 16807 10455
rect 10609 10217 10643 10251
rect 12449 10217 12483 10251
rect 14105 10217 14139 10251
rect 16589 10217 16623 10251
rect 18429 10217 18463 10251
rect 28549 10217 28583 10251
rect 15945 10149 15979 10183
rect 11253 10081 11287 10115
rect 12909 10081 12943 10115
rect 13001 10081 13035 10115
rect 14749 10081 14783 10115
rect 21649 10081 21683 10115
rect 21741 10081 21775 10115
rect 24961 10081 24995 10115
rect 10977 10013 11011 10047
rect 12817 10013 12851 10047
rect 15301 10013 15335 10047
rect 15449 10013 15483 10047
rect 15766 10013 15800 10047
rect 16497 10013 16531 10047
rect 17141 10013 17175 10047
rect 17234 10013 17268 10047
rect 17417 10013 17451 10047
rect 17647 10013 17681 10047
rect 19257 10013 19291 10047
rect 19524 10013 19558 10047
rect 21373 10013 21407 10047
rect 21557 10013 21591 10047
rect 21925 10013 21959 10047
rect 25237 10013 25271 10047
rect 26341 10013 26375 10047
rect 27169 10013 27203 10047
rect 30113 10013 30147 10047
rect 11069 9945 11103 9979
rect 14473 9945 14507 9979
rect 15577 9945 15611 9979
rect 15669 9945 15703 9979
rect 17509 9945 17543 9979
rect 18337 9945 18371 9979
rect 27436 9945 27470 9979
rect 14565 9877 14599 9911
rect 17785 9877 17819 9911
rect 20637 9877 20671 9911
rect 22109 9877 22143 9911
rect 26433 9877 26467 9911
rect 29929 9877 29963 9911
rect 10241 9673 10275 9707
rect 12633 9673 12667 9707
rect 15853 9673 15887 9707
rect 18061 9673 18095 9707
rect 25329 9673 25363 9707
rect 14381 9605 14415 9639
rect 16948 9605 16982 9639
rect 26249 9605 26283 9639
rect 10609 9537 10643 9571
rect 12173 9537 12207 9571
rect 13001 9537 13035 9571
rect 14013 9537 14047 9571
rect 14197 9537 14231 9571
rect 15117 9537 15151 9571
rect 15301 9537 15335 9571
rect 15393 9537 15427 9571
rect 16037 9537 16071 9571
rect 18521 9537 18555 9571
rect 18614 9537 18648 9571
rect 18797 9537 18831 9571
rect 18889 9537 18923 9571
rect 19027 9537 19061 9571
rect 19901 9537 19935 9571
rect 20168 9537 20202 9571
rect 22017 9537 22051 9571
rect 22284 9537 22318 9571
rect 23949 9537 23983 9571
rect 24205 9537 24239 9571
rect 27445 9537 27479 9571
rect 27721 9537 27755 9571
rect 29000 9537 29034 9571
rect 10701 9469 10735 9503
rect 10793 9469 10827 9503
rect 13093 9469 13127 9503
rect 13277 9469 13311 9503
rect 16681 9469 16715 9503
rect 28733 9469 28767 9503
rect 11989 9401 12023 9435
rect 14933 9401 14967 9435
rect 26433 9401 26467 9435
rect 30113 9401 30147 9435
rect 19165 9333 19199 9367
rect 21281 9333 21315 9367
rect 23397 9333 23431 9367
rect 10977 9129 11011 9163
rect 13185 9129 13219 9163
rect 14197 9129 14231 9163
rect 15669 9129 15703 9163
rect 16865 9129 16899 9163
rect 19809 9129 19843 9163
rect 22569 9129 22603 9163
rect 28641 9129 28675 9163
rect 21373 9061 21407 9095
rect 11621 8993 11655 9027
rect 14841 8993 14875 9027
rect 17417 8993 17451 9027
rect 17693 8993 17727 9027
rect 23397 8993 23431 9027
rect 25697 8993 25731 9027
rect 26801 8993 26835 9027
rect 27353 8993 27387 9027
rect 27629 8993 27663 9027
rect 1409 8925 1443 8959
rect 13001 8925 13035 8959
rect 15577 8925 15611 8959
rect 15761 8925 15795 8959
rect 16773 8925 16807 8959
rect 19717 8925 19751 8959
rect 20729 8925 20763 8959
rect 20877 8925 20911 8959
rect 21005 8925 21039 8959
rect 21235 8925 21269 8959
rect 21925 8925 21959 8959
rect 22018 8925 22052 8959
rect 22390 8925 22424 8959
rect 23121 8925 23155 8959
rect 23305 8925 23339 8959
rect 23489 8925 23523 8959
rect 23673 8925 23707 8959
rect 25421 8925 25455 8959
rect 26709 8925 26743 8959
rect 28825 8925 28859 8959
rect 30113 8925 30147 8959
rect 12817 8857 12851 8891
rect 21097 8857 21131 8891
rect 22201 8857 22235 8891
rect 22293 8857 22327 8891
rect 1593 8789 1627 8823
rect 11345 8789 11379 8823
rect 11437 8789 11471 8823
rect 14565 8789 14599 8823
rect 14657 8789 14691 8823
rect 23857 8789 23891 8823
rect 29929 8789 29963 8823
rect 10793 8585 10827 8619
rect 13829 8585 13863 8619
rect 15393 8585 15427 8619
rect 19441 8585 19475 8619
rect 20545 8585 20579 8619
rect 23581 8585 23615 8619
rect 30113 8585 30147 8619
rect 11713 8517 11747 8551
rect 14841 8517 14875 8551
rect 16865 8517 16899 8551
rect 18328 8517 18362 8551
rect 20453 8517 20487 8551
rect 22109 8517 22143 8551
rect 24286 8517 24320 8551
rect 10977 8449 11011 8483
rect 11529 8449 11563 8483
rect 12541 8449 12575 8483
rect 14013 8449 14047 8483
rect 14473 8449 14507 8483
rect 14657 8449 14691 8483
rect 15761 8449 15795 8483
rect 15853 8449 15887 8483
rect 16681 8449 16715 8483
rect 21925 8449 21959 8483
rect 22845 8449 22879 8483
rect 23029 8449 23063 8483
rect 23121 8449 23155 8483
rect 23397 8449 23431 8483
rect 24041 8449 24075 8483
rect 27261 8449 27295 8483
rect 29000 8449 29034 8483
rect 11897 8381 11931 8415
rect 15945 8381 15979 8415
rect 18061 8381 18095 8415
rect 23213 8381 23247 8415
rect 26985 8381 27019 8415
rect 28733 8381 28767 8415
rect 12357 8313 12391 8347
rect 25421 8313 25455 8347
rect 17049 8245 17083 8279
rect 12633 8041 12667 8075
rect 16037 8041 16071 8075
rect 18613 8041 18647 8075
rect 19625 8041 19659 8075
rect 20269 8041 20303 8075
rect 23489 8041 23523 8075
rect 24501 8041 24535 8075
rect 26709 8041 26743 8075
rect 28365 8041 28399 8075
rect 21097 7905 21131 7939
rect 25329 7905 25363 7939
rect 12265 7837 12299 7871
rect 13093 7837 13127 7871
rect 14289 7837 14323 7871
rect 16221 7837 16255 7871
rect 17325 7837 17359 7871
rect 17473 7837 17507 7871
rect 17693 7837 17727 7871
rect 17831 7837 17865 7871
rect 19441 7837 19475 7871
rect 19717 7837 19751 7871
rect 20177 7837 20211 7871
rect 20821 7837 20855 7871
rect 22098 7837 22132 7871
rect 22257 7837 22291 7871
rect 22615 7837 22649 7871
rect 23397 7837 23431 7871
rect 24409 7837 24443 7871
rect 25585 7837 25619 7871
rect 27629 7837 27663 7871
rect 27813 7837 27847 7871
rect 27905 7837 27939 7871
rect 27997 7837 28031 7871
rect 28181 7837 28215 7871
rect 30113 7837 30147 7871
rect 12449 7769 12483 7803
rect 17601 7769 17635 7803
rect 18521 7769 18555 7803
rect 22385 7769 22419 7803
rect 22477 7769 22511 7803
rect 13277 7701 13311 7735
rect 14289 7701 14323 7735
rect 17969 7701 18003 7735
rect 19257 7701 19291 7735
rect 22753 7701 22787 7735
rect 29929 7701 29963 7735
rect 14657 7497 14691 7531
rect 24133 7497 24167 7531
rect 28365 7497 28399 7531
rect 29561 7497 29595 7531
rect 14197 7429 14231 7463
rect 17040 7429 17074 7463
rect 1409 7361 1443 7395
rect 12357 7361 12391 7395
rect 12541 7361 12575 7395
rect 13277 7361 13311 7395
rect 14841 7361 14875 7395
rect 16773 7361 16807 7395
rect 19349 7361 19383 7395
rect 19616 7361 19650 7395
rect 21833 7361 21867 7395
rect 22753 7361 22787 7395
rect 23020 7361 23054 7395
rect 25329 7361 25363 7395
rect 27252 7361 27286 7395
rect 28825 7361 28859 7395
rect 29009 7361 29043 7395
rect 29377 7361 29411 7395
rect 13394 7293 13428 7327
rect 13553 7293 13587 7327
rect 25053 7293 25087 7327
rect 26985 7293 27019 7327
rect 29101 7293 29135 7327
rect 29193 7293 29227 7327
rect 13001 7225 13035 7259
rect 1593 7157 1627 7191
rect 18153 7157 18187 7191
rect 20729 7157 20763 7191
rect 21925 7157 21959 7191
rect 15485 6953 15519 6987
rect 20453 6953 20487 6987
rect 22293 6953 22327 6987
rect 23397 6953 23431 6987
rect 27169 6953 27203 6987
rect 11253 6885 11287 6919
rect 10609 6817 10643 6851
rect 11529 6817 11563 6851
rect 11805 6817 11839 6851
rect 13277 6817 13311 6851
rect 16129 6817 16163 6851
rect 17141 6817 17175 6851
rect 18337 6817 18371 6851
rect 25513 6817 25547 6851
rect 25605 6817 25639 6851
rect 26801 6817 26835 6851
rect 10793 6749 10827 6783
rect 11667 6749 11701 6783
rect 12909 6749 12943 6783
rect 13093 6749 13127 6783
rect 16681 6749 16715 6783
rect 16865 6749 16899 6783
rect 16957 6749 16991 6783
rect 17233 6749 17267 6783
rect 17969 6749 18003 6783
rect 18153 6747 18187 6781
rect 18248 6749 18282 6783
rect 18521 6749 18555 6783
rect 19809 6749 19843 6783
rect 19957 6749 19991 6783
rect 20315 6749 20349 6783
rect 20913 6749 20947 6783
rect 22753 6749 22787 6783
rect 22846 6749 22880 6783
rect 23029 6749 23063 6783
rect 23218 6749 23252 6783
rect 25237 6749 25271 6783
rect 25421 6749 25455 6783
rect 25789 6749 25823 6783
rect 26433 6749 26467 6783
rect 26617 6749 26651 6783
rect 26709 6749 26743 6783
rect 26985 6749 27019 6783
rect 27629 6749 27663 6783
rect 30113 6749 30147 6783
rect 15945 6681 15979 6715
rect 20085 6681 20119 6715
rect 20177 6681 20211 6715
rect 21180 6681 21214 6715
rect 23121 6681 23155 6715
rect 27896 6681 27930 6715
rect 12449 6613 12483 6647
rect 15853 6613 15887 6647
rect 16681 6613 16715 6647
rect 18705 6613 18739 6647
rect 25973 6613 26007 6647
rect 29009 6613 29043 6647
rect 29929 6613 29963 6647
rect 11989 6409 12023 6443
rect 12449 6409 12483 6443
rect 13277 6409 13311 6443
rect 15945 6409 15979 6443
rect 21925 6409 21959 6443
rect 25697 6409 25731 6443
rect 27905 6409 27939 6443
rect 29101 6409 29135 6443
rect 29929 6409 29963 6443
rect 17693 6341 17727 6375
rect 12357 6273 12391 6307
rect 13185 6273 13219 6307
rect 17417 6273 17451 6307
rect 17510 6273 17544 6307
rect 17785 6273 17819 6307
rect 17882 6273 17916 6307
rect 18705 6273 18739 6307
rect 18889 6273 18923 6307
rect 18981 6273 19015 6307
rect 19257 6273 19291 6307
rect 20453 6273 20487 6307
rect 21833 6273 21867 6307
rect 22477 6273 22511 6307
rect 22744 6273 22778 6307
rect 24317 6273 24351 6307
rect 24584 6273 24618 6307
rect 27077 6273 27111 6307
rect 27169 6273 27203 6307
rect 27353 6273 27387 6307
rect 27721 6273 27755 6307
rect 28365 6273 28399 6307
rect 28549 6273 28583 6307
rect 28917 6273 28951 6307
rect 30113 6273 30147 6307
rect 12633 6205 12667 6239
rect 14105 6205 14139 6239
rect 14289 6205 14323 6239
rect 15025 6205 15059 6239
rect 15142 6205 15176 6239
rect 15301 6205 15335 6239
rect 19073 6205 19107 6239
rect 20729 6205 20763 6239
rect 14749 6137 14783 6171
rect 27445 6205 27479 6239
rect 27537 6205 27571 6239
rect 28641 6205 28675 6239
rect 28733 6205 28767 6239
rect 18061 6069 18095 6103
rect 19441 6069 19475 6103
rect 23857 6069 23891 6103
rect 27077 6069 27111 6103
rect 12449 5865 12483 5899
rect 15945 5865 15979 5899
rect 19441 5865 19475 5899
rect 22661 5865 22695 5899
rect 26709 5865 26743 5899
rect 28549 5865 28583 5899
rect 9965 5797 9999 5831
rect 19717 5797 19751 5831
rect 19809 5797 19843 5831
rect 10793 5729 10827 5763
rect 11253 5729 11287 5763
rect 11529 5729 11563 5763
rect 11646 5729 11680 5763
rect 11805 5729 11839 5763
rect 13553 5729 13587 5763
rect 14749 5729 14783 5763
rect 15142 5729 15176 5763
rect 15301 5729 15335 5763
rect 21189 5729 21223 5763
rect 25329 5729 25363 5763
rect 10149 5661 10183 5695
rect 10609 5661 10643 5695
rect 13277 5661 13311 5695
rect 13369 5661 13403 5695
rect 14105 5661 14139 5695
rect 14289 5661 14323 5695
rect 15025 5661 15059 5695
rect 16405 5661 16439 5695
rect 19625 5661 19659 5695
rect 19901 5661 19935 5695
rect 20821 5661 20855 5695
rect 20993 5661 21027 5695
rect 21097 5661 21131 5695
rect 21373 5661 21407 5695
rect 22017 5661 22051 5695
rect 22110 5661 22144 5695
rect 22293 5661 22327 5695
rect 22521 5661 22555 5695
rect 27169 5661 27203 5695
rect 22385 5593 22419 5627
rect 25596 5593 25630 5627
rect 27414 5593 27448 5627
rect 29929 5593 29963 5627
rect 13553 5525 13587 5559
rect 16497 5525 16531 5559
rect 21557 5525 21591 5559
rect 30021 5525 30055 5559
rect 11897 5321 11931 5355
rect 14841 5321 14875 5355
rect 18429 5321 18463 5355
rect 20361 5321 20395 5355
rect 25789 5321 25823 5355
rect 19248 5253 19282 5287
rect 1409 5185 1443 5219
rect 11713 5185 11747 5219
rect 13185 5185 13219 5219
rect 13645 5185 13679 5219
rect 15025 5185 15059 5219
rect 15117 5185 15151 5219
rect 15393 5185 15427 5219
rect 17049 5185 17083 5219
rect 17316 5185 17350 5219
rect 18981 5185 19015 5219
rect 21833 5185 21867 5219
rect 22017 5185 22051 5219
rect 22109 5185 22143 5219
rect 22385 5185 22419 5219
rect 25053 5185 25087 5219
rect 25237 5185 25271 5219
rect 25605 5185 25639 5219
rect 29929 5185 29963 5219
rect 11529 5117 11563 5151
rect 13737 5117 13771 5151
rect 22201 5117 22235 5151
rect 25329 5117 25363 5151
rect 25421 5117 25455 5151
rect 13001 5049 13035 5083
rect 14013 5049 14047 5083
rect 1593 4981 1627 5015
rect 13829 4981 13863 5015
rect 15301 4981 15335 5015
rect 22569 4981 22603 5015
rect 30021 4981 30055 5015
rect 12725 4777 12759 4811
rect 21373 4777 21407 4811
rect 23213 4777 23247 4811
rect 26157 4777 26191 4811
rect 14105 4709 14139 4743
rect 13369 4641 13403 4675
rect 14473 4641 14507 4675
rect 16129 4641 16163 4675
rect 25789 4641 25823 4675
rect 14289 4573 14323 4607
rect 14565 4573 14599 4607
rect 15025 4573 15059 4607
rect 16396 4573 16430 4607
rect 19993 4573 20027 4607
rect 21833 4573 21867 4607
rect 22100 4573 22134 4607
rect 25421 4573 25455 4607
rect 25605 4573 25639 4607
rect 25697 4573 25731 4607
rect 25973 4573 26007 4607
rect 20260 4505 20294 4539
rect 29929 4505 29963 4539
rect 13093 4437 13127 4471
rect 13185 4437 13219 4471
rect 15117 4437 15151 4471
rect 17509 4437 17543 4471
rect 30021 4437 30055 4471
rect 11713 4097 11747 4131
rect 12541 4097 12575 4131
rect 13553 4097 13587 4131
rect 14381 4097 14415 4131
rect 15209 4097 15243 4131
rect 15393 4097 15427 4131
rect 17049 4097 17083 4131
rect 18245 4097 18279 4131
rect 18512 4097 18546 4131
rect 29837 4097 29871 4131
rect 13001 4029 13035 4063
rect 13645 4029 13679 4063
rect 14197 4029 14231 4063
rect 14749 4029 14783 4063
rect 17141 4029 17175 4063
rect 17233 4029 17267 4063
rect 12357 3961 12391 3995
rect 13277 3961 13311 3995
rect 14657 3961 14691 3995
rect 16681 3961 16715 3995
rect 30021 3961 30055 3995
rect 11529 3893 11563 3927
rect 15301 3893 15335 3927
rect 19625 3893 19659 3927
rect 10517 3689 10551 3723
rect 13001 3689 13035 3723
rect 16221 3689 16255 3723
rect 11805 3621 11839 3655
rect 15025 3621 15059 3655
rect 11161 3553 11195 3587
rect 11345 3553 11379 3587
rect 12081 3553 12115 3587
rect 12219 3553 12253 3587
rect 14565 3553 14599 3587
rect 15301 3553 15335 3587
rect 10701 3485 10735 3519
rect 12357 3485 12391 3519
rect 14381 3485 14415 3519
rect 15418 3485 15452 3519
rect 15577 3485 15611 3519
rect 29837 3485 29871 3519
rect 30021 3349 30055 3383
rect 13369 3145 13403 3179
rect 16129 3145 16163 3179
rect 29837 3145 29871 3179
rect 1409 3009 1443 3043
rect 11529 3009 11563 3043
rect 11713 3009 11747 3043
rect 12566 3009 12600 3043
rect 14289 3009 14323 3043
rect 14473 3009 14507 3043
rect 15209 3009 15243 3043
rect 15347 3009 15381 3043
rect 29745 3009 29779 3043
rect 12449 2941 12483 2975
rect 12725 2941 12759 2975
rect 15485 2941 15519 2975
rect 1593 2873 1627 2907
rect 12173 2873 12207 2907
rect 14933 2873 14967 2907
rect 13277 2601 13311 2635
rect 14105 2601 14139 2635
rect 28917 2601 28951 2635
rect 29837 2601 29871 2635
rect 1409 2397 1443 2431
rect 12909 2397 12943 2431
rect 13093 2397 13127 2431
rect 14105 2397 14139 2431
rect 14289 2397 14323 2431
rect 28733 2397 28767 2431
rect 29745 2329 29779 2363
rect 1593 2261 1627 2295
<< metal1 >>
rect 14182 45772 14188 45824
rect 14240 45812 14246 45824
rect 15562 45812 15568 45824
rect 14240 45784 15568 45812
rect 14240 45772 14246 45784
rect 15562 45772 15568 45784
rect 15620 45772 15626 45824
rect 23290 45772 23296 45824
rect 23348 45812 23354 45824
rect 27062 45812 27068 45824
rect 23348 45784 27068 45812
rect 23348 45772 23354 45784
rect 27062 45772 27068 45784
rect 27120 45772 27126 45824
rect 1104 45722 30820 45744
rect 1104 45670 10880 45722
rect 10932 45670 10944 45722
rect 10996 45670 11008 45722
rect 11060 45670 11072 45722
rect 11124 45670 11136 45722
rect 11188 45670 20811 45722
rect 20863 45670 20875 45722
rect 20927 45670 20939 45722
rect 20991 45670 21003 45722
rect 21055 45670 21067 45722
rect 21119 45670 30820 45722
rect 1104 45648 30820 45670
rect 6365 45611 6423 45617
rect 6365 45577 6377 45611
rect 6411 45608 6423 45611
rect 8021 45611 8079 45617
rect 6411 45580 6445 45608
rect 6411 45577 6423 45580
rect 6365 45571 6423 45577
rect 8021 45577 8033 45611
rect 8067 45608 8079 45611
rect 16666 45608 16672 45620
rect 8067 45580 8101 45608
rect 9646 45580 16672 45608
rect 8067 45577 8079 45580
rect 8021 45571 8079 45577
rect 6380 45540 6408 45571
rect 8036 45540 8064 45571
rect 9646 45540 9674 45580
rect 16666 45568 16672 45580
rect 16724 45568 16730 45620
rect 16761 45611 16819 45617
rect 16761 45577 16773 45611
rect 16807 45608 16819 45611
rect 17494 45608 17500 45620
rect 16807 45580 17500 45608
rect 16807 45577 16819 45580
rect 16761 45571 16819 45577
rect 17494 45568 17500 45580
rect 17552 45568 17558 45620
rect 21085 45611 21143 45617
rect 21085 45577 21097 45611
rect 21131 45608 21143 45611
rect 23842 45608 23848 45620
rect 21131 45580 23848 45608
rect 21131 45577 21143 45580
rect 21085 45571 21143 45577
rect 23842 45568 23848 45580
rect 23900 45568 23906 45620
rect 30006 45608 30012 45620
rect 29967 45580 30012 45608
rect 30006 45568 30012 45580
rect 30064 45568 30070 45620
rect 16390 45540 16396 45552
rect 6380 45512 7880 45540
rect 8036 45512 9076 45540
rect 1578 45472 1584 45484
rect 1539 45444 1584 45472
rect 1578 45432 1584 45444
rect 1636 45432 1642 45484
rect 2409 45475 2467 45481
rect 2409 45441 2421 45475
rect 2455 45472 2467 45475
rect 2590 45472 2596 45484
rect 2455 45444 2596 45472
rect 2455 45441 2467 45444
rect 2409 45435 2467 45441
rect 2590 45432 2596 45444
rect 2648 45432 2654 45484
rect 3418 45432 3424 45484
rect 3476 45472 3482 45484
rect 3789 45475 3847 45481
rect 3789 45472 3801 45475
rect 3476 45444 3801 45472
rect 3476 45432 3482 45444
rect 3789 45441 3801 45444
rect 3835 45441 3847 45475
rect 3789 45435 3847 45441
rect 4154 45432 4160 45484
rect 4212 45472 4218 45484
rect 5077 45475 5135 45481
rect 5077 45472 5089 45475
rect 4212 45444 5089 45472
rect 4212 45432 4218 45444
rect 5077 45441 5089 45444
rect 5123 45441 5135 45475
rect 5077 45435 5135 45441
rect 5718 45432 5724 45484
rect 5776 45472 5782 45484
rect 6549 45475 6607 45481
rect 6549 45472 6561 45475
rect 5776 45444 6561 45472
rect 5776 45432 5782 45444
rect 6549 45441 6561 45444
rect 6595 45441 6607 45475
rect 6549 45435 6607 45441
rect 6914 45432 6920 45484
rect 6972 45472 6978 45484
rect 7193 45475 7251 45481
rect 7193 45472 7205 45475
rect 6972 45444 7205 45472
rect 6972 45432 6978 45444
rect 7193 45441 7205 45444
rect 7239 45441 7251 45475
rect 7193 45435 7251 45441
rect 2682 45404 2688 45416
rect 2643 45376 2688 45404
rect 2682 45364 2688 45376
rect 2740 45364 2746 45416
rect 4065 45407 4123 45413
rect 4065 45373 4077 45407
rect 4111 45373 4123 45407
rect 5350 45404 5356 45416
rect 5311 45376 5356 45404
rect 4065 45367 4123 45373
rect 4080 45336 4108 45367
rect 5350 45364 5356 45376
rect 5408 45364 5414 45416
rect 7852 45404 7880 45512
rect 7926 45432 7932 45484
rect 7984 45472 7990 45484
rect 8205 45475 8263 45481
rect 8205 45472 8217 45475
rect 7984 45444 8217 45472
rect 7984 45432 7990 45444
rect 8205 45441 8217 45444
rect 8251 45441 8263 45475
rect 8205 45435 8263 45441
rect 8754 45432 8760 45484
rect 8812 45472 8818 45484
rect 8941 45475 8999 45481
rect 8941 45472 8953 45475
rect 8812 45444 8953 45472
rect 8812 45432 8818 45444
rect 8941 45441 8953 45444
rect 8987 45441 8999 45475
rect 8941 45435 8999 45441
rect 8846 45404 8852 45416
rect 7852 45376 8852 45404
rect 8846 45364 8852 45376
rect 8904 45364 8910 45416
rect 8938 45336 8944 45348
rect 4080 45308 8944 45336
rect 8938 45296 8944 45308
rect 8996 45296 9002 45348
rect 9048 45336 9076 45512
rect 9232 45512 9674 45540
rect 14660 45512 16396 45540
rect 9232 45481 9260 45512
rect 9217 45475 9275 45481
rect 9217 45441 9229 45475
rect 9263 45441 9275 45475
rect 9217 45435 9275 45441
rect 9490 45432 9496 45484
rect 9548 45472 9554 45484
rect 10229 45475 10287 45481
rect 10229 45472 10241 45475
rect 9548 45444 10241 45472
rect 9548 45432 9554 45444
rect 10229 45441 10241 45444
rect 10275 45441 10287 45475
rect 10229 45435 10287 45441
rect 11238 45432 11244 45484
rect 11296 45472 11302 45484
rect 11517 45475 11575 45481
rect 11517 45472 11529 45475
rect 11296 45444 11529 45472
rect 11296 45432 11302 45444
rect 11517 45441 11529 45444
rect 11563 45441 11575 45475
rect 11517 45435 11575 45441
rect 12621 45475 12679 45481
rect 12621 45441 12633 45475
rect 12667 45472 12679 45475
rect 12897 45475 12955 45481
rect 12897 45472 12909 45475
rect 12667 45470 12756 45472
rect 12820 45470 12909 45472
rect 12667 45444 12909 45470
rect 12667 45441 12679 45444
rect 12728 45442 12848 45444
rect 12621 45435 12679 45441
rect 12897 45441 12909 45444
rect 12943 45472 12955 45475
rect 13446 45472 13452 45484
rect 12943 45444 13452 45472
rect 12943 45441 12955 45444
rect 12897 45435 12955 45441
rect 13446 45432 13452 45444
rect 13504 45432 13510 45484
rect 13541 45475 13599 45481
rect 13541 45441 13553 45475
rect 13587 45472 13599 45475
rect 13814 45472 13820 45484
rect 13587 45444 13820 45472
rect 13587 45441 13599 45444
rect 13541 45435 13599 45441
rect 13814 45432 13820 45444
rect 13872 45432 13878 45484
rect 14660 45481 14688 45512
rect 16390 45500 16396 45512
rect 16448 45500 16454 45552
rect 20990 45540 20996 45552
rect 16776 45512 20996 45540
rect 14645 45475 14703 45481
rect 14645 45441 14657 45475
rect 14691 45441 14703 45475
rect 15286 45472 15292 45484
rect 15247 45444 15292 45472
rect 14645 45435 14703 45441
rect 15286 45432 15292 45444
rect 15344 45432 15350 45484
rect 16776 45472 16804 45512
rect 20990 45500 20996 45512
rect 21048 45500 21054 45552
rect 21450 45540 21456 45552
rect 21292 45512 21456 45540
rect 16942 45472 16948 45484
rect 15488 45444 16804 45472
rect 16903 45444 16948 45472
rect 15488 45404 15516 45444
rect 16942 45432 16948 45444
rect 17000 45432 17006 45484
rect 17773 45475 17831 45481
rect 17773 45441 17785 45475
rect 17819 45441 17831 45475
rect 18414 45472 18420 45484
rect 18375 45444 18420 45472
rect 17773 45435 17831 45441
rect 12636 45376 15516 45404
rect 15565 45407 15623 45413
rect 12636 45336 12664 45376
rect 15565 45373 15577 45407
rect 15611 45404 15623 45407
rect 16666 45404 16672 45416
rect 15611 45376 16672 45404
rect 15611 45373 15623 45376
rect 15565 45367 15623 45373
rect 16666 45364 16672 45376
rect 16724 45404 16730 45416
rect 17221 45407 17279 45413
rect 17221 45404 17233 45407
rect 16724 45376 17233 45404
rect 16724 45364 16730 45376
rect 17221 45373 17233 45376
rect 17267 45404 17279 45407
rect 17402 45404 17408 45416
rect 17267 45376 17408 45404
rect 17267 45373 17279 45376
rect 17221 45367 17279 45373
rect 17402 45364 17408 45376
rect 17460 45364 17466 45416
rect 12713 45339 12771 45345
rect 12713 45336 12725 45339
rect 9048 45308 12434 45336
rect 12636 45308 12725 45336
rect 1394 45268 1400 45280
rect 1355 45240 1400 45268
rect 1394 45228 1400 45240
rect 1452 45228 1458 45280
rect 7006 45268 7012 45280
rect 6967 45240 7012 45268
rect 7006 45228 7012 45240
rect 7064 45228 7070 45280
rect 9858 45228 9864 45280
rect 9916 45268 9922 45280
rect 10413 45271 10471 45277
rect 10413 45268 10425 45271
rect 9916 45240 10425 45268
rect 9916 45228 9922 45240
rect 10413 45237 10425 45240
rect 10459 45237 10471 45271
rect 11698 45268 11704 45280
rect 11659 45240 11704 45268
rect 10413 45231 10471 45237
rect 11698 45228 11704 45240
rect 11756 45228 11762 45280
rect 12406 45268 12434 45308
rect 12713 45305 12725 45308
rect 12759 45305 12771 45339
rect 16574 45336 16580 45348
rect 12713 45299 12771 45305
rect 12820 45308 16580 45336
rect 12820 45268 12848 45308
rect 16574 45296 16580 45308
rect 16632 45296 16638 45348
rect 17788 45336 17816 45435
rect 18414 45432 18420 45444
rect 18472 45432 18478 45484
rect 18506 45432 18512 45484
rect 18564 45472 18570 45484
rect 19245 45475 19303 45481
rect 19245 45472 19257 45475
rect 18564 45444 19257 45472
rect 18564 45432 18570 45444
rect 19245 45441 19257 45444
rect 19291 45472 19303 45475
rect 20530 45472 20536 45484
rect 19291 45444 20536 45472
rect 19291 45441 19303 45444
rect 19245 45435 19303 45441
rect 20530 45432 20536 45444
rect 20588 45432 20594 45484
rect 20625 45475 20683 45481
rect 20625 45441 20637 45475
rect 20671 45472 20683 45475
rect 21082 45472 21088 45484
rect 20671 45444 21088 45472
rect 20671 45441 20683 45444
rect 20625 45435 20683 45441
rect 21082 45432 21088 45444
rect 21140 45432 21146 45484
rect 21292 45481 21320 45512
rect 21450 45500 21456 45512
rect 21508 45500 21514 45552
rect 21269 45475 21327 45481
rect 21269 45441 21281 45475
rect 21315 45441 21327 45475
rect 21269 45435 21327 45441
rect 21726 45432 21732 45484
rect 21784 45472 21790 45484
rect 21821 45475 21879 45481
rect 21821 45472 21833 45475
rect 21784 45444 21833 45472
rect 21784 45432 21790 45444
rect 21821 45441 21833 45444
rect 21867 45441 21879 45475
rect 21821 45435 21879 45441
rect 23842 45432 23848 45484
rect 23900 45472 23906 45484
rect 26142 45472 26148 45484
rect 23900 45444 23945 45472
rect 26103 45444 26148 45472
rect 23900 45432 23906 45444
rect 26142 45432 26148 45444
rect 26200 45432 26206 45484
rect 27430 45472 27436 45484
rect 27391 45444 27436 45472
rect 27430 45432 27436 45444
rect 27488 45432 27494 45484
rect 27614 45432 27620 45484
rect 27672 45472 27678 45484
rect 27709 45475 27767 45481
rect 27709 45472 27721 45475
rect 27672 45444 27721 45472
rect 27672 45432 27678 45444
rect 27709 45441 27721 45444
rect 27755 45441 27767 45475
rect 28353 45475 28411 45481
rect 28353 45472 28365 45475
rect 27709 45435 27767 45441
rect 27908 45444 28365 45472
rect 18693 45407 18751 45413
rect 18693 45373 18705 45407
rect 18739 45404 18751 45407
rect 19334 45404 19340 45416
rect 18739 45376 19340 45404
rect 18739 45373 18751 45376
rect 18693 45367 18751 45373
rect 19334 45364 19340 45376
rect 19392 45364 19398 45416
rect 20438 45364 20444 45416
rect 20496 45404 20502 45416
rect 22097 45407 22155 45413
rect 22097 45404 22109 45407
rect 20496 45376 22109 45404
rect 20496 45364 20502 45376
rect 22097 45373 22109 45376
rect 22143 45373 22155 45407
rect 22097 45367 22155 45373
rect 23198 45364 23204 45416
rect 23256 45404 23262 45416
rect 24397 45407 24455 45413
rect 24397 45404 24409 45407
rect 23256 45376 24409 45404
rect 23256 45364 23262 45376
rect 24397 45373 24409 45376
rect 24443 45373 24455 45407
rect 24397 45367 24455 45373
rect 24673 45407 24731 45413
rect 24673 45373 24685 45407
rect 24719 45373 24731 45407
rect 27522 45404 27528 45416
rect 27483 45376 27528 45404
rect 24673 45367 24731 45373
rect 16684 45308 17816 45336
rect 17865 45339 17923 45345
rect 12406 45240 12848 45268
rect 13357 45271 13415 45277
rect 13357 45237 13369 45271
rect 13403 45268 13415 45271
rect 14274 45268 14280 45280
rect 13403 45240 14280 45268
rect 13403 45237 13415 45240
rect 13357 45231 13415 45237
rect 14274 45228 14280 45240
rect 14332 45228 14338 45280
rect 14458 45268 14464 45280
rect 14419 45240 14464 45268
rect 14458 45228 14464 45240
rect 14516 45228 14522 45280
rect 15102 45268 15108 45280
rect 15063 45240 15108 45268
rect 15102 45228 15108 45240
rect 15160 45228 15166 45280
rect 15194 45228 15200 45280
rect 15252 45268 15258 45280
rect 15473 45271 15531 45277
rect 15473 45268 15485 45271
rect 15252 45240 15485 45268
rect 15252 45228 15258 45240
rect 15473 45237 15485 45240
rect 15519 45237 15531 45271
rect 15473 45231 15531 45237
rect 15654 45228 15660 45280
rect 15712 45268 15718 45280
rect 16684 45268 16712 45308
rect 17865 45305 17877 45339
rect 17911 45336 17923 45339
rect 18509 45339 18567 45345
rect 18509 45336 18521 45339
rect 17911 45308 18521 45336
rect 17911 45305 17923 45308
rect 17865 45299 17923 45305
rect 18509 45305 18521 45308
rect 18555 45336 18567 45339
rect 24688 45336 24716 45367
rect 27522 45364 27528 45376
rect 27580 45364 27586 45416
rect 18555 45308 19288 45336
rect 18555 45305 18567 45308
rect 18509 45299 18567 45305
rect 15712 45240 16712 45268
rect 15712 45228 15718 45240
rect 17034 45228 17040 45280
rect 17092 45268 17098 45280
rect 17129 45271 17187 45277
rect 17129 45268 17141 45271
rect 17092 45240 17141 45268
rect 17092 45228 17098 45240
rect 17129 45237 17141 45240
rect 17175 45237 17187 45271
rect 17129 45231 17187 45237
rect 17586 45228 17592 45280
rect 17644 45268 17650 45280
rect 19260 45277 19288 45308
rect 23216 45308 24716 45336
rect 26329 45339 26387 45345
rect 18417 45271 18475 45277
rect 18417 45268 18429 45271
rect 17644 45240 18429 45268
rect 17644 45228 17650 45240
rect 18417 45237 18429 45240
rect 18463 45237 18475 45271
rect 18417 45231 18475 45237
rect 19245 45271 19303 45277
rect 19245 45237 19257 45271
rect 19291 45268 19303 45271
rect 19426 45268 19432 45280
rect 19291 45240 19432 45268
rect 19291 45237 19303 45240
rect 19245 45231 19303 45237
rect 19426 45228 19432 45240
rect 19484 45228 19490 45280
rect 19610 45268 19616 45280
rect 19571 45240 19616 45268
rect 19610 45228 19616 45240
rect 19668 45228 19674 45280
rect 20441 45271 20499 45277
rect 20441 45237 20453 45271
rect 20487 45268 20499 45271
rect 20622 45268 20628 45280
rect 20487 45240 20628 45268
rect 20487 45237 20499 45240
rect 20441 45231 20499 45237
rect 20622 45228 20628 45240
rect 20680 45228 20686 45280
rect 20990 45228 20996 45280
rect 21048 45268 21054 45280
rect 23216 45268 23244 45308
rect 26329 45305 26341 45339
rect 26375 45336 26387 45339
rect 27706 45336 27712 45348
rect 26375 45308 27712 45336
rect 26375 45305 26387 45308
rect 26329 45299 26387 45305
rect 27706 45296 27712 45308
rect 27764 45296 27770 45348
rect 27908 45345 27936 45444
rect 28353 45441 28365 45444
rect 28399 45441 28411 45475
rect 28534 45472 28540 45484
rect 28495 45444 28540 45472
rect 28353 45435 28411 45441
rect 28534 45432 28540 45444
rect 28592 45432 28598 45484
rect 29178 45432 29184 45484
rect 29236 45472 29242 45484
rect 29825 45475 29883 45481
rect 29825 45472 29837 45475
rect 29236 45444 29837 45472
rect 29236 45432 29242 45444
rect 29825 45441 29837 45444
rect 29871 45441 29883 45475
rect 29825 45435 29883 45441
rect 27893 45339 27951 45345
rect 27893 45305 27905 45339
rect 27939 45305 27951 45339
rect 27893 45299 27951 45305
rect 21048 45240 23244 45268
rect 23661 45271 23719 45277
rect 21048 45228 21054 45240
rect 23661 45237 23673 45271
rect 23707 45268 23719 45271
rect 27154 45268 27160 45280
rect 23707 45240 27160 45268
rect 23707 45237 23719 45240
rect 23661 45231 23719 45237
rect 27154 45228 27160 45240
rect 27212 45228 27218 45280
rect 27246 45228 27252 45280
rect 27304 45268 27310 45280
rect 27433 45271 27491 45277
rect 27433 45268 27445 45271
rect 27304 45240 27445 45268
rect 27304 45228 27310 45240
rect 27433 45237 27445 45240
rect 27479 45237 27491 45271
rect 27433 45231 27491 45237
rect 27522 45228 27528 45280
rect 27580 45268 27586 45280
rect 28721 45271 28779 45277
rect 28721 45268 28733 45271
rect 27580 45240 28733 45268
rect 27580 45228 27586 45240
rect 28721 45237 28733 45240
rect 28767 45237 28779 45271
rect 28721 45231 28779 45237
rect 1104 45178 30820 45200
rect 1104 45126 5915 45178
rect 5967 45126 5979 45178
rect 6031 45126 6043 45178
rect 6095 45126 6107 45178
rect 6159 45126 6171 45178
rect 6223 45126 15846 45178
rect 15898 45126 15910 45178
rect 15962 45126 15974 45178
rect 16026 45126 16038 45178
rect 16090 45126 16102 45178
rect 16154 45126 25776 45178
rect 25828 45126 25840 45178
rect 25892 45126 25904 45178
rect 25956 45126 25968 45178
rect 26020 45126 26032 45178
rect 26084 45126 30820 45178
rect 1104 45104 30820 45126
rect 8938 45024 8944 45076
rect 8996 45064 9002 45076
rect 11885 45067 11943 45073
rect 8996 45036 11376 45064
rect 8996 45024 9002 45036
rect 9766 44956 9772 45008
rect 9824 44996 9830 45008
rect 10505 44999 10563 45005
rect 10505 44996 10517 44999
rect 9824 44968 10517 44996
rect 9824 44956 9830 44968
rect 10505 44965 10517 44968
rect 10551 44965 10563 44999
rect 10505 44959 10563 44965
rect 1394 44888 1400 44940
rect 1452 44928 1458 44940
rect 11238 44928 11244 44940
rect 1452 44900 11244 44928
rect 1452 44888 1458 44900
rect 11238 44888 11244 44900
rect 11296 44888 11302 44940
rect 11348 44928 11376 45036
rect 11885 45033 11897 45067
rect 11931 45064 11943 45067
rect 13906 45064 13912 45076
rect 11931 45036 13912 45064
rect 11931 45033 11943 45036
rect 11885 45027 11943 45033
rect 13906 45024 13912 45036
rect 13964 45024 13970 45076
rect 14734 45024 14740 45076
rect 14792 45064 14798 45076
rect 15010 45064 15016 45076
rect 14792 45036 15016 45064
rect 14792 45024 14798 45036
rect 15010 45024 15016 45036
rect 15068 45064 15074 45076
rect 15473 45067 15531 45073
rect 15473 45064 15485 45067
rect 15068 45036 15485 45064
rect 15068 45024 15074 45036
rect 15473 45033 15485 45036
rect 15519 45033 15531 45067
rect 16574 45064 16580 45076
rect 16535 45036 16580 45064
rect 15473 45027 15531 45033
rect 16574 45024 16580 45036
rect 16632 45024 16638 45076
rect 16942 45024 16948 45076
rect 17000 45064 17006 45076
rect 17589 45067 17647 45073
rect 17589 45064 17601 45067
rect 17000 45036 17601 45064
rect 17000 45024 17006 45036
rect 17589 45033 17601 45036
rect 17635 45033 17647 45067
rect 20714 45064 20720 45076
rect 20675 45036 20720 45064
rect 17589 45027 17647 45033
rect 20714 45024 20720 45036
rect 20772 45024 20778 45076
rect 21082 45024 21088 45076
rect 21140 45064 21146 45076
rect 21140 45036 22324 45064
rect 21140 45024 21146 45036
rect 12621 44999 12679 45005
rect 12621 44965 12633 44999
rect 12667 44996 12679 44999
rect 14366 44996 14372 45008
rect 12667 44968 14372 44996
rect 12667 44965 12679 44968
rect 12621 44959 12679 44965
rect 14366 44956 14372 44968
rect 14424 44956 14430 45008
rect 14458 44956 14464 45008
rect 14516 44996 14522 45008
rect 15933 44999 15991 45005
rect 14516 44968 15608 44996
rect 14516 44956 14522 44968
rect 15580 44937 15608 44968
rect 15933 44965 15945 44999
rect 15979 44996 15991 44999
rect 18049 44999 18107 45005
rect 18049 44996 18061 44999
rect 15979 44968 16712 44996
rect 15979 44965 15991 44968
rect 15933 44959 15991 44965
rect 15565 44931 15623 44937
rect 11348 44900 15516 44928
rect 1854 44820 1860 44872
rect 1912 44860 1918 44872
rect 2041 44863 2099 44869
rect 2041 44860 2053 44863
rect 1912 44832 2053 44860
rect 1912 44820 1918 44832
rect 2041 44829 2053 44832
rect 2087 44829 2099 44863
rect 2041 44823 2099 44829
rect 4890 44820 4896 44872
rect 4948 44860 4954 44872
rect 5077 44863 5135 44869
rect 5077 44860 5089 44863
rect 4948 44832 5089 44860
rect 4948 44820 4954 44832
rect 5077 44829 5089 44832
rect 5123 44829 5135 44863
rect 5077 44823 5135 44829
rect 7190 44820 7196 44872
rect 7248 44860 7254 44872
rect 7469 44863 7527 44869
rect 7469 44860 7481 44863
rect 7248 44832 7481 44860
rect 7248 44820 7254 44832
rect 7469 44829 7481 44832
rect 7515 44829 7527 44863
rect 7469 44823 7527 44829
rect 10226 44820 10232 44872
rect 10284 44860 10290 44872
rect 10321 44863 10379 44869
rect 10321 44860 10333 44863
rect 10284 44832 10333 44860
rect 10284 44820 10290 44832
rect 10321 44829 10333 44832
rect 10367 44829 10379 44863
rect 10321 44823 10379 44829
rect 11790 44820 11796 44872
rect 11848 44860 11854 44872
rect 12069 44863 12127 44869
rect 12069 44860 12081 44863
rect 11848 44832 12081 44860
rect 11848 44820 11854 44832
rect 12069 44829 12081 44832
rect 12115 44829 12127 44863
rect 12069 44823 12127 44829
rect 12526 44820 12532 44872
rect 12584 44860 12590 44872
rect 12805 44863 12863 44869
rect 12805 44860 12817 44863
rect 12584 44832 12817 44860
rect 12584 44820 12590 44832
rect 12805 44829 12817 44832
rect 12851 44829 12863 44863
rect 13538 44860 13544 44872
rect 13499 44832 13544 44860
rect 12805 44823 12863 44829
rect 13538 44820 13544 44832
rect 13596 44820 13602 44872
rect 14734 44860 14740 44872
rect 14695 44832 14740 44860
rect 14734 44820 14740 44832
rect 14792 44820 14798 44872
rect 14918 44860 14924 44872
rect 14879 44832 14924 44860
rect 14918 44820 14924 44832
rect 14976 44820 14982 44872
rect 15013 44863 15071 44869
rect 15013 44829 15025 44863
rect 15059 44862 15071 44863
rect 15059 44860 15148 44862
rect 15488 44860 15516 44900
rect 15565 44897 15577 44931
rect 15611 44928 15623 44931
rect 16206 44928 16212 44940
rect 15611 44900 16212 44928
rect 15611 44897 15623 44900
rect 15565 44891 15623 44897
rect 16206 44888 16212 44900
rect 16264 44888 16270 44940
rect 16684 44937 16712 44968
rect 16776 44968 18061 44996
rect 16669 44931 16727 44937
rect 16669 44897 16681 44931
rect 16715 44897 16727 44931
rect 16669 44891 16727 44897
rect 15746 44860 15752 44872
rect 15059 44834 15240 44860
rect 15059 44829 15071 44834
rect 15120 44832 15240 44834
rect 15488 44832 15608 44860
rect 15707 44832 15752 44860
rect 15013 44823 15071 44829
rect 2406 44792 2412 44804
rect 2367 44764 2412 44792
rect 2406 44752 2412 44764
rect 2464 44752 2470 44804
rect 14642 44792 14648 44804
rect 13372 44764 14648 44792
rect 5166 44724 5172 44736
rect 5127 44696 5172 44724
rect 5166 44684 5172 44696
rect 5224 44684 5230 44736
rect 7285 44727 7343 44733
rect 7285 44693 7297 44727
rect 7331 44724 7343 44727
rect 10042 44724 10048 44736
rect 7331 44696 10048 44724
rect 7331 44693 7343 44696
rect 7285 44687 7343 44693
rect 10042 44684 10048 44696
rect 10100 44684 10106 44736
rect 13372 44733 13400 44764
rect 14642 44752 14648 44764
rect 14700 44752 14706 44804
rect 13357 44727 13415 44733
rect 13357 44693 13369 44727
rect 13403 44693 13415 44727
rect 13357 44687 13415 44693
rect 13446 44684 13452 44736
rect 13504 44724 13510 44736
rect 14458 44724 14464 44736
rect 13504 44696 14464 44724
rect 13504 44684 13510 44696
rect 14458 44684 14464 44696
rect 14516 44684 14522 44736
rect 14553 44727 14611 44733
rect 14553 44693 14565 44727
rect 14599 44724 14611 44727
rect 14918 44724 14924 44736
rect 14599 44696 14924 44724
rect 14599 44693 14611 44696
rect 14553 44687 14611 44693
rect 14918 44684 14924 44696
rect 14976 44684 14982 44736
rect 15212 44724 15240 44832
rect 15286 44752 15292 44804
rect 15344 44792 15350 44804
rect 15473 44795 15531 44801
rect 15473 44792 15485 44795
rect 15344 44764 15485 44792
rect 15344 44752 15350 44764
rect 15473 44761 15485 44764
rect 15519 44761 15531 44795
rect 15580 44792 15608 44832
rect 15746 44820 15752 44832
rect 15804 44820 15810 44872
rect 16577 44863 16635 44869
rect 16577 44829 16589 44863
rect 16623 44860 16635 44863
rect 16776 44860 16804 44968
rect 18049 44965 18061 44968
rect 18095 44965 18107 44999
rect 18049 44959 18107 44965
rect 19242 44956 19248 45008
rect 19300 44996 19306 45008
rect 22186 44996 22192 45008
rect 19300 44968 22192 44996
rect 19300 44956 19306 44968
rect 22186 44956 22192 44968
rect 22244 44956 22250 45008
rect 22296 44996 22324 45036
rect 22370 45024 22376 45076
rect 22428 45064 22434 45076
rect 27522 45064 27528 45076
rect 22428 45036 27528 45064
rect 22428 45024 22434 45036
rect 27522 45024 27528 45036
rect 27580 45024 27586 45076
rect 28258 45064 28264 45076
rect 28219 45036 28264 45064
rect 28258 45024 28264 45036
rect 28316 45024 28322 45076
rect 28445 44999 28503 45005
rect 28445 44996 28457 44999
rect 22296 44968 25268 44996
rect 17218 44888 17224 44940
rect 17276 44928 17282 44940
rect 17681 44931 17739 44937
rect 17681 44928 17693 44931
rect 17276 44900 17693 44928
rect 17276 44888 17282 44900
rect 17681 44897 17693 44900
rect 17727 44928 17739 44931
rect 17727 44900 18092 44928
rect 17727 44897 17739 44900
rect 17681 44891 17739 44897
rect 18064 44872 18092 44900
rect 18414 44888 18420 44940
rect 18472 44928 18478 44940
rect 19705 44931 19763 44937
rect 19705 44928 19717 44931
rect 18472 44900 19717 44928
rect 18472 44888 18478 44900
rect 19705 44897 19717 44900
rect 19751 44928 19763 44931
rect 19978 44928 19984 44940
rect 19751 44900 19984 44928
rect 19751 44897 19763 44900
rect 19705 44891 19763 44897
rect 19978 44888 19984 44900
rect 20036 44888 20042 44940
rect 21450 44928 21456 44940
rect 20640 44900 21456 44928
rect 16623 44832 16804 44860
rect 16623 44829 16635 44832
rect 16577 44823 16635 44829
rect 16850 44820 16856 44872
rect 16908 44860 16914 44872
rect 16908 44832 16953 44860
rect 17052 44832 17724 44860
rect 16908 44820 16914 44832
rect 17052 44792 17080 44832
rect 15580 44764 17080 44792
rect 15473 44755 15531 44761
rect 17310 44752 17316 44804
rect 17368 44792 17374 44804
rect 17589 44795 17647 44801
rect 17589 44792 17601 44795
rect 17368 44764 17601 44792
rect 17368 44752 17374 44764
rect 17589 44761 17601 44764
rect 17635 44761 17647 44795
rect 17696 44792 17724 44832
rect 17770 44820 17776 44872
rect 17828 44860 17834 44872
rect 17865 44863 17923 44869
rect 17865 44860 17877 44863
rect 17828 44832 17877 44860
rect 17828 44820 17834 44832
rect 17865 44829 17877 44832
rect 17911 44829 17923 44863
rect 17865 44823 17923 44829
rect 18046 44820 18052 44872
rect 18104 44820 18110 44872
rect 18509 44863 18567 44869
rect 18509 44829 18521 44863
rect 18555 44829 18567 44863
rect 19886 44860 19892 44872
rect 19847 44832 19892 44860
rect 18509 44823 18567 44829
rect 18524 44792 18552 44823
rect 19886 44820 19892 44832
rect 19944 44820 19950 44872
rect 20640 44869 20668 44900
rect 21450 44888 21456 44900
rect 21508 44888 21514 44940
rect 22370 44928 22376 44940
rect 21744 44900 22376 44928
rect 20625 44863 20683 44869
rect 20625 44829 20637 44863
rect 20671 44829 20683 44863
rect 20990 44860 20996 44872
rect 20951 44832 20996 44860
rect 20625 44823 20683 44829
rect 20990 44820 20996 44832
rect 21048 44820 21054 44872
rect 21085 44863 21143 44869
rect 21085 44829 21097 44863
rect 21131 44856 21143 44863
rect 21131 44829 21146 44856
rect 21085 44823 21146 44829
rect 17696 44764 18552 44792
rect 21118 44792 21146 44823
rect 21450 44792 21456 44804
rect 21118 44764 21456 44792
rect 17589 44755 17647 44761
rect 21450 44752 21456 44764
rect 21508 44752 21514 44804
rect 21634 44752 21640 44804
rect 21692 44792 21698 44804
rect 21744 44792 21772 44900
rect 22370 44888 22376 44900
rect 22428 44888 22434 44940
rect 22462 44888 22468 44940
rect 22520 44928 22526 44940
rect 22557 44931 22615 44937
rect 22557 44928 22569 44931
rect 22520 44900 22569 44928
rect 22520 44888 22526 44900
rect 22557 44897 22569 44900
rect 22603 44897 22615 44931
rect 22557 44891 22615 44897
rect 23934 44888 23940 44940
rect 23992 44928 23998 44940
rect 24397 44931 24455 44937
rect 24397 44928 24409 44931
rect 23992 44900 24409 44928
rect 23992 44888 23998 44900
rect 24397 44897 24409 44900
rect 24443 44897 24455 44931
rect 25240 44928 25268 44968
rect 26896 44968 28457 44996
rect 25240 44900 26004 44928
rect 24397 44891 24455 44897
rect 21910 44869 21916 44872
rect 21905 44823 21916 44869
rect 21968 44860 21974 44872
rect 22830 44860 22836 44872
rect 21968 44832 22005 44860
rect 22791 44832 22836 44860
rect 21910 44820 21916 44823
rect 21968 44820 21974 44832
rect 22830 44820 22836 44832
rect 22888 44820 22894 44872
rect 24673 44863 24731 44869
rect 24673 44829 24685 44863
rect 24719 44829 24731 44863
rect 24673 44823 24731 44829
rect 21692 44764 21772 44792
rect 21692 44752 21698 44764
rect 22186 44752 22192 44804
rect 22244 44792 22250 44804
rect 24688 44792 24716 44823
rect 25038 44820 25044 44872
rect 25096 44860 25102 44872
rect 25869 44863 25927 44869
rect 25869 44860 25881 44863
rect 25096 44832 25881 44860
rect 25096 44820 25102 44832
rect 25869 44829 25881 44832
rect 25915 44829 25927 44863
rect 25976 44860 26004 44900
rect 26896 44860 26924 44968
rect 28445 44965 28457 44968
rect 28491 44965 28503 44999
rect 28445 44959 28503 44965
rect 27154 44888 27160 44940
rect 27212 44928 27218 44940
rect 27212 44900 29868 44928
rect 27212 44888 27218 44900
rect 25976 44832 26924 44860
rect 27893 44863 27951 44869
rect 25869 44823 25927 44829
rect 27893 44829 27905 44863
rect 27939 44860 27951 44863
rect 28074 44860 28080 44872
rect 27939 44832 28080 44860
rect 27939 44829 27951 44832
rect 27893 44823 27951 44829
rect 28074 44820 28080 44832
rect 28132 44820 28138 44872
rect 29840 44869 29868 44900
rect 29825 44863 29883 44869
rect 29825 44829 29837 44863
rect 29871 44829 29883 44863
rect 29825 44823 29883 44829
rect 22244 44764 24716 44792
rect 26136 44795 26194 44801
rect 22244 44752 22250 44764
rect 26136 44761 26148 44795
rect 26182 44792 26194 44795
rect 26326 44792 26332 44804
rect 26182 44764 26332 44792
rect 26182 44761 26194 44764
rect 26136 44755 26194 44761
rect 26326 44752 26332 44764
rect 26384 44752 26390 44804
rect 28261 44795 28319 44801
rect 28261 44792 28273 44795
rect 26436 44764 28273 44792
rect 16666 44724 16672 44736
rect 15212 44696 16672 44724
rect 16666 44684 16672 44696
rect 16724 44684 16730 44736
rect 17037 44727 17095 44733
rect 17037 44693 17049 44727
rect 17083 44724 17095 44727
rect 17862 44724 17868 44736
rect 17083 44696 17868 44724
rect 17083 44693 17095 44696
rect 17037 44687 17095 44693
rect 17862 44684 17868 44696
rect 17920 44684 17926 44736
rect 18601 44727 18659 44733
rect 18601 44693 18613 44727
rect 18647 44724 18659 44727
rect 19334 44724 19340 44736
rect 18647 44696 19340 44724
rect 18647 44693 18659 44696
rect 18601 44687 18659 44693
rect 19334 44684 19340 44696
rect 19392 44684 19398 44736
rect 20070 44724 20076 44736
rect 20031 44696 20076 44724
rect 20070 44684 20076 44696
rect 20128 44684 20134 44736
rect 21266 44724 21272 44736
rect 21227 44696 21272 44724
rect 21266 44684 21272 44696
rect 21324 44684 21330 44736
rect 21729 44727 21787 44733
rect 21729 44693 21741 44727
rect 21775 44724 21787 44727
rect 22094 44724 22100 44736
rect 21775 44696 22100 44724
rect 21775 44693 21787 44696
rect 21729 44687 21787 44693
rect 22094 44684 22100 44696
rect 22152 44684 22158 44736
rect 25314 44684 25320 44736
rect 25372 44724 25378 44736
rect 26436 44724 26464 44764
rect 28261 44761 28273 44764
rect 28307 44761 28319 44795
rect 28261 44755 28319 44761
rect 25372 44696 26464 44724
rect 25372 44684 25378 44696
rect 26786 44684 26792 44736
rect 26844 44724 26850 44736
rect 27249 44727 27307 44733
rect 27249 44724 27261 44727
rect 26844 44696 27261 44724
rect 26844 44684 26850 44696
rect 27249 44693 27261 44696
rect 27295 44724 27307 44727
rect 27522 44724 27528 44736
rect 27295 44696 27528 44724
rect 27295 44693 27307 44696
rect 27249 44687 27307 44693
rect 27522 44684 27528 44696
rect 27580 44684 27586 44736
rect 30006 44724 30012 44736
rect 29967 44696 30012 44724
rect 30006 44684 30012 44696
rect 30064 44684 30070 44736
rect 1104 44634 30820 44656
rect 1104 44582 10880 44634
rect 10932 44582 10944 44634
rect 10996 44582 11008 44634
rect 11060 44582 11072 44634
rect 11124 44582 11136 44634
rect 11188 44582 20811 44634
rect 20863 44582 20875 44634
rect 20927 44582 20939 44634
rect 20991 44582 21003 44634
rect 21055 44582 21067 44634
rect 21119 44582 30820 44634
rect 1104 44560 30820 44582
rect 5166 44480 5172 44532
rect 5224 44520 5230 44532
rect 12618 44520 12624 44532
rect 5224 44492 12624 44520
rect 5224 44480 5230 44492
rect 12618 44480 12624 44492
rect 12676 44480 12682 44532
rect 15654 44520 15660 44532
rect 13096 44492 15660 44520
rect 2774 44452 2780 44464
rect 1596 44424 2780 44452
rect 1596 44393 1624 44424
rect 2774 44412 2780 44424
rect 2832 44412 2838 44464
rect 1581 44387 1639 44393
rect 1581 44353 1593 44387
rect 1627 44353 1639 44387
rect 2038 44384 2044 44396
rect 1999 44356 2044 44384
rect 1581 44347 1639 44353
rect 2038 44344 2044 44356
rect 2096 44344 2102 44396
rect 2225 44387 2283 44393
rect 2225 44353 2237 44387
rect 2271 44384 2283 44387
rect 2406 44384 2412 44396
rect 2271 44356 2412 44384
rect 2271 44353 2283 44356
rect 2225 44347 2283 44353
rect 2406 44344 2412 44356
rect 2464 44344 2470 44396
rect 2590 44316 2596 44328
rect 2551 44288 2596 44316
rect 2590 44276 2596 44288
rect 2648 44276 2654 44328
rect 2682 44276 2688 44328
rect 2740 44316 2746 44328
rect 13096 44316 13124 44492
rect 15654 44480 15660 44492
rect 15712 44480 15718 44532
rect 15933 44523 15991 44529
rect 15933 44489 15945 44523
rect 15979 44489 15991 44523
rect 15933 44483 15991 44489
rect 17037 44523 17095 44529
rect 17037 44489 17049 44523
rect 17083 44520 17095 44523
rect 17494 44520 17500 44532
rect 17083 44492 17500 44520
rect 17083 44489 17095 44492
rect 17037 44483 17095 44489
rect 14918 44452 14924 44464
rect 14879 44424 14924 44452
rect 14918 44412 14924 44424
rect 14976 44412 14982 44464
rect 15948 44452 15976 44483
rect 17494 44480 17500 44492
rect 17552 44480 17558 44532
rect 27341 44523 27399 44529
rect 17696 44492 27200 44520
rect 17696 44452 17724 44492
rect 17862 44452 17868 44464
rect 15948 44424 17724 44452
rect 17823 44424 17868 44452
rect 17862 44412 17868 44424
rect 17920 44412 17926 44464
rect 18049 44455 18107 44461
rect 18049 44421 18061 44455
rect 18095 44452 18107 44455
rect 18506 44452 18512 44464
rect 18095 44424 18512 44452
rect 18095 44421 18107 44424
rect 18049 44415 18107 44421
rect 18506 44412 18512 44424
rect 18564 44412 18570 44464
rect 18690 44412 18696 44464
rect 18748 44452 18754 44464
rect 18748 44424 19840 44452
rect 18748 44412 18754 44424
rect 13173 44387 13231 44393
rect 13173 44353 13185 44387
rect 13219 44384 13231 44387
rect 13449 44387 13507 44393
rect 13449 44384 13461 44387
rect 13219 44356 13461 44384
rect 13219 44353 13231 44356
rect 13173 44347 13231 44353
rect 13449 44353 13461 44356
rect 13495 44384 13507 44387
rect 13998 44384 14004 44396
rect 13495 44356 14004 44384
rect 13495 44353 13507 44356
rect 13449 44347 13507 44353
rect 13998 44344 14004 44356
rect 14056 44344 14062 44396
rect 14093 44387 14151 44393
rect 14093 44353 14105 44387
rect 14139 44384 14151 44387
rect 14182 44384 14188 44396
rect 14139 44356 14188 44384
rect 14139 44353 14151 44356
rect 14093 44347 14151 44353
rect 14182 44344 14188 44356
rect 14240 44344 14246 44396
rect 16117 44387 16175 44393
rect 16117 44353 16129 44387
rect 16163 44384 16175 44387
rect 16390 44384 16396 44396
rect 16163 44356 16396 44384
rect 16163 44353 16175 44356
rect 16117 44347 16175 44353
rect 16390 44344 16396 44356
rect 16448 44344 16454 44396
rect 16482 44344 16488 44396
rect 16540 44384 16546 44396
rect 18969 44387 19027 44393
rect 16540 44356 17356 44384
rect 16540 44344 16546 44356
rect 2740 44288 13124 44316
rect 2740 44276 2746 44288
rect 15010 44276 15016 44328
rect 15068 44316 15074 44328
rect 15068 44288 15113 44316
rect 15068 44276 15074 44288
rect 15194 44276 15200 44328
rect 15252 44316 15258 44328
rect 15252 44288 15297 44316
rect 15252 44276 15258 44288
rect 16758 44276 16764 44328
rect 16816 44316 16822 44328
rect 16942 44316 16948 44328
rect 16816 44288 16948 44316
rect 16816 44276 16822 44288
rect 16942 44276 16948 44288
rect 17000 44316 17006 44328
rect 17328 44325 17356 44356
rect 18969 44353 18981 44387
rect 19015 44384 19027 44387
rect 19334 44384 19340 44396
rect 19015 44356 19340 44384
rect 19015 44353 19027 44356
rect 18969 44347 19027 44353
rect 19334 44344 19340 44356
rect 19392 44344 19398 44396
rect 19521 44387 19579 44393
rect 19521 44353 19533 44387
rect 19567 44384 19579 44387
rect 19702 44384 19708 44396
rect 19567 44356 19708 44384
rect 19567 44353 19579 44356
rect 19521 44347 19579 44353
rect 19702 44344 19708 44356
rect 19760 44344 19766 44396
rect 17129 44319 17187 44325
rect 17129 44316 17141 44319
rect 17000 44288 17141 44316
rect 17000 44276 17006 44288
rect 17129 44285 17141 44288
rect 17175 44285 17187 44319
rect 17129 44279 17187 44285
rect 17313 44319 17371 44325
rect 17313 44285 17325 44319
rect 17359 44316 17371 44319
rect 19426 44316 19432 44328
rect 17359 44288 19288 44316
rect 19387 44288 19432 44316
rect 17359 44285 17371 44288
rect 17313 44279 17371 44285
rect 1397 44251 1455 44257
rect 1397 44217 1409 44251
rect 1443 44248 1455 44251
rect 10870 44248 10876 44260
rect 1443 44220 10876 44248
rect 1443 44217 1455 44220
rect 1397 44211 1455 44217
rect 10870 44208 10876 44220
rect 10928 44208 10934 44260
rect 13265 44251 13323 44257
rect 13265 44217 13277 44251
rect 13311 44248 13323 44251
rect 18690 44248 18696 44260
rect 13311 44220 18696 44248
rect 13311 44217 13323 44220
rect 13265 44211 13323 44217
rect 18690 44208 18696 44220
rect 18748 44208 18754 44260
rect 19260 44248 19288 44288
rect 19426 44276 19432 44288
rect 19484 44276 19490 44328
rect 19521 44251 19579 44257
rect 19521 44248 19533 44251
rect 19260 44220 19533 44248
rect 19521 44217 19533 44220
rect 19567 44217 19579 44251
rect 19812 44248 19840 44424
rect 19886 44412 19892 44464
rect 19944 44452 19950 44464
rect 22189 44455 22247 44461
rect 22189 44452 22201 44455
rect 19944 44424 22201 44452
rect 19944 44412 19950 44424
rect 22189 44421 22201 44424
rect 22235 44421 22247 44455
rect 22189 44415 22247 44421
rect 20254 44384 20260 44396
rect 20215 44356 20260 44384
rect 20254 44344 20260 44356
rect 20312 44344 20318 44396
rect 20717 44387 20775 44393
rect 20717 44353 20729 44387
rect 20763 44353 20775 44387
rect 20717 44347 20775 44353
rect 20346 44276 20352 44328
rect 20404 44316 20410 44328
rect 20533 44319 20591 44325
rect 20533 44316 20545 44319
rect 20404 44288 20545 44316
rect 20404 44276 20410 44288
rect 20533 44285 20545 44288
rect 20579 44285 20591 44319
rect 20732 44316 20760 44347
rect 21174 44344 21180 44396
rect 21232 44384 21238 44396
rect 21634 44384 21640 44396
rect 21232 44356 21640 44384
rect 21232 44344 21238 44356
rect 21634 44344 21640 44356
rect 21692 44384 21698 44396
rect 21821 44387 21879 44393
rect 21821 44384 21833 44387
rect 21692 44356 21833 44384
rect 21692 44344 21698 44356
rect 21821 44353 21833 44356
rect 21867 44353 21879 44387
rect 22002 44384 22008 44396
rect 21963 44356 22008 44384
rect 21821 44347 21879 44353
rect 22002 44344 22008 44356
rect 22060 44344 22066 44396
rect 22922 44384 22928 44396
rect 22883 44356 22928 44384
rect 22922 44344 22928 44356
rect 22980 44344 22986 44396
rect 23836 44387 23894 44393
rect 23836 44353 23848 44387
rect 23882 44384 23894 44387
rect 23882 44356 24808 44384
rect 23882 44353 23894 44356
rect 23836 44347 23894 44353
rect 20806 44316 20812 44328
rect 20719 44288 20812 44316
rect 20533 44279 20591 44285
rect 20806 44276 20812 44288
rect 20864 44316 20870 44328
rect 21726 44316 21732 44328
rect 20864 44288 21732 44316
rect 20864 44276 20870 44288
rect 21726 44276 21732 44288
rect 21784 44276 21790 44328
rect 22094 44276 22100 44328
rect 22152 44316 22158 44328
rect 23382 44316 23388 44328
rect 22152 44288 23388 44316
rect 22152 44276 22158 44288
rect 23382 44276 23388 44288
rect 23440 44276 23446 44328
rect 23566 44316 23572 44328
rect 23527 44288 23572 44316
rect 23566 44276 23572 44288
rect 23624 44276 23630 44328
rect 24780 44316 24808 44356
rect 24854 44344 24860 44396
rect 24912 44384 24918 44396
rect 25409 44387 25467 44393
rect 25409 44384 25421 44387
rect 24912 44356 25421 44384
rect 24912 44344 24918 44356
rect 25409 44353 25421 44356
rect 25455 44353 25467 44387
rect 25682 44384 25688 44396
rect 25643 44356 25688 44384
rect 25409 44347 25467 44353
rect 25682 44344 25688 44356
rect 25740 44344 25746 44396
rect 27172 44393 27200 44492
rect 27341 44489 27353 44523
rect 27387 44489 27399 44523
rect 27341 44483 27399 44489
rect 27356 44452 27384 44483
rect 27522 44480 27528 44532
rect 27580 44520 27586 44532
rect 28261 44523 28319 44529
rect 28261 44520 28273 44523
rect 27580 44492 28273 44520
rect 27580 44480 27586 44492
rect 28261 44489 28273 44492
rect 28307 44489 28319 44523
rect 28442 44520 28448 44532
rect 28403 44492 28448 44520
rect 28261 44483 28319 44489
rect 28442 44480 28448 44492
rect 28500 44480 28506 44532
rect 28534 44480 28540 44532
rect 28592 44520 28598 44532
rect 30101 44523 30159 44529
rect 30101 44520 30113 44523
rect 28592 44492 30113 44520
rect 28592 44480 28598 44492
rect 30101 44489 30113 44492
rect 30147 44489 30159 44523
rect 30101 44483 30159 44489
rect 27890 44452 27896 44464
rect 27356 44424 27896 44452
rect 27890 44412 27896 44424
rect 27948 44412 27954 44464
rect 27157 44387 27215 44393
rect 27157 44353 27169 44387
rect 27203 44353 27215 44387
rect 29546 44384 29552 44396
rect 29507 44356 29552 44384
rect 27157 44347 27215 44353
rect 29546 44344 29552 44356
rect 29604 44344 29610 44396
rect 29914 44384 29920 44396
rect 29875 44356 29920 44384
rect 29914 44344 29920 44356
rect 29972 44344 29978 44396
rect 25130 44316 25136 44328
rect 24780 44288 25136 44316
rect 25130 44276 25136 44288
rect 25188 44276 25194 44328
rect 29457 44319 29515 44325
rect 29457 44316 29469 44319
rect 25792 44288 29469 44316
rect 25792 44248 25820 44288
rect 29457 44285 29469 44288
rect 29503 44285 29515 44319
rect 29457 44279 29515 44285
rect 19812 44220 23612 44248
rect 19521 44211 19579 44217
rect 13909 44183 13967 44189
rect 13909 44149 13921 44183
rect 13955 44180 13967 44183
rect 14182 44180 14188 44192
rect 13955 44152 14188 44180
rect 13955 44149 13967 44152
rect 13909 44143 13967 44149
rect 14182 44140 14188 44152
rect 14240 44140 14246 44192
rect 14553 44183 14611 44189
rect 14553 44149 14565 44183
rect 14599 44180 14611 44183
rect 14734 44180 14740 44192
rect 14599 44152 14740 44180
rect 14599 44149 14611 44152
rect 14553 44143 14611 44149
rect 14734 44140 14740 44152
rect 14792 44140 14798 44192
rect 16298 44140 16304 44192
rect 16356 44180 16362 44192
rect 16669 44183 16727 44189
rect 16669 44180 16681 44183
rect 16356 44152 16681 44180
rect 16356 44140 16362 44152
rect 16669 44149 16681 44152
rect 16715 44149 16727 44183
rect 16669 44143 16727 44149
rect 17310 44140 17316 44192
rect 17368 44180 17374 44192
rect 17954 44180 17960 44192
rect 17368 44152 17960 44180
rect 17368 44140 17374 44152
rect 17954 44140 17960 44152
rect 18012 44140 18018 44192
rect 18141 44183 18199 44189
rect 18141 44149 18153 44183
rect 18187 44180 18199 44183
rect 18966 44180 18972 44192
rect 18187 44152 18972 44180
rect 18187 44149 18199 44152
rect 18141 44143 18199 44149
rect 18966 44140 18972 44152
rect 19024 44140 19030 44192
rect 20438 44180 20444 44192
rect 20399 44152 20444 44180
rect 20438 44140 20444 44152
rect 20496 44140 20502 44192
rect 20714 44140 20720 44192
rect 20772 44180 20778 44192
rect 20901 44183 20959 44189
rect 20901 44180 20913 44183
rect 20772 44152 20913 44180
rect 20772 44140 20778 44152
rect 20901 44149 20913 44152
rect 20947 44149 20959 44183
rect 20901 44143 20959 44149
rect 21726 44140 21732 44192
rect 21784 44180 21790 44192
rect 22830 44180 22836 44192
rect 21784 44152 22836 44180
rect 21784 44140 21790 44152
rect 22830 44140 22836 44152
rect 22888 44140 22894 44192
rect 23106 44180 23112 44192
rect 23067 44152 23112 44180
rect 23106 44140 23112 44152
rect 23164 44140 23170 44192
rect 23584 44180 23612 44220
rect 24504 44220 25820 44248
rect 27893 44251 27951 44257
rect 24504 44180 24532 44220
rect 27893 44217 27905 44251
rect 27939 44248 27951 44251
rect 28074 44248 28080 44260
rect 27939 44220 28080 44248
rect 27939 44217 27951 44220
rect 27893 44211 27951 44217
rect 28074 44208 28080 44220
rect 28132 44208 28138 44260
rect 28994 44248 29000 44260
rect 28184 44220 29000 44248
rect 24946 44180 24952 44192
rect 23584 44152 24532 44180
rect 24907 44152 24952 44180
rect 24946 44140 24952 44152
rect 25004 44140 25010 44192
rect 25222 44140 25228 44192
rect 25280 44180 25286 44192
rect 28184 44180 28212 44220
rect 28994 44208 29000 44220
rect 29052 44208 29058 44260
rect 25280 44152 28212 44180
rect 25280 44140 25286 44152
rect 28258 44140 28264 44192
rect 28316 44180 28322 44192
rect 28316 44152 28361 44180
rect 28316 44140 28322 44152
rect 29638 44140 29644 44192
rect 29696 44180 29702 44192
rect 29825 44183 29883 44189
rect 29825 44180 29837 44183
rect 29696 44152 29837 44180
rect 29696 44140 29702 44152
rect 29825 44149 29837 44152
rect 29871 44149 29883 44183
rect 29825 44143 29883 44149
rect 31570 44112 31576 44124
rect 1104 44090 30820 44112
rect 1104 44038 5915 44090
rect 5967 44038 5979 44090
rect 6031 44038 6043 44090
rect 6095 44038 6107 44090
rect 6159 44038 6171 44090
rect 6223 44038 15846 44090
rect 15898 44038 15910 44090
rect 15962 44038 15974 44090
rect 16026 44038 16038 44090
rect 16090 44038 16102 44090
rect 16154 44038 25776 44090
rect 25828 44038 25840 44090
rect 25892 44038 25904 44090
rect 25956 44038 25968 44090
rect 26020 44038 26032 44090
rect 26084 44038 30820 44090
rect 31531 44084 31576 44112
rect 31570 44072 31576 44084
rect 31628 44072 31634 44124
rect 1104 44016 30820 44038
rect 1397 43979 1455 43985
rect 1397 43945 1409 43979
rect 1443 43976 1455 43979
rect 2038 43976 2044 43988
rect 1443 43948 2044 43976
rect 1443 43945 1455 43948
rect 1397 43939 1455 43945
rect 2038 43936 2044 43948
rect 2096 43936 2102 43988
rect 13814 43936 13820 43988
rect 13872 43976 13878 43988
rect 18598 43976 18604 43988
rect 13872 43948 18604 43976
rect 13872 43936 13878 43948
rect 18598 43936 18604 43948
rect 18656 43936 18662 43988
rect 19426 43976 19432 43988
rect 19387 43948 19432 43976
rect 19426 43936 19432 43948
rect 19484 43936 19490 43988
rect 20438 43976 20444 43988
rect 20399 43948 20444 43976
rect 20438 43936 20444 43948
rect 20496 43936 20502 43988
rect 20625 43979 20683 43985
rect 20625 43945 20637 43979
rect 20671 43976 20683 43979
rect 21085 43979 21143 43985
rect 21085 43976 21097 43979
rect 20671 43948 21097 43976
rect 20671 43945 20683 43948
rect 20625 43939 20683 43945
rect 21085 43945 21097 43948
rect 21131 43945 21143 43979
rect 21085 43939 21143 43945
rect 22649 43979 22707 43985
rect 22649 43945 22661 43979
rect 22695 43976 22707 43979
rect 23566 43976 23572 43988
rect 22695 43948 23572 43976
rect 22695 43945 22707 43948
rect 22649 43939 22707 43945
rect 23566 43936 23572 43948
rect 23624 43936 23630 43988
rect 23658 43936 23664 43988
rect 23716 43976 23722 43988
rect 28258 43976 28264 43988
rect 23716 43948 28120 43976
rect 28219 43948 28264 43976
rect 23716 43936 23722 43948
rect 22830 43908 22836 43920
rect 12406 43880 22836 43908
rect 10870 43840 10876 43852
rect 10831 43812 10876 43840
rect 10870 43800 10876 43812
rect 10928 43800 10934 43852
rect 11238 43800 11244 43852
rect 11296 43840 11302 43852
rect 11793 43843 11851 43849
rect 11793 43840 11805 43843
rect 11296 43812 11805 43840
rect 11296 43800 11302 43812
rect 11793 43809 11805 43812
rect 11839 43809 11851 43843
rect 11793 43803 11851 43809
rect 12161 43843 12219 43849
rect 12161 43809 12173 43843
rect 12207 43840 12219 43843
rect 12406 43840 12434 43880
rect 22830 43868 22836 43880
rect 22888 43908 22894 43920
rect 25130 43908 25136 43920
rect 22888 43880 23336 43908
rect 22888 43868 22894 43880
rect 12207 43812 12434 43840
rect 12207 43809 12219 43812
rect 12161 43803 12219 43809
rect 14458 43800 14464 43852
rect 14516 43840 14522 43852
rect 15010 43840 15016 43852
rect 14516 43812 15016 43840
rect 14516 43800 14522 43812
rect 15010 43800 15016 43812
rect 15068 43800 15074 43852
rect 15194 43800 15200 43852
rect 15252 43840 15258 43852
rect 15289 43843 15347 43849
rect 15289 43840 15301 43843
rect 15252 43812 15301 43840
rect 15252 43800 15258 43812
rect 15289 43809 15301 43812
rect 15335 43840 15347 43843
rect 15335 43812 16160 43840
rect 15335 43809 15347 43812
rect 15289 43803 15347 43809
rect 382 43732 388 43784
rect 440 43772 446 43784
rect 1581 43775 1639 43781
rect 1581 43772 1593 43775
rect 440 43744 1593 43772
rect 440 43732 446 43744
rect 1581 43741 1593 43744
rect 1627 43741 1639 43775
rect 1581 43735 1639 43741
rect 11057 43775 11115 43781
rect 11057 43741 11069 43775
rect 11103 43772 11115 43775
rect 11330 43772 11336 43784
rect 11103 43744 11336 43772
rect 11103 43741 11115 43744
rect 11057 43735 11115 43741
rect 11330 43732 11336 43744
rect 11388 43772 11394 43784
rect 11977 43775 12035 43781
rect 11977 43772 11989 43775
rect 11388 43744 11989 43772
rect 11388 43732 11394 43744
rect 11977 43741 11989 43744
rect 12023 43741 12035 43775
rect 11977 43735 12035 43741
rect 13262 43732 13268 43784
rect 13320 43772 13326 43784
rect 13449 43775 13507 43781
rect 13449 43772 13461 43775
rect 13320 43744 13461 43772
rect 13320 43732 13326 43744
rect 13449 43741 13461 43744
rect 13495 43741 13507 43775
rect 13449 43735 13507 43741
rect 13538 43732 13544 43784
rect 13596 43772 13602 43784
rect 15105 43775 15163 43781
rect 15105 43772 15117 43775
rect 13596 43744 15117 43772
rect 13596 43732 13602 43744
rect 15105 43741 15117 43744
rect 15151 43772 15163 43775
rect 15746 43772 15752 43784
rect 15151 43744 15752 43772
rect 15151 43741 15163 43744
rect 15105 43735 15163 43741
rect 15746 43732 15752 43744
rect 15804 43732 15810 43784
rect 14182 43664 14188 43716
rect 14240 43704 14246 43716
rect 14918 43704 14924 43716
rect 14240 43676 14924 43704
rect 14240 43664 14246 43676
rect 14918 43664 14924 43676
rect 14976 43664 14982 43716
rect 15013 43707 15071 43713
rect 15013 43673 15025 43707
rect 15059 43704 15071 43707
rect 15470 43704 15476 43716
rect 15059 43676 15476 43704
rect 15059 43673 15071 43676
rect 15013 43667 15071 43673
rect 15470 43664 15476 43676
rect 15528 43664 15534 43716
rect 16132 43704 16160 43812
rect 16206 43800 16212 43852
rect 16264 43840 16270 43852
rect 16301 43843 16359 43849
rect 16301 43840 16313 43843
rect 16264 43812 16313 43840
rect 16264 43800 16270 43812
rect 16301 43809 16313 43812
rect 16347 43809 16359 43843
rect 16301 43803 16359 43809
rect 16393 43843 16451 43849
rect 16393 43809 16405 43843
rect 16439 43840 16451 43843
rect 16574 43840 16580 43852
rect 16439 43812 16580 43840
rect 16439 43809 16451 43812
rect 16393 43803 16451 43809
rect 16316 43772 16344 43803
rect 16574 43800 16580 43812
rect 16632 43800 16638 43852
rect 17402 43840 17408 43852
rect 17363 43812 17408 43840
rect 17402 43800 17408 43812
rect 17460 43800 17466 43852
rect 19334 43840 19340 43852
rect 19295 43812 19340 43840
rect 19334 43800 19340 43812
rect 19392 43800 19398 43852
rect 22646 43840 22652 43852
rect 20180 43812 22652 43840
rect 16482 43772 16488 43784
rect 16316 43744 16488 43772
rect 16482 43732 16488 43744
rect 16540 43732 16546 43784
rect 16592 43704 16620 43800
rect 16942 43732 16948 43784
rect 17000 43772 17006 43784
rect 17129 43775 17187 43781
rect 17129 43772 17141 43775
rect 17000 43744 17141 43772
rect 17000 43732 17006 43744
rect 17129 43741 17141 43744
rect 17175 43772 17187 43775
rect 17586 43772 17592 43784
rect 17175 43744 17592 43772
rect 17175 43741 17187 43744
rect 17129 43735 17187 43741
rect 17586 43732 17592 43744
rect 17644 43732 17650 43784
rect 18417 43775 18475 43781
rect 18417 43741 18429 43775
rect 18463 43741 18475 43775
rect 18417 43735 18475 43741
rect 19245 43775 19303 43781
rect 19245 43741 19257 43775
rect 19291 43772 19303 43775
rect 20070 43772 20076 43784
rect 19291 43744 20076 43772
rect 19291 43741 19303 43744
rect 19245 43735 19303 43741
rect 16132 43676 16620 43704
rect 18432 43704 18460 43735
rect 20070 43732 20076 43744
rect 20128 43772 20134 43784
rect 20180 43772 20208 43812
rect 22646 43800 22652 43812
rect 22704 43800 22710 43852
rect 20346 43772 20352 43784
rect 20128 43744 20208 43772
rect 20307 43744 20352 43772
rect 20128 43732 20134 43744
rect 20346 43732 20352 43744
rect 20404 43732 20410 43784
rect 20441 43775 20499 43781
rect 20441 43741 20453 43775
rect 20487 43772 20499 43775
rect 20806 43772 20812 43784
rect 20487 43744 20812 43772
rect 20487 43741 20499 43744
rect 20441 43735 20499 43741
rect 20806 43732 20812 43744
rect 20864 43732 20870 43784
rect 21082 43772 21088 43784
rect 21043 43744 21088 43772
rect 21082 43732 21088 43744
rect 21140 43732 21146 43784
rect 21266 43772 21272 43784
rect 21227 43744 21272 43772
rect 21266 43732 21272 43744
rect 21324 43732 21330 43784
rect 22462 43772 22468 43784
rect 22423 43744 22468 43772
rect 22462 43732 22468 43744
rect 22520 43732 22526 43784
rect 22554 43732 22560 43784
rect 22612 43772 22618 43784
rect 23109 43775 23167 43781
rect 23109 43772 23121 43775
rect 22612 43744 23121 43772
rect 22612 43732 22618 43744
rect 23109 43741 23121 43744
rect 23155 43772 23167 43775
rect 23198 43772 23204 43784
rect 23155 43744 23204 43772
rect 23155 43741 23167 43744
rect 23109 43735 23167 43741
rect 23198 43732 23204 43744
rect 23256 43732 23262 43784
rect 23308 43781 23336 43880
rect 23492 43880 24808 43908
rect 25091 43880 25136 43908
rect 23492 43849 23520 43880
rect 23477 43843 23535 43849
rect 23477 43809 23489 43843
rect 23523 43809 23535 43843
rect 24486 43840 24492 43852
rect 23477 43803 23535 43809
rect 23676 43812 24492 43840
rect 23293 43775 23351 43781
rect 23293 43741 23305 43775
rect 23339 43741 23351 43775
rect 23293 43735 23351 43741
rect 23385 43775 23443 43781
rect 23385 43741 23397 43775
rect 23431 43772 23443 43775
rect 23566 43772 23572 43784
rect 23431 43744 23572 43772
rect 23431 43741 23443 43744
rect 23385 43735 23443 43741
rect 23566 43732 23572 43744
rect 23624 43732 23630 43784
rect 23676 43781 23704 43812
rect 24486 43800 24492 43812
rect 24544 43800 24550 43852
rect 24780 43849 24808 43880
rect 25130 43868 25136 43880
rect 25188 43868 25194 43920
rect 24765 43843 24823 43849
rect 24765 43809 24777 43843
rect 24811 43840 24823 43843
rect 25406 43840 25412 43852
rect 24811 43812 25412 43840
rect 24811 43809 24823 43812
rect 24765 43803 24823 43809
rect 25406 43800 25412 43812
rect 25464 43840 25470 43852
rect 25866 43840 25872 43852
rect 25464 43812 25872 43840
rect 25464 43800 25470 43812
rect 25866 43800 25872 43812
rect 25924 43800 25930 43852
rect 28092 43840 28120 43948
rect 28258 43936 28264 43948
rect 28316 43936 28322 43988
rect 30834 43936 30840 43988
rect 30892 43976 30898 43988
rect 30929 43979 30987 43985
rect 30929 43976 30941 43979
rect 30892 43948 30941 43976
rect 30892 43936 30898 43948
rect 30929 43945 30941 43948
rect 30975 43945 30987 43979
rect 30929 43939 30987 43945
rect 30006 43908 30012 43920
rect 29967 43880 30012 43908
rect 30006 43868 30012 43880
rect 30064 43868 30070 43920
rect 29086 43840 29092 43852
rect 28092 43812 29092 43840
rect 29086 43800 29092 43812
rect 29144 43800 29150 43852
rect 23661 43775 23719 43781
rect 23661 43741 23673 43775
rect 23707 43741 23719 43775
rect 24394 43772 24400 43784
rect 24355 43744 24400 43772
rect 23661 43735 23719 43741
rect 24394 43732 24400 43744
rect 24452 43732 24458 43784
rect 24578 43779 24584 43784
rect 24569 43773 24584 43779
rect 24569 43739 24581 43773
rect 24569 43733 24584 43739
rect 24578 43732 24584 43733
rect 24636 43732 24642 43784
rect 24670 43732 24676 43784
rect 24728 43772 24734 43784
rect 24946 43772 24952 43784
rect 24728 43744 24773 43772
rect 24907 43744 24952 43772
rect 24728 43732 24734 43744
rect 24946 43732 24952 43744
rect 25004 43732 25010 43784
rect 25961 43775 26019 43781
rect 25961 43741 25973 43775
rect 26007 43772 26019 43775
rect 26050 43772 26056 43784
rect 26007 43744 26056 43772
rect 26007 43741 26019 43744
rect 25961 43735 26019 43741
rect 26050 43732 26056 43744
rect 26108 43732 26114 43784
rect 27062 43772 27068 43784
rect 26160 43744 27068 43772
rect 20165 43707 20223 43713
rect 18432 43676 19656 43704
rect 11238 43636 11244 43648
rect 11199 43608 11244 43636
rect 11238 43596 11244 43608
rect 11296 43596 11302 43648
rect 13265 43639 13323 43645
rect 13265 43605 13277 43639
rect 13311 43636 13323 43639
rect 14458 43636 14464 43648
rect 13311 43608 14464 43636
rect 13311 43605 13323 43608
rect 13265 43599 13323 43605
rect 14458 43596 14464 43608
rect 14516 43596 14522 43648
rect 14550 43596 14556 43648
rect 14608 43636 14614 43648
rect 14645 43639 14703 43645
rect 14645 43636 14657 43639
rect 14608 43608 14657 43636
rect 14608 43596 14614 43608
rect 14645 43605 14657 43608
rect 14691 43605 14703 43639
rect 14645 43599 14703 43605
rect 15378 43596 15384 43648
rect 15436 43636 15442 43648
rect 15841 43639 15899 43645
rect 15841 43636 15853 43639
rect 15436 43608 15853 43636
rect 15436 43596 15442 43608
rect 15841 43605 15853 43608
rect 15887 43605 15899 43639
rect 16206 43636 16212 43648
rect 16167 43608 16212 43636
rect 15841 43599 15899 43605
rect 16206 43596 16212 43608
rect 16264 43596 16270 43648
rect 16390 43596 16396 43648
rect 16448 43636 16454 43648
rect 17586 43636 17592 43648
rect 16448 43608 17592 43636
rect 16448 43596 16454 43608
rect 17586 43596 17592 43608
rect 17644 43596 17650 43648
rect 18601 43639 18659 43645
rect 18601 43605 18613 43639
rect 18647 43636 18659 43639
rect 18782 43636 18788 43648
rect 18647 43608 18788 43636
rect 18647 43605 18659 43608
rect 18601 43599 18659 43605
rect 18782 43596 18788 43608
rect 18840 43596 18846 43648
rect 19628 43645 19656 43676
rect 20165 43673 20177 43707
rect 20211 43704 20223 43707
rect 20254 43704 20260 43716
rect 20211 43676 20260 43704
rect 20211 43673 20223 43676
rect 20165 43667 20223 43673
rect 20254 43664 20260 43676
rect 20312 43664 20318 43716
rect 20622 43664 20628 43716
rect 20680 43704 20686 43716
rect 24118 43704 24124 43716
rect 20680 43676 24124 43704
rect 20680 43664 20686 43676
rect 24118 43664 24124 43676
rect 24176 43664 24182 43716
rect 24302 43664 24308 43716
rect 24360 43704 24366 43716
rect 26160 43704 26188 43744
rect 27062 43732 27068 43744
rect 27120 43732 27126 43784
rect 27893 43775 27951 43781
rect 27893 43741 27905 43775
rect 27939 43772 27951 43775
rect 28074 43772 28080 43784
rect 27939 43744 28080 43772
rect 27939 43741 27951 43744
rect 27893 43735 27951 43741
rect 28074 43732 28080 43744
rect 28132 43732 28138 43784
rect 28994 43732 29000 43784
rect 29052 43772 29058 43784
rect 29825 43775 29883 43781
rect 29825 43772 29837 43775
rect 29052 43744 29837 43772
rect 29052 43732 29058 43744
rect 29825 43741 29837 43744
rect 29871 43741 29883 43775
rect 29825 43735 29883 43741
rect 26234 43713 26240 43716
rect 24360 43676 26188 43704
rect 24360 43664 24366 43676
rect 26228 43667 26240 43713
rect 26292 43704 26298 43716
rect 26292 43676 26328 43704
rect 26436 43676 28488 43704
rect 26234 43664 26240 43667
rect 26292 43664 26298 43676
rect 19613 43639 19671 43645
rect 19613 43605 19625 43639
rect 19659 43605 19671 43639
rect 19613 43599 19671 43605
rect 19978 43596 19984 43648
rect 20036 43636 20042 43648
rect 21453 43639 21511 43645
rect 21453 43636 21465 43639
rect 20036 43608 21465 43636
rect 20036 43596 20042 43608
rect 21453 43605 21465 43608
rect 21499 43605 21511 43639
rect 21453 43599 21511 43605
rect 22370 43596 22376 43648
rect 22428 43636 22434 43648
rect 23382 43636 23388 43648
rect 22428 43608 23388 43636
rect 22428 43596 22434 43608
rect 23382 43596 23388 43608
rect 23440 43596 23446 43648
rect 23842 43636 23848 43648
rect 23803 43608 23848 43636
rect 23842 43596 23848 43608
rect 23900 43596 23906 43648
rect 23934 43596 23940 43648
rect 23992 43636 23998 43648
rect 26436 43636 26464 43676
rect 23992 43608 26464 43636
rect 23992 43596 23998 43608
rect 26602 43596 26608 43648
rect 26660 43636 26666 43648
rect 28460 43645 28488 43676
rect 27341 43639 27399 43645
rect 27341 43636 27353 43639
rect 26660 43608 27353 43636
rect 26660 43596 26666 43608
rect 27341 43605 27353 43608
rect 27387 43636 27399 43639
rect 28261 43639 28319 43645
rect 28261 43636 28273 43639
rect 27387 43608 28273 43636
rect 27387 43605 27399 43608
rect 27341 43599 27399 43605
rect 28261 43605 28273 43608
rect 28307 43605 28319 43639
rect 28261 43599 28319 43605
rect 28445 43639 28503 43645
rect 28445 43605 28457 43639
rect 28491 43605 28503 43639
rect 28445 43599 28503 43605
rect 1104 43546 30820 43568
rect 1104 43494 10880 43546
rect 10932 43494 10944 43546
rect 10996 43494 11008 43546
rect 11060 43494 11072 43546
rect 11124 43494 11136 43546
rect 11188 43494 20811 43546
rect 20863 43494 20875 43546
rect 20927 43494 20939 43546
rect 20991 43494 21003 43546
rect 21055 43494 21067 43546
rect 21119 43494 30820 43546
rect 1104 43472 30820 43494
rect 13357 43435 13415 43441
rect 13357 43401 13369 43435
rect 13403 43432 13415 43435
rect 13538 43432 13544 43444
rect 13403 43404 13544 43432
rect 13403 43401 13415 43404
rect 13357 43395 13415 43401
rect 13538 43392 13544 43404
rect 13596 43392 13602 43444
rect 14182 43432 14188 43444
rect 14143 43404 14188 43432
rect 14182 43392 14188 43404
rect 14240 43392 14246 43444
rect 15102 43392 15108 43444
rect 15160 43432 15166 43444
rect 15197 43435 15255 43441
rect 15197 43432 15209 43435
rect 15160 43404 15209 43432
rect 15160 43392 15166 43404
rect 15197 43401 15209 43404
rect 15243 43401 15255 43435
rect 15197 43395 15255 43401
rect 15286 43392 15292 43444
rect 15344 43432 15350 43444
rect 16758 43432 16764 43444
rect 15344 43404 15389 43432
rect 16719 43404 16764 43432
rect 15344 43392 15350 43404
rect 16758 43392 16764 43404
rect 16816 43392 16822 43444
rect 17586 43392 17592 43444
rect 17644 43432 17650 43444
rect 21174 43432 21180 43444
rect 17644 43404 19748 43432
rect 17644 43392 17650 43404
rect 14826 43364 14832 43376
rect 13556 43336 14832 43364
rect 1578 43296 1584 43308
rect 1539 43268 1584 43296
rect 1578 43256 1584 43268
rect 1636 43256 1642 43308
rect 13556 43305 13584 43336
rect 14826 43324 14832 43336
rect 14884 43324 14890 43376
rect 17218 43324 17224 43376
rect 17276 43364 17282 43376
rect 19518 43364 19524 43376
rect 17276 43336 19524 43364
rect 17276 43324 17282 43336
rect 19518 43324 19524 43336
rect 19576 43324 19582 43376
rect 13541 43299 13599 43305
rect 13541 43265 13553 43299
rect 13587 43265 13599 43299
rect 13541 43259 13599 43265
rect 14090 43256 14096 43308
rect 14148 43296 14154 43308
rect 14369 43299 14427 43305
rect 14369 43296 14381 43299
rect 14148 43268 14381 43296
rect 14148 43256 14154 43268
rect 14369 43265 14381 43268
rect 14415 43265 14427 43299
rect 14369 43259 14427 43265
rect 16945 43299 17003 43305
rect 16945 43265 16957 43299
rect 16991 43296 17003 43299
rect 17126 43296 17132 43308
rect 16991 43268 17132 43296
rect 16991 43265 17003 43268
rect 16945 43259 17003 43265
rect 17126 43256 17132 43268
rect 17184 43256 17190 43308
rect 17681 43299 17739 43305
rect 17681 43296 17693 43299
rect 17236 43268 17693 43296
rect 15194 43188 15200 43240
rect 15252 43228 15258 43240
rect 15381 43231 15439 43237
rect 15381 43228 15393 43231
rect 15252 43200 15393 43228
rect 15252 43188 15258 43200
rect 15381 43197 15393 43200
rect 15427 43197 15439 43231
rect 15381 43191 15439 43197
rect 17034 43188 17040 43240
rect 17092 43228 17098 43240
rect 17236 43228 17264 43268
rect 17681 43265 17693 43268
rect 17727 43265 17739 43299
rect 17681 43259 17739 43265
rect 17954 43256 17960 43308
rect 18012 43296 18018 43308
rect 18138 43296 18144 43308
rect 18012 43268 18144 43296
rect 18012 43256 18018 43268
rect 18138 43256 18144 43268
rect 18196 43296 18202 43308
rect 18877 43299 18935 43305
rect 18877 43296 18889 43299
rect 18196 43268 18889 43296
rect 18196 43256 18202 43268
rect 18877 43265 18889 43268
rect 18923 43265 18935 43299
rect 19610 43296 19616 43308
rect 19571 43268 19616 43296
rect 18877 43259 18935 43265
rect 19610 43256 19616 43268
rect 19668 43256 19674 43308
rect 17402 43228 17408 43240
rect 17092 43200 17264 43228
rect 17363 43200 17408 43228
rect 17092 43188 17098 43200
rect 17402 43188 17408 43200
rect 17460 43188 17466 43240
rect 18598 43188 18604 43240
rect 18656 43228 18662 43240
rect 19153 43231 19211 43237
rect 19153 43228 19165 43231
rect 18656 43200 19165 43228
rect 18656 43188 18662 43200
rect 19153 43197 19165 43200
rect 19199 43197 19211 43231
rect 19720 43228 19748 43404
rect 20272 43404 21180 43432
rect 20272 43305 20300 43404
rect 21174 43392 21180 43404
rect 21232 43392 21238 43444
rect 22462 43392 22468 43444
rect 22520 43432 22526 43444
rect 22925 43435 22983 43441
rect 22925 43432 22937 43435
rect 22520 43404 22937 43432
rect 22520 43392 22526 43404
rect 22925 43401 22937 43404
rect 22971 43401 22983 43435
rect 22925 43395 22983 43401
rect 23198 43392 23204 43444
rect 23256 43432 23262 43444
rect 24394 43432 24400 43444
rect 23256 43404 24400 43432
rect 23256 43392 23262 43404
rect 24394 43392 24400 43404
rect 24452 43392 24458 43444
rect 24486 43392 24492 43444
rect 24544 43432 24550 43444
rect 24765 43435 24823 43441
rect 24765 43432 24777 43435
rect 24544 43404 24777 43432
rect 24544 43392 24550 43404
rect 24765 43401 24777 43404
rect 24811 43432 24823 43435
rect 25314 43432 25320 43444
rect 24811 43404 25320 43432
rect 24811 43401 24823 43404
rect 24765 43395 24823 43401
rect 25314 43392 25320 43404
rect 25372 43392 25378 43444
rect 26237 43435 26295 43441
rect 26237 43401 26249 43435
rect 26283 43432 26295 43435
rect 26326 43432 26332 43444
rect 26283 43404 26332 43432
rect 26283 43401 26295 43404
rect 26237 43395 26295 43401
rect 26326 43392 26332 43404
rect 26384 43392 26390 43444
rect 26510 43392 26516 43444
rect 26568 43432 26574 43444
rect 26568 43404 28396 43432
rect 26568 43392 26574 43404
rect 23652 43367 23710 43373
rect 20364 43336 23612 43364
rect 20257 43299 20315 43305
rect 20257 43265 20269 43299
rect 20303 43265 20315 43299
rect 20257 43259 20315 43265
rect 20364 43228 20392 43336
rect 20441 43299 20499 43305
rect 20441 43265 20453 43299
rect 20487 43296 20499 43299
rect 21174 43296 21180 43308
rect 20487 43268 21180 43296
rect 20487 43265 20499 43268
rect 20441 43259 20499 43265
rect 21174 43256 21180 43268
rect 21232 43256 21238 43308
rect 21269 43299 21327 43305
rect 21269 43265 21281 43299
rect 21315 43296 21327 43299
rect 21928 43296 22048 43300
rect 22186 43296 22192 43308
rect 21315 43272 22192 43296
rect 21315 43268 21956 43272
rect 22020 43268 22192 43272
rect 21315 43265 21327 43268
rect 21269 43259 21327 43265
rect 22186 43256 22192 43268
rect 22244 43256 22250 43308
rect 22281 43299 22339 43305
rect 22281 43265 22293 43299
rect 22327 43265 22339 43299
rect 22738 43296 22744 43308
rect 22699 43268 22744 43296
rect 22281 43259 22339 43265
rect 21910 43228 21916 43240
rect 19720 43200 20392 43228
rect 20456 43200 21916 43228
rect 19153 43191 19211 43197
rect 11238 43120 11244 43172
rect 11296 43160 11302 43172
rect 20456 43160 20484 43200
rect 21910 43188 21916 43200
rect 21968 43188 21974 43240
rect 22296 43228 22324 43259
rect 22738 43256 22744 43268
rect 22796 43256 22802 43308
rect 23106 43256 23112 43308
rect 23164 43296 23170 43308
rect 23385 43299 23443 43305
rect 23385 43296 23397 43299
rect 23164 43268 23397 43296
rect 23164 43256 23170 43268
rect 23385 43265 23397 43268
rect 23431 43265 23443 43299
rect 23385 43259 23443 43265
rect 23474 43256 23480 43308
rect 23532 43256 23538 43308
rect 23584 43296 23612 43336
rect 23652 43333 23664 43367
rect 23698 43364 23710 43367
rect 23842 43364 23848 43376
rect 23698 43336 23848 43364
rect 23698 43333 23710 43336
rect 23652 43327 23710 43333
rect 23842 43324 23848 43336
rect 23900 43324 23906 43376
rect 24412 43364 24440 43392
rect 24412 43336 24808 43364
rect 24780 43296 24808 43336
rect 24946 43324 24952 43376
rect 25004 43364 25010 43376
rect 28261 43367 28319 43373
rect 28261 43364 28273 43367
rect 25004 43336 28273 43364
rect 25004 43324 25010 43336
rect 28261 43333 28273 43336
rect 28307 43333 28319 43367
rect 28368 43364 28396 43404
rect 28902 43392 28908 43444
rect 28960 43432 28966 43444
rect 29273 43435 29331 43441
rect 29273 43432 29285 43435
rect 28960 43404 29285 43432
rect 28960 43392 28966 43404
rect 29273 43401 29285 43404
rect 29319 43401 29331 43435
rect 29273 43395 29331 43401
rect 28368 43336 29868 43364
rect 28261 43327 28319 43333
rect 25314 43296 25320 43308
rect 23584 43268 24440 43296
rect 24780 43268 25320 43296
rect 23492 43228 23520 43256
rect 22296 43200 23520 43228
rect 20714 43160 20720 43172
rect 11296 43132 20484 43160
rect 20548 43132 20720 43160
rect 11296 43120 11302 43132
rect 1397 43095 1455 43101
rect 1397 43061 1409 43095
rect 1443 43092 1455 43095
rect 10870 43092 10876 43104
rect 1443 43064 10876 43092
rect 1443 43061 1455 43064
rect 1397 43055 1455 43061
rect 10870 43052 10876 43064
rect 10928 43052 10934 43104
rect 14829 43095 14887 43101
rect 14829 43061 14841 43095
rect 14875 43092 14887 43095
rect 14918 43092 14924 43104
rect 14875 43064 14924 43092
rect 14875 43061 14887 43064
rect 14829 43055 14887 43061
rect 14918 43052 14924 43064
rect 14976 43052 14982 43104
rect 15010 43052 15016 43104
rect 15068 43092 15074 43104
rect 18506 43092 18512 43104
rect 15068 43064 18512 43092
rect 15068 43052 15074 43064
rect 18506 43052 18512 43064
rect 18564 43052 18570 43104
rect 18690 43092 18696 43104
rect 18651 43064 18696 43092
rect 18690 43052 18696 43064
rect 18748 43052 18754 43104
rect 19058 43092 19064 43104
rect 19019 43064 19064 43092
rect 19058 43052 19064 43064
rect 19116 43052 19122 43104
rect 19702 43092 19708 43104
rect 19663 43064 19708 43092
rect 19702 43052 19708 43064
rect 19760 43052 19766 43104
rect 20441 43095 20499 43101
rect 20441 43061 20453 43095
rect 20487 43092 20499 43095
rect 20548 43092 20576 43132
rect 20714 43120 20720 43132
rect 20772 43120 20778 43172
rect 21085 43163 21143 43169
rect 21085 43129 21097 43163
rect 21131 43160 21143 43163
rect 23382 43160 23388 43172
rect 21131 43132 23388 43160
rect 21131 43129 21143 43132
rect 21085 43123 21143 43129
rect 23382 43120 23388 43132
rect 23440 43120 23446 43172
rect 24412 43160 24440 43268
rect 25314 43256 25320 43268
rect 25372 43256 25378 43308
rect 25501 43299 25559 43305
rect 25501 43265 25513 43299
rect 25547 43265 25559 43299
rect 25682 43296 25688 43308
rect 25643 43268 25688 43296
rect 25501 43259 25559 43265
rect 25332 43228 25360 43256
rect 25516 43228 25544 43259
rect 25682 43256 25688 43268
rect 25740 43256 25746 43308
rect 25866 43296 25872 43308
rect 25827 43268 25872 43296
rect 25866 43256 25872 43268
rect 25924 43256 25930 43308
rect 26053 43299 26111 43305
rect 26053 43265 26065 43299
rect 26099 43296 26111 43299
rect 26786 43296 26792 43308
rect 26099 43268 26792 43296
rect 26099 43265 26111 43268
rect 26053 43259 26111 43265
rect 26786 43256 26792 43268
rect 26844 43256 26850 43308
rect 26970 43296 26976 43308
rect 26931 43268 26976 43296
rect 26970 43256 26976 43268
rect 27028 43256 27034 43308
rect 27062 43256 27068 43308
rect 27120 43296 27126 43308
rect 29840 43305 29868 43336
rect 29089 43299 29147 43305
rect 29089 43296 29101 43299
rect 27120 43268 29101 43296
rect 27120 43256 27126 43268
rect 29089 43265 29101 43268
rect 29135 43265 29147 43299
rect 29089 43259 29147 43265
rect 29825 43299 29883 43305
rect 29825 43265 29837 43299
rect 29871 43265 29883 43299
rect 29825 43259 29883 43265
rect 25332 43200 25544 43228
rect 25590 43188 25596 43240
rect 25648 43228 25654 43240
rect 25777 43231 25835 43237
rect 25777 43228 25789 43231
rect 25648 43200 25789 43228
rect 25648 43188 25654 43200
rect 25777 43197 25789 43200
rect 25823 43197 25835 43231
rect 25777 43191 25835 43197
rect 25976 43200 28488 43228
rect 25976 43160 26004 43200
rect 24412 43132 26004 43160
rect 26326 43120 26332 43172
rect 26384 43160 26390 43172
rect 27798 43160 27804 43172
rect 26384 43132 27804 43160
rect 26384 43120 26390 43132
rect 27798 43120 27804 43132
rect 27856 43120 27862 43172
rect 27893 43163 27951 43169
rect 27893 43129 27905 43163
rect 27939 43160 27951 43163
rect 28074 43160 28080 43172
rect 27939 43132 28080 43160
rect 27939 43129 27951 43132
rect 27893 43123 27951 43129
rect 28074 43120 28080 43132
rect 28132 43120 28138 43172
rect 28460 43169 28488 43200
rect 28445 43163 28503 43169
rect 28445 43129 28457 43163
rect 28491 43129 28503 43163
rect 28445 43123 28503 43129
rect 20487 43064 20576 43092
rect 20487 43061 20499 43064
rect 20441 43055 20499 43061
rect 20622 43052 20628 43104
rect 20680 43092 20686 43104
rect 22094 43092 22100 43104
rect 20680 43064 20725 43092
rect 22055 43064 22100 43092
rect 20680 43052 20686 43064
rect 22094 43052 22100 43064
rect 22152 43052 22158 43104
rect 22278 43052 22284 43104
rect 22336 43092 22342 43104
rect 24578 43092 24584 43104
rect 22336 43064 24584 43092
rect 22336 43052 22342 43064
rect 24578 43052 24584 43064
rect 24636 43052 24642 43104
rect 25498 43052 25504 43104
rect 25556 43092 25562 43104
rect 25682 43092 25688 43104
rect 25556 43064 25688 43092
rect 25556 43052 25562 43064
rect 25682 43052 25688 43064
rect 25740 43052 25746 43104
rect 27154 43092 27160 43104
rect 27115 43064 27160 43092
rect 27154 43052 27160 43064
rect 27212 43052 27218 43104
rect 27706 43052 27712 43104
rect 27764 43092 27770 43104
rect 28258 43092 28264 43104
rect 27764 43064 28264 43092
rect 27764 43052 27770 43064
rect 28258 43052 28264 43064
rect 28316 43052 28322 43104
rect 30006 43092 30012 43104
rect 29967 43064 30012 43092
rect 30006 43052 30012 43064
rect 30064 43052 30070 43104
rect 1104 43002 30820 43024
rect 1104 42950 5915 43002
rect 5967 42950 5979 43002
rect 6031 42950 6043 43002
rect 6095 42950 6107 43002
rect 6159 42950 6171 43002
rect 6223 42950 15846 43002
rect 15898 42950 15910 43002
rect 15962 42950 15974 43002
rect 16026 42950 16038 43002
rect 16090 42950 16102 43002
rect 16154 42950 25776 43002
rect 25828 42950 25840 43002
rect 25892 42950 25904 43002
rect 25956 42950 25968 43002
rect 26020 42950 26032 43002
rect 26084 42950 30820 43002
rect 1104 42928 30820 42950
rect 16206 42848 16212 42900
rect 16264 42888 16270 42900
rect 16393 42891 16451 42897
rect 16393 42888 16405 42891
rect 16264 42860 16405 42888
rect 16264 42848 16270 42860
rect 16393 42857 16405 42860
rect 16439 42857 16451 42891
rect 16393 42851 16451 42857
rect 16761 42891 16819 42897
rect 16761 42857 16773 42891
rect 16807 42888 16819 42891
rect 17034 42888 17040 42900
rect 16807 42860 17040 42888
rect 16807 42857 16819 42860
rect 16761 42851 16819 42857
rect 17034 42848 17040 42860
rect 17092 42848 17098 42900
rect 17402 42848 17408 42900
rect 17460 42888 17466 42900
rect 19702 42888 19708 42900
rect 17460 42860 19708 42888
rect 17460 42848 17466 42860
rect 17678 42780 17684 42832
rect 17736 42820 17742 42832
rect 17736 42792 18552 42820
rect 17736 42780 17742 42792
rect 10870 42752 10876 42764
rect 10831 42724 10876 42752
rect 10870 42712 10876 42724
rect 10928 42712 10934 42764
rect 15470 42752 15476 42764
rect 15431 42724 15476 42752
rect 15470 42712 15476 42724
rect 15528 42712 15534 42764
rect 15933 42755 15991 42761
rect 15933 42721 15945 42755
rect 15979 42752 15991 42755
rect 16853 42755 16911 42761
rect 16853 42752 16865 42755
rect 15979 42724 16865 42752
rect 15979 42721 15991 42724
rect 15933 42715 15991 42721
rect 16853 42721 16865 42724
rect 16899 42752 16911 42755
rect 17310 42752 17316 42764
rect 16899 42724 17316 42752
rect 16899 42721 16911 42724
rect 16853 42715 16911 42721
rect 17310 42712 17316 42724
rect 17368 42712 17374 42764
rect 17770 42752 17776 42764
rect 17731 42724 17776 42752
rect 17770 42712 17776 42724
rect 17828 42712 17834 42764
rect 17957 42755 18015 42761
rect 17957 42721 17969 42755
rect 18003 42752 18015 42755
rect 18414 42752 18420 42764
rect 18003 42724 18420 42752
rect 18003 42721 18015 42724
rect 17957 42715 18015 42721
rect 18414 42712 18420 42724
rect 18472 42712 18478 42764
rect 11057 42687 11115 42693
rect 11057 42653 11069 42687
rect 11103 42684 11115 42687
rect 11330 42684 11336 42696
rect 11103 42656 11336 42684
rect 11103 42653 11115 42656
rect 11057 42647 11115 42653
rect 11330 42644 11336 42656
rect 11388 42644 11394 42696
rect 14458 42644 14464 42696
rect 14516 42684 14522 42696
rect 14737 42687 14795 42693
rect 14737 42684 14749 42687
rect 14516 42656 14749 42684
rect 14516 42644 14522 42656
rect 14737 42653 14749 42656
rect 14783 42653 14795 42687
rect 14737 42647 14795 42653
rect 14921 42687 14979 42693
rect 14921 42653 14933 42687
rect 14967 42653 14979 42687
rect 14921 42647 14979 42653
rect 15013 42687 15071 42693
rect 15013 42653 15025 42687
rect 15059 42684 15071 42687
rect 15102 42684 15108 42696
rect 15059 42656 15108 42684
rect 15059 42653 15071 42656
rect 15013 42647 15071 42653
rect 14936 42616 14964 42647
rect 15102 42644 15108 42656
rect 15160 42644 15166 42696
rect 15657 42687 15715 42693
rect 15657 42653 15669 42687
rect 15703 42684 15715 42687
rect 15746 42684 15752 42696
rect 15703 42656 15752 42684
rect 15703 42653 15715 42656
rect 15657 42647 15715 42653
rect 15746 42644 15752 42656
rect 15804 42644 15810 42696
rect 15841 42687 15899 42693
rect 15841 42653 15853 42687
rect 15887 42653 15899 42687
rect 15841 42647 15899 42653
rect 15194 42616 15200 42628
rect 14936 42588 15200 42616
rect 15194 42576 15200 42588
rect 15252 42576 15258 42628
rect 15856 42616 15884 42647
rect 16482 42644 16488 42696
rect 16540 42684 16546 42696
rect 16577 42687 16635 42693
rect 16577 42684 16589 42687
rect 16540 42656 16589 42684
rect 16540 42644 16546 42656
rect 16577 42653 16589 42656
rect 16623 42653 16635 42687
rect 18524 42684 18552 42792
rect 19628 42693 19656 42860
rect 19702 42848 19708 42860
rect 19760 42848 19766 42900
rect 25041 42891 25099 42897
rect 25041 42857 25053 42891
rect 25087 42857 25099 42891
rect 25041 42851 25099 42857
rect 25056 42764 25084 42851
rect 25130 42780 25136 42832
rect 25188 42820 25194 42832
rect 25406 42820 25412 42832
rect 25188 42792 25412 42820
rect 25188 42780 25194 42792
rect 25406 42780 25412 42792
rect 25464 42820 25470 42832
rect 25866 42820 25872 42832
rect 25464 42792 25872 42820
rect 25464 42780 25470 42792
rect 25866 42780 25872 42792
rect 25924 42780 25930 42832
rect 25038 42712 25044 42764
rect 25096 42712 25102 42764
rect 27154 42752 27160 42764
rect 25148 42724 27160 42752
rect 18693 42687 18751 42693
rect 18693 42684 18705 42687
rect 18524 42656 18705 42684
rect 16577 42647 16635 42653
rect 18693 42653 18705 42656
rect 18739 42653 18751 42687
rect 18693 42647 18751 42653
rect 19521 42687 19579 42693
rect 19521 42653 19533 42687
rect 19567 42653 19579 42687
rect 19521 42647 19579 42653
rect 19613 42687 19671 42693
rect 19613 42653 19625 42687
rect 19659 42653 19671 42687
rect 19613 42647 19671 42653
rect 17034 42616 17040 42628
rect 15856 42588 17040 42616
rect 17034 42576 17040 42588
rect 17092 42576 17098 42628
rect 19536 42616 19564 42647
rect 20070 42644 20076 42696
rect 20128 42684 20134 42696
rect 20533 42687 20591 42693
rect 20533 42684 20545 42687
rect 20128 42656 20545 42684
rect 20128 42644 20134 42656
rect 20533 42653 20545 42656
rect 20579 42653 20591 42687
rect 20533 42647 20591 42653
rect 20622 42644 20628 42696
rect 20680 42684 20686 42696
rect 22738 42684 22744 42696
rect 20680 42656 22094 42684
rect 22699 42656 22744 42684
rect 20680 42644 20686 42656
rect 20800 42619 20858 42625
rect 19536 42588 20024 42616
rect 11238 42548 11244 42560
rect 11199 42520 11244 42548
rect 11238 42508 11244 42520
rect 11296 42508 11302 42560
rect 14553 42551 14611 42557
rect 14553 42517 14565 42551
rect 14599 42548 14611 42551
rect 14642 42548 14648 42560
rect 14599 42520 14648 42548
rect 14599 42517 14611 42520
rect 14553 42511 14611 42517
rect 14642 42508 14648 42520
rect 14700 42508 14706 42560
rect 17218 42508 17224 42560
rect 17276 42548 17282 42560
rect 17313 42551 17371 42557
rect 17313 42548 17325 42551
rect 17276 42520 17325 42548
rect 17276 42508 17282 42520
rect 17313 42517 17325 42520
rect 17359 42517 17371 42551
rect 17678 42548 17684 42560
rect 17639 42520 17684 42548
rect 17313 42511 17371 42517
rect 17678 42508 17684 42520
rect 17736 42508 17742 42560
rect 17770 42508 17776 42560
rect 17828 42548 17834 42560
rect 18509 42551 18567 42557
rect 18509 42548 18521 42551
rect 17828 42520 18521 42548
rect 17828 42508 17834 42520
rect 18509 42517 18521 42520
rect 18555 42517 18567 42551
rect 19794 42548 19800 42560
rect 19755 42520 19800 42548
rect 18509 42511 18567 42517
rect 19794 42508 19800 42520
rect 19852 42508 19858 42560
rect 19996 42548 20024 42588
rect 20800 42585 20812 42619
rect 20846 42616 20858 42619
rect 21174 42616 21180 42628
rect 20846 42588 21180 42616
rect 20846 42585 20858 42588
rect 20800 42579 20858 42585
rect 21174 42576 21180 42588
rect 21232 42576 21238 42628
rect 22066 42616 22094 42656
rect 22738 42644 22744 42656
rect 22796 42644 22802 42696
rect 23569 42687 23627 42693
rect 23569 42653 23581 42687
rect 23615 42653 23627 42687
rect 23569 42647 23627 42653
rect 24857 42687 24915 42693
rect 24857 42653 24869 42687
rect 24903 42684 24915 42687
rect 25148 42684 25176 42724
rect 27154 42712 27160 42724
rect 27212 42712 27218 42764
rect 27430 42712 27436 42764
rect 27488 42752 27494 42764
rect 27488 42724 29868 42752
rect 27488 42712 27494 42724
rect 24903 42656 25176 42684
rect 24903 42653 24915 42656
rect 24857 42647 24915 42653
rect 23584 42616 23612 42647
rect 25314 42644 25320 42696
rect 25372 42684 25378 42696
rect 25501 42687 25559 42693
rect 25501 42684 25513 42687
rect 25372 42656 25513 42684
rect 25372 42644 25378 42656
rect 25501 42653 25513 42656
rect 25547 42653 25559 42687
rect 25501 42647 25559 42653
rect 25590 42644 25596 42696
rect 25648 42684 25654 42696
rect 25685 42687 25743 42693
rect 25685 42684 25697 42687
rect 25648 42656 25697 42684
rect 25648 42644 25654 42656
rect 25685 42653 25697 42656
rect 25731 42653 25743 42687
rect 25685 42647 25743 42653
rect 25777 42687 25835 42693
rect 25777 42653 25789 42687
rect 25823 42653 25835 42687
rect 25777 42647 25835 42653
rect 24946 42616 24952 42628
rect 22066 42588 23520 42616
rect 23584 42588 24952 42616
rect 21913 42551 21971 42557
rect 21913 42548 21925 42551
rect 19996 42520 21925 42548
rect 21913 42517 21925 42520
rect 21959 42517 21971 42551
rect 22922 42548 22928 42560
rect 22883 42520 22928 42548
rect 21913 42511 21971 42517
rect 22922 42508 22928 42520
rect 22980 42508 22986 42560
rect 23382 42548 23388 42560
rect 23343 42520 23388 42548
rect 23382 42508 23388 42520
rect 23440 42508 23446 42560
rect 23492 42548 23520 42588
rect 24946 42576 24952 42588
rect 25004 42576 25010 42628
rect 24670 42548 24676 42560
rect 23492 42520 24676 42548
rect 24670 42508 24676 42520
rect 24728 42508 24734 42560
rect 24762 42508 24768 42560
rect 24820 42548 24826 42560
rect 25682 42548 25688 42560
rect 24820 42520 25688 42548
rect 24820 42508 24826 42520
rect 25682 42508 25688 42520
rect 25740 42548 25746 42560
rect 25792 42548 25820 42647
rect 25866 42644 25872 42696
rect 25924 42684 25930 42696
rect 26053 42687 26111 42693
rect 25924 42656 25969 42684
rect 25924 42644 25930 42656
rect 26053 42653 26065 42687
rect 26099 42653 26111 42687
rect 26053 42647 26111 42653
rect 25740 42520 25820 42548
rect 26068 42548 26096 42647
rect 26234 42644 26240 42696
rect 26292 42684 26298 42696
rect 26694 42684 26700 42696
rect 26292 42656 26337 42684
rect 26655 42656 26700 42684
rect 26292 42644 26298 42656
rect 26694 42644 26700 42656
rect 26752 42644 26758 42696
rect 27338 42684 27344 42696
rect 27299 42656 27344 42684
rect 27338 42644 27344 42656
rect 27396 42644 27402 42696
rect 28169 42687 28227 42693
rect 28169 42653 28181 42687
rect 28215 42684 28227 42687
rect 28442 42684 28448 42696
rect 28215 42656 28448 42684
rect 28215 42653 28227 42656
rect 28169 42647 28227 42653
rect 28442 42644 28448 42656
rect 28500 42644 28506 42696
rect 28813 42687 28871 42693
rect 28813 42653 28825 42687
rect 28859 42684 28871 42687
rect 28902 42684 28908 42696
rect 28859 42656 28908 42684
rect 28859 42653 28871 42656
rect 28813 42647 28871 42653
rect 28902 42644 28908 42656
rect 28960 42644 28966 42696
rect 29840 42693 29868 42724
rect 29825 42687 29883 42693
rect 29825 42653 29837 42687
rect 29871 42653 29883 42687
rect 29825 42647 29883 42653
rect 26142 42576 26148 42628
rect 26200 42616 26206 42628
rect 29730 42616 29736 42628
rect 26200 42588 26924 42616
rect 26200 42576 26206 42588
rect 26602 42548 26608 42560
rect 26068 42520 26608 42548
rect 25740 42508 25746 42520
rect 26602 42508 26608 42520
rect 26660 42508 26666 42560
rect 26896 42557 26924 42588
rect 28000 42588 29736 42616
rect 26881 42551 26939 42557
rect 26881 42517 26893 42551
rect 26927 42517 26939 42551
rect 27522 42548 27528 42560
rect 27483 42520 27528 42548
rect 26881 42511 26939 42517
rect 27522 42508 27528 42520
rect 27580 42508 27586 42560
rect 28000 42557 28028 42588
rect 29730 42576 29736 42588
rect 29788 42576 29794 42628
rect 27985 42551 28043 42557
rect 27985 42517 27997 42551
rect 28031 42517 28043 42551
rect 28626 42548 28632 42560
rect 28587 42520 28632 42548
rect 27985 42511 28043 42517
rect 28626 42508 28632 42520
rect 28684 42508 28690 42560
rect 30006 42548 30012 42560
rect 29967 42520 30012 42548
rect 30006 42508 30012 42520
rect 30064 42508 30070 42560
rect 1104 42458 30820 42480
rect 1104 42406 10880 42458
rect 10932 42406 10944 42458
rect 10996 42406 11008 42458
rect 11060 42406 11072 42458
rect 11124 42406 11136 42458
rect 11188 42406 20811 42458
rect 20863 42406 20875 42458
rect 20927 42406 20939 42458
rect 20991 42406 21003 42458
rect 21055 42406 21067 42458
rect 21119 42406 30820 42458
rect 1104 42384 30820 42406
rect 17678 42304 17684 42356
rect 17736 42344 17742 42356
rect 18233 42347 18291 42353
rect 18233 42344 18245 42347
rect 17736 42316 18245 42344
rect 17736 42304 17742 42316
rect 18233 42313 18245 42316
rect 18279 42313 18291 42347
rect 18233 42307 18291 42313
rect 18506 42304 18512 42356
rect 18564 42344 18570 42356
rect 19058 42344 19064 42356
rect 18564 42316 19064 42344
rect 18564 42304 18570 42316
rect 19058 42304 19064 42316
rect 19116 42304 19122 42356
rect 19153 42347 19211 42353
rect 19153 42313 19165 42347
rect 19199 42344 19211 42347
rect 20622 42344 20628 42356
rect 19199 42316 20628 42344
rect 19199 42313 19211 42316
rect 19153 42307 19211 42313
rect 20622 42304 20628 42316
rect 20680 42304 20686 42356
rect 21174 42344 21180 42356
rect 21135 42316 21180 42344
rect 21174 42304 21180 42316
rect 21232 42304 21238 42356
rect 23842 42344 23848 42356
rect 23803 42316 23848 42344
rect 23842 42304 23848 42316
rect 23900 42304 23906 42356
rect 25961 42347 26019 42353
rect 25961 42313 25973 42347
rect 26007 42344 26019 42347
rect 26694 42344 26700 42356
rect 26007 42316 26700 42344
rect 26007 42313 26019 42316
rect 25961 42307 26019 42313
rect 26694 42304 26700 42316
rect 26752 42304 26758 42356
rect 26786 42304 26792 42356
rect 26844 42344 26850 42356
rect 29089 42347 29147 42353
rect 29089 42344 29101 42347
rect 26844 42316 29101 42344
rect 26844 42304 26850 42316
rect 29089 42313 29101 42316
rect 29135 42313 29147 42347
rect 29089 42307 29147 42313
rect 11238 42236 11244 42288
rect 11296 42276 11302 42288
rect 15933 42279 15991 42285
rect 11296 42248 12434 42276
rect 11296 42236 11302 42248
rect 12406 42072 12434 42248
rect 15933 42245 15945 42279
rect 15979 42276 15991 42279
rect 17402 42276 17408 42288
rect 15979 42248 17408 42276
rect 15979 42245 15991 42248
rect 15933 42239 15991 42245
rect 17402 42236 17408 42248
rect 17460 42236 17466 42288
rect 19426 42276 19432 42288
rect 18708 42248 19432 42276
rect 14366 42168 14372 42220
rect 14424 42208 14430 42220
rect 15010 42208 15016 42220
rect 14424 42180 15016 42208
rect 14424 42168 14430 42180
rect 15010 42168 15016 42180
rect 15068 42168 15074 42220
rect 15194 42208 15200 42220
rect 15155 42180 15200 42208
rect 15194 42168 15200 42180
rect 15252 42168 15258 42220
rect 15289 42211 15347 42217
rect 15289 42177 15301 42211
rect 15335 42208 15347 42211
rect 15335 42180 17172 42208
rect 15335 42177 15347 42180
rect 15289 42171 15347 42177
rect 15102 42100 15108 42152
rect 15160 42140 15166 42152
rect 15304 42140 15332 42171
rect 17144 42152 17172 42180
rect 17770 42168 17776 42220
rect 17828 42208 17834 42220
rect 18417 42211 18475 42217
rect 18417 42208 18429 42211
rect 17828 42180 18429 42208
rect 17828 42168 17834 42180
rect 18417 42177 18429 42180
rect 18463 42177 18475 42211
rect 18417 42171 18475 42177
rect 16942 42140 16948 42152
rect 15160 42112 15332 42140
rect 16903 42112 16948 42140
rect 15160 42100 15166 42112
rect 16942 42100 16948 42112
rect 17000 42100 17006 42152
rect 17126 42100 17132 42152
rect 17184 42140 17190 42152
rect 17221 42143 17279 42149
rect 17221 42140 17233 42143
rect 17184 42112 17233 42140
rect 17184 42100 17190 42112
rect 17221 42109 17233 42112
rect 17267 42109 17279 42143
rect 17221 42103 17279 42109
rect 18598 42100 18604 42152
rect 18656 42140 18662 42152
rect 18708 42149 18736 42248
rect 19426 42236 19432 42248
rect 19484 42236 19490 42288
rect 19613 42279 19671 42285
rect 19613 42245 19625 42279
rect 19659 42276 19671 42279
rect 19702 42276 19708 42288
rect 19659 42248 19708 42276
rect 19659 42245 19671 42248
rect 19613 42239 19671 42245
rect 19702 42236 19708 42248
rect 19760 42236 19766 42288
rect 19794 42236 19800 42288
rect 19852 42276 19858 42288
rect 19852 42248 22048 42276
rect 19852 42236 19858 42248
rect 19518 42208 19524 42220
rect 19479 42180 19524 42208
rect 19518 42168 19524 42180
rect 19576 42168 19582 42220
rect 19886 42208 19892 42220
rect 19812 42180 19892 42208
rect 18693 42143 18751 42149
rect 18693 42140 18705 42143
rect 18656 42112 18705 42140
rect 18656 42100 18662 42112
rect 18693 42109 18705 42112
rect 18739 42109 18751 42143
rect 18693 42103 18751 42109
rect 18782 42100 18788 42152
rect 18840 42140 18846 42152
rect 19334 42140 19340 42152
rect 18840 42112 19340 42140
rect 18840 42100 18846 42112
rect 19334 42100 19340 42112
rect 19392 42100 19398 42152
rect 19812 42149 19840 42180
rect 19886 42168 19892 42180
rect 19944 42168 19950 42220
rect 19978 42168 19984 42220
rect 20036 42208 20042 42220
rect 20441 42211 20499 42217
rect 20441 42208 20453 42211
rect 20036 42180 20453 42208
rect 20036 42168 20042 42180
rect 20441 42177 20453 42180
rect 20487 42177 20499 42211
rect 20622 42208 20628 42220
rect 20583 42180 20628 42208
rect 20441 42171 20499 42177
rect 20622 42168 20628 42180
rect 20680 42168 20686 42220
rect 21085 42211 21143 42217
rect 21085 42177 21097 42211
rect 21131 42177 21143 42211
rect 21266 42208 21272 42220
rect 21227 42180 21272 42208
rect 21085 42171 21143 42177
rect 19797 42143 19855 42149
rect 19797 42109 19809 42143
rect 19843 42109 19855 42143
rect 21100 42140 21128 42171
rect 21266 42168 21272 42180
rect 21324 42168 21330 42220
rect 22020 42217 22048 42248
rect 22646 42236 22652 42288
rect 22704 42276 22710 42288
rect 22704 42248 23244 42276
rect 22704 42236 22710 42248
rect 22005 42211 22063 42217
rect 22005 42177 22017 42211
rect 22051 42177 22063 42211
rect 22005 42171 22063 42177
rect 23014 42168 23020 42220
rect 23072 42208 23078 42220
rect 23216 42208 23244 42248
rect 23382 42236 23388 42288
rect 23440 42276 23446 42288
rect 23440 42248 27108 42276
rect 23440 42236 23446 42248
rect 24026 42208 24032 42220
rect 23072 42180 23117 42208
rect 23216 42180 24032 42208
rect 23072 42168 23078 42180
rect 24026 42168 24032 42180
rect 24084 42168 24090 42220
rect 24118 42168 24124 42220
rect 24176 42208 24182 42220
rect 25777 42211 25835 42217
rect 25777 42208 25789 42211
rect 24176 42180 25789 42208
rect 24176 42168 24182 42180
rect 25777 42177 25789 42180
rect 25823 42208 25835 42211
rect 26970 42208 26976 42220
rect 25823 42180 26976 42208
rect 25823 42177 25835 42180
rect 25777 42171 25835 42177
rect 26970 42168 26976 42180
rect 27028 42168 27034 42220
rect 21542 42140 21548 42152
rect 21100 42112 21548 42140
rect 19797 42103 19855 42109
rect 21542 42100 21548 42112
rect 21600 42100 21606 42152
rect 24210 42100 24216 42152
rect 24268 42140 24274 42152
rect 24489 42143 24547 42149
rect 24489 42140 24501 42143
rect 24268 42112 24501 42140
rect 24268 42100 24274 42112
rect 24489 42109 24501 42112
rect 24535 42109 24547 42143
rect 24762 42140 24768 42152
rect 24723 42112 24768 42140
rect 24489 42103 24547 42109
rect 24762 42100 24768 42112
rect 24820 42100 24826 42152
rect 27080 42140 27108 42248
rect 27430 42236 27436 42288
rect 27488 42276 27494 42288
rect 27488 42248 27568 42276
rect 27488 42236 27494 42248
rect 27540 42217 27568 42248
rect 27706 42236 27712 42288
rect 27764 42276 27770 42288
rect 27893 42279 27951 42285
rect 27893 42276 27905 42279
rect 27764 42248 27905 42276
rect 27764 42236 27770 42248
rect 27893 42245 27905 42248
rect 27939 42245 27951 42279
rect 27893 42239 27951 42245
rect 27982 42236 27988 42288
rect 28040 42276 28046 42288
rect 28905 42279 28963 42285
rect 28905 42276 28917 42279
rect 28040 42248 28917 42276
rect 28040 42236 28046 42248
rect 28905 42245 28917 42248
rect 28951 42245 28963 42279
rect 28905 42239 28963 42245
rect 27525 42211 27583 42217
rect 27525 42177 27537 42211
rect 27571 42208 27583 42211
rect 28534 42208 28540 42220
rect 27571 42180 28540 42208
rect 27571 42177 27583 42180
rect 27525 42171 27583 42177
rect 28534 42168 28540 42180
rect 28592 42168 28598 42220
rect 29825 42211 29883 42217
rect 29825 42208 29837 42211
rect 28966 42180 29837 42208
rect 28966 42140 28994 42180
rect 29825 42177 29837 42180
rect 29871 42177 29883 42211
rect 29825 42171 29883 42177
rect 27080 42112 28994 42140
rect 12406 42044 18736 42072
rect 14826 42004 14832 42016
rect 14787 41976 14832 42004
rect 14826 41964 14832 41976
rect 14884 41964 14890 42016
rect 16025 42007 16083 42013
rect 16025 41973 16037 42007
rect 16071 42004 16083 42007
rect 18506 42004 18512 42016
rect 16071 41976 18512 42004
rect 16071 41973 16083 41976
rect 16025 41967 16083 41973
rect 18506 41964 18512 41976
rect 18564 42004 18570 42016
rect 18601 42007 18659 42013
rect 18601 42004 18613 42007
rect 18564 41976 18613 42004
rect 18564 41964 18570 41976
rect 18601 41973 18613 41976
rect 18647 41973 18659 42007
rect 18708 42004 18736 42044
rect 19886 42032 19892 42084
rect 19944 42072 19950 42084
rect 21821 42075 21879 42081
rect 21821 42072 21833 42075
rect 19944 42044 21833 42072
rect 19944 42032 19950 42044
rect 21821 42041 21833 42044
rect 21867 42041 21879 42075
rect 21821 42035 21879 42041
rect 22833 42075 22891 42081
rect 22833 42041 22845 42075
rect 22879 42072 22891 42075
rect 26970 42072 26976 42084
rect 22879 42044 26976 42072
rect 22879 42041 22891 42044
rect 22833 42035 22891 42041
rect 26970 42032 26976 42044
rect 27028 42032 27034 42084
rect 28077 42075 28135 42081
rect 28077 42072 28089 42075
rect 27448 42044 28089 42072
rect 21082 42004 21088 42016
rect 18708 41976 21088 42004
rect 18601 41967 18659 41973
rect 21082 41964 21088 41976
rect 21140 41964 21146 42016
rect 25038 41964 25044 42016
rect 25096 42004 25102 42016
rect 27448 42004 27476 42044
rect 28077 42041 28089 42044
rect 28123 42041 28135 42075
rect 28077 42035 28135 42041
rect 25096 41976 27476 42004
rect 27893 42007 27951 42013
rect 25096 41964 25102 41976
rect 27893 41973 27905 42007
rect 27939 42004 27951 42007
rect 28258 42004 28264 42016
rect 27939 41976 28264 42004
rect 27939 41973 27951 41976
rect 27893 41967 27951 41973
rect 28258 41964 28264 41976
rect 28316 41964 28322 42016
rect 28626 41964 28632 42016
rect 28684 42004 28690 42016
rect 28905 42007 28963 42013
rect 28905 42004 28917 42007
rect 28684 41976 28917 42004
rect 28684 41964 28690 41976
rect 28905 41973 28917 41976
rect 28951 41973 28963 42007
rect 30006 42004 30012 42016
rect 29967 41976 30012 42004
rect 28905 41967 28963 41973
rect 30006 41964 30012 41976
rect 30064 41964 30070 42016
rect 1104 41914 30820 41936
rect 1104 41862 5915 41914
rect 5967 41862 5979 41914
rect 6031 41862 6043 41914
rect 6095 41862 6107 41914
rect 6159 41862 6171 41914
rect 6223 41862 15846 41914
rect 15898 41862 15910 41914
rect 15962 41862 15974 41914
rect 16026 41862 16038 41914
rect 16090 41862 16102 41914
rect 16154 41862 25776 41914
rect 25828 41862 25840 41914
rect 25892 41862 25904 41914
rect 25956 41862 25968 41914
rect 26020 41862 26032 41914
rect 26084 41862 30820 41914
rect 1104 41840 30820 41862
rect 19061 41803 19119 41809
rect 19061 41769 19073 41803
rect 19107 41800 19119 41803
rect 21266 41800 21272 41812
rect 19107 41772 21272 41800
rect 19107 41769 19119 41772
rect 19061 41763 19119 41769
rect 21266 41760 21272 41772
rect 21324 41760 21330 41812
rect 23845 41803 23903 41809
rect 23845 41769 23857 41803
rect 23891 41800 23903 41803
rect 27338 41800 27344 41812
rect 23891 41772 27344 41800
rect 23891 41769 23903 41772
rect 23845 41763 23903 41769
rect 27338 41760 27344 41772
rect 27396 41760 27402 41812
rect 28626 41760 28632 41812
rect 28684 41800 28690 41812
rect 28810 41800 28816 41812
rect 28684 41772 28816 41800
rect 28684 41760 28690 41772
rect 28810 41760 28816 41772
rect 28868 41760 28874 41812
rect 28997 41803 29055 41809
rect 28997 41769 29009 41803
rect 29043 41800 29055 41803
rect 29086 41800 29092 41812
rect 29043 41772 29092 41800
rect 29043 41769 29055 41772
rect 28997 41763 29055 41769
rect 29086 41760 29092 41772
rect 29144 41760 29150 41812
rect 16942 41692 16948 41744
rect 17000 41732 17006 41744
rect 19978 41732 19984 41744
rect 17000 41704 19984 41732
rect 17000 41692 17006 41704
rect 19978 41692 19984 41704
rect 20036 41692 20042 41744
rect 21082 41692 21088 41744
rect 21140 41732 21146 41744
rect 21140 41704 23980 41732
rect 21140 41692 21146 41704
rect 14458 41624 14464 41676
rect 14516 41664 14522 41676
rect 14737 41667 14795 41673
rect 14737 41664 14749 41667
rect 14516 41636 14749 41664
rect 14516 41624 14522 41636
rect 14737 41633 14749 41636
rect 14783 41633 14795 41667
rect 14737 41627 14795 41633
rect 14921 41667 14979 41673
rect 14921 41633 14933 41667
rect 14967 41664 14979 41667
rect 15286 41664 15292 41676
rect 14967 41636 15292 41664
rect 14967 41633 14979 41636
rect 14921 41627 14979 41633
rect 15286 41624 15292 41636
rect 15344 41624 15350 41676
rect 16482 41624 16488 41676
rect 16540 41664 16546 41676
rect 16577 41667 16635 41673
rect 16577 41664 16589 41667
rect 16540 41636 16589 41664
rect 16540 41624 16546 41636
rect 16577 41633 16589 41636
rect 16623 41633 16635 41667
rect 19705 41667 19763 41673
rect 19705 41664 19717 41667
rect 16577 41627 16635 41633
rect 17144 41636 19717 41664
rect 14642 41596 14648 41608
rect 14603 41568 14648 41596
rect 14642 41556 14648 41568
rect 14700 41556 14706 41608
rect 17144 41596 17172 41636
rect 16316 41568 17172 41596
rect 17221 41599 17279 41605
rect 2590 41488 2596 41540
rect 2648 41528 2654 41540
rect 16316 41528 16344 41568
rect 17221 41565 17233 41599
rect 17267 41565 17279 41599
rect 17494 41596 17500 41608
rect 17455 41568 17500 41596
rect 17221 41559 17279 41565
rect 2648 41500 16344 41528
rect 16393 41531 16451 41537
rect 2648 41488 2654 41500
rect 16393 41497 16405 41531
rect 16439 41528 16451 41531
rect 16666 41528 16672 41540
rect 16439 41500 16672 41528
rect 16439 41497 16451 41500
rect 16393 41491 16451 41497
rect 16666 41488 16672 41500
rect 16724 41488 16730 41540
rect 17236 41528 17264 41559
rect 17494 41556 17500 41568
rect 17552 41556 17558 41608
rect 18892 41605 18920 41636
rect 19705 41633 19717 41636
rect 19751 41633 19763 41667
rect 20070 41664 20076 41676
rect 20031 41636 20076 41664
rect 19705 41627 19763 41633
rect 20070 41624 20076 41636
rect 20128 41624 20134 41676
rect 23842 41664 23848 41676
rect 21100 41636 23848 41664
rect 18877 41599 18935 41605
rect 18877 41565 18889 41599
rect 18923 41596 18935 41599
rect 19058 41596 19064 41608
rect 18923 41568 19064 41596
rect 18923 41565 18935 41568
rect 18877 41559 18935 41565
rect 19058 41556 19064 41568
rect 19116 41556 19122 41608
rect 19429 41599 19487 41605
rect 19429 41565 19441 41599
rect 19475 41596 19487 41599
rect 21100 41596 21128 41636
rect 23842 41624 23848 41636
rect 23900 41624 23906 41676
rect 23952 41664 23980 41704
rect 24026 41692 24032 41744
rect 24084 41732 24090 41744
rect 25222 41732 25228 41744
rect 24084 41704 25228 41732
rect 24084 41692 24090 41704
rect 25222 41692 25228 41704
rect 25280 41692 25286 41744
rect 28445 41735 28503 41741
rect 28445 41701 28457 41735
rect 28491 41732 28503 41735
rect 28534 41732 28540 41744
rect 28491 41704 28540 41732
rect 28491 41701 28503 41704
rect 28445 41695 28503 41701
rect 28534 41692 28540 41704
rect 28592 41692 28598 41744
rect 24949 41667 25007 41673
rect 23952 41636 24900 41664
rect 19475 41568 21128 41596
rect 19475 41565 19487 41568
rect 19429 41559 19487 41565
rect 21266 41556 21272 41608
rect 21324 41596 21330 41608
rect 21913 41599 21971 41605
rect 21913 41596 21925 41599
rect 21324 41568 21925 41596
rect 21324 41556 21330 41568
rect 21913 41565 21925 41568
rect 21959 41565 21971 41599
rect 21913 41559 21971 41565
rect 23017 41599 23075 41605
rect 23017 41565 23029 41599
rect 23063 41596 23075 41599
rect 23382 41596 23388 41608
rect 23063 41568 23388 41596
rect 23063 41565 23075 41568
rect 23017 41559 23075 41565
rect 23382 41556 23388 41568
rect 23440 41596 23446 41608
rect 23661 41599 23719 41605
rect 23661 41596 23673 41599
rect 23440 41568 23673 41596
rect 23440 41556 23446 41568
rect 23661 41565 23673 41568
rect 23707 41596 23719 41599
rect 24118 41596 24124 41608
rect 23707 41568 24124 41596
rect 23707 41565 23719 41568
rect 23661 41559 23719 41565
rect 24118 41556 24124 41568
rect 24176 41556 24182 41608
rect 24302 41556 24308 41608
rect 24360 41596 24366 41608
rect 24673 41599 24731 41605
rect 24673 41596 24685 41599
rect 24360 41568 24685 41596
rect 24360 41556 24366 41568
rect 24673 41565 24685 41568
rect 24719 41565 24731 41599
rect 24872 41596 24900 41636
rect 24949 41633 24961 41667
rect 24995 41664 25007 41667
rect 25130 41664 25136 41676
rect 24995 41636 25136 41664
rect 24995 41633 25007 41636
rect 24949 41627 25007 41633
rect 25130 41624 25136 41636
rect 25188 41624 25194 41676
rect 26970 41624 26976 41676
rect 27028 41664 27034 41676
rect 27028 41636 29868 41664
rect 27028 41624 27034 41636
rect 25498 41596 25504 41608
rect 24872 41568 25504 41596
rect 24673 41559 24731 41565
rect 25498 41556 25504 41568
rect 25556 41556 25562 41608
rect 25961 41599 26019 41605
rect 25961 41565 25973 41599
rect 26007 41596 26019 41599
rect 27522 41596 27528 41608
rect 26007 41568 27528 41596
rect 26007 41565 26019 41568
rect 25961 41559 26019 41565
rect 27522 41556 27528 41568
rect 27580 41556 27586 41608
rect 27982 41596 27988 41608
rect 27943 41568 27988 41596
rect 27982 41556 27988 41568
rect 28040 41556 28046 41608
rect 29840 41605 29868 41636
rect 29825 41599 29883 41605
rect 29825 41565 29837 41599
rect 29871 41565 29883 41599
rect 29825 41559 29883 41565
rect 18506 41528 18512 41540
rect 17236 41500 18512 41528
rect 18506 41488 18512 41500
rect 18564 41488 18570 41540
rect 18693 41531 18751 41537
rect 18693 41497 18705 41531
rect 18739 41528 18751 41531
rect 19610 41528 19616 41540
rect 18739 41500 19616 41528
rect 18739 41497 18751 41500
rect 18693 41491 18751 41497
rect 19610 41488 19616 41500
rect 19668 41488 19674 41540
rect 20340 41531 20398 41537
rect 20340 41497 20352 41531
rect 20386 41528 20398 41531
rect 22189 41531 22247 41537
rect 22189 41528 22201 41531
rect 20386 41500 22201 41528
rect 20386 41497 20398 41500
rect 20340 41491 20398 41497
rect 22189 41497 22201 41500
rect 22235 41497 22247 41531
rect 25038 41528 25044 41540
rect 22189 41491 22247 41497
rect 23124 41500 25044 41528
rect 14274 41460 14280 41472
rect 14235 41432 14280 41460
rect 14274 41420 14280 41432
rect 14332 41420 14338 41472
rect 15562 41420 15568 41472
rect 15620 41460 15626 41472
rect 16025 41463 16083 41469
rect 16025 41460 16037 41463
rect 15620 41432 16037 41460
rect 15620 41420 15626 41432
rect 16025 41429 16037 41432
rect 16071 41429 16083 41463
rect 16025 41423 16083 41429
rect 16485 41463 16543 41469
rect 16485 41429 16497 41463
rect 16531 41460 16543 41463
rect 16850 41460 16856 41472
rect 16531 41432 16856 41460
rect 16531 41429 16543 41432
rect 16485 41423 16543 41429
rect 16850 41420 16856 41432
rect 16908 41420 16914 41472
rect 19242 41460 19248 41472
rect 19203 41432 19248 41460
rect 19242 41420 19248 41432
rect 19300 41420 19306 41472
rect 19628 41460 19656 41488
rect 20714 41460 20720 41472
rect 19628 41432 20720 41460
rect 20714 41420 20720 41432
rect 20772 41420 20778 41472
rect 21450 41460 21456 41472
rect 21411 41432 21456 41460
rect 21450 41420 21456 41432
rect 21508 41420 21514 41472
rect 21818 41420 21824 41472
rect 21876 41460 21882 41472
rect 23124 41460 23152 41500
rect 25038 41488 25044 41500
rect 25096 41488 25102 41540
rect 26234 41537 26240 41540
rect 26228 41491 26240 41537
rect 26292 41528 26298 41540
rect 26292 41500 26328 41528
rect 26234 41488 26240 41491
rect 26292 41488 26298 41500
rect 27154 41488 27160 41540
rect 27212 41528 27218 41540
rect 28813 41531 28871 41537
rect 28813 41528 28825 41531
rect 27212 41500 28825 41528
rect 27212 41488 27218 41500
rect 28813 41497 28825 41500
rect 28859 41497 28871 41531
rect 28813 41491 28871 41497
rect 21876 41432 23152 41460
rect 23201 41463 23259 41469
rect 21876 41420 21882 41432
rect 23201 41429 23213 41463
rect 23247 41460 23259 41463
rect 23566 41460 23572 41472
rect 23247 41432 23572 41460
rect 23247 41429 23259 41432
rect 23201 41423 23259 41429
rect 23566 41420 23572 41432
rect 23624 41420 23630 41472
rect 24578 41420 24584 41472
rect 24636 41460 24642 41472
rect 24762 41460 24768 41472
rect 24636 41432 24768 41460
rect 24636 41420 24642 41432
rect 24762 41420 24768 41432
rect 24820 41420 24826 41472
rect 26970 41420 26976 41472
rect 27028 41460 27034 41472
rect 27341 41463 27399 41469
rect 27341 41460 27353 41463
rect 27028 41432 27353 41460
rect 27028 41420 27034 41432
rect 27341 41429 27353 41432
rect 27387 41460 27399 41463
rect 27706 41460 27712 41472
rect 27387 41432 27712 41460
rect 27387 41429 27399 41432
rect 27341 41423 27399 41429
rect 27706 41420 27712 41432
rect 27764 41420 27770 41472
rect 27801 41463 27859 41469
rect 27801 41429 27813 41463
rect 27847 41460 27859 41463
rect 28718 41460 28724 41472
rect 27847 41432 28724 41460
rect 27847 41429 27859 41432
rect 27801 41423 27859 41429
rect 28718 41420 28724 41432
rect 28776 41420 28782 41472
rect 30006 41460 30012 41472
rect 29967 41432 30012 41460
rect 30006 41420 30012 41432
rect 30064 41420 30070 41472
rect 1104 41370 30820 41392
rect 1104 41318 10880 41370
rect 10932 41318 10944 41370
rect 10996 41318 11008 41370
rect 11060 41318 11072 41370
rect 11124 41318 11136 41370
rect 11188 41318 20811 41370
rect 20863 41318 20875 41370
rect 20927 41318 20939 41370
rect 20991 41318 21003 41370
rect 21055 41318 21067 41370
rect 21119 41318 30820 41370
rect 1104 41296 30820 41318
rect 13906 41216 13912 41268
rect 13964 41256 13970 41268
rect 14366 41256 14372 41268
rect 13964 41228 14372 41256
rect 13964 41216 13970 41228
rect 14366 41216 14372 41228
rect 14424 41256 14430 41268
rect 14829 41259 14887 41265
rect 14829 41256 14841 41259
rect 14424 41228 14841 41256
rect 14424 41216 14430 41228
rect 14829 41225 14841 41228
rect 14875 41225 14887 41259
rect 16666 41256 16672 41268
rect 16627 41228 16672 41256
rect 14829 41219 14887 41225
rect 14844 41188 14872 41219
rect 16666 41216 16672 41228
rect 16724 41216 16730 41268
rect 18138 41256 18144 41268
rect 18099 41228 18144 41256
rect 18138 41216 18144 41228
rect 18196 41216 18202 41268
rect 26234 41256 26240 41268
rect 26195 41228 26240 41256
rect 26234 41216 26240 41228
rect 26292 41216 26298 41268
rect 26418 41216 26424 41268
rect 26476 41256 26482 41268
rect 29365 41259 29423 41265
rect 29365 41256 29377 41259
rect 26476 41228 29377 41256
rect 26476 41216 26482 41228
rect 29365 41225 29377 41228
rect 29411 41225 29423 41259
rect 29365 41219 29423 41225
rect 18049 41191 18107 41197
rect 14844 41160 15700 41188
rect 1578 41120 1584 41132
rect 1539 41092 1584 41120
rect 1578 41080 1584 41092
rect 1636 41080 1642 41132
rect 14642 41080 14648 41132
rect 14700 41120 14706 41132
rect 14737 41123 14795 41129
rect 14737 41120 14749 41123
rect 14700 41092 14749 41120
rect 14700 41080 14706 41092
rect 14737 41089 14749 41092
rect 14783 41089 14795 41123
rect 14737 41083 14795 41089
rect 15010 41080 15016 41132
rect 15068 41120 15074 41132
rect 15672 41129 15700 41160
rect 18049 41157 18061 41191
rect 18095 41188 18107 41191
rect 18690 41188 18696 41200
rect 18095 41160 18696 41188
rect 18095 41157 18107 41160
rect 18049 41151 18107 41157
rect 18690 41148 18696 41160
rect 18748 41148 18754 41200
rect 19076 41160 19380 41188
rect 15565 41123 15623 41129
rect 15565 41120 15577 41123
rect 15068 41092 15577 41120
rect 15068 41080 15074 41092
rect 15565 41089 15577 41092
rect 15611 41089 15623 41123
rect 15565 41083 15623 41089
rect 15657 41123 15715 41129
rect 15657 41089 15669 41123
rect 15703 41089 15715 41123
rect 16850 41120 16856 41132
rect 16811 41092 16856 41120
rect 15657 41083 15715 41089
rect 16850 41080 16856 41092
rect 16908 41080 16914 41132
rect 19076 41120 19104 41160
rect 19242 41120 19248 41132
rect 18432 41092 19104 41120
rect 19203 41092 19248 41120
rect 18432 41064 18460 41092
rect 19242 41080 19248 41092
rect 19300 41080 19306 41132
rect 19352 41120 19380 41160
rect 23842 41148 23848 41200
rect 23900 41188 23906 41200
rect 26970 41188 26976 41200
rect 23900 41160 24707 41188
rect 23900 41148 23906 41160
rect 19352 41092 19472 41120
rect 14921 41055 14979 41061
rect 14921 41021 14933 41055
rect 14967 41052 14979 41055
rect 15286 41052 15292 41064
rect 14967 41024 15292 41052
rect 14967 41021 14979 41024
rect 14921 41015 14979 41021
rect 15286 41012 15292 41024
rect 15344 41012 15350 41064
rect 17126 41052 17132 41064
rect 17087 41024 17132 41052
rect 17126 41012 17132 41024
rect 17184 41012 17190 41064
rect 18325 41055 18383 41061
rect 18325 41021 18337 41055
rect 18371 41052 18383 41055
rect 18414 41052 18420 41064
rect 18371 41024 18420 41052
rect 18371 41021 18383 41024
rect 18325 41015 18383 41021
rect 18414 41012 18420 41024
rect 18472 41012 18478 41064
rect 19444 41061 19472 41092
rect 21818 41080 21824 41132
rect 21876 41120 21882 41132
rect 22281 41123 22339 41129
rect 22281 41120 22293 41123
rect 21876 41092 22293 41120
rect 21876 41080 21882 41092
rect 22281 41089 22293 41092
rect 22327 41089 22339 41123
rect 22281 41083 22339 41089
rect 23744 41123 23802 41129
rect 23744 41089 23756 41123
rect 23790 41120 23802 41123
rect 24578 41120 24584 41132
rect 23790 41092 24584 41120
rect 23790 41089 23802 41092
rect 23744 41083 23802 41089
rect 24578 41080 24584 41092
rect 24636 41080 24642 41132
rect 19337 41055 19395 41061
rect 19337 41052 19349 41055
rect 18616 41024 19349 41052
rect 14458 40944 14464 40996
rect 14516 40984 14522 40996
rect 14516 40956 15608 40984
rect 14516 40944 14522 40956
rect 1397 40919 1455 40925
rect 1397 40885 1409 40919
rect 1443 40916 1455 40919
rect 12066 40916 12072 40928
rect 1443 40888 12072 40916
rect 1443 40885 1455 40888
rect 1397 40879 1455 40885
rect 12066 40876 12072 40888
rect 12124 40876 12130 40928
rect 14182 40876 14188 40928
rect 14240 40916 14246 40928
rect 15580 40925 15608 40956
rect 18046 40944 18052 40996
rect 18104 40984 18110 40996
rect 18616 40984 18644 41024
rect 19337 41021 19349 41024
rect 19383 41021 19395 41055
rect 19337 41015 19395 41021
rect 19429 41055 19487 41061
rect 19429 41021 19441 41055
rect 19475 41021 19487 41055
rect 19429 41015 19487 41021
rect 20714 41012 20720 41064
rect 20772 41052 20778 41064
rect 20901 41055 20959 41061
rect 20901 41052 20913 41055
rect 20772 41024 20913 41052
rect 20772 41012 20778 41024
rect 20901 41021 20913 41024
rect 20947 41021 20959 41055
rect 20901 41015 20959 41021
rect 21174 41012 21180 41064
rect 21232 41052 21238 41064
rect 21634 41052 21640 41064
rect 21232 41024 21640 41052
rect 21232 41012 21238 41024
rect 21634 41012 21640 41024
rect 21692 41012 21698 41064
rect 23474 41052 23480 41064
rect 23435 41024 23480 41052
rect 23474 41012 23480 41024
rect 23532 41012 23538 41064
rect 24679 41052 24707 41160
rect 26528 41160 26976 41188
rect 25501 41123 25559 41129
rect 25501 41120 25513 41123
rect 24955 41092 25513 41120
rect 24955 41052 24983 41092
rect 25501 41089 25513 41092
rect 25547 41089 25559 41123
rect 25673 41123 25731 41129
rect 25673 41120 25685 41123
rect 25501 41083 25559 41089
rect 25608 41092 25685 41120
rect 24679 41024 24983 41052
rect 25038 41012 25044 41064
rect 25096 41052 25102 41064
rect 25608 41052 25636 41092
rect 25673 41089 25685 41092
rect 25719 41089 25731 41123
rect 25673 41083 25731 41089
rect 25774 41080 25780 41132
rect 25832 41120 25838 41132
rect 26053 41123 26111 41129
rect 25832 41092 25877 41120
rect 25832 41080 25838 41092
rect 26053 41089 26065 41123
rect 26099 41120 26111 41123
rect 26528 41120 26556 41160
rect 26970 41148 26976 41160
rect 27028 41148 27034 41200
rect 28350 41148 28356 41200
rect 28408 41188 28414 41200
rect 29181 41191 29239 41197
rect 29181 41188 29193 41191
rect 28408 41160 29193 41188
rect 28408 41148 28414 41160
rect 29181 41157 29193 41160
rect 29227 41157 29239 41191
rect 29181 41151 29239 41157
rect 26099 41092 26556 41120
rect 26099 41089 26111 41092
rect 26053 41083 26111 41089
rect 26602 41080 26608 41132
rect 26660 41120 26666 41132
rect 27229 41123 27287 41129
rect 27229 41120 27241 41123
rect 26660 41092 27241 41120
rect 26660 41080 26666 41092
rect 27229 41089 27241 41092
rect 27275 41089 27287 41123
rect 27229 41083 27287 41089
rect 28534 41080 28540 41132
rect 28592 41120 28598 41132
rect 28813 41123 28871 41129
rect 28813 41120 28825 41123
rect 28592 41092 28825 41120
rect 28592 41080 28598 41092
rect 28813 41089 28825 41092
rect 28859 41089 28871 41123
rect 28813 41083 28871 41089
rect 29730 41080 29736 41132
rect 29788 41120 29794 41132
rect 29825 41123 29883 41129
rect 29825 41120 29837 41123
rect 29788 41092 29837 41120
rect 29788 41080 29794 41092
rect 29825 41089 29837 41092
rect 29871 41089 29883 41123
rect 29825 41083 29883 41089
rect 25096 41024 25636 41052
rect 25869 41055 25927 41061
rect 25096 41012 25102 41024
rect 25869 41021 25881 41055
rect 25915 41021 25927 41055
rect 25869 41015 25927 41021
rect 18104 40956 18644 40984
rect 18104 40944 18110 40956
rect 19518 40944 19524 40996
rect 19576 40984 19582 40996
rect 20349 40987 20407 40993
rect 20349 40984 20361 40987
rect 19576 40956 20361 40984
rect 19576 40944 19582 40956
rect 20349 40953 20361 40956
rect 20395 40953 20407 40987
rect 20349 40947 20407 40953
rect 20809 40987 20867 40993
rect 20809 40953 20821 40987
rect 20855 40984 20867 40987
rect 21450 40984 21456 40996
rect 20855 40956 21456 40984
rect 20855 40953 20867 40956
rect 20809 40947 20867 40953
rect 21450 40944 21456 40956
rect 21508 40944 21514 40996
rect 22186 40944 22192 40996
rect 22244 40984 22250 40996
rect 22465 40987 22523 40993
rect 22465 40984 22477 40987
rect 22244 40956 22477 40984
rect 22244 40944 22250 40956
rect 22465 40953 22477 40956
rect 22511 40984 22523 40987
rect 23106 40984 23112 40996
rect 22511 40956 23112 40984
rect 22511 40953 22523 40956
rect 22465 40947 22523 40953
rect 23106 40944 23112 40956
rect 23164 40944 23170 40996
rect 25130 40944 25136 40996
rect 25188 40984 25194 40996
rect 25884 40984 25912 41015
rect 26418 41012 26424 41064
rect 26476 41052 26482 41064
rect 26973 41055 27031 41061
rect 26973 41052 26985 41055
rect 26476 41024 26985 41052
rect 26476 41012 26482 41024
rect 26973 41021 26985 41024
rect 27019 41021 27031 41055
rect 26973 41015 27031 41021
rect 28258 41012 28264 41064
rect 28316 41052 28322 41064
rect 29546 41052 29552 41064
rect 28316 41024 29552 41052
rect 28316 41012 28322 41024
rect 29546 41012 29552 41024
rect 29604 41012 29610 41064
rect 25188 40956 25912 40984
rect 25188 40944 25194 40956
rect 28166 40944 28172 40996
rect 28224 40984 28230 40996
rect 31573 40987 31631 40993
rect 31573 40984 31585 40987
rect 28224 40956 31585 40984
rect 28224 40944 28230 40956
rect 31573 40953 31585 40956
rect 31619 40953 31631 40987
rect 31573 40947 31631 40953
rect 14369 40919 14427 40925
rect 14369 40916 14381 40919
rect 14240 40888 14381 40916
rect 14240 40876 14246 40888
rect 14369 40885 14381 40888
rect 14415 40885 14427 40919
rect 14369 40879 14427 40885
rect 15565 40919 15623 40925
rect 15565 40885 15577 40919
rect 15611 40885 15623 40919
rect 15565 40879 15623 40885
rect 15933 40919 15991 40925
rect 15933 40885 15945 40919
rect 15979 40916 15991 40919
rect 16390 40916 16396 40928
rect 15979 40888 16396 40916
rect 15979 40885 15991 40888
rect 15933 40879 15991 40885
rect 16390 40876 16396 40888
rect 16448 40876 16454 40928
rect 17034 40916 17040 40928
rect 16995 40888 17040 40916
rect 17034 40876 17040 40888
rect 17092 40916 17098 40928
rect 17494 40916 17500 40928
rect 17092 40888 17500 40916
rect 17092 40876 17098 40888
rect 17494 40876 17500 40888
rect 17552 40876 17558 40928
rect 17681 40919 17739 40925
rect 17681 40885 17693 40919
rect 17727 40916 17739 40919
rect 17862 40916 17868 40928
rect 17727 40888 17868 40916
rect 17727 40885 17739 40888
rect 17681 40879 17739 40885
rect 17862 40876 17868 40888
rect 17920 40876 17926 40928
rect 18138 40876 18144 40928
rect 18196 40916 18202 40928
rect 18877 40919 18935 40925
rect 18877 40916 18889 40919
rect 18196 40888 18889 40916
rect 18196 40876 18202 40888
rect 18877 40885 18889 40888
rect 18923 40885 18935 40919
rect 20714 40916 20720 40928
rect 20675 40888 20720 40916
rect 18877 40879 18935 40885
rect 20714 40876 20720 40888
rect 20772 40876 20778 40928
rect 21177 40919 21235 40925
rect 21177 40885 21189 40919
rect 21223 40916 21235 40919
rect 21726 40916 21732 40928
rect 21223 40888 21732 40916
rect 21223 40885 21235 40888
rect 21177 40879 21235 40885
rect 21726 40876 21732 40888
rect 21784 40876 21790 40928
rect 24394 40876 24400 40928
rect 24452 40916 24458 40928
rect 24857 40919 24915 40925
rect 24857 40916 24869 40919
rect 24452 40888 24869 40916
rect 24452 40876 24458 40888
rect 24857 40885 24869 40888
rect 24903 40916 24915 40919
rect 27890 40916 27896 40928
rect 24903 40888 27896 40916
rect 24903 40885 24915 40888
rect 24857 40879 24915 40885
rect 27890 40876 27896 40888
rect 27948 40876 27954 40928
rect 28350 40916 28356 40928
rect 28311 40888 28356 40916
rect 28350 40876 28356 40888
rect 28408 40876 28414 40928
rect 29178 40916 29184 40928
rect 29139 40888 29184 40916
rect 29178 40876 29184 40888
rect 29236 40876 29242 40928
rect 30009 40919 30067 40925
rect 30009 40885 30021 40919
rect 30055 40916 30067 40919
rect 30098 40916 30104 40928
rect 30055 40888 30104 40916
rect 30055 40885 30067 40888
rect 30009 40879 30067 40885
rect 30098 40876 30104 40888
rect 30156 40876 30162 40928
rect 1104 40826 30820 40848
rect 1104 40774 5915 40826
rect 5967 40774 5979 40826
rect 6031 40774 6043 40826
rect 6095 40774 6107 40826
rect 6159 40774 6171 40826
rect 6223 40774 15846 40826
rect 15898 40774 15910 40826
rect 15962 40774 15974 40826
rect 16026 40774 16038 40826
rect 16090 40774 16102 40826
rect 16154 40774 25776 40826
rect 25828 40774 25840 40826
rect 25892 40774 25904 40826
rect 25956 40774 25968 40826
rect 26020 40774 26032 40826
rect 26084 40774 30820 40826
rect 1104 40752 30820 40774
rect 12618 40672 12624 40724
rect 12676 40712 12682 40724
rect 18233 40715 18291 40721
rect 12676 40684 17172 40712
rect 12676 40672 12682 40684
rect 5350 40604 5356 40656
rect 5408 40644 5414 40656
rect 5408 40616 14964 40644
rect 5408 40604 5414 40616
rect 11698 40536 11704 40588
rect 11756 40576 11762 40588
rect 14550 40576 14556 40588
rect 11756 40548 14556 40576
rect 11756 40536 11762 40548
rect 14550 40536 14556 40548
rect 14608 40536 14614 40588
rect 14936 40576 14964 40616
rect 15010 40604 15016 40656
rect 15068 40644 15074 40656
rect 16209 40647 16267 40653
rect 15068 40616 15148 40644
rect 15068 40604 15074 40616
rect 15120 40585 15148 40616
rect 16209 40613 16221 40647
rect 16255 40644 16267 40647
rect 16850 40644 16856 40656
rect 16255 40616 16856 40644
rect 16255 40613 16267 40616
rect 16209 40607 16267 40613
rect 16850 40604 16856 40616
rect 16908 40604 16914 40656
rect 17144 40644 17172 40684
rect 18233 40681 18245 40715
rect 18279 40712 18291 40715
rect 19242 40712 19248 40724
rect 18279 40684 19248 40712
rect 18279 40681 18291 40684
rect 18233 40675 18291 40681
rect 19242 40672 19248 40684
rect 19300 40672 19306 40724
rect 19702 40672 19708 40724
rect 19760 40712 19766 40724
rect 20254 40712 20260 40724
rect 19760 40684 20260 40712
rect 19760 40672 19766 40684
rect 20254 40672 20260 40684
rect 20312 40672 20318 40724
rect 20714 40672 20720 40724
rect 20772 40712 20778 40724
rect 21818 40712 21824 40724
rect 20772 40684 21824 40712
rect 20772 40672 20778 40684
rect 21818 40672 21824 40684
rect 21876 40672 21882 40724
rect 23474 40672 23480 40724
rect 23532 40712 23538 40724
rect 23753 40715 23811 40721
rect 23753 40712 23765 40715
rect 23532 40684 23765 40712
rect 23532 40672 23538 40684
rect 23753 40681 23765 40684
rect 23799 40681 23811 40715
rect 23753 40675 23811 40681
rect 24213 40715 24271 40721
rect 24213 40681 24225 40715
rect 24259 40712 24271 40715
rect 26510 40712 26516 40724
rect 24259 40684 26516 40712
rect 24259 40681 24271 40684
rect 24213 40675 24271 40681
rect 26510 40672 26516 40684
rect 26568 40672 26574 40724
rect 28810 40712 28816 40724
rect 28723 40684 28816 40712
rect 28810 40672 28816 40684
rect 28868 40712 28874 40724
rect 29178 40712 29184 40724
rect 28868 40684 29184 40712
rect 28868 40672 28874 40684
rect 29178 40672 29184 40684
rect 29236 40672 29242 40724
rect 19518 40644 19524 40656
rect 17144 40616 19524 40644
rect 19518 40604 19524 40616
rect 19576 40604 19582 40656
rect 20346 40604 20352 40656
rect 20404 40644 20410 40656
rect 20993 40647 21051 40653
rect 20993 40644 21005 40647
rect 20404 40616 21005 40644
rect 20404 40604 20410 40616
rect 20993 40613 21005 40616
rect 21039 40644 21051 40647
rect 21174 40644 21180 40656
rect 21039 40616 21180 40644
rect 21039 40613 21051 40616
rect 20993 40607 21051 40613
rect 21174 40604 21180 40616
rect 21232 40604 21238 40656
rect 23109 40647 23167 40653
rect 23109 40613 23121 40647
rect 23155 40644 23167 40647
rect 23155 40616 24440 40644
rect 23155 40613 23167 40616
rect 23109 40607 23167 40613
rect 15105 40579 15163 40585
rect 14936 40548 15056 40576
rect 14826 40468 14832 40520
rect 14884 40508 14890 40520
rect 15028 40508 15056 40548
rect 15105 40545 15117 40579
rect 15151 40545 15163 40579
rect 15105 40539 15163 40545
rect 15286 40536 15292 40588
rect 15344 40576 15350 40588
rect 16482 40576 16488 40588
rect 15344 40548 16488 40576
rect 15344 40536 15350 40548
rect 16482 40536 16488 40548
rect 16540 40576 16546 40588
rect 16761 40579 16819 40585
rect 16761 40576 16773 40579
rect 16540 40548 16773 40576
rect 16540 40536 16546 40548
rect 16761 40545 16773 40548
rect 16807 40576 16819 40579
rect 16807 40548 17172 40576
rect 16807 40545 16819 40548
rect 16761 40539 16819 40545
rect 14884 40480 14964 40508
rect 15028 40480 17080 40508
rect 14884 40468 14890 40480
rect 14936 40440 14964 40480
rect 15013 40443 15071 40449
rect 15013 40440 15025 40443
rect 14936 40412 15025 40440
rect 15013 40409 15025 40412
rect 15059 40409 15071 40443
rect 15013 40403 15071 40409
rect 14645 40375 14703 40381
rect 14645 40341 14657 40375
rect 14691 40372 14703 40375
rect 15286 40372 15292 40384
rect 14691 40344 15292 40372
rect 14691 40341 14703 40344
rect 14645 40335 14703 40341
rect 15286 40332 15292 40344
rect 15344 40332 15350 40384
rect 16574 40372 16580 40384
rect 16535 40344 16580 40372
rect 16574 40332 16580 40344
rect 16632 40332 16638 40384
rect 16669 40375 16727 40381
rect 16669 40341 16681 40375
rect 16715 40372 16727 40375
rect 16942 40372 16948 40384
rect 16715 40344 16948 40372
rect 16715 40341 16727 40344
rect 16669 40335 16727 40341
rect 16942 40332 16948 40344
rect 17000 40332 17006 40384
rect 17052 40372 17080 40480
rect 17144 40440 17172 40548
rect 17954 40536 17960 40588
rect 18012 40576 18018 40588
rect 18506 40576 18512 40588
rect 18012 40548 18512 40576
rect 18012 40536 18018 40548
rect 18506 40536 18512 40548
rect 18564 40576 18570 40588
rect 18601 40579 18659 40585
rect 18601 40576 18613 40579
rect 18564 40548 18613 40576
rect 18564 40536 18570 40548
rect 18601 40545 18613 40548
rect 18647 40545 18659 40579
rect 18601 40539 18659 40545
rect 22554 40536 22560 40588
rect 22612 40576 22618 40588
rect 24412 40585 24440 40616
rect 25406 40604 25412 40656
rect 25464 40644 25470 40656
rect 25777 40647 25835 40653
rect 25777 40644 25789 40647
rect 25464 40616 25789 40644
rect 25464 40604 25470 40616
rect 25777 40613 25789 40616
rect 25823 40644 25835 40647
rect 27154 40644 27160 40656
rect 25823 40616 27160 40644
rect 25823 40613 25835 40616
rect 25777 40607 25835 40613
rect 27154 40604 27160 40616
rect 27212 40604 27218 40656
rect 28445 40647 28503 40653
rect 28445 40613 28457 40647
rect 28491 40644 28503 40647
rect 28534 40644 28540 40656
rect 28491 40616 28540 40644
rect 28491 40613 28503 40616
rect 28445 40607 28503 40613
rect 28534 40604 28540 40616
rect 28592 40604 28598 40656
rect 28997 40647 29055 40653
rect 28997 40613 29009 40647
rect 29043 40613 29055 40647
rect 28997 40607 29055 40613
rect 24213 40579 24271 40585
rect 24213 40576 24225 40579
rect 22612 40548 24225 40576
rect 22612 40536 22618 40548
rect 24213 40545 24225 40548
rect 24259 40545 24271 40579
rect 24213 40539 24271 40545
rect 24397 40579 24455 40585
rect 24397 40545 24409 40579
rect 24443 40545 24455 40579
rect 24397 40539 24455 40545
rect 25498 40536 25504 40588
rect 25556 40576 25562 40588
rect 29012 40576 29040 40607
rect 25556 40548 29040 40576
rect 25556 40536 25562 40548
rect 18046 40468 18052 40520
rect 18104 40508 18110 40520
rect 18417 40511 18475 40517
rect 18417 40508 18429 40511
rect 18104 40480 18429 40508
rect 18104 40468 18110 40480
rect 18417 40477 18429 40480
rect 18463 40477 18475 40511
rect 18417 40471 18475 40477
rect 18693 40511 18751 40517
rect 18693 40477 18705 40511
rect 18739 40477 18751 40511
rect 18693 40471 18751 40477
rect 19521 40511 19579 40517
rect 19521 40477 19533 40511
rect 19567 40508 19579 40511
rect 19794 40508 19800 40520
rect 19567 40480 19800 40508
rect 19567 40477 19579 40480
rect 19521 40471 19579 40477
rect 18230 40440 18236 40452
rect 17144 40412 18236 40440
rect 18230 40400 18236 40412
rect 18288 40400 18294 40452
rect 18322 40400 18328 40452
rect 18380 40440 18386 40452
rect 18598 40440 18604 40452
rect 18380 40412 18604 40440
rect 18380 40400 18386 40412
rect 18598 40400 18604 40412
rect 18656 40440 18662 40452
rect 18708 40440 18736 40471
rect 19794 40468 19800 40480
rect 19852 40468 19858 40520
rect 20162 40468 20168 40520
rect 20220 40508 20226 40520
rect 20441 40511 20499 40517
rect 20441 40508 20453 40511
rect 20220 40480 20453 40508
rect 20220 40468 20226 40480
rect 20441 40477 20453 40480
rect 20487 40477 20499 40511
rect 20441 40471 20499 40477
rect 21177 40511 21235 40517
rect 21177 40477 21189 40511
rect 21223 40508 21235 40511
rect 21358 40508 21364 40520
rect 21223 40480 21364 40508
rect 21223 40477 21235 40480
rect 21177 40471 21235 40477
rect 21358 40468 21364 40480
rect 21416 40468 21422 40520
rect 21637 40511 21695 40517
rect 21637 40477 21649 40511
rect 21683 40508 21695 40511
rect 21729 40511 21787 40517
rect 21729 40508 21741 40511
rect 21683 40480 21741 40508
rect 21683 40477 21695 40480
rect 21637 40471 21695 40477
rect 21729 40477 21741 40480
rect 21775 40477 21787 40511
rect 22922 40508 22928 40520
rect 22883 40480 22928 40508
rect 21729 40471 21787 40477
rect 22922 40468 22928 40480
rect 22980 40468 22986 40520
rect 23566 40508 23572 40520
rect 23527 40480 23572 40508
rect 23566 40468 23572 40480
rect 23624 40468 23630 40520
rect 24596 40480 25452 40508
rect 18656 40412 18736 40440
rect 18800 40412 19748 40440
rect 18656 40400 18662 40412
rect 18800 40372 18828 40412
rect 19610 40372 19616 40384
rect 17052 40344 18828 40372
rect 19571 40344 19616 40372
rect 19610 40332 19616 40344
rect 19668 40332 19674 40384
rect 19720 40372 19748 40412
rect 21266 40400 21272 40452
rect 21324 40440 21330 40452
rect 23198 40440 23204 40452
rect 21324 40412 23204 40440
rect 21324 40400 21330 40412
rect 23198 40400 23204 40412
rect 23256 40400 23262 40452
rect 23290 40400 23296 40452
rect 23348 40440 23354 40452
rect 24596 40440 24624 40480
rect 23348 40412 24624 40440
rect 24664 40443 24722 40449
rect 23348 40400 23354 40412
rect 24664 40409 24676 40443
rect 24710 40440 24722 40443
rect 25130 40440 25136 40452
rect 24710 40412 25136 40440
rect 24710 40409 24722 40412
rect 24664 40403 24722 40409
rect 25130 40400 25136 40412
rect 25188 40400 25194 40452
rect 21358 40372 21364 40384
rect 19720 40344 21364 40372
rect 21358 40332 21364 40344
rect 21416 40372 21422 40384
rect 21637 40375 21695 40381
rect 21637 40372 21649 40375
rect 21416 40344 21649 40372
rect 21416 40332 21422 40344
rect 21637 40341 21649 40344
rect 21683 40341 21695 40375
rect 21637 40335 21695 40341
rect 22094 40332 22100 40384
rect 22152 40372 22158 40384
rect 24854 40372 24860 40384
rect 22152 40344 24860 40372
rect 22152 40332 22158 40344
rect 24854 40332 24860 40344
rect 24912 40332 24918 40384
rect 25424 40372 25452 40480
rect 25866 40468 25872 40520
rect 25924 40508 25930 40520
rect 26237 40511 26295 40517
rect 26237 40508 26249 40511
rect 25924 40480 26249 40508
rect 25924 40468 25930 40480
rect 26237 40477 26249 40480
rect 26283 40477 26295 40511
rect 26237 40471 26295 40477
rect 26418 40468 26424 40520
rect 26476 40468 26482 40520
rect 26878 40508 26884 40520
rect 26839 40480 26884 40508
rect 26878 40468 26884 40480
rect 26936 40468 26942 40520
rect 27985 40511 28043 40517
rect 27985 40477 27997 40511
rect 28031 40508 28043 40511
rect 28902 40508 28908 40520
rect 28031 40480 28908 40508
rect 28031 40477 28043 40480
rect 27985 40471 28043 40477
rect 28902 40468 28908 40480
rect 28960 40468 28966 40520
rect 29086 40468 29092 40520
rect 29144 40508 29150 40520
rect 29825 40511 29883 40517
rect 29825 40508 29837 40511
rect 29144 40480 29837 40508
rect 29144 40468 29150 40480
rect 29825 40477 29837 40480
rect 29871 40477 29883 40511
rect 29825 40471 29883 40477
rect 26234 40372 26240 40384
rect 25424 40344 26240 40372
rect 26234 40332 26240 40344
rect 26292 40332 26298 40384
rect 26436 40381 26464 40468
rect 26510 40400 26516 40452
rect 26568 40440 26574 40452
rect 28813 40443 28871 40449
rect 28813 40440 28825 40443
rect 26568 40412 28825 40440
rect 26568 40400 26574 40412
rect 28813 40409 28825 40412
rect 28859 40409 28871 40443
rect 28813 40403 28871 40409
rect 26421 40375 26479 40381
rect 26421 40341 26433 40375
rect 26467 40341 26479 40375
rect 27062 40372 27068 40384
rect 27023 40344 27068 40372
rect 26421 40335 26479 40341
rect 27062 40332 27068 40344
rect 27120 40332 27126 40384
rect 27801 40375 27859 40381
rect 27801 40341 27813 40375
rect 27847 40372 27859 40375
rect 28626 40372 28632 40384
rect 27847 40344 28632 40372
rect 27847 40341 27859 40344
rect 27801 40335 27859 40341
rect 28626 40332 28632 40344
rect 28684 40332 28690 40384
rect 30006 40372 30012 40384
rect 29967 40344 30012 40372
rect 30006 40332 30012 40344
rect 30064 40332 30070 40384
rect 1104 40282 30820 40304
rect 1104 40230 10880 40282
rect 10932 40230 10944 40282
rect 10996 40230 11008 40282
rect 11060 40230 11072 40282
rect 11124 40230 11136 40282
rect 11188 40230 20811 40282
rect 20863 40230 20875 40282
rect 20927 40230 20939 40282
rect 20991 40230 21003 40282
rect 21055 40230 21067 40282
rect 21119 40230 30820 40282
rect 1104 40208 30820 40230
rect 14642 40168 14648 40180
rect 14603 40140 14648 40168
rect 14642 40128 14648 40140
rect 14700 40128 14706 40180
rect 16574 40128 16580 40180
rect 16632 40168 16638 40180
rect 16669 40171 16727 40177
rect 16669 40168 16681 40171
rect 16632 40140 16681 40168
rect 16632 40128 16638 40140
rect 16669 40137 16681 40140
rect 16715 40137 16727 40171
rect 16669 40131 16727 40137
rect 17126 40128 17132 40180
rect 17184 40128 17190 40180
rect 21085 40171 21143 40177
rect 21085 40137 21097 40171
rect 21131 40168 21143 40171
rect 21450 40168 21456 40180
rect 21131 40140 21456 40168
rect 21131 40137 21143 40140
rect 21085 40131 21143 40137
rect 21450 40128 21456 40140
rect 21508 40128 21514 40180
rect 21913 40171 21971 40177
rect 21913 40137 21925 40171
rect 21959 40168 21971 40171
rect 22002 40168 22008 40180
rect 21959 40140 22008 40168
rect 21959 40137 21971 40140
rect 21913 40131 21971 40137
rect 22002 40128 22008 40140
rect 22060 40128 22066 40180
rect 22554 40168 22560 40180
rect 22515 40140 22560 40168
rect 22554 40128 22560 40140
rect 22612 40128 22618 40180
rect 22922 40128 22928 40180
rect 22980 40168 22986 40180
rect 25225 40171 25283 40177
rect 25225 40168 25237 40171
rect 22980 40140 25237 40168
rect 22980 40128 22986 40140
rect 25225 40137 25237 40140
rect 25271 40137 25283 40171
rect 25866 40168 25872 40180
rect 25827 40140 25872 40168
rect 25225 40131 25283 40137
rect 25866 40128 25872 40140
rect 25924 40128 25930 40180
rect 26234 40128 26240 40180
rect 26292 40168 26298 40180
rect 26786 40168 26792 40180
rect 26292 40140 26792 40168
rect 26292 40128 26298 40140
rect 26786 40128 26792 40140
rect 26844 40128 26850 40180
rect 27154 40128 27160 40180
rect 27212 40168 27218 40180
rect 27212 40140 27257 40168
rect 27212 40128 27218 40140
rect 27338 40128 27344 40180
rect 27396 40168 27402 40180
rect 29454 40168 29460 40180
rect 27396 40140 29460 40168
rect 27396 40128 27402 40140
rect 29454 40128 29460 40140
rect 29512 40128 29518 40180
rect 14550 40060 14556 40112
rect 14608 40100 14614 40112
rect 14608 40072 16896 40100
rect 14608 40060 14614 40072
rect 12066 40032 12072 40044
rect 12027 40004 12072 40032
rect 12066 39992 12072 40004
rect 12124 39992 12130 40044
rect 12250 40032 12256 40044
rect 12211 40004 12256 40032
rect 12250 39992 12256 40004
rect 12308 39992 12314 40044
rect 14366 39992 14372 40044
rect 14424 40032 14430 40044
rect 14829 40035 14887 40041
rect 14829 40032 14841 40035
rect 14424 40004 14841 40032
rect 14424 39992 14430 40004
rect 14829 40001 14841 40004
rect 14875 40001 14887 40035
rect 15102 40032 15108 40044
rect 15063 40004 15108 40032
rect 14829 39995 14887 40001
rect 15102 39992 15108 40004
rect 15160 39992 15166 40044
rect 16868 40041 16896 40072
rect 16853 40035 16911 40041
rect 16853 40001 16865 40035
rect 16899 40032 16911 40035
rect 16942 40032 16948 40044
rect 16899 40004 16948 40032
rect 16899 40001 16911 40004
rect 16853 39995 16911 40001
rect 16942 39992 16948 40004
rect 17000 39992 17006 40044
rect 17144 40041 17172 40128
rect 19702 40100 19708 40112
rect 19628 40072 19708 40100
rect 17129 40035 17187 40041
rect 17129 40001 17141 40035
rect 17175 40001 17187 40035
rect 17129 39995 17187 40001
rect 17678 39992 17684 40044
rect 17736 40032 17742 40044
rect 19429 40035 19487 40041
rect 19429 40032 19441 40035
rect 17736 40004 19441 40032
rect 17736 39992 17742 40004
rect 19429 40001 19441 40004
rect 19475 40032 19487 40035
rect 19518 40032 19524 40044
rect 19475 40004 19524 40032
rect 19475 40001 19487 40004
rect 19429 39995 19487 40001
rect 19518 39992 19524 40004
rect 19576 39992 19582 40044
rect 19628 40041 19656 40072
rect 19702 40060 19708 40072
rect 19760 40060 19766 40112
rect 20898 40100 20904 40112
rect 19996 40072 20904 40100
rect 19996 40041 20024 40072
rect 20898 40060 20904 40072
rect 20956 40060 20962 40112
rect 23290 40100 23296 40112
rect 22756 40072 23296 40100
rect 19613 40035 19671 40041
rect 19613 40001 19625 40035
rect 19659 40001 19671 40035
rect 19613 39995 19671 40001
rect 19981 40035 20039 40041
rect 19981 40001 19993 40035
rect 20027 40001 20039 40035
rect 20530 40032 20536 40044
rect 19981 39995 20039 40001
rect 20088 40004 20536 40032
rect 15013 39967 15071 39973
rect 15013 39933 15025 39967
rect 15059 39964 15071 39967
rect 15194 39964 15200 39976
rect 15059 39936 15200 39964
rect 15059 39933 15071 39936
rect 15013 39927 15071 39933
rect 15194 39924 15200 39936
rect 15252 39964 15258 39976
rect 17034 39964 17040 39976
rect 15252 39936 17040 39964
rect 15252 39924 15258 39936
rect 17034 39924 17040 39936
rect 17092 39924 17098 39976
rect 19702 39964 19708 39976
rect 19663 39936 19708 39964
rect 19702 39924 19708 39936
rect 19760 39924 19766 39976
rect 19797 39967 19855 39973
rect 19797 39933 19809 39967
rect 19843 39964 19855 39967
rect 20088 39964 20116 40004
rect 20530 39992 20536 40004
rect 20588 39992 20594 40044
rect 21266 40032 21272 40044
rect 21227 40004 21272 40032
rect 21266 39992 21272 40004
rect 21324 39992 21330 40044
rect 22094 39992 22100 40044
rect 22152 40032 22158 40044
rect 22756 40041 22784 40072
rect 23290 40060 23296 40072
rect 23348 40060 23354 40112
rect 23382 40060 23388 40112
rect 23440 40100 23446 40112
rect 26510 40100 26516 40112
rect 23440 40072 24707 40100
rect 23440 40060 23446 40072
rect 22741 40035 22799 40041
rect 22152 40004 22197 40032
rect 22152 39992 22158 40004
rect 22741 40001 22753 40035
rect 22787 40001 22799 40035
rect 22741 39995 22799 40001
rect 22830 39992 22836 40044
rect 22888 40032 22894 40044
rect 23201 40035 23259 40041
rect 23201 40032 23213 40035
rect 22888 40004 23213 40032
rect 22888 39992 22894 40004
rect 23201 40001 23213 40004
rect 23247 40001 23259 40035
rect 23842 40032 23848 40044
rect 23803 40004 23848 40032
rect 23201 39995 23259 40001
rect 23842 39992 23848 40004
rect 23900 39992 23906 40044
rect 24029 40035 24087 40041
rect 24029 40032 24041 40035
rect 23952 40004 24041 40032
rect 19843 39936 20116 39964
rect 19843 39933 19855 39936
rect 19797 39927 19855 39933
rect 23290 39924 23296 39976
rect 23348 39964 23354 39976
rect 23952 39964 23980 40004
rect 24029 40001 24041 40004
rect 24075 40001 24087 40035
rect 24029 39995 24087 40001
rect 24394 39992 24400 40044
rect 24452 40032 24458 40044
rect 24578 40032 24584 40044
rect 24452 40004 24497 40032
rect 24539 40004 24584 40032
rect 24452 39992 24458 40004
rect 24578 39992 24584 40004
rect 24636 39992 24642 40044
rect 24679 40032 24707 40072
rect 25700 40072 26516 40100
rect 25700 40041 25728 40072
rect 26510 40060 26516 40072
rect 26568 40060 26574 40112
rect 26694 40060 26700 40112
rect 26752 40100 26758 40112
rect 29086 40100 29092 40112
rect 26752 40072 29092 40100
rect 26752 40060 26758 40072
rect 29086 40060 29092 40072
rect 29144 40060 29150 40112
rect 25041 40035 25099 40041
rect 25041 40032 25053 40035
rect 24679 40004 25053 40032
rect 25041 40001 25053 40004
rect 25087 40001 25099 40035
rect 25041 39995 25099 40001
rect 25685 40035 25743 40041
rect 25685 40001 25697 40035
rect 25731 40001 25743 40035
rect 26970 40032 26976 40044
rect 26931 40004 26976 40032
rect 25685 39995 25743 40001
rect 26970 39992 26976 40004
rect 27028 39992 27034 40044
rect 28353 40035 28411 40041
rect 28353 40001 28365 40035
rect 28399 40032 28411 40035
rect 28442 40032 28448 40044
rect 28399 40004 28448 40032
rect 28399 40001 28411 40004
rect 28353 39995 28411 40001
rect 28442 39992 28448 40004
rect 28500 39992 28506 40044
rect 28810 39992 28816 40044
rect 28868 40032 28874 40044
rect 28997 40035 29055 40041
rect 28997 40032 29009 40035
rect 28868 40004 29009 40032
rect 28868 39992 28874 40004
rect 28997 40001 29009 40004
rect 29043 40001 29055 40035
rect 28997 39995 29055 40001
rect 29825 40035 29883 40041
rect 29825 40001 29837 40035
rect 29871 40001 29883 40035
rect 29825 39995 29883 40001
rect 24118 39964 24124 39976
rect 23348 39936 23980 39964
rect 24079 39936 24124 39964
rect 23348 39924 23354 39936
rect 24118 39924 24124 39936
rect 24176 39924 24182 39976
rect 24213 39967 24271 39973
rect 24213 39933 24225 39967
rect 24259 39964 24271 39967
rect 24302 39964 24308 39976
rect 24259 39936 24308 39964
rect 24259 39933 24271 39936
rect 24213 39927 24271 39933
rect 24302 39924 24308 39936
rect 24360 39924 24366 39976
rect 24486 39924 24492 39976
rect 24544 39964 24550 39976
rect 29638 39964 29644 39976
rect 24544 39936 29644 39964
rect 24544 39924 24550 39936
rect 29638 39924 29644 39936
rect 29696 39924 29702 39976
rect 12437 39899 12495 39905
rect 12437 39865 12449 39899
rect 12483 39896 12495 39899
rect 23198 39896 23204 39908
rect 12483 39868 23204 39896
rect 12483 39865 12495 39868
rect 12437 39859 12495 39865
rect 23198 39856 23204 39868
rect 23256 39856 23262 39908
rect 23382 39896 23388 39908
rect 23343 39868 23388 39896
rect 23382 39856 23388 39868
rect 23440 39856 23446 39908
rect 29840 39896 29868 39995
rect 24423 39868 29868 39896
rect 16942 39788 16948 39840
rect 17000 39828 17006 39840
rect 17586 39828 17592 39840
rect 17000 39800 17592 39828
rect 17000 39788 17006 39800
rect 17586 39788 17592 39800
rect 17644 39788 17650 39840
rect 20162 39828 20168 39840
rect 20123 39800 20168 39828
rect 20162 39788 20168 39800
rect 20220 39788 20226 39840
rect 20898 39788 20904 39840
rect 20956 39828 20962 39840
rect 21266 39828 21272 39840
rect 20956 39800 21272 39828
rect 20956 39788 20962 39800
rect 21266 39788 21272 39800
rect 21324 39788 21330 39840
rect 23658 39788 23664 39840
rect 23716 39828 23722 39840
rect 24423 39828 24451 39868
rect 23716 39800 24451 39828
rect 23716 39788 23722 39800
rect 24762 39788 24768 39840
rect 24820 39828 24826 39840
rect 25314 39828 25320 39840
rect 24820 39800 25320 39828
rect 24820 39788 24826 39800
rect 25314 39788 25320 39800
rect 25372 39788 25378 39840
rect 26234 39788 26240 39840
rect 26292 39828 26298 39840
rect 27246 39828 27252 39840
rect 26292 39800 27252 39828
rect 26292 39788 26298 39800
rect 27246 39788 27252 39800
rect 27304 39788 27310 39840
rect 28166 39828 28172 39840
rect 28127 39800 28172 39828
rect 28166 39788 28172 39800
rect 28224 39788 28230 39840
rect 28813 39831 28871 39837
rect 28813 39797 28825 39831
rect 28859 39828 28871 39831
rect 29362 39828 29368 39840
rect 28859 39800 29368 39828
rect 28859 39797 28871 39800
rect 28813 39791 28871 39797
rect 29362 39788 29368 39800
rect 29420 39788 29426 39840
rect 30009 39831 30067 39837
rect 30009 39797 30021 39831
rect 30055 39828 30067 39831
rect 30098 39828 30104 39840
rect 30055 39800 30104 39828
rect 30055 39797 30067 39800
rect 30009 39791 30067 39797
rect 30098 39788 30104 39800
rect 30156 39788 30162 39840
rect 1104 39738 30820 39760
rect 1104 39686 5915 39738
rect 5967 39686 5979 39738
rect 6031 39686 6043 39738
rect 6095 39686 6107 39738
rect 6159 39686 6171 39738
rect 6223 39686 15846 39738
rect 15898 39686 15910 39738
rect 15962 39686 15974 39738
rect 16026 39686 16038 39738
rect 16090 39686 16102 39738
rect 16154 39686 25776 39738
rect 25828 39686 25840 39738
rect 25892 39686 25904 39738
rect 25956 39686 25968 39738
rect 26020 39686 26032 39738
rect 26084 39686 30820 39738
rect 1104 39664 30820 39686
rect 19610 39624 19616 39636
rect 19571 39596 19616 39624
rect 19610 39584 19616 39596
rect 19668 39584 19674 39636
rect 22738 39584 22744 39636
rect 22796 39624 22802 39636
rect 22925 39627 22983 39633
rect 22925 39624 22937 39627
rect 22796 39596 22937 39624
rect 22796 39584 22802 39596
rect 22925 39593 22937 39596
rect 22971 39593 22983 39627
rect 22925 39587 22983 39593
rect 23198 39584 23204 39636
rect 23256 39624 23262 39636
rect 24854 39624 24860 39636
rect 23256 39596 24860 39624
rect 23256 39584 23262 39596
rect 24854 39584 24860 39596
rect 24912 39584 24918 39636
rect 25130 39624 25136 39636
rect 25091 39596 25136 39624
rect 25130 39584 25136 39596
rect 25188 39584 25194 39636
rect 27614 39624 27620 39636
rect 25240 39596 27620 39624
rect 19702 39556 19708 39568
rect 17972 39528 19708 39556
rect 16574 39488 16580 39500
rect 15212 39460 16580 39488
rect 1578 39420 1584 39432
rect 1539 39392 1584 39420
rect 1578 39380 1584 39392
rect 1636 39380 1642 39432
rect 15212 39429 15240 39460
rect 16574 39448 16580 39460
rect 16632 39448 16638 39500
rect 17770 39448 17776 39500
rect 17828 39488 17834 39500
rect 17972 39497 18000 39528
rect 19702 39516 19708 39528
rect 19760 39516 19766 39568
rect 22097 39559 22155 39565
rect 22097 39525 22109 39559
rect 22143 39556 22155 39559
rect 25240 39556 25268 39596
rect 27614 39584 27620 39596
rect 27672 39584 27678 39636
rect 29178 39584 29184 39636
rect 29236 39624 29242 39636
rect 29917 39627 29975 39633
rect 29917 39624 29929 39627
rect 29236 39596 29929 39624
rect 29236 39584 29242 39596
rect 29917 39593 29929 39596
rect 29963 39593 29975 39627
rect 29917 39587 29975 39593
rect 22143 39528 25268 39556
rect 22143 39525 22155 39528
rect 22097 39519 22155 39525
rect 25314 39516 25320 39568
rect 25372 39556 25378 39568
rect 25958 39556 25964 39568
rect 25372 39528 25964 39556
rect 25372 39516 25378 39528
rect 25958 39516 25964 39528
rect 26016 39516 26022 39568
rect 26252 39528 27476 39556
rect 17957 39491 18015 39497
rect 17957 39488 17969 39491
rect 17828 39460 17969 39488
rect 17828 39448 17834 39460
rect 17957 39457 17969 39460
rect 18003 39457 18015 39491
rect 17957 39451 18015 39457
rect 18506 39448 18512 39500
rect 18564 39488 18570 39500
rect 20257 39491 20315 39497
rect 20257 39488 20269 39491
rect 18564 39460 20269 39488
rect 18564 39448 18570 39460
rect 20257 39457 20269 39460
rect 20303 39457 20315 39491
rect 20257 39451 20315 39457
rect 21450 39448 21456 39500
rect 21508 39488 21514 39500
rect 21634 39488 21640 39500
rect 21508 39460 21640 39488
rect 21508 39448 21514 39460
rect 21634 39448 21640 39460
rect 21692 39448 21698 39500
rect 23474 39488 23480 39500
rect 22066 39460 23480 39488
rect 15197 39423 15255 39429
rect 15197 39389 15209 39423
rect 15243 39389 15255 39423
rect 15378 39420 15384 39432
rect 15339 39392 15384 39420
rect 15197 39383 15255 39389
rect 15378 39380 15384 39392
rect 15436 39380 15442 39432
rect 15470 39380 15476 39432
rect 15528 39420 15534 39432
rect 15654 39429 15660 39432
rect 15611 39423 15660 39429
rect 15528 39392 15573 39420
rect 15528 39380 15534 39392
rect 15611 39389 15623 39423
rect 15657 39389 15660 39423
rect 15611 39383 15660 39389
rect 15654 39380 15660 39383
rect 15712 39380 15718 39432
rect 15760 39423 15818 39429
rect 15760 39389 15772 39423
rect 15806 39420 15818 39423
rect 16022 39420 16028 39432
rect 15806 39392 16028 39420
rect 15806 39389 15818 39392
rect 15760 39383 15818 39389
rect 16022 39380 16028 39392
rect 16080 39380 16086 39432
rect 17678 39420 17684 39432
rect 17639 39392 17684 39420
rect 17678 39380 17684 39392
rect 17736 39380 17742 39432
rect 17862 39420 17868 39432
rect 17823 39392 17868 39420
rect 17862 39380 17868 39392
rect 17920 39380 17926 39432
rect 18049 39423 18107 39429
rect 18049 39389 18061 39423
rect 18095 39389 18107 39423
rect 18230 39420 18236 39432
rect 18191 39392 18236 39420
rect 18049 39383 18107 39389
rect 15672 39352 15700 39380
rect 18064 39352 18092 39383
rect 18230 39380 18236 39392
rect 18288 39380 18294 39432
rect 19797 39423 19855 39429
rect 19797 39389 19809 39423
rect 19843 39420 19855 39423
rect 22066 39420 22094 39460
rect 23474 39448 23480 39460
rect 23532 39448 23538 39500
rect 23753 39491 23811 39497
rect 23753 39457 23765 39491
rect 23799 39488 23811 39491
rect 24762 39488 24768 39500
rect 23799 39460 24768 39488
rect 23799 39457 23811 39460
rect 23753 39451 23811 39457
rect 24762 39448 24768 39460
rect 24820 39448 24826 39500
rect 25590 39448 25596 39500
rect 25648 39488 25654 39500
rect 26252 39497 26280 39528
rect 26237 39491 26295 39497
rect 26237 39488 26249 39491
rect 25648 39460 26249 39488
rect 25648 39448 25654 39460
rect 26237 39457 26249 39460
rect 26283 39457 26295 39491
rect 26786 39488 26792 39500
rect 26237 39451 26295 39457
rect 26436 39460 26792 39488
rect 22278 39420 22284 39432
rect 19843 39392 22094 39420
rect 22239 39392 22284 39420
rect 19843 39389 19855 39392
rect 19797 39383 19855 39389
rect 22278 39380 22284 39392
rect 22336 39380 22342 39432
rect 22741 39423 22799 39429
rect 22741 39389 22753 39423
rect 22787 39420 22799 39423
rect 22830 39420 22836 39432
rect 22787 39392 22836 39420
rect 22787 39389 22799 39392
rect 22741 39383 22799 39389
rect 22830 39380 22836 39392
rect 22888 39380 22894 39432
rect 23661 39423 23719 39429
rect 23661 39389 23673 39423
rect 23707 39389 23719 39423
rect 23661 39383 23719 39389
rect 18782 39352 18788 39364
rect 15672 39324 18788 39352
rect 18782 39312 18788 39324
rect 18840 39312 18846 39364
rect 20524 39355 20582 39361
rect 20524 39321 20536 39355
rect 20570 39352 20582 39355
rect 20714 39352 20720 39364
rect 20570 39324 20720 39352
rect 20570 39321 20582 39324
rect 20524 39315 20582 39321
rect 20714 39312 20720 39324
rect 20772 39312 20778 39364
rect 23566 39312 23572 39364
rect 23624 39352 23630 39364
rect 23676 39352 23704 39383
rect 23842 39380 23848 39432
rect 23900 39420 23906 39432
rect 24302 39420 24308 39432
rect 23900 39392 24308 39420
rect 23900 39380 23906 39392
rect 24302 39380 24308 39392
rect 24360 39420 24366 39432
rect 24397 39423 24455 39429
rect 24397 39420 24409 39423
rect 24360 39392 24409 39420
rect 24360 39380 24366 39392
rect 24397 39389 24409 39392
rect 24443 39389 24455 39423
rect 24397 39383 24455 39389
rect 24486 39380 24492 39432
rect 24544 39420 24550 39432
rect 24581 39423 24639 39429
rect 24581 39420 24593 39423
rect 24544 39392 24593 39420
rect 24544 39380 24550 39392
rect 24581 39389 24593 39392
rect 24627 39389 24639 39423
rect 24581 39383 24639 39389
rect 24673 39423 24731 39429
rect 24673 39389 24685 39423
rect 24719 39389 24731 39423
rect 24673 39383 24731 39389
rect 24949 39423 25007 39429
rect 24949 39389 24961 39423
rect 24995 39420 25007 39423
rect 25406 39420 25412 39432
rect 24995 39392 25412 39420
rect 24995 39389 25007 39392
rect 24949 39383 25007 39389
rect 24210 39352 24216 39364
rect 23624 39324 24216 39352
rect 23624 39312 23630 39324
rect 24210 39312 24216 39324
rect 24268 39352 24274 39364
rect 24688 39352 24716 39383
rect 25406 39380 25412 39392
rect 25464 39380 25470 39432
rect 25869 39423 25927 39429
rect 25869 39389 25881 39423
rect 25915 39389 25927 39423
rect 25869 39383 25927 39389
rect 24268 39324 24716 39352
rect 24268 39312 24274 39324
rect 24854 39312 24860 39364
rect 24912 39352 24918 39364
rect 25498 39352 25504 39364
rect 24912 39324 25504 39352
rect 24912 39312 24918 39324
rect 25498 39312 25504 39324
rect 25556 39312 25562 39364
rect 25682 39312 25688 39364
rect 25740 39352 25746 39364
rect 25884 39352 25912 39383
rect 25958 39380 25964 39432
rect 26016 39420 26022 39432
rect 26053 39423 26111 39429
rect 26053 39420 26065 39423
rect 26016 39392 26065 39420
rect 26016 39380 26022 39392
rect 26053 39389 26065 39392
rect 26099 39389 26111 39423
rect 26053 39383 26111 39389
rect 26142 39380 26148 39432
rect 26200 39420 26206 39432
rect 26436 39429 26464 39460
rect 26786 39448 26792 39460
rect 26844 39448 26850 39500
rect 27448 39497 27476 39528
rect 27522 39516 27528 39568
rect 27580 39556 27586 39568
rect 27580 39528 28488 39556
rect 27580 39516 27586 39528
rect 27433 39491 27491 39497
rect 27433 39457 27445 39491
rect 27479 39457 27491 39491
rect 28460 39488 28488 39528
rect 28534 39516 28540 39568
rect 28592 39556 28598 39568
rect 30101 39559 30159 39565
rect 30101 39556 30113 39559
rect 28592 39528 30113 39556
rect 28592 39516 28598 39528
rect 30101 39525 30113 39528
rect 30147 39525 30159 39559
rect 30101 39519 30159 39525
rect 30929 39491 30987 39497
rect 30929 39488 30941 39491
rect 28460 39460 30941 39488
rect 27433 39451 27491 39457
rect 30929 39457 30941 39460
rect 30975 39457 30987 39491
rect 30929 39451 30987 39457
rect 26421 39423 26479 39429
rect 26200 39392 26245 39420
rect 26200 39380 26206 39392
rect 26421 39389 26433 39423
rect 26467 39389 26479 39423
rect 26602 39420 26608 39432
rect 26563 39392 26608 39420
rect 26421 39383 26479 39389
rect 26602 39380 26608 39392
rect 26660 39380 26666 39432
rect 27065 39423 27123 39429
rect 27065 39389 27077 39423
rect 27111 39389 27123 39423
rect 27246 39420 27252 39432
rect 27207 39392 27252 39420
rect 27065 39383 27123 39389
rect 27080 39352 27108 39383
rect 27246 39380 27252 39392
rect 27304 39380 27310 39432
rect 27341 39423 27399 39429
rect 27341 39389 27353 39423
rect 27387 39389 27399 39423
rect 27341 39383 27399 39389
rect 27617 39423 27675 39429
rect 27617 39389 27629 39423
rect 27663 39420 27675 39423
rect 28534 39420 28540 39432
rect 27663 39392 28540 39420
rect 27663 39389 27675 39392
rect 27617 39383 27675 39389
rect 25740 39324 27108 39352
rect 25740 39312 25746 39324
rect 1397 39287 1455 39293
rect 1397 39253 1409 39287
rect 1443 39284 1455 39287
rect 12066 39284 12072 39296
rect 1443 39256 12072 39284
rect 1443 39253 1455 39256
rect 1397 39247 1455 39253
rect 12066 39244 12072 39256
rect 12124 39244 12130 39296
rect 15930 39284 15936 39296
rect 15891 39256 15936 39284
rect 15930 39244 15936 39256
rect 15988 39244 15994 39296
rect 18414 39284 18420 39296
rect 18375 39256 18420 39284
rect 18414 39244 18420 39256
rect 18472 39244 18478 39296
rect 19150 39244 19156 39296
rect 19208 39284 19214 39296
rect 20346 39284 20352 39296
rect 19208 39256 20352 39284
rect 19208 39244 19214 39256
rect 20346 39244 20352 39256
rect 20404 39244 20410 39296
rect 21634 39284 21640 39296
rect 21595 39256 21640 39284
rect 21634 39244 21640 39256
rect 21692 39244 21698 39296
rect 22094 39244 22100 39296
rect 22152 39284 22158 39296
rect 26050 39284 26056 39296
rect 22152 39256 26056 39284
rect 22152 39244 22158 39256
rect 26050 39244 26056 39256
rect 26108 39244 26114 39296
rect 26142 39244 26148 39296
rect 26200 39284 26206 39296
rect 27356 39284 27384 39383
rect 28534 39380 28540 39392
rect 28592 39380 28598 39432
rect 28718 39420 28724 39432
rect 28679 39392 28724 39420
rect 28718 39380 28724 39392
rect 28776 39380 28782 39432
rect 29086 39380 29092 39432
rect 29144 39420 29150 39432
rect 29549 39423 29607 39429
rect 29549 39420 29561 39423
rect 29144 39392 29561 39420
rect 29144 39380 29150 39392
rect 29549 39389 29561 39392
rect 29595 39389 29607 39423
rect 29549 39383 29607 39389
rect 28350 39312 28356 39364
rect 28408 39352 28414 39364
rect 29917 39355 29975 39361
rect 29917 39352 29929 39355
rect 28408 39324 29929 39352
rect 28408 39312 28414 39324
rect 29917 39321 29929 39324
rect 29963 39321 29975 39355
rect 29917 39315 29975 39321
rect 27798 39284 27804 39296
rect 26200 39256 27384 39284
rect 27759 39256 27804 39284
rect 26200 39244 26206 39256
rect 27798 39244 27804 39256
rect 27856 39244 27862 39296
rect 28902 39284 28908 39296
rect 28863 39256 28908 39284
rect 28902 39244 28908 39256
rect 28960 39244 28966 39296
rect 1104 39194 30820 39216
rect 1104 39142 10880 39194
rect 10932 39142 10944 39194
rect 10996 39142 11008 39194
rect 11060 39142 11072 39194
rect 11124 39142 11136 39194
rect 11188 39142 20811 39194
rect 20863 39142 20875 39194
rect 20927 39142 20939 39194
rect 20991 39142 21003 39194
rect 21055 39142 21067 39194
rect 21119 39142 30820 39194
rect 1104 39120 30820 39142
rect 15746 39040 15752 39092
rect 15804 39080 15810 39092
rect 16022 39080 16028 39092
rect 15804 39052 16028 39080
rect 15804 39040 15810 39052
rect 16022 39040 16028 39052
rect 16080 39040 16086 39092
rect 20714 39040 20720 39092
rect 20772 39080 20778 39092
rect 21085 39083 21143 39089
rect 21085 39080 21097 39083
rect 20772 39052 21097 39080
rect 20772 39040 20778 39052
rect 21085 39049 21097 39052
rect 21131 39049 21143 39083
rect 21085 39043 21143 39049
rect 22094 39040 22100 39092
rect 22152 39080 22158 39092
rect 23014 39080 23020 39092
rect 22152 39052 22197 39080
rect 22975 39052 23020 39080
rect 22152 39040 22158 39052
rect 23014 39040 23020 39052
rect 23072 39040 23078 39092
rect 23658 39080 23664 39092
rect 23619 39052 23664 39080
rect 23658 39040 23664 39052
rect 23716 39040 23722 39092
rect 23750 39040 23756 39092
rect 23808 39080 23814 39092
rect 28534 39080 28540 39092
rect 23808 39052 27936 39080
rect 28495 39052 28540 39080
rect 23808 39040 23814 39052
rect 14660 38984 16712 39012
rect 12066 38944 12072 38956
rect 12027 38916 12072 38944
rect 12066 38904 12072 38916
rect 12124 38904 12130 38956
rect 12250 38944 12256 38956
rect 12211 38916 12256 38944
rect 12250 38904 12256 38916
rect 12308 38904 12314 38956
rect 14090 38836 14096 38888
rect 14148 38876 14154 38888
rect 14660 38885 14688 38984
rect 16684 38956 16712 38984
rect 18414 38972 18420 39024
rect 18472 39012 18478 39024
rect 18754 39015 18812 39021
rect 18754 39012 18766 39015
rect 18472 38984 18766 39012
rect 18472 38972 18478 38984
rect 18754 38981 18766 38984
rect 18800 38981 18812 39015
rect 21174 39012 21180 39024
rect 18754 38975 18812 38981
rect 20548 38984 21180 39012
rect 14912 38947 14970 38953
rect 14912 38913 14924 38947
rect 14958 38944 14970 38947
rect 15930 38944 15936 38956
rect 14958 38916 15936 38944
rect 14958 38913 14970 38916
rect 14912 38907 14970 38913
rect 15930 38904 15936 38916
rect 15988 38904 15994 38956
rect 16666 38944 16672 38956
rect 16579 38916 16672 38944
rect 16666 38904 16672 38916
rect 16724 38904 16730 38956
rect 16942 38953 16948 38956
rect 16936 38907 16948 38953
rect 17000 38944 17006 38956
rect 18506 38944 18512 38956
rect 17000 38916 17036 38944
rect 18467 38916 18512 38944
rect 16942 38904 16948 38907
rect 17000 38904 17006 38916
rect 18506 38904 18512 38916
rect 18564 38904 18570 38956
rect 19150 38944 19156 38956
rect 18616 38916 19156 38944
rect 14645 38879 14703 38885
rect 14645 38876 14657 38879
rect 14148 38848 14657 38876
rect 14148 38836 14154 38848
rect 14645 38845 14657 38848
rect 14691 38845 14703 38879
rect 18616 38876 18644 38916
rect 19150 38904 19156 38916
rect 19208 38904 19214 38956
rect 19518 38904 19524 38956
rect 19576 38944 19582 38956
rect 19978 38944 19984 38956
rect 19576 38916 19984 38944
rect 19576 38904 19582 38916
rect 19978 38904 19984 38916
rect 20036 38944 20042 38956
rect 20548 38953 20576 38984
rect 21174 38972 21180 38984
rect 21232 38972 21238 39024
rect 26326 39012 26332 39024
rect 22296 38984 26332 39012
rect 20349 38947 20407 38953
rect 20349 38944 20361 38947
rect 20036 38916 20361 38944
rect 20036 38904 20042 38916
rect 20349 38913 20361 38916
rect 20395 38913 20407 38947
rect 20349 38907 20407 38913
rect 20533 38947 20591 38953
rect 20533 38913 20545 38947
rect 20579 38913 20591 38947
rect 20533 38907 20591 38913
rect 20901 38947 20959 38953
rect 20901 38913 20913 38947
rect 20947 38944 20959 38947
rect 21634 38944 21640 38956
rect 20947 38916 21640 38944
rect 20947 38913 20959 38916
rect 20901 38907 20959 38913
rect 21634 38904 21640 38916
rect 21692 38904 21698 38956
rect 22296 38953 22324 38984
rect 26326 38972 26332 38984
rect 26384 38972 26390 39024
rect 27424 39015 27482 39021
rect 27424 38981 27436 39015
rect 27470 39012 27482 39015
rect 27798 39012 27804 39024
rect 27470 38984 27804 39012
rect 27470 38981 27482 38984
rect 27424 38975 27482 38981
rect 27798 38972 27804 38984
rect 27856 38972 27862 39024
rect 27908 39012 27936 39052
rect 28534 39040 28540 39052
rect 28592 39080 28598 39092
rect 29365 39083 29423 39089
rect 29365 39080 29377 39083
rect 28592 39052 29377 39080
rect 28592 39040 28598 39052
rect 29365 39049 29377 39052
rect 29411 39049 29423 39083
rect 29365 39043 29423 39049
rect 29549 39083 29607 39089
rect 29549 39049 29561 39083
rect 29595 39049 29607 39083
rect 29549 39043 29607 39049
rect 29564 39012 29592 39043
rect 27908 38984 29592 39012
rect 22281 38947 22339 38953
rect 22281 38913 22293 38947
rect 22327 38913 22339 38947
rect 22281 38907 22339 38913
rect 23201 38947 23259 38953
rect 23201 38913 23213 38947
rect 23247 38944 23259 38947
rect 23750 38944 23756 38956
rect 23247 38916 23756 38944
rect 23247 38913 23259 38916
rect 23201 38907 23259 38913
rect 23750 38904 23756 38916
rect 23808 38904 23814 38956
rect 23845 38947 23903 38953
rect 23845 38913 23857 38947
rect 23891 38913 23903 38947
rect 24302 38944 24308 38956
rect 24263 38916 24308 38944
rect 23845 38907 23903 38913
rect 14645 38839 14703 38845
rect 17696 38848 18644 38876
rect 12437 38743 12495 38749
rect 12437 38709 12449 38743
rect 12483 38740 12495 38743
rect 17696 38740 17724 38848
rect 19702 38836 19708 38888
rect 19760 38876 19766 38888
rect 20625 38879 20683 38885
rect 20625 38876 20637 38879
rect 19760 38848 20637 38876
rect 19760 38836 19766 38848
rect 20625 38845 20637 38848
rect 20671 38845 20683 38879
rect 20625 38839 20683 38845
rect 20717 38879 20775 38885
rect 20717 38845 20729 38879
rect 20763 38845 20775 38879
rect 20717 38839 20775 38845
rect 20530 38768 20536 38820
rect 20588 38808 20594 38820
rect 20732 38808 20760 38839
rect 20588 38780 20760 38808
rect 23860 38808 23888 38907
rect 24302 38904 24308 38916
rect 24360 38904 24366 38956
rect 24394 38904 24400 38956
rect 24452 38944 24458 38956
rect 24489 38947 24547 38953
rect 24489 38944 24501 38947
rect 24452 38916 24501 38944
rect 24452 38904 24458 38916
rect 24489 38913 24501 38916
rect 24535 38913 24547 38947
rect 24670 38944 24676 38956
rect 24631 38916 24676 38944
rect 24489 38907 24547 38913
rect 24670 38904 24676 38916
rect 24728 38904 24734 38956
rect 24857 38947 24915 38953
rect 24857 38913 24869 38947
rect 24903 38944 24915 38947
rect 25498 38944 25504 38956
rect 24903 38916 25504 38944
rect 24903 38913 24915 38916
rect 24857 38907 24915 38913
rect 25498 38904 25504 38916
rect 25556 38904 25562 38956
rect 25682 38944 25688 38956
rect 25643 38916 25688 38944
rect 25682 38904 25688 38916
rect 25740 38904 25746 38956
rect 25774 38904 25780 38956
rect 25832 38944 25838 38956
rect 25869 38947 25927 38953
rect 25869 38944 25881 38947
rect 25832 38916 25881 38944
rect 25832 38904 25838 38916
rect 25869 38913 25881 38916
rect 25915 38913 25927 38947
rect 25869 38907 25927 38913
rect 25961 38947 26019 38953
rect 25961 38913 25973 38947
rect 26007 38944 26019 38947
rect 26142 38944 26148 38956
rect 26007 38916 26148 38944
rect 26007 38913 26019 38916
rect 25961 38907 26019 38913
rect 26142 38904 26148 38916
rect 26200 38904 26206 38956
rect 26237 38947 26295 38953
rect 26237 38913 26249 38947
rect 26283 38913 26295 38947
rect 26237 38907 26295 38913
rect 24210 38836 24216 38888
rect 24268 38876 24274 38888
rect 24581 38879 24639 38885
rect 24581 38876 24593 38879
rect 24268 38848 24593 38876
rect 24268 38836 24274 38848
rect 24581 38845 24593 38848
rect 24627 38845 24639 38879
rect 24581 38839 24639 38845
rect 25590 38836 25596 38888
rect 25648 38876 25654 38888
rect 26053 38879 26111 38885
rect 26053 38876 26065 38879
rect 25648 38848 26065 38876
rect 25648 38836 25654 38848
rect 26053 38845 26065 38848
rect 26099 38845 26111 38879
rect 26252 38876 26280 38907
rect 27062 38904 27068 38956
rect 27120 38944 27126 38956
rect 27157 38947 27215 38953
rect 27157 38944 27169 38947
rect 27120 38916 27169 38944
rect 27120 38904 27126 38916
rect 27157 38913 27169 38916
rect 27203 38913 27215 38947
rect 28350 38944 28356 38956
rect 27157 38907 27215 38913
rect 27264 38916 28356 38944
rect 27264 38876 27292 38916
rect 28350 38904 28356 38916
rect 28408 38904 28414 38956
rect 26252 38848 27292 38876
rect 26053 38839 26111 38845
rect 25406 38808 25412 38820
rect 23860 38780 25412 38808
rect 20588 38768 20594 38780
rect 25406 38768 25412 38780
rect 25464 38768 25470 38820
rect 25774 38768 25780 38820
rect 25832 38808 25838 38820
rect 26326 38808 26332 38820
rect 25832 38780 26332 38808
rect 25832 38768 25838 38780
rect 26326 38768 26332 38780
rect 26384 38768 26390 38820
rect 28997 38811 29055 38817
rect 28997 38777 29009 38811
rect 29043 38808 29055 38811
rect 29086 38808 29092 38820
rect 29043 38780 29092 38808
rect 29043 38777 29055 38780
rect 28997 38771 29055 38777
rect 29086 38768 29092 38780
rect 29144 38768 29150 38820
rect 18046 38740 18052 38752
rect 12483 38712 17724 38740
rect 18007 38712 18052 38740
rect 12483 38709 12495 38712
rect 12437 38703 12495 38709
rect 18046 38700 18052 38712
rect 18104 38700 18110 38752
rect 18230 38700 18236 38752
rect 18288 38740 18294 38752
rect 19889 38743 19947 38749
rect 19889 38740 19901 38743
rect 18288 38712 19901 38740
rect 18288 38700 18294 38712
rect 19889 38709 19901 38712
rect 19935 38709 19947 38743
rect 19889 38703 19947 38709
rect 24946 38700 24952 38752
rect 25004 38740 25010 38752
rect 25041 38743 25099 38749
rect 25041 38740 25053 38743
rect 25004 38712 25053 38740
rect 25004 38700 25010 38712
rect 25041 38709 25053 38712
rect 25087 38709 25099 38743
rect 25041 38703 25099 38709
rect 26421 38743 26479 38749
rect 26421 38709 26433 38743
rect 26467 38740 26479 38743
rect 27062 38740 27068 38752
rect 26467 38712 27068 38740
rect 26467 38709 26479 38712
rect 26421 38703 26479 38709
rect 27062 38700 27068 38712
rect 27120 38700 27126 38752
rect 29362 38740 29368 38752
rect 29323 38712 29368 38740
rect 29362 38700 29368 38712
rect 29420 38700 29426 38752
rect 1104 38650 30820 38672
rect 1104 38598 5915 38650
rect 5967 38598 5979 38650
rect 6031 38598 6043 38650
rect 6095 38598 6107 38650
rect 6159 38598 6171 38650
rect 6223 38598 15846 38650
rect 15898 38598 15910 38650
rect 15962 38598 15974 38650
rect 16026 38598 16038 38650
rect 16090 38598 16102 38650
rect 16154 38598 25776 38650
rect 25828 38598 25840 38650
rect 25892 38598 25904 38650
rect 25956 38598 25968 38650
rect 26020 38598 26032 38650
rect 26084 38598 30820 38650
rect 1104 38576 30820 38598
rect 16853 38539 16911 38545
rect 16853 38505 16865 38539
rect 16899 38536 16911 38539
rect 16942 38536 16948 38548
rect 16899 38508 16948 38536
rect 16899 38505 16911 38508
rect 16853 38499 16911 38505
rect 16942 38496 16948 38508
rect 17000 38496 17006 38548
rect 20070 38536 20076 38548
rect 19812 38508 20076 38536
rect 15654 38428 15660 38480
rect 15712 38468 15718 38480
rect 19610 38468 19616 38480
rect 15712 38440 16528 38468
rect 15712 38428 15718 38440
rect 15194 38360 15200 38412
rect 15252 38400 15258 38412
rect 15470 38400 15476 38412
rect 15252 38372 15476 38400
rect 15252 38360 15258 38372
rect 15470 38360 15476 38372
rect 15528 38400 15534 38412
rect 16500 38409 16528 38440
rect 18524 38440 19616 38468
rect 16393 38403 16451 38409
rect 16393 38400 16405 38403
rect 15528 38372 16405 38400
rect 15528 38360 15534 38372
rect 16393 38369 16405 38372
rect 16439 38369 16451 38403
rect 16393 38363 16451 38369
rect 16485 38403 16543 38409
rect 16485 38369 16497 38403
rect 16531 38369 16543 38403
rect 18046 38400 18052 38412
rect 16485 38363 16543 38369
rect 17328 38372 18052 38400
rect 10134 38332 10140 38344
rect 10095 38304 10140 38332
rect 10134 38292 10140 38304
rect 10192 38292 10198 38344
rect 14090 38332 14096 38344
rect 14051 38304 14096 38332
rect 14090 38292 14096 38304
rect 14148 38292 14154 38344
rect 16117 38335 16175 38341
rect 16117 38301 16129 38335
rect 16163 38301 16175 38335
rect 16298 38332 16304 38344
rect 16259 38304 16304 38332
rect 16117 38295 16175 38301
rect 10404 38267 10462 38273
rect 10404 38233 10416 38267
rect 10450 38264 10462 38267
rect 10594 38264 10600 38276
rect 10450 38236 10600 38264
rect 10450 38233 10462 38236
rect 10404 38227 10462 38233
rect 10594 38224 10600 38236
rect 10652 38224 10658 38276
rect 14360 38267 14418 38273
rect 14360 38233 14372 38267
rect 14406 38264 14418 38267
rect 15378 38264 15384 38276
rect 14406 38236 15384 38264
rect 14406 38233 14418 38236
rect 14360 38227 14418 38233
rect 15378 38224 15384 38236
rect 15436 38224 15442 38276
rect 16132 38264 16160 38295
rect 16298 38292 16304 38304
rect 16356 38292 16362 38344
rect 17328 38341 17356 38372
rect 18046 38360 18052 38372
rect 18104 38360 18110 38412
rect 16669 38335 16727 38341
rect 16669 38301 16681 38335
rect 16715 38332 16727 38335
rect 17313 38335 17371 38341
rect 17313 38332 17325 38335
rect 16715 38304 17325 38332
rect 16715 38301 16727 38304
rect 16669 38295 16727 38301
rect 17313 38301 17325 38304
rect 17359 38301 17371 38335
rect 17313 38295 17371 38301
rect 17678 38292 17684 38344
rect 17736 38332 17742 38344
rect 17957 38335 18015 38341
rect 17957 38332 17969 38335
rect 17736 38304 17969 38332
rect 17736 38292 17742 38304
rect 17957 38301 17969 38304
rect 18003 38301 18015 38335
rect 18138 38332 18144 38344
rect 18099 38304 18144 38332
rect 17957 38295 18015 38301
rect 18138 38292 18144 38304
rect 18196 38292 18202 38344
rect 18524 38341 18552 38440
rect 19610 38428 19616 38440
rect 19668 38428 19674 38480
rect 19812 38409 19840 38508
rect 20070 38496 20076 38508
rect 20128 38496 20134 38548
rect 26053 38539 26111 38545
rect 26053 38505 26065 38539
rect 26099 38536 26111 38539
rect 26418 38536 26424 38548
rect 26099 38508 26424 38536
rect 26099 38505 26111 38508
rect 26053 38499 26111 38505
rect 19797 38403 19855 38409
rect 19797 38369 19809 38403
rect 19843 38369 19855 38403
rect 19797 38363 19855 38369
rect 18233 38335 18291 38341
rect 18233 38301 18245 38335
rect 18279 38301 18291 38335
rect 18233 38295 18291 38301
rect 18325 38335 18383 38341
rect 18325 38301 18337 38335
rect 18371 38301 18383 38335
rect 18325 38295 18383 38301
rect 18509 38335 18567 38341
rect 18509 38301 18521 38335
rect 18555 38301 18567 38335
rect 20530 38332 20536 38344
rect 18509 38295 18567 38301
rect 18616 38304 20536 38332
rect 16574 38264 16580 38276
rect 16132 38236 16580 38264
rect 16574 38224 16580 38236
rect 16632 38224 16638 38276
rect 17770 38224 17776 38276
rect 17828 38264 17834 38276
rect 18046 38264 18052 38276
rect 17828 38236 18052 38264
rect 17828 38224 17834 38236
rect 18046 38224 18052 38236
rect 18104 38264 18110 38276
rect 18248 38264 18276 38295
rect 18104 38236 18276 38264
rect 18340 38264 18368 38295
rect 18616 38264 18644 38304
rect 20530 38292 20536 38304
rect 20588 38292 20594 38344
rect 21634 38332 21640 38344
rect 21595 38304 21640 38332
rect 21634 38292 21640 38304
rect 21692 38292 21698 38344
rect 22094 38292 22100 38344
rect 22152 38332 22158 38344
rect 22649 38335 22707 38341
rect 22649 38332 22661 38335
rect 22152 38304 22661 38332
rect 22152 38292 22158 38304
rect 22649 38301 22661 38304
rect 22695 38301 22707 38335
rect 22649 38295 22707 38301
rect 23293 38335 23351 38341
rect 23293 38301 23305 38335
rect 23339 38332 23351 38335
rect 24486 38332 24492 38344
rect 23339 38304 24492 38332
rect 23339 38301 23351 38304
rect 23293 38295 23351 38301
rect 24486 38292 24492 38304
rect 24544 38292 24550 38344
rect 24670 38332 24676 38344
rect 24631 38304 24676 38332
rect 24670 38292 24676 38304
rect 24728 38292 24734 38344
rect 24946 38341 24952 38344
rect 24940 38332 24952 38341
rect 24907 38304 24952 38332
rect 24940 38295 24952 38304
rect 24946 38292 24952 38295
rect 25004 38292 25010 38344
rect 25498 38292 25504 38344
rect 25556 38332 25562 38344
rect 26068 38332 26096 38499
rect 26418 38496 26424 38508
rect 26476 38496 26482 38548
rect 26697 38539 26755 38545
rect 26697 38505 26709 38539
rect 26743 38536 26755 38539
rect 26970 38536 26976 38548
rect 26743 38508 26976 38536
rect 26743 38505 26755 38508
rect 26697 38499 26755 38505
rect 26970 38496 26976 38508
rect 27028 38496 27034 38548
rect 28350 38496 28356 38548
rect 28408 38536 28414 38548
rect 28537 38539 28595 38545
rect 28537 38536 28549 38539
rect 28408 38508 28549 38536
rect 28408 38496 28414 38508
rect 28537 38505 28549 38508
rect 28583 38505 28595 38539
rect 28537 38499 28595 38505
rect 27154 38400 27160 38412
rect 27115 38372 27160 38400
rect 27154 38360 27160 38372
rect 27212 38360 27218 38412
rect 26510 38332 26516 38344
rect 25556 38304 26096 38332
rect 26471 38304 26516 38332
rect 25556 38292 25562 38304
rect 26510 38292 26516 38304
rect 26568 38292 26574 38344
rect 27062 38292 27068 38344
rect 27120 38332 27126 38344
rect 27413 38335 27471 38341
rect 27413 38332 27425 38335
rect 27120 38304 27425 38332
rect 27120 38292 27126 38304
rect 27413 38301 27425 38304
rect 27459 38301 27471 38335
rect 27413 38295 27471 38301
rect 28626 38292 28632 38344
rect 28684 38332 28690 38344
rect 29825 38335 29883 38341
rect 29825 38332 29837 38335
rect 28684 38304 29837 38332
rect 28684 38292 28690 38304
rect 29825 38301 29837 38304
rect 29871 38301 29883 38335
rect 29825 38295 29883 38301
rect 18340 38236 18644 38264
rect 20064 38267 20122 38273
rect 18104 38224 18110 38236
rect 20064 38233 20076 38267
rect 20110 38264 20122 38267
rect 20162 38264 20168 38276
rect 20110 38236 20168 38264
rect 20110 38233 20122 38236
rect 20064 38227 20122 38233
rect 20162 38224 20168 38236
rect 20220 38224 20226 38276
rect 11238 38156 11244 38208
rect 11296 38196 11302 38208
rect 11517 38199 11575 38205
rect 11517 38196 11529 38199
rect 11296 38168 11529 38196
rect 11296 38156 11302 38168
rect 11517 38165 11529 38168
rect 11563 38165 11575 38199
rect 11517 38159 11575 38165
rect 15473 38199 15531 38205
rect 15473 38165 15485 38199
rect 15519 38196 15531 38199
rect 16022 38196 16028 38208
rect 15519 38168 16028 38196
rect 15519 38165 15531 38168
rect 15473 38159 15531 38165
rect 16022 38156 16028 38168
rect 16080 38156 16086 38208
rect 17405 38199 17463 38205
rect 17405 38165 17417 38199
rect 17451 38196 17463 38199
rect 17494 38196 17500 38208
rect 17451 38168 17500 38196
rect 17451 38165 17463 38168
rect 17405 38159 17463 38165
rect 17494 38156 17500 38168
rect 17552 38156 17558 38208
rect 18690 38196 18696 38208
rect 18651 38168 18696 38196
rect 18690 38156 18696 38168
rect 18748 38156 18754 38208
rect 21177 38199 21235 38205
rect 21177 38165 21189 38199
rect 21223 38196 21235 38199
rect 21266 38196 21272 38208
rect 21223 38168 21272 38196
rect 21223 38165 21235 38168
rect 21177 38159 21235 38165
rect 21266 38156 21272 38168
rect 21324 38156 21330 38208
rect 21358 38156 21364 38208
rect 21416 38196 21422 38208
rect 21634 38196 21640 38208
rect 21416 38168 21640 38196
rect 21416 38156 21422 38168
rect 21634 38156 21640 38168
rect 21692 38156 21698 38208
rect 21729 38199 21787 38205
rect 21729 38165 21741 38199
rect 21775 38196 21787 38199
rect 21910 38196 21916 38208
rect 21775 38168 21916 38196
rect 21775 38165 21787 38168
rect 21729 38159 21787 38165
rect 21910 38156 21916 38168
rect 21968 38156 21974 38208
rect 22554 38156 22560 38208
rect 22612 38196 22618 38208
rect 22833 38199 22891 38205
rect 22833 38196 22845 38199
rect 22612 38168 22845 38196
rect 22612 38156 22618 38168
rect 22833 38165 22845 38168
rect 22879 38165 22891 38199
rect 23474 38196 23480 38208
rect 23435 38168 23480 38196
rect 22833 38159 22891 38165
rect 23474 38156 23480 38168
rect 23532 38156 23538 38208
rect 30006 38196 30012 38208
rect 29967 38168 30012 38196
rect 30006 38156 30012 38168
rect 30064 38156 30070 38208
rect 1104 38106 30820 38128
rect 1104 38054 10880 38106
rect 10932 38054 10944 38106
rect 10996 38054 11008 38106
rect 11060 38054 11072 38106
rect 11124 38054 11136 38106
rect 11188 38054 20811 38106
rect 20863 38054 20875 38106
rect 20927 38054 20939 38106
rect 20991 38054 21003 38106
rect 21055 38054 21067 38106
rect 21119 38054 30820 38106
rect 1104 38032 30820 38054
rect 15654 37992 15660 38004
rect 15212 37964 15660 37992
rect 7006 37884 7012 37936
rect 7064 37924 7070 37936
rect 14090 37924 14096 37936
rect 7064 37896 10272 37924
rect 7064 37884 7070 37896
rect 9950 37816 9956 37868
rect 10008 37856 10014 37868
rect 10244 37865 10272 37896
rect 12406 37896 14096 37924
rect 10045 37859 10103 37865
rect 10045 37856 10057 37859
rect 10008 37828 10057 37856
rect 10008 37816 10014 37828
rect 10045 37825 10057 37828
rect 10091 37825 10103 37859
rect 10045 37819 10103 37825
rect 10229 37859 10287 37865
rect 10229 37825 10241 37859
rect 10275 37825 10287 37859
rect 10229 37819 10287 37825
rect 10597 37859 10655 37865
rect 10597 37825 10609 37859
rect 10643 37856 10655 37859
rect 10778 37856 10784 37868
rect 10643 37828 10784 37856
rect 10643 37825 10655 37828
rect 10597 37819 10655 37825
rect 10778 37816 10784 37828
rect 10836 37816 10842 37868
rect 12253 37859 12311 37865
rect 12253 37825 12265 37859
rect 12299 37856 12311 37859
rect 12406 37856 12434 37896
rect 14090 37884 14096 37896
rect 14148 37884 14154 37936
rect 15102 37924 15108 37936
rect 15028 37896 15108 37924
rect 12299 37828 12434 37856
rect 12520 37859 12578 37865
rect 12299 37825 12311 37828
rect 12253 37819 12311 37825
rect 12520 37825 12532 37859
rect 12566 37856 12578 37859
rect 13078 37856 13084 37868
rect 12566 37828 13084 37856
rect 12566 37825 12578 37828
rect 12520 37819 12578 37825
rect 13078 37816 13084 37828
rect 13136 37816 13142 37868
rect 14737 37859 14795 37865
rect 14737 37825 14749 37859
rect 14783 37825 14795 37859
rect 14918 37856 14924 37868
rect 14879 37828 14924 37856
rect 14737 37819 14795 37825
rect 10318 37788 10324 37800
rect 10279 37760 10324 37788
rect 10318 37748 10324 37760
rect 10376 37748 10382 37800
rect 10413 37791 10471 37797
rect 10413 37757 10425 37791
rect 10459 37788 10471 37791
rect 10502 37788 10508 37800
rect 10459 37760 10508 37788
rect 10459 37757 10471 37760
rect 10413 37751 10471 37757
rect 10502 37748 10508 37760
rect 10560 37748 10566 37800
rect 14752 37788 14780 37819
rect 14918 37816 14924 37828
rect 14976 37816 14982 37868
rect 15028 37797 15056 37896
rect 15102 37884 15108 37896
rect 15160 37884 15166 37936
rect 15013 37791 15071 37797
rect 14752 37760 14872 37788
rect 14844 37720 14872 37760
rect 15013 37757 15025 37791
rect 15059 37757 15071 37791
rect 15013 37751 15071 37757
rect 15105 37791 15163 37797
rect 15105 37757 15117 37791
rect 15151 37788 15163 37791
rect 15212 37788 15240 37964
rect 15654 37952 15660 37964
rect 15712 37952 15718 38004
rect 18506 37952 18512 38004
rect 18564 37952 18570 38004
rect 22094 37952 22100 38004
rect 22152 37992 22158 38004
rect 22152 37964 22197 37992
rect 22152 37952 22158 37964
rect 22738 37952 22744 38004
rect 22796 37952 22802 38004
rect 26878 37952 26884 38004
rect 26936 37992 26942 38004
rect 27157 37995 27215 38001
rect 27157 37992 27169 37995
rect 26936 37964 27169 37992
rect 26936 37952 26942 37964
rect 27157 37961 27169 37964
rect 27203 37961 27215 37995
rect 29549 37995 29607 38001
rect 29549 37992 29561 37995
rect 27157 37955 27215 37961
rect 27264 37964 29561 37992
rect 18524 37924 18552 37952
rect 15304 37896 16068 37924
rect 15304 37865 15332 37896
rect 16040 37868 16068 37896
rect 18248 37896 18552 37924
rect 15289 37859 15347 37865
rect 15289 37825 15301 37859
rect 15335 37825 15347 37859
rect 15289 37819 15347 37825
rect 15746 37816 15752 37868
rect 15804 37856 15810 37868
rect 15933 37859 15991 37865
rect 15933 37856 15945 37859
rect 15804 37828 15945 37856
rect 15804 37816 15810 37828
rect 15933 37825 15945 37828
rect 15979 37825 15991 37859
rect 15933 37819 15991 37825
rect 16022 37816 16028 37868
rect 16080 37856 16086 37868
rect 16669 37859 16727 37865
rect 16669 37856 16681 37859
rect 16080 37828 16681 37856
rect 16080 37816 16086 37828
rect 16669 37825 16681 37828
rect 16715 37825 16727 37859
rect 16669 37819 16727 37825
rect 17589 37859 17647 37865
rect 17589 37825 17601 37859
rect 17635 37856 17647 37859
rect 18138 37856 18144 37868
rect 17635 37828 18144 37856
rect 17635 37825 17647 37828
rect 17589 37819 17647 37825
rect 18138 37816 18144 37828
rect 18196 37816 18202 37868
rect 18248 37865 18276 37896
rect 18690 37884 18696 37936
rect 18748 37884 18754 37936
rect 20438 37884 20444 37936
rect 20496 37884 20502 37936
rect 22756 37924 22784 37952
rect 22066 37896 22784 37924
rect 18233 37859 18291 37865
rect 18233 37825 18245 37859
rect 18279 37825 18291 37859
rect 18233 37819 18291 37825
rect 18500 37859 18558 37865
rect 18500 37825 18512 37859
rect 18546 37856 18558 37859
rect 18708 37856 18736 37884
rect 18546 37828 18736 37856
rect 18546 37825 18558 37828
rect 18500 37819 18558 37825
rect 19978 37816 19984 37868
rect 20036 37856 20042 37868
rect 20073 37859 20131 37865
rect 20073 37856 20085 37859
rect 20036 37828 20085 37856
rect 20036 37816 20042 37828
rect 20073 37825 20085 37828
rect 20119 37825 20131 37859
rect 20073 37819 20131 37825
rect 20257 37859 20315 37865
rect 20257 37825 20269 37859
rect 20303 37856 20315 37859
rect 20456 37856 20484 37884
rect 22066 37868 22094 37896
rect 25406 37884 25412 37936
rect 25464 37924 25470 37936
rect 27264 37924 27292 37964
rect 29549 37961 29561 37964
rect 29595 37961 29607 37995
rect 29549 37955 29607 37961
rect 25464 37896 27292 37924
rect 25464 37884 25470 37896
rect 28258 37884 28264 37936
rect 28316 37924 28322 37936
rect 29365 37927 29423 37933
rect 29365 37924 29377 37927
rect 28316 37896 29377 37924
rect 28316 37884 28322 37896
rect 29365 37893 29377 37896
rect 29411 37893 29423 37927
rect 29365 37887 29423 37893
rect 20622 37856 20628 37868
rect 20303 37828 20484 37856
rect 20583 37828 20628 37856
rect 20303 37825 20315 37828
rect 20257 37819 20315 37825
rect 20622 37816 20628 37828
rect 20680 37816 20686 37868
rect 21913 37859 21971 37865
rect 21913 37825 21925 37859
rect 21959 37856 21971 37859
rect 22066 37856 22100 37868
rect 21959 37828 22100 37856
rect 21959 37825 21971 37828
rect 21913 37819 21971 37825
rect 22094 37816 22100 37828
rect 22152 37816 22158 37868
rect 22554 37856 22560 37868
rect 22515 37828 22560 37856
rect 22554 37816 22560 37828
rect 22612 37816 22618 37868
rect 22824 37859 22882 37865
rect 22824 37825 22836 37859
rect 22870 37856 22882 37859
rect 23750 37856 23756 37868
rect 22870 37828 23756 37856
rect 22870 37825 22882 37828
rect 22824 37819 22882 37825
rect 23750 37816 23756 37828
rect 23808 37816 23814 37868
rect 24762 37856 24768 37868
rect 24723 37828 24768 37856
rect 24762 37816 24768 37828
rect 24820 37816 24826 37868
rect 25501 37859 25559 37865
rect 25501 37825 25513 37859
rect 25547 37856 25559 37859
rect 25682 37856 25688 37868
rect 25547 37828 25688 37856
rect 25547 37825 25559 37828
rect 25501 37819 25559 37825
rect 25682 37816 25688 37828
rect 25740 37816 25746 37868
rect 26510 37816 26516 37868
rect 26568 37856 26574 37868
rect 26973 37859 27031 37865
rect 26973 37856 26985 37859
rect 26568 37828 26985 37856
rect 26568 37816 26574 37828
rect 26973 37825 26985 37828
rect 27019 37825 27031 37859
rect 27890 37856 27896 37868
rect 27851 37828 27896 37856
rect 26973 37819 27031 37825
rect 27890 37816 27896 37828
rect 27948 37816 27954 37868
rect 28534 37856 28540 37868
rect 28495 37828 28540 37856
rect 28534 37816 28540 37828
rect 28592 37816 28598 37868
rect 15151 37760 15240 37788
rect 15151 37757 15163 37760
rect 15105 37751 15163 37757
rect 15378 37748 15384 37800
rect 15436 37788 15442 37800
rect 15473 37791 15531 37797
rect 15473 37788 15485 37791
rect 15436 37760 15485 37788
rect 15436 37748 15442 37760
rect 15473 37757 15485 37760
rect 15519 37757 15531 37791
rect 20346 37788 20352 37800
rect 20307 37760 20352 37788
rect 15473 37751 15531 37757
rect 20346 37748 20352 37760
rect 20404 37748 20410 37800
rect 20438 37748 20444 37800
rect 20496 37788 20502 37800
rect 25225 37791 25283 37797
rect 20496 37760 20541 37788
rect 20496 37748 20502 37760
rect 25225 37757 25237 37791
rect 25271 37757 25283 37791
rect 28997 37791 29055 37797
rect 28997 37788 29009 37791
rect 25225 37751 25283 37757
rect 27632 37760 29009 37788
rect 16574 37720 16580 37732
rect 14844 37692 16580 37720
rect 16574 37680 16580 37692
rect 16632 37720 16638 37732
rect 17126 37720 17132 37732
rect 16632 37692 17132 37720
rect 16632 37680 16638 37692
rect 17126 37680 17132 37692
rect 17184 37680 17190 37732
rect 25240 37720 25268 37751
rect 23492 37692 25268 37720
rect 10686 37612 10692 37664
rect 10744 37652 10750 37664
rect 10781 37655 10839 37661
rect 10781 37652 10793 37655
rect 10744 37624 10793 37652
rect 10744 37612 10750 37624
rect 10781 37621 10793 37624
rect 10827 37621 10839 37655
rect 13630 37652 13636 37664
rect 13591 37624 13636 37652
rect 10781 37615 10839 37621
rect 13630 37612 13636 37624
rect 13688 37612 13694 37664
rect 16025 37655 16083 37661
rect 16025 37621 16037 37655
rect 16071 37652 16083 37655
rect 16482 37652 16488 37664
rect 16071 37624 16488 37652
rect 16071 37621 16083 37624
rect 16025 37615 16083 37621
rect 16482 37612 16488 37624
rect 16540 37612 16546 37664
rect 16761 37655 16819 37661
rect 16761 37621 16773 37655
rect 16807 37652 16819 37655
rect 16942 37652 16948 37664
rect 16807 37624 16948 37652
rect 16807 37621 16819 37624
rect 16761 37615 16819 37621
rect 16942 37612 16948 37624
rect 17000 37612 17006 37664
rect 17681 37655 17739 37661
rect 17681 37621 17693 37655
rect 17727 37652 17739 37655
rect 18414 37652 18420 37664
rect 17727 37624 18420 37652
rect 17727 37621 17739 37624
rect 17681 37615 17739 37621
rect 18414 37612 18420 37624
rect 18472 37612 18478 37664
rect 19610 37652 19616 37664
rect 19523 37624 19616 37652
rect 19610 37612 19616 37624
rect 19668 37652 19674 37664
rect 20530 37652 20536 37664
rect 19668 37624 20536 37652
rect 19668 37612 19674 37624
rect 20530 37612 20536 37624
rect 20588 37612 20594 37664
rect 20809 37655 20867 37661
rect 20809 37621 20821 37655
rect 20855 37652 20867 37655
rect 21174 37652 21180 37664
rect 20855 37624 21180 37652
rect 20855 37621 20867 37624
rect 20809 37615 20867 37621
rect 21174 37612 21180 37624
rect 21232 37612 21238 37664
rect 22922 37612 22928 37664
rect 22980 37652 22986 37664
rect 23492 37652 23520 37692
rect 23934 37652 23940 37664
rect 22980 37624 23520 37652
rect 23895 37624 23940 37652
rect 22980 37612 22986 37624
rect 23934 37612 23940 37624
rect 23992 37612 23998 37664
rect 24581 37655 24639 37661
rect 24581 37621 24593 37655
rect 24627 37652 24639 37655
rect 27632 37652 27660 37760
rect 28997 37757 29009 37760
rect 29043 37788 29055 37791
rect 29086 37788 29092 37800
rect 29043 37760 29092 37788
rect 29043 37757 29055 37760
rect 28997 37751 29055 37757
rect 29086 37748 29092 37760
rect 29144 37748 29150 37800
rect 27709 37723 27767 37729
rect 27709 37689 27721 37723
rect 27755 37720 27767 37723
rect 27755 37692 28948 37720
rect 27755 37689 27767 37692
rect 27709 37683 27767 37689
rect 24627 37624 27660 37652
rect 28353 37655 28411 37661
rect 24627 37621 24639 37624
rect 24581 37615 24639 37621
rect 28353 37621 28365 37655
rect 28399 37652 28411 37655
rect 28718 37652 28724 37664
rect 28399 37624 28724 37652
rect 28399 37621 28411 37624
rect 28353 37615 28411 37621
rect 28718 37612 28724 37624
rect 28776 37612 28782 37664
rect 28920 37652 28948 37692
rect 29270 37652 29276 37664
rect 28920 37624 29276 37652
rect 29270 37612 29276 37624
rect 29328 37612 29334 37664
rect 29362 37612 29368 37664
rect 29420 37652 29426 37664
rect 29420 37624 29465 37652
rect 29420 37612 29426 37624
rect 1104 37562 30820 37584
rect 1104 37510 5915 37562
rect 5967 37510 5979 37562
rect 6031 37510 6043 37562
rect 6095 37510 6107 37562
rect 6159 37510 6171 37562
rect 6223 37510 15846 37562
rect 15898 37510 15910 37562
rect 15962 37510 15974 37562
rect 16026 37510 16038 37562
rect 16090 37510 16102 37562
rect 16154 37510 25776 37562
rect 25828 37510 25840 37562
rect 25892 37510 25904 37562
rect 25956 37510 25968 37562
rect 26020 37510 26032 37562
rect 26084 37510 30820 37562
rect 1104 37488 30820 37510
rect 13078 37408 13084 37460
rect 13136 37448 13142 37460
rect 13173 37451 13231 37457
rect 13173 37448 13185 37451
rect 13136 37420 13185 37448
rect 13136 37408 13142 37420
rect 13173 37417 13185 37420
rect 13219 37417 13231 37451
rect 13173 37411 13231 37417
rect 15102 37408 15108 37460
rect 15160 37448 15166 37460
rect 21266 37448 21272 37460
rect 15160 37420 21272 37448
rect 15160 37408 15166 37420
rect 21266 37408 21272 37420
rect 21324 37408 21330 37460
rect 23750 37448 23756 37460
rect 23711 37420 23756 37448
rect 23750 37408 23756 37420
rect 23808 37408 23814 37460
rect 24486 37408 24492 37460
rect 24544 37448 24550 37460
rect 24581 37451 24639 37457
rect 24581 37448 24593 37451
rect 24544 37420 24593 37448
rect 24544 37408 24550 37420
rect 24581 37417 24593 37420
rect 24627 37417 24639 37451
rect 28258 37448 28264 37460
rect 24581 37411 24639 37417
rect 27632 37420 28264 37448
rect 12618 37340 12624 37392
rect 12676 37340 12682 37392
rect 16669 37383 16727 37389
rect 16669 37380 16681 37383
rect 15028 37352 16681 37380
rect 1578 37244 1584 37256
rect 1539 37216 1584 37244
rect 1578 37204 1584 37216
rect 1636 37204 1642 37256
rect 10134 37204 10140 37256
rect 10192 37244 10198 37256
rect 10410 37244 10416 37256
rect 10192 37216 10416 37244
rect 10192 37204 10198 37216
rect 10410 37204 10416 37216
rect 10468 37204 10474 37256
rect 10686 37253 10692 37256
rect 10680 37244 10692 37253
rect 10647 37216 10692 37244
rect 10680 37207 10692 37216
rect 10686 37204 10692 37207
rect 10744 37204 10750 37256
rect 12636 37253 12664 37340
rect 12805 37315 12863 37321
rect 12805 37281 12817 37315
rect 12851 37312 12863 37315
rect 13262 37312 13268 37324
rect 12851 37284 13268 37312
rect 12851 37281 12863 37284
rect 12805 37275 12863 37281
rect 13262 37272 13268 37284
rect 13320 37272 13326 37324
rect 15028 37256 15056 37352
rect 16669 37349 16681 37352
rect 16715 37349 16727 37383
rect 16669 37343 16727 37349
rect 18417 37383 18475 37389
rect 18417 37349 18429 37383
rect 18463 37380 18475 37383
rect 18782 37380 18788 37392
rect 18463 37352 18788 37380
rect 18463 37349 18475 37352
rect 18417 37343 18475 37349
rect 18782 37340 18788 37352
rect 18840 37340 18846 37392
rect 23198 37340 23204 37392
rect 23256 37340 23262 37392
rect 27632 37380 27660 37420
rect 28258 37408 28264 37420
rect 28316 37408 28322 37460
rect 28813 37451 28871 37457
rect 28813 37417 28825 37451
rect 28859 37448 28871 37451
rect 29362 37448 29368 37460
rect 28859 37420 29368 37448
rect 28859 37417 28871 37420
rect 28813 37411 28871 37417
rect 29362 37408 29368 37420
rect 29420 37448 29426 37460
rect 29917 37451 29975 37457
rect 29917 37448 29929 37451
rect 29420 37420 29929 37448
rect 29420 37408 29426 37420
rect 29917 37417 29929 37420
rect 29963 37417 29975 37451
rect 29917 37411 29975 37417
rect 27080 37352 27660 37380
rect 15194 37312 15200 37324
rect 15155 37284 15200 37312
rect 15194 37272 15200 37284
rect 15252 37272 15258 37324
rect 15654 37312 15660 37324
rect 15615 37284 15660 37312
rect 15654 37272 15660 37284
rect 15712 37272 15718 37324
rect 19521 37315 19579 37321
rect 19521 37281 19533 37315
rect 19567 37312 19579 37315
rect 19978 37312 19984 37324
rect 19567 37284 19984 37312
rect 19567 37281 19579 37284
rect 19521 37275 19579 37281
rect 19978 37272 19984 37284
rect 20036 37272 20042 37324
rect 20070 37272 20076 37324
rect 20128 37312 20134 37324
rect 20625 37315 20683 37321
rect 20625 37312 20637 37315
rect 20128 37284 20637 37312
rect 20128 37272 20134 37284
rect 20625 37281 20637 37284
rect 20671 37281 20683 37315
rect 20625 37275 20683 37281
rect 23204 37274 23232 37340
rect 12437 37247 12495 37253
rect 12437 37213 12449 37247
rect 12483 37244 12495 37247
rect 12621 37247 12679 37253
rect 12483 37216 12517 37244
rect 12483 37213 12495 37216
rect 12437 37207 12495 37213
rect 12621 37213 12633 37247
rect 12667 37213 12679 37247
rect 12621 37207 12679 37213
rect 12713 37247 12771 37253
rect 12713 37213 12725 37247
rect 12759 37213 12771 37247
rect 12713 37207 12771 37213
rect 9950 37136 9956 37188
rect 10008 37176 10014 37188
rect 12452 37176 12480 37207
rect 12526 37176 12532 37188
rect 10008 37148 12532 37176
rect 10008 37136 10014 37148
rect 12526 37136 12532 37148
rect 12584 37136 12590 37188
rect 1397 37111 1455 37117
rect 1397 37077 1409 37111
rect 1443 37108 1455 37111
rect 10686 37108 10692 37120
rect 1443 37080 10692 37108
rect 1443 37077 1455 37080
rect 1397 37071 1455 37077
rect 10686 37068 10692 37080
rect 10744 37068 10750 37120
rect 10778 37068 10784 37120
rect 10836 37108 10842 37120
rect 11793 37111 11851 37117
rect 11793 37108 11805 37111
rect 10836 37080 11805 37108
rect 10836 37068 10842 37080
rect 11793 37077 11805 37080
rect 11839 37077 11851 37111
rect 11793 37071 11851 37077
rect 12158 37068 12164 37120
rect 12216 37108 12222 37120
rect 12728 37108 12756 37207
rect 12894 37204 12900 37256
rect 12952 37244 12958 37256
rect 12989 37247 13047 37253
rect 12989 37244 13001 37247
rect 12952 37216 13001 37244
rect 12952 37204 12958 37216
rect 12989 37213 13001 37216
rect 13035 37244 13047 37247
rect 13630 37244 13636 37256
rect 13035 37216 13636 37244
rect 13035 37213 13047 37216
rect 12989 37207 13047 37213
rect 13630 37204 13636 37216
rect 13688 37204 13694 37256
rect 14921 37247 14979 37253
rect 14921 37213 14933 37247
rect 14967 37244 14979 37247
rect 15010 37244 15016 37256
rect 14967 37216 15016 37244
rect 14967 37213 14979 37216
rect 14921 37207 14979 37213
rect 15010 37204 15016 37216
rect 15068 37204 15074 37256
rect 15105 37247 15163 37253
rect 15105 37213 15117 37247
rect 15151 37213 15163 37247
rect 15105 37207 15163 37213
rect 15289 37247 15347 37253
rect 15289 37213 15301 37247
rect 15335 37244 15347 37247
rect 15378 37244 15384 37256
rect 15335 37216 15384 37244
rect 15335 37213 15347 37216
rect 15289 37207 15347 37213
rect 14734 37136 14740 37188
rect 14792 37176 14798 37188
rect 15120 37176 15148 37207
rect 15378 37204 15384 37216
rect 15436 37204 15442 37256
rect 15473 37247 15531 37253
rect 15473 37213 15485 37247
rect 15519 37213 15531 37247
rect 15473 37207 15531 37213
rect 16485 37247 16543 37253
rect 16485 37213 16497 37247
rect 16531 37244 16543 37247
rect 16574 37244 16580 37256
rect 16531 37216 16580 37244
rect 16531 37213 16543 37216
rect 16485 37207 16543 37213
rect 14792 37148 15148 37176
rect 15488 37176 15516 37207
rect 16574 37204 16580 37216
rect 16632 37204 16638 37256
rect 17129 37247 17187 37253
rect 17129 37213 17141 37247
rect 17175 37244 17187 37247
rect 17175 37216 19196 37244
rect 17175 37213 17187 37216
rect 17129 37207 17187 37213
rect 16758 37176 16764 37188
rect 15488 37148 16764 37176
rect 14792 37136 14798 37148
rect 16758 37136 16764 37148
rect 16816 37136 16822 37188
rect 18233 37179 18291 37185
rect 18233 37145 18245 37179
rect 18279 37176 18291 37179
rect 18690 37176 18696 37188
rect 18279 37148 18696 37176
rect 18279 37145 18291 37148
rect 18233 37139 18291 37145
rect 18690 37136 18696 37148
rect 18748 37136 18754 37188
rect 19168 37176 19196 37216
rect 19242 37204 19248 37256
rect 19300 37244 19306 37256
rect 22186 37244 22192 37256
rect 19300 37216 22192 37244
rect 19300 37204 19306 37216
rect 22186 37204 22192 37216
rect 22244 37244 22250 37256
rect 22922 37244 22928 37256
rect 22244 37216 22928 37244
rect 22244 37204 22250 37216
rect 22922 37204 22928 37216
rect 22980 37204 22986 37256
rect 23014 37204 23020 37256
rect 23072 37244 23078 37256
rect 23204 37253 23244 37274
rect 23290 37272 23296 37324
rect 23348 37312 23354 37324
rect 23934 37312 23940 37324
rect 23348 37284 23393 37312
rect 23584 37284 23940 37312
rect 23348 37272 23354 37284
rect 23189 37247 23247 37253
rect 23072 37216 23117 37244
rect 23072 37204 23078 37216
rect 23189 37213 23201 37247
rect 23235 37213 23247 37247
rect 23189 37207 23247 37213
rect 23382 37204 23388 37256
rect 23440 37244 23446 37256
rect 23584 37253 23612 37284
rect 23934 37272 23940 37284
rect 23992 37312 23998 37324
rect 26142 37312 26148 37324
rect 23992 37284 24532 37312
rect 23992 37272 23998 37284
rect 24504 37256 24532 37284
rect 25608 37284 26148 37312
rect 23569 37247 23627 37253
rect 23440 37216 23485 37244
rect 23440 37204 23446 37216
rect 23569 37213 23581 37247
rect 23615 37244 23627 37247
rect 24397 37247 24455 37253
rect 23615 37216 23649 37244
rect 23615 37213 23627 37216
rect 23569 37207 23627 37213
rect 24397 37213 24409 37247
rect 24443 37213 24455 37247
rect 24397 37207 24455 37213
rect 20622 37176 20628 37188
rect 19168 37148 20628 37176
rect 20622 37136 20628 37148
rect 20680 37136 20686 37188
rect 20898 37185 20904 37188
rect 20892 37176 20904 37185
rect 20859 37148 20904 37176
rect 20892 37139 20904 37148
rect 20898 37136 20904 37139
rect 20956 37136 20962 37188
rect 22094 37136 22100 37188
rect 22152 37176 22158 37188
rect 24412 37176 24440 37207
rect 24486 37204 24492 37256
rect 24544 37204 24550 37256
rect 24946 37204 24952 37256
rect 25004 37244 25010 37256
rect 25608 37253 25636 37284
rect 26142 37272 26148 37284
rect 26200 37312 26206 37324
rect 26973 37315 27031 37321
rect 26200 37284 26924 37312
rect 26200 37272 26206 37284
rect 25317 37247 25375 37253
rect 25317 37244 25329 37247
rect 25004 37216 25329 37244
rect 25004 37204 25010 37216
rect 25317 37213 25329 37216
rect 25363 37213 25375 37247
rect 25317 37207 25375 37213
rect 25593 37247 25651 37253
rect 25593 37213 25605 37247
rect 25639 37244 25651 37247
rect 25639 37216 25673 37244
rect 25639 37213 25651 37216
rect 25593 37207 25651 37213
rect 25774 37204 25780 37256
rect 25832 37244 25838 37256
rect 26605 37247 26663 37253
rect 26605 37244 26617 37247
rect 25832 37216 26617 37244
rect 25832 37204 25838 37216
rect 26605 37213 26617 37216
rect 26651 37213 26663 37247
rect 26605 37207 26663 37213
rect 26694 37204 26700 37256
rect 26752 37244 26758 37256
rect 26896 37253 26924 37284
rect 26973 37281 26985 37315
rect 27019 37281 27031 37315
rect 26973 37275 27031 37281
rect 26789 37247 26847 37253
rect 26789 37244 26801 37247
rect 26752 37216 26801 37244
rect 26752 37204 26758 37216
rect 26789 37213 26801 37216
rect 26835 37213 26847 37247
rect 26789 37207 26847 37213
rect 26875 37247 26933 37253
rect 26875 37213 26887 37247
rect 26921 37213 26933 37247
rect 26875 37207 26933 37213
rect 26988 37176 27016 37275
rect 27080 37260 27108 37352
rect 27982 37340 27988 37392
rect 28040 37380 28046 37392
rect 28997 37383 29055 37389
rect 28997 37380 29009 37383
rect 28040 37352 29009 37380
rect 28040 37340 28046 37352
rect 28997 37349 29009 37352
rect 29043 37349 29055 37383
rect 28997 37343 29055 37349
rect 28445 37315 28503 37321
rect 27632 37284 27936 37312
rect 27080 37253 27183 37260
rect 27080 37247 27215 37253
rect 27080 37232 27169 37247
rect 27155 37216 27169 37232
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 27157 37207 27215 37213
rect 27338 37204 27344 37256
rect 27396 37244 27402 37256
rect 27632 37244 27660 37284
rect 27798 37244 27804 37256
rect 27396 37216 27660 37244
rect 27759 37216 27804 37244
rect 27396 37204 27402 37216
rect 27798 37204 27804 37216
rect 27856 37204 27862 37256
rect 27908 37244 27936 37284
rect 28445 37281 28457 37315
rect 28491 37312 28503 37315
rect 29086 37312 29092 37324
rect 28491 37284 29092 37312
rect 28491 37281 28503 37284
rect 28445 37275 28503 37281
rect 29086 37272 29092 37284
rect 29144 37312 29150 37324
rect 29549 37315 29607 37321
rect 29549 37312 29561 37315
rect 29144 37284 29561 37312
rect 29144 37272 29150 37284
rect 29549 37281 29561 37284
rect 29595 37281 29607 37315
rect 29549 37275 29607 37281
rect 27908 37216 29960 37244
rect 29932 37185 29960 37216
rect 22152 37148 24440 37176
rect 25792 37148 27016 37176
rect 29917 37179 29975 37185
rect 22152 37136 22158 37148
rect 25792 37120 25820 37148
rect 29917 37145 29929 37179
rect 29963 37145 29975 37179
rect 29917 37139 29975 37145
rect 12216 37080 12756 37108
rect 12216 37068 12222 37080
rect 17034 37068 17040 37120
rect 17092 37108 17098 37120
rect 17221 37111 17279 37117
rect 17221 37108 17233 37111
rect 17092 37080 17233 37108
rect 17092 37068 17098 37080
rect 17221 37077 17233 37080
rect 17267 37077 17279 37111
rect 17221 37071 17279 37077
rect 21358 37068 21364 37120
rect 21416 37108 21422 37120
rect 22005 37111 22063 37117
rect 22005 37108 22017 37111
rect 21416 37080 22017 37108
rect 21416 37068 21422 37080
rect 22005 37077 22017 37080
rect 22051 37077 22063 37111
rect 22005 37071 22063 37077
rect 22922 37068 22928 37120
rect 22980 37108 22986 37120
rect 23290 37108 23296 37120
rect 22980 37080 23296 37108
rect 22980 37068 22986 37080
rect 23290 37068 23296 37080
rect 23348 37068 23354 37120
rect 25774 37068 25780 37120
rect 25832 37068 25838 37120
rect 27338 37108 27344 37120
rect 27299 37080 27344 37108
rect 27338 37068 27344 37080
rect 27396 37068 27402 37120
rect 27982 37108 27988 37120
rect 27943 37080 27988 37108
rect 27982 37068 27988 37080
rect 28040 37068 28046 37120
rect 28810 37108 28816 37120
rect 28771 37080 28816 37108
rect 28810 37068 28816 37080
rect 28868 37068 28874 37120
rect 28902 37068 28908 37120
rect 28960 37108 28966 37120
rect 30101 37111 30159 37117
rect 30101 37108 30113 37111
rect 28960 37080 30113 37108
rect 28960 37068 28966 37080
rect 30101 37077 30113 37080
rect 30147 37077 30159 37111
rect 30101 37071 30159 37077
rect 1104 37018 30820 37040
rect 1104 36966 10880 37018
rect 10932 36966 10944 37018
rect 10996 36966 11008 37018
rect 11060 36966 11072 37018
rect 11124 36966 11136 37018
rect 11188 36966 20811 37018
rect 20863 36966 20875 37018
rect 20927 36966 20939 37018
rect 20991 36966 21003 37018
rect 21055 36966 21067 37018
rect 21119 36966 30820 37018
rect 1104 36944 30820 36966
rect 10594 36904 10600 36916
rect 10555 36876 10600 36904
rect 10594 36864 10600 36876
rect 10652 36864 10658 36916
rect 10686 36864 10692 36916
rect 10744 36904 10750 36916
rect 12066 36904 12072 36916
rect 10744 36876 12072 36904
rect 10744 36864 10750 36876
rect 12066 36864 12072 36876
rect 12124 36864 12130 36916
rect 19426 36904 19432 36916
rect 14936 36876 19432 36904
rect 9950 36836 9956 36848
rect 8680 36808 9956 36836
rect 8680 36777 8708 36808
rect 8665 36771 8723 36777
rect 8665 36737 8677 36771
rect 8711 36737 8723 36771
rect 8846 36768 8852 36780
rect 8807 36740 8852 36768
rect 8665 36731 8723 36737
rect 8846 36728 8852 36740
rect 8904 36728 8910 36780
rect 8941 36771 8999 36777
rect 8941 36737 8953 36771
rect 8987 36768 8999 36771
rect 9217 36771 9275 36777
rect 8987 36740 9168 36768
rect 8987 36737 8999 36740
rect 8941 36731 8999 36737
rect 9033 36703 9091 36709
rect 9033 36669 9045 36703
rect 9079 36669 9091 36703
rect 9140 36700 9168 36740
rect 9217 36737 9229 36771
rect 9263 36768 9275 36771
rect 9674 36768 9680 36780
rect 9263 36740 9680 36768
rect 9263 36737 9275 36740
rect 9217 36731 9275 36737
rect 9674 36728 9680 36740
rect 9732 36728 9738 36780
rect 9876 36777 9904 36808
rect 9950 36796 9956 36808
rect 10008 36796 10014 36848
rect 14936 36836 14964 36876
rect 19426 36864 19432 36876
rect 19484 36864 19490 36916
rect 23290 36904 23296 36916
rect 23124 36876 23296 36904
rect 19242 36836 19248 36848
rect 13648 36808 14964 36836
rect 9861 36771 9919 36777
rect 9861 36737 9873 36771
rect 9907 36737 9919 36771
rect 10042 36768 10048 36780
rect 10003 36740 10048 36768
rect 9861 36731 9919 36737
rect 10042 36728 10048 36740
rect 10100 36728 10106 36780
rect 10318 36768 10324 36780
rect 10152 36740 10324 36768
rect 10152 36709 10180 36740
rect 10318 36728 10324 36740
rect 10376 36728 10382 36780
rect 10413 36771 10471 36777
rect 10413 36737 10425 36771
rect 10459 36768 10471 36771
rect 11238 36768 11244 36780
rect 10459 36740 11244 36768
rect 10459 36737 10471 36740
rect 10413 36731 10471 36737
rect 11238 36728 11244 36740
rect 11296 36728 11302 36780
rect 11701 36771 11759 36777
rect 11701 36737 11713 36771
rect 11747 36768 11759 36771
rect 13170 36768 13176 36780
rect 11747 36740 13176 36768
rect 11747 36737 11759 36740
rect 11701 36731 11759 36737
rect 13170 36728 13176 36740
rect 13228 36728 13234 36780
rect 13648 36777 13676 36808
rect 14936 36777 14964 36808
rect 16960 36808 19248 36836
rect 13633 36771 13691 36777
rect 13633 36737 13645 36771
rect 13679 36737 13691 36771
rect 14921 36771 14979 36777
rect 13633 36731 13691 36737
rect 13832 36740 14872 36768
rect 10137 36703 10195 36709
rect 10137 36700 10149 36703
rect 9140 36672 10149 36700
rect 9033 36663 9091 36669
rect 10137 36669 10149 36672
rect 10183 36669 10195 36703
rect 10137 36663 10195 36669
rect 10229 36703 10287 36709
rect 10229 36669 10241 36703
rect 10275 36669 10287 36703
rect 10336 36700 10364 36728
rect 12158 36700 12164 36712
rect 10336 36672 12164 36700
rect 10229 36663 10287 36669
rect 9048 36632 9076 36663
rect 10244 36632 10272 36663
rect 12158 36660 12164 36672
rect 12216 36700 12222 36712
rect 12345 36703 12403 36709
rect 12216 36672 12296 36700
rect 12216 36660 12222 36672
rect 9048 36604 10364 36632
rect 9306 36524 9312 36576
rect 9364 36564 9370 36576
rect 9401 36567 9459 36573
rect 9401 36564 9413 36567
rect 9364 36536 9413 36564
rect 9364 36524 9370 36536
rect 9401 36533 9413 36536
rect 9447 36533 9459 36567
rect 10336 36564 10364 36604
rect 10410 36592 10416 36644
rect 10468 36632 10474 36644
rect 10468 36604 11836 36632
rect 10468 36592 10474 36604
rect 11808 36576 11836 36604
rect 10502 36564 10508 36576
rect 10336 36536 10508 36564
rect 9401 36527 9459 36533
rect 10502 36524 10508 36536
rect 10560 36524 10566 36576
rect 11790 36564 11796 36576
rect 11751 36536 11796 36564
rect 11790 36524 11796 36536
rect 11848 36524 11854 36576
rect 12268 36564 12296 36672
rect 12345 36669 12357 36703
rect 12391 36669 12403 36703
rect 12618 36700 12624 36712
rect 12579 36672 12624 36700
rect 12345 36663 12403 36669
rect 12360 36632 12388 36663
rect 12618 36660 12624 36672
rect 12676 36660 12682 36712
rect 13832 36632 13860 36740
rect 13909 36703 13967 36709
rect 13909 36669 13921 36703
rect 13955 36669 13967 36703
rect 14844 36700 14872 36740
rect 14921 36737 14933 36771
rect 14967 36737 14979 36771
rect 15194 36768 15200 36780
rect 15155 36740 15200 36768
rect 14921 36731 14979 36737
rect 15194 36728 15200 36740
rect 15252 36768 15258 36780
rect 15378 36768 15384 36780
rect 15252 36740 15384 36768
rect 15252 36728 15258 36740
rect 15378 36728 15384 36740
rect 15436 36728 15442 36780
rect 16960 36700 16988 36808
rect 17037 36771 17095 36777
rect 17037 36737 17049 36771
rect 17083 36737 17095 36771
rect 17218 36768 17224 36780
rect 17179 36740 17224 36768
rect 17037 36731 17095 36737
rect 14844 36672 16988 36700
rect 17052 36700 17080 36731
rect 17218 36728 17224 36740
rect 17276 36728 17282 36780
rect 17313 36771 17371 36777
rect 17313 36737 17325 36771
rect 17359 36768 17371 36771
rect 17589 36771 17647 36777
rect 17359 36740 17540 36768
rect 17359 36737 17371 36740
rect 17313 36731 17371 36737
rect 17405 36703 17463 36709
rect 17052 36672 17264 36700
rect 13909 36663 13967 36669
rect 12360 36604 13860 36632
rect 13924 36564 13952 36663
rect 17236 36644 17264 36672
rect 17405 36669 17417 36703
rect 17451 36669 17463 36703
rect 17512 36700 17540 36740
rect 17589 36737 17601 36771
rect 17635 36768 17647 36771
rect 17678 36768 17684 36780
rect 17635 36740 17684 36768
rect 17635 36737 17647 36740
rect 17589 36731 17647 36737
rect 17678 36728 17684 36740
rect 17736 36728 17742 36780
rect 18800 36777 18828 36808
rect 19242 36796 19248 36808
rect 19300 36796 19306 36848
rect 18785 36771 18843 36777
rect 18785 36737 18797 36771
rect 18831 36737 18843 36771
rect 20349 36771 20407 36777
rect 20349 36768 20361 36771
rect 18785 36731 18843 36737
rect 18984 36740 20361 36768
rect 18046 36700 18052 36712
rect 17512 36672 18052 36700
rect 17405 36663 17463 36669
rect 17218 36592 17224 36644
rect 17276 36592 17282 36644
rect 17420 36632 17448 36663
rect 18046 36660 18052 36672
rect 18104 36700 18110 36712
rect 18984 36700 19012 36740
rect 20349 36737 20361 36740
rect 20395 36737 20407 36771
rect 20349 36731 20407 36737
rect 22005 36771 22063 36777
rect 22005 36737 22017 36771
rect 22051 36768 22063 36771
rect 22094 36768 22100 36780
rect 22051 36740 22100 36768
rect 22051 36737 22063 36740
rect 22005 36731 22063 36737
rect 22094 36728 22100 36740
rect 22152 36728 22158 36780
rect 22646 36768 22652 36780
rect 22607 36740 22652 36768
rect 22646 36728 22652 36740
rect 22704 36728 22710 36780
rect 22833 36771 22891 36777
rect 22833 36737 22845 36771
rect 22879 36737 22891 36771
rect 22833 36731 22891 36737
rect 18104 36672 19012 36700
rect 19061 36703 19119 36709
rect 18104 36660 18110 36672
rect 19061 36669 19073 36703
rect 19107 36669 19119 36703
rect 19061 36663 19119 36669
rect 18782 36632 18788 36644
rect 17420 36604 18788 36632
rect 18782 36592 18788 36604
rect 18840 36592 18846 36644
rect 19076 36632 19104 36663
rect 19426 36660 19432 36712
rect 19484 36700 19490 36712
rect 20073 36703 20131 36709
rect 20073 36700 20085 36703
rect 19484 36672 20085 36700
rect 19484 36660 19490 36672
rect 20073 36669 20085 36672
rect 20119 36669 20131 36703
rect 20073 36663 20131 36669
rect 22370 36660 22376 36712
rect 22428 36700 22434 36712
rect 22848 36700 22876 36731
rect 22922 36728 22928 36780
rect 22980 36768 22986 36780
rect 22980 36740 23025 36768
rect 22980 36728 22986 36740
rect 22428 36672 22876 36700
rect 23017 36703 23075 36709
rect 22428 36660 22434 36672
rect 23017 36669 23029 36703
rect 23063 36700 23075 36703
rect 23124 36700 23152 36876
rect 23290 36864 23296 36876
rect 23348 36904 23354 36916
rect 24486 36904 24492 36916
rect 23348 36876 24492 36904
rect 23348 36864 23354 36876
rect 24486 36864 24492 36876
rect 24544 36864 24550 36916
rect 28353 36907 28411 36913
rect 28353 36904 28365 36907
rect 26252 36876 28365 36904
rect 23385 36839 23443 36845
rect 23385 36805 23397 36839
rect 23431 36836 23443 36839
rect 24090 36839 24148 36845
rect 24090 36836 24102 36839
rect 23431 36808 24102 36836
rect 23431 36805 23443 36808
rect 23385 36799 23443 36805
rect 24090 36805 24102 36808
rect 24136 36805 24148 36839
rect 24090 36799 24148 36805
rect 24854 36796 24860 36848
rect 24912 36836 24918 36848
rect 26050 36836 26056 36848
rect 24912 36808 26056 36836
rect 24912 36796 24918 36808
rect 23201 36771 23259 36777
rect 23201 36737 23213 36771
rect 23247 36737 23259 36771
rect 23201 36731 23259 36737
rect 23063 36672 23152 36700
rect 23063 36669 23075 36672
rect 23017 36663 23075 36669
rect 19518 36632 19524 36644
rect 19076 36604 19524 36632
rect 19518 36592 19524 36604
rect 19576 36592 19582 36644
rect 12268 36536 13952 36564
rect 17126 36524 17132 36576
rect 17184 36564 17190 36576
rect 17773 36567 17831 36573
rect 17773 36564 17785 36567
rect 17184 36536 17785 36564
rect 17184 36524 17190 36536
rect 17773 36533 17785 36536
rect 17819 36533 17831 36567
rect 17773 36527 17831 36533
rect 22189 36567 22247 36573
rect 22189 36533 22201 36567
rect 22235 36564 22247 36567
rect 22738 36564 22744 36576
rect 22235 36536 22744 36564
rect 22235 36533 22247 36536
rect 22189 36527 22247 36533
rect 22738 36524 22744 36536
rect 22796 36524 22802 36576
rect 23216 36564 23244 36731
rect 23474 36728 23480 36780
rect 23532 36768 23538 36780
rect 23845 36771 23903 36777
rect 23845 36768 23857 36771
rect 23532 36740 23857 36768
rect 23532 36728 23538 36740
rect 23845 36737 23857 36740
rect 23891 36737 23903 36771
rect 25682 36768 25688 36780
rect 25643 36740 25688 36768
rect 23845 36731 23903 36737
rect 25682 36728 25688 36740
rect 25740 36728 25746 36780
rect 25884 36777 25912 36808
rect 26050 36796 26056 36808
rect 26108 36796 26114 36848
rect 25869 36771 25927 36777
rect 25869 36737 25881 36771
rect 25915 36737 25927 36771
rect 25869 36731 25927 36737
rect 25961 36771 26019 36777
rect 25961 36737 25973 36771
rect 26007 36768 26019 36771
rect 26142 36768 26148 36780
rect 26007 36740 26148 36768
rect 26007 36737 26019 36740
rect 25961 36731 26019 36737
rect 26142 36728 26148 36740
rect 26200 36728 26206 36780
rect 26252 36777 26280 36876
rect 28353 36873 28365 36876
rect 28399 36904 28411 36907
rect 28810 36904 28816 36916
rect 28399 36876 28816 36904
rect 28399 36873 28411 36876
rect 28353 36867 28411 36873
rect 28810 36864 28816 36876
rect 28868 36864 28874 36916
rect 29641 36907 29699 36913
rect 29641 36904 29653 36907
rect 29012 36876 29653 36904
rect 26421 36839 26479 36845
rect 26421 36805 26433 36839
rect 26467 36836 26479 36839
rect 27218 36839 27276 36845
rect 27218 36836 27230 36839
rect 26467 36808 27230 36836
rect 26467 36805 26479 36808
rect 26421 36799 26479 36805
rect 27218 36805 27230 36808
rect 27264 36805 27276 36839
rect 27218 36799 27276 36805
rect 28442 36796 28448 36848
rect 28500 36836 28506 36848
rect 29012 36836 29040 36876
rect 29641 36873 29653 36876
rect 29687 36873 29699 36907
rect 29641 36867 29699 36873
rect 28500 36808 29040 36836
rect 29457 36839 29515 36845
rect 28500 36796 28506 36808
rect 29457 36805 29469 36839
rect 29503 36805 29515 36839
rect 29457 36799 29515 36805
rect 26237 36771 26295 36777
rect 26237 36737 26249 36771
rect 26283 36737 26295 36771
rect 29472 36768 29500 36799
rect 26237 36731 26295 36737
rect 26344 36740 29500 36768
rect 25774 36660 25780 36712
rect 25832 36700 25838 36712
rect 26053 36703 26111 36709
rect 26053 36700 26065 36703
rect 25832 36672 26065 36700
rect 25832 36660 25838 36672
rect 26053 36669 26065 36672
rect 26099 36669 26111 36703
rect 26053 36663 26111 36669
rect 25225 36635 25283 36641
rect 25225 36601 25237 36635
rect 25271 36632 25283 36635
rect 26344 36632 26372 36740
rect 26970 36700 26976 36712
rect 26931 36672 26976 36700
rect 26970 36660 26976 36672
rect 27028 36660 27034 36712
rect 29086 36632 29092 36644
rect 25271 36604 26372 36632
rect 29047 36604 29092 36632
rect 25271 36601 25283 36604
rect 25225 36595 25283 36601
rect 25240 36564 25268 36595
rect 29086 36592 29092 36604
rect 29144 36592 29150 36644
rect 23216 36536 25268 36564
rect 29362 36524 29368 36576
rect 29420 36564 29426 36576
rect 29457 36567 29515 36573
rect 29457 36564 29469 36567
rect 29420 36536 29469 36564
rect 29420 36524 29426 36536
rect 29457 36533 29469 36536
rect 29503 36533 29515 36567
rect 29457 36527 29515 36533
rect 1104 36474 30820 36496
rect 1104 36422 5915 36474
rect 5967 36422 5979 36474
rect 6031 36422 6043 36474
rect 6095 36422 6107 36474
rect 6159 36422 6171 36474
rect 6223 36422 15846 36474
rect 15898 36422 15910 36474
rect 15962 36422 15974 36474
rect 16026 36422 16038 36474
rect 16090 36422 16102 36474
rect 16154 36422 25776 36474
rect 25828 36422 25840 36474
rect 25892 36422 25904 36474
rect 25956 36422 25968 36474
rect 26020 36422 26032 36474
rect 26084 36422 30820 36474
rect 1104 36400 30820 36422
rect 13262 36320 13268 36372
rect 13320 36360 13326 36372
rect 19150 36360 19156 36372
rect 13320 36332 19156 36360
rect 13320 36320 13326 36332
rect 19150 36320 19156 36332
rect 19208 36360 19214 36372
rect 19705 36363 19763 36369
rect 19705 36360 19717 36363
rect 19208 36332 19717 36360
rect 19208 36320 19214 36332
rect 19705 36329 19717 36332
rect 19751 36329 19763 36363
rect 19705 36323 19763 36329
rect 19794 36320 19800 36372
rect 19852 36360 19858 36372
rect 22370 36360 22376 36372
rect 19852 36332 22376 36360
rect 19852 36320 19858 36332
rect 22370 36320 22376 36332
rect 22428 36360 22434 36372
rect 24578 36360 24584 36372
rect 22428 36332 24584 36360
rect 22428 36320 22434 36332
rect 24578 36320 24584 36332
rect 24636 36320 24642 36372
rect 28258 36360 28264 36372
rect 28219 36332 28264 36360
rect 28258 36320 28264 36332
rect 28316 36320 28322 36372
rect 28902 36360 28908 36372
rect 28863 36332 28908 36360
rect 28902 36320 28908 36332
rect 28960 36320 28966 36372
rect 13814 36292 13820 36304
rect 12406 36264 13820 36292
rect 12406 36224 12434 36264
rect 13814 36252 13820 36264
rect 13872 36252 13878 36304
rect 22281 36295 22339 36301
rect 22281 36261 22293 36295
rect 22327 36292 22339 36295
rect 22646 36292 22652 36304
rect 22327 36264 22652 36292
rect 22327 36261 22339 36264
rect 22281 36255 22339 36261
rect 22646 36252 22652 36264
rect 22704 36292 22710 36304
rect 23014 36292 23020 36304
rect 22704 36264 23020 36292
rect 22704 36252 22710 36264
rect 23014 36252 23020 36264
rect 23072 36292 23078 36304
rect 23290 36292 23296 36304
rect 23072 36264 23296 36292
rect 23072 36252 23078 36264
rect 23290 36252 23296 36264
rect 23348 36252 23354 36304
rect 25038 36252 25044 36304
rect 25096 36292 25102 36304
rect 26694 36292 26700 36304
rect 25096 36264 26700 36292
rect 25096 36252 25102 36264
rect 26694 36252 26700 36264
rect 26752 36252 26758 36304
rect 11822 36196 12434 36224
rect 13004 36196 14688 36224
rect 11057 36159 11115 36165
rect 11057 36125 11069 36159
rect 11103 36156 11115 36159
rect 11238 36156 11244 36168
rect 11103 36128 11244 36156
rect 11103 36125 11115 36128
rect 11057 36119 11115 36125
rect 11238 36116 11244 36128
rect 11296 36116 11302 36168
rect 11606 36156 11612 36168
rect 11440 36128 11612 36156
rect 10778 36088 10784 36100
rect 10739 36060 10784 36088
rect 10778 36048 10784 36060
rect 10836 36048 10842 36100
rect 11149 36091 11207 36097
rect 11149 36057 11161 36091
rect 11195 36088 11207 36091
rect 11440 36088 11468 36128
rect 11606 36116 11612 36128
rect 11664 36116 11670 36168
rect 12618 36116 12624 36168
rect 12676 36156 12682 36168
rect 13004 36165 13032 36196
rect 12805 36159 12863 36165
rect 12805 36156 12817 36159
rect 12676 36128 12817 36156
rect 12676 36116 12682 36128
rect 12805 36125 12817 36128
rect 12851 36125 12863 36159
rect 12805 36119 12863 36125
rect 12989 36159 13047 36165
rect 12989 36125 13001 36159
rect 13035 36125 13047 36159
rect 12989 36119 13047 36125
rect 13081 36159 13139 36165
rect 13081 36125 13093 36159
rect 13127 36125 13139 36159
rect 13081 36119 13139 36125
rect 13173 36159 13231 36165
rect 13173 36125 13185 36159
rect 13219 36156 13231 36159
rect 13262 36156 13268 36168
rect 13219 36128 13268 36156
rect 13219 36125 13231 36128
rect 13173 36119 13231 36125
rect 11195 36060 11468 36088
rect 11517 36091 11575 36097
rect 11195 36057 11207 36060
rect 11149 36051 11207 36057
rect 11517 36057 11529 36091
rect 11563 36057 11575 36091
rect 11517 36051 11575 36057
rect 11885 36091 11943 36097
rect 11885 36057 11897 36091
rect 11931 36088 11943 36091
rect 12894 36088 12900 36100
rect 11931 36060 12900 36088
rect 11931 36057 11943 36060
rect 11885 36051 11943 36057
rect 9674 35980 9680 36032
rect 9732 36020 9738 36032
rect 11532 36020 11560 36051
rect 12894 36048 12900 36060
rect 12952 36048 12958 36100
rect 9732 35992 11560 36020
rect 9732 35980 9738 35992
rect 11974 35980 11980 36032
rect 12032 36020 12038 36032
rect 12069 36023 12127 36029
rect 12069 36020 12081 36023
rect 12032 35992 12081 36020
rect 12032 35980 12038 35992
rect 12069 35989 12081 35992
rect 12115 35989 12127 36023
rect 12069 35983 12127 35989
rect 12158 35980 12164 36032
rect 12216 36020 12222 36032
rect 13096 36020 13124 36119
rect 13262 36116 13268 36128
rect 13320 36116 13326 36168
rect 13357 36159 13415 36165
rect 13357 36125 13369 36159
rect 13403 36125 13415 36159
rect 13357 36119 13415 36125
rect 13372 36088 13400 36119
rect 13538 36116 13544 36168
rect 13596 36156 13602 36168
rect 14553 36159 14611 36165
rect 14553 36156 14565 36159
rect 13596 36128 14565 36156
rect 13596 36116 13602 36128
rect 14553 36125 14565 36128
rect 14599 36125 14611 36159
rect 14660 36156 14688 36196
rect 16666 36184 16672 36236
rect 16724 36224 16730 36236
rect 16853 36227 16911 36233
rect 16853 36224 16865 36227
rect 16724 36196 16865 36224
rect 16724 36184 16730 36196
rect 16853 36193 16865 36196
rect 16899 36193 16911 36227
rect 16853 36187 16911 36193
rect 19610 36184 19616 36236
rect 19668 36224 19674 36236
rect 20070 36224 20076 36236
rect 19668 36196 20076 36224
rect 19668 36184 19674 36196
rect 20070 36184 20076 36196
rect 20128 36224 20134 36236
rect 20257 36227 20315 36233
rect 20257 36224 20269 36227
rect 20128 36196 20269 36224
rect 20128 36184 20134 36196
rect 20257 36193 20269 36196
rect 20303 36193 20315 36227
rect 20257 36187 20315 36193
rect 22922 36184 22928 36236
rect 22980 36224 22986 36236
rect 24673 36227 24731 36233
rect 24673 36224 24685 36227
rect 22980 36196 24685 36224
rect 22980 36184 22986 36196
rect 24673 36193 24685 36196
rect 24719 36224 24731 36227
rect 24854 36224 24860 36236
rect 24719 36196 24860 36224
rect 24719 36193 24731 36196
rect 24673 36187 24731 36193
rect 24854 36184 24860 36196
rect 24912 36184 24918 36236
rect 25682 36224 25688 36236
rect 25643 36196 25688 36224
rect 25682 36184 25688 36196
rect 25740 36184 25746 36236
rect 17126 36165 17132 36168
rect 17120 36156 17132 36165
rect 14660 36128 16988 36156
rect 17087 36128 17132 36156
rect 14553 36119 14611 36125
rect 13906 36088 13912 36100
rect 13372 36060 13912 36088
rect 13906 36048 13912 36060
rect 13964 36048 13970 36100
rect 14820 36091 14878 36097
rect 14820 36057 14832 36091
rect 14866 36088 14878 36091
rect 15838 36088 15844 36100
rect 14866 36060 15844 36088
rect 14866 36057 14878 36060
rect 14820 36051 14878 36057
rect 15838 36048 15844 36060
rect 15896 36048 15902 36100
rect 16960 36088 16988 36128
rect 17120 36119 17132 36128
rect 17126 36116 17132 36119
rect 17184 36116 17190 36168
rect 18598 36116 18604 36168
rect 18656 36156 18662 36168
rect 19058 36156 19064 36168
rect 18656 36128 19064 36156
rect 18656 36116 18662 36128
rect 19058 36116 19064 36128
rect 19116 36116 19122 36168
rect 19536 36128 21404 36156
rect 19536 36088 19564 36128
rect 16960 36060 19564 36088
rect 19613 36091 19671 36097
rect 19613 36057 19625 36091
rect 19659 36057 19671 36091
rect 19613 36051 19671 36057
rect 20524 36091 20582 36097
rect 20524 36057 20536 36091
rect 20570 36088 20582 36091
rect 21266 36088 21272 36100
rect 20570 36060 21272 36088
rect 20570 36057 20582 36060
rect 20524 36051 20582 36057
rect 12216 35992 13124 36020
rect 12216 35980 12222 35992
rect 13262 35980 13268 36032
rect 13320 36020 13326 36032
rect 13541 36023 13599 36029
rect 13541 36020 13553 36023
rect 13320 35992 13553 36020
rect 13320 35980 13326 35992
rect 13541 35989 13553 35992
rect 13587 35989 13599 36023
rect 13541 35983 13599 35989
rect 15194 35980 15200 36032
rect 15252 36020 15258 36032
rect 15746 36020 15752 36032
rect 15252 35992 15752 36020
rect 15252 35980 15258 35992
rect 15746 35980 15752 35992
rect 15804 36020 15810 36032
rect 15933 36023 15991 36029
rect 15933 36020 15945 36023
rect 15804 35992 15945 36020
rect 15804 35980 15810 35992
rect 15933 35989 15945 35992
rect 15979 35989 15991 36023
rect 15933 35983 15991 35989
rect 17678 35980 17684 36032
rect 17736 36020 17742 36032
rect 18233 36023 18291 36029
rect 18233 36020 18245 36023
rect 17736 35992 18245 36020
rect 17736 35980 17742 35992
rect 18233 35989 18245 35992
rect 18279 35989 18291 36023
rect 18233 35983 18291 35989
rect 18690 35980 18696 36032
rect 18748 36020 18754 36032
rect 19058 36020 19064 36032
rect 18748 35992 19064 36020
rect 18748 35980 18754 35992
rect 19058 35980 19064 35992
rect 19116 36020 19122 36032
rect 19628 36020 19656 36051
rect 21266 36048 21272 36060
rect 21324 36048 21330 36100
rect 21376 36088 21404 36128
rect 22094 36116 22100 36168
rect 22152 36156 22158 36168
rect 22152 36128 22197 36156
rect 22152 36116 22158 36128
rect 22738 36116 22744 36168
rect 22796 36156 22802 36168
rect 23569 36159 23627 36165
rect 23569 36156 23581 36159
rect 22796 36128 23581 36156
rect 22796 36116 22802 36128
rect 23569 36125 23581 36128
rect 23615 36125 23627 36159
rect 23569 36119 23627 36125
rect 24486 36116 24492 36168
rect 24544 36156 24550 36168
rect 24581 36159 24639 36165
rect 24581 36156 24593 36159
rect 24544 36128 24593 36156
rect 24544 36116 24550 36128
rect 24581 36125 24593 36128
rect 24627 36156 24639 36159
rect 25409 36159 25467 36165
rect 25409 36156 25421 36159
rect 24627 36128 25421 36156
rect 24627 36125 24639 36128
rect 24581 36119 24639 36125
rect 25409 36125 25421 36128
rect 25455 36125 25467 36159
rect 25409 36119 25467 36125
rect 26881 36159 26939 36165
rect 26881 36125 26893 36159
rect 26927 36156 26939 36159
rect 27982 36156 27988 36168
rect 26927 36128 27988 36156
rect 26927 36125 26939 36128
rect 26881 36119 26939 36125
rect 27982 36116 27988 36128
rect 28040 36116 28046 36168
rect 28166 36116 28172 36168
rect 28224 36156 28230 36168
rect 28721 36159 28779 36165
rect 28721 36156 28733 36159
rect 28224 36128 28733 36156
rect 28224 36116 28230 36128
rect 28721 36125 28733 36128
rect 28767 36125 28779 36159
rect 28721 36119 28779 36125
rect 29270 36116 29276 36168
rect 29328 36156 29334 36168
rect 29825 36159 29883 36165
rect 29825 36156 29837 36159
rect 29328 36128 29837 36156
rect 29328 36116 29334 36128
rect 29825 36125 29837 36128
rect 29871 36125 29883 36159
rect 29825 36119 29883 36125
rect 22925 36091 22983 36097
rect 21376 36060 22692 36088
rect 19116 35992 19656 36020
rect 19116 35980 19122 35992
rect 21358 35980 21364 36032
rect 21416 36020 21422 36032
rect 21637 36023 21695 36029
rect 21637 36020 21649 36023
rect 21416 35992 21649 36020
rect 21416 35980 21422 35992
rect 21637 35989 21649 35992
rect 21683 35989 21695 36023
rect 22664 36020 22692 36060
rect 22925 36057 22937 36091
rect 22971 36088 22983 36091
rect 23106 36088 23112 36100
rect 22971 36060 23112 36088
rect 22971 36057 22983 36060
rect 22925 36051 22983 36057
rect 23106 36048 23112 36060
rect 23164 36088 23170 36100
rect 27148 36091 27206 36097
rect 23164 36060 23888 36088
rect 23164 36048 23170 36060
rect 23014 36020 23020 36032
rect 22664 35992 23020 36020
rect 21637 35983 21695 35989
rect 23014 35980 23020 35992
rect 23072 35980 23078 36032
rect 23750 36020 23756 36032
rect 23711 35992 23756 36020
rect 23750 35980 23756 35992
rect 23808 35980 23814 36032
rect 23860 36020 23888 36060
rect 27148 36057 27160 36091
rect 27194 36088 27206 36091
rect 27338 36088 27344 36100
rect 27194 36060 27344 36088
rect 27194 36057 27206 36060
rect 27148 36051 27206 36057
rect 27338 36048 27344 36060
rect 27396 36048 27402 36100
rect 27706 36020 27712 36032
rect 23860 35992 27712 36020
rect 27706 35980 27712 35992
rect 27764 35980 27770 36032
rect 30006 36020 30012 36032
rect 29967 35992 30012 36020
rect 30006 35980 30012 35992
rect 30064 35980 30070 36032
rect 1104 35930 30820 35952
rect 1104 35878 10880 35930
rect 10932 35878 10944 35930
rect 10996 35878 11008 35930
rect 11060 35878 11072 35930
rect 11124 35878 11136 35930
rect 11188 35878 20811 35930
rect 20863 35878 20875 35930
rect 20927 35878 20939 35930
rect 20991 35878 21003 35930
rect 21055 35878 21067 35930
rect 21119 35878 30820 35930
rect 1104 35856 30820 35878
rect 12437 35819 12495 35825
rect 12437 35785 12449 35819
rect 12483 35816 12495 35819
rect 20622 35816 20628 35828
rect 12483 35788 15884 35816
rect 12483 35785 12495 35788
rect 12437 35779 12495 35785
rect 10410 35748 10416 35760
rect 9048 35720 10416 35748
rect 9048 35689 9076 35720
rect 10410 35708 10416 35720
rect 10468 35708 10474 35760
rect 11790 35708 11796 35760
rect 11848 35748 11854 35760
rect 15746 35748 15752 35760
rect 11848 35720 12434 35748
rect 11848 35708 11854 35720
rect 9306 35689 9312 35692
rect 9033 35683 9091 35689
rect 9033 35649 9045 35683
rect 9079 35649 9091 35683
rect 9300 35680 9312 35689
rect 9267 35652 9312 35680
rect 9033 35643 9091 35649
rect 9300 35643 9312 35652
rect 9306 35640 9312 35643
rect 9364 35640 9370 35692
rect 12066 35680 12072 35692
rect 12027 35652 12072 35680
rect 12066 35640 12072 35652
rect 12124 35640 12130 35692
rect 12250 35680 12256 35692
rect 12211 35652 12256 35680
rect 12250 35640 12256 35652
rect 12308 35640 12314 35692
rect 12406 35680 12434 35720
rect 15120 35720 15608 35748
rect 12989 35683 13047 35689
rect 12989 35680 13001 35683
rect 12406 35652 13001 35680
rect 12989 35649 13001 35652
rect 13035 35680 13047 35683
rect 13538 35680 13544 35692
rect 13035 35652 13544 35680
rect 13035 35649 13047 35652
rect 12989 35643 13047 35649
rect 13538 35640 13544 35652
rect 13596 35640 13602 35692
rect 15120 35689 15148 35720
rect 15105 35683 15163 35689
rect 15105 35649 15117 35683
rect 15151 35649 15163 35683
rect 15105 35643 15163 35649
rect 15289 35683 15347 35689
rect 15289 35649 15301 35683
rect 15335 35649 15347 35683
rect 15289 35643 15347 35649
rect 13262 35612 13268 35624
rect 13223 35584 13268 35612
rect 13262 35572 13268 35584
rect 13320 35572 13326 35624
rect 14458 35572 14464 35624
rect 14516 35612 14522 35624
rect 15304 35612 15332 35643
rect 15378 35640 15384 35692
rect 15436 35680 15442 35692
rect 15436 35652 15481 35680
rect 15436 35640 15442 35652
rect 15470 35612 15476 35624
rect 14516 35584 15332 35612
rect 15431 35584 15476 35612
rect 14516 35572 14522 35584
rect 15470 35572 15476 35584
rect 15528 35572 15534 35624
rect 15580 35612 15608 35720
rect 15672 35720 15752 35748
rect 15672 35689 15700 35720
rect 15746 35708 15752 35720
rect 15804 35708 15810 35760
rect 15856 35748 15884 35788
rect 20456 35788 20628 35816
rect 19978 35748 19984 35760
rect 15856 35720 19984 35748
rect 19978 35708 19984 35720
rect 20036 35708 20042 35760
rect 20156 35751 20214 35757
rect 20156 35717 20168 35751
rect 20202 35748 20214 35751
rect 20456 35748 20484 35788
rect 20622 35776 20628 35788
rect 20680 35776 20686 35828
rect 22922 35816 22928 35828
rect 22066 35788 22928 35816
rect 20202 35720 20484 35748
rect 20202 35717 20214 35720
rect 20156 35711 20214 35717
rect 20806 35708 20812 35760
rect 20864 35748 20870 35760
rect 22066 35748 22094 35788
rect 22922 35776 22928 35788
rect 22980 35816 22986 35828
rect 23198 35816 23204 35828
rect 22980 35788 23204 35816
rect 22980 35776 22986 35788
rect 23198 35776 23204 35788
rect 23256 35776 23262 35828
rect 25961 35819 26019 35825
rect 25961 35785 25973 35819
rect 26007 35816 26019 35819
rect 26510 35816 26516 35828
rect 26007 35788 26516 35816
rect 26007 35785 26019 35788
rect 25961 35779 26019 35785
rect 26510 35776 26516 35788
rect 26568 35776 26574 35828
rect 27798 35816 27804 35828
rect 27759 35788 27804 35816
rect 27798 35776 27804 35788
rect 27856 35776 27862 35828
rect 27890 35776 27896 35828
rect 27948 35816 27954 35828
rect 29641 35819 29699 35825
rect 29641 35816 29653 35819
rect 27948 35788 29653 35816
rect 27948 35776 27954 35788
rect 29641 35785 29653 35788
rect 29687 35785 29699 35819
rect 29641 35779 29699 35785
rect 22646 35748 22652 35760
rect 20864 35720 22094 35748
rect 22204 35720 22652 35748
rect 20864 35708 20870 35720
rect 15657 35683 15715 35689
rect 15657 35649 15669 35683
rect 15703 35649 15715 35683
rect 16945 35683 17003 35689
rect 16945 35680 16957 35683
rect 15657 35643 15715 35649
rect 15764 35652 16957 35680
rect 15764 35612 15792 35652
rect 16945 35649 16957 35652
rect 16991 35680 17003 35683
rect 17126 35680 17132 35692
rect 16991 35652 17132 35680
rect 16991 35649 17003 35652
rect 16945 35643 17003 35649
rect 17126 35640 17132 35652
rect 17184 35640 17190 35692
rect 17954 35680 17960 35692
rect 17915 35652 17960 35680
rect 17954 35640 17960 35652
rect 18012 35640 18018 35692
rect 18141 35683 18199 35689
rect 18141 35649 18153 35683
rect 18187 35680 18199 35683
rect 18322 35680 18328 35692
rect 18187 35652 18328 35680
rect 18187 35649 18199 35652
rect 18141 35643 18199 35649
rect 18322 35640 18328 35652
rect 18380 35640 18386 35692
rect 18601 35683 18659 35689
rect 18601 35649 18613 35683
rect 18647 35680 18659 35683
rect 19426 35680 19432 35692
rect 18647 35652 19432 35680
rect 18647 35649 18659 35652
rect 18601 35643 18659 35649
rect 19426 35640 19432 35652
rect 19484 35640 19490 35692
rect 19610 35640 19616 35692
rect 19668 35680 19674 35692
rect 19889 35683 19947 35689
rect 19889 35680 19901 35683
rect 19668 35652 19901 35680
rect 19668 35640 19674 35652
rect 19889 35649 19901 35652
rect 19935 35649 19947 35683
rect 22204 35680 22232 35720
rect 22646 35708 22652 35720
rect 22704 35748 22710 35760
rect 22704 35720 25820 35748
rect 22704 35708 22710 35720
rect 19889 35643 19947 35649
rect 19996 35652 22232 35680
rect 22557 35683 22615 35689
rect 15580 35584 15792 35612
rect 15838 35572 15844 35624
rect 15896 35612 15902 35624
rect 15896 35584 15941 35612
rect 15896 35572 15902 35584
rect 16574 35572 16580 35624
rect 16632 35612 16638 35624
rect 16669 35615 16727 35621
rect 16669 35612 16681 35615
rect 16632 35584 16681 35612
rect 16632 35572 16638 35584
rect 16669 35581 16681 35584
rect 16715 35581 16727 35615
rect 18874 35612 18880 35624
rect 18835 35584 18880 35612
rect 16669 35575 16727 35581
rect 18874 35572 18880 35584
rect 18932 35572 18938 35624
rect 19702 35572 19708 35624
rect 19760 35612 19766 35624
rect 19996 35612 20024 35652
rect 22557 35649 22569 35683
rect 22603 35680 22615 35683
rect 23201 35683 23259 35689
rect 22603 35652 23152 35680
rect 22603 35649 22615 35652
rect 22557 35643 22615 35649
rect 19760 35584 20024 35612
rect 19760 35572 19766 35584
rect 22094 35572 22100 35624
rect 22152 35612 22158 35624
rect 22741 35615 22799 35621
rect 22741 35612 22753 35615
rect 22152 35584 22753 35612
rect 22152 35572 22158 35584
rect 22741 35581 22753 35584
rect 22787 35581 22799 35615
rect 23124 35612 23152 35652
rect 23201 35649 23213 35683
rect 23247 35680 23259 35683
rect 23382 35680 23388 35692
rect 23247 35652 23388 35680
rect 23247 35649 23259 35652
rect 23201 35643 23259 35649
rect 23382 35640 23388 35652
rect 23440 35640 23446 35692
rect 23750 35640 23756 35692
rect 23808 35680 23814 35692
rect 23937 35683 23995 35689
rect 23937 35680 23949 35683
rect 23808 35652 23949 35680
rect 23808 35640 23814 35652
rect 23937 35649 23949 35652
rect 23983 35649 23995 35683
rect 23937 35643 23995 35649
rect 24204 35683 24262 35689
rect 24204 35649 24216 35683
rect 24250 35680 24262 35683
rect 25130 35680 25136 35692
rect 24250 35652 25136 35680
rect 24250 35649 24262 35652
rect 24204 35643 24262 35649
rect 25130 35640 25136 35652
rect 25188 35640 25194 35692
rect 25792 35689 25820 35720
rect 25777 35683 25835 35689
rect 25777 35649 25789 35683
rect 25823 35649 25835 35683
rect 26528 35680 26556 35776
rect 29457 35751 29515 35757
rect 29457 35717 29469 35751
rect 29503 35717 29515 35751
rect 29457 35711 29515 35717
rect 26973 35683 27031 35689
rect 26973 35680 26985 35683
rect 26528 35652 26985 35680
rect 25777 35643 25835 35649
rect 26973 35649 26985 35652
rect 27019 35680 27031 35683
rect 27617 35683 27675 35689
rect 27617 35680 27629 35683
rect 27019 35652 27629 35680
rect 27019 35649 27031 35652
rect 26973 35643 27031 35649
rect 27617 35649 27629 35652
rect 27663 35649 27675 35683
rect 27617 35643 27675 35649
rect 27706 35640 27712 35692
rect 27764 35680 27770 35692
rect 28626 35680 28632 35692
rect 27764 35652 28632 35680
rect 27764 35640 27770 35652
rect 28626 35640 28632 35652
rect 28684 35640 28690 35692
rect 29086 35680 29092 35692
rect 29047 35652 29092 35680
rect 29086 35640 29092 35652
rect 29144 35640 29150 35692
rect 23842 35612 23848 35624
rect 23124 35584 23848 35612
rect 22741 35575 22799 35581
rect 23842 35572 23848 35584
rect 23900 35572 23906 35624
rect 29472 35612 29500 35711
rect 25332 35584 29500 35612
rect 19794 35544 19800 35556
rect 17328 35516 19800 35544
rect 9674 35436 9680 35488
rect 9732 35476 9738 35488
rect 10413 35479 10471 35485
rect 10413 35476 10425 35479
rect 9732 35448 10425 35476
rect 9732 35436 9738 35448
rect 10413 35445 10425 35448
rect 10459 35445 10471 35479
rect 10413 35439 10471 35445
rect 13906 35436 13912 35488
rect 13964 35476 13970 35488
rect 14369 35479 14427 35485
rect 14369 35476 14381 35479
rect 13964 35448 14381 35476
rect 13964 35436 13970 35448
rect 14369 35445 14381 35448
rect 14415 35445 14427 35479
rect 14369 35439 14427 35445
rect 14458 35436 14464 35488
rect 14516 35476 14522 35488
rect 17328 35476 17356 35516
rect 19794 35504 19800 35516
rect 19852 35504 19858 35556
rect 24946 35504 24952 35556
rect 25004 35544 25010 35556
rect 25332 35553 25360 35584
rect 25317 35547 25375 35553
rect 25317 35544 25329 35547
rect 25004 35516 25329 35544
rect 25004 35504 25010 35516
rect 25317 35513 25329 35516
rect 25363 35513 25375 35547
rect 25317 35507 25375 35513
rect 14516 35448 17356 35476
rect 17957 35479 18015 35485
rect 14516 35436 14522 35448
rect 17957 35445 17969 35479
rect 18003 35476 18015 35479
rect 18046 35476 18052 35488
rect 18003 35448 18052 35476
rect 18003 35445 18015 35448
rect 17957 35439 18015 35445
rect 18046 35436 18052 35448
rect 18104 35436 18110 35488
rect 20254 35436 20260 35488
rect 20312 35476 20318 35488
rect 21269 35479 21327 35485
rect 21269 35476 21281 35479
rect 20312 35448 21281 35476
rect 20312 35436 20318 35448
rect 21269 35445 21281 35448
rect 21315 35445 21327 35479
rect 21269 35439 21327 35445
rect 22830 35436 22836 35488
rect 22888 35476 22894 35488
rect 23385 35479 23443 35485
rect 23385 35476 23397 35479
rect 22888 35448 23397 35476
rect 22888 35436 22894 35448
rect 23385 35445 23397 35448
rect 23431 35476 23443 35479
rect 23566 35476 23572 35488
rect 23431 35448 23572 35476
rect 23431 35445 23443 35448
rect 23385 35439 23443 35445
rect 23566 35436 23572 35448
rect 23624 35436 23630 35488
rect 26418 35436 26424 35488
rect 26476 35476 26482 35488
rect 27157 35479 27215 35485
rect 27157 35476 27169 35479
rect 26476 35448 27169 35476
rect 26476 35436 26482 35448
rect 27157 35445 27169 35448
rect 27203 35445 27215 35479
rect 27157 35439 27215 35445
rect 28445 35479 28503 35485
rect 28445 35445 28457 35479
rect 28491 35476 28503 35479
rect 29457 35479 29515 35485
rect 29457 35476 29469 35479
rect 28491 35448 29469 35476
rect 28491 35445 28503 35448
rect 28445 35439 28503 35445
rect 29457 35445 29469 35448
rect 29503 35476 29515 35479
rect 29914 35476 29920 35488
rect 29503 35448 29920 35476
rect 29503 35445 29515 35448
rect 29457 35439 29515 35445
rect 29914 35436 29920 35448
rect 29972 35436 29978 35488
rect 1104 35386 30820 35408
rect 1104 35334 5915 35386
rect 5967 35334 5979 35386
rect 6031 35334 6043 35386
rect 6095 35334 6107 35386
rect 6159 35334 6171 35386
rect 6223 35334 15846 35386
rect 15898 35334 15910 35386
rect 15962 35334 15974 35386
rect 16026 35334 16038 35386
rect 16090 35334 16102 35386
rect 16154 35334 25776 35386
rect 25828 35334 25840 35386
rect 25892 35334 25904 35386
rect 25956 35334 25968 35386
rect 26020 35334 26032 35386
rect 26084 35334 30820 35386
rect 1104 35312 30820 35334
rect 12437 35275 12495 35281
rect 12437 35241 12449 35275
rect 12483 35272 12495 35275
rect 14458 35272 14464 35284
rect 12483 35244 14464 35272
rect 12483 35241 12495 35244
rect 12437 35235 12495 35241
rect 14458 35232 14464 35244
rect 14516 35232 14522 35284
rect 14645 35275 14703 35281
rect 14645 35241 14657 35275
rect 14691 35272 14703 35275
rect 15381 35275 15439 35281
rect 15381 35272 15393 35275
rect 14691 35244 15393 35272
rect 14691 35241 14703 35244
rect 14645 35235 14703 35241
rect 15381 35241 15393 35244
rect 15427 35272 15439 35275
rect 16666 35272 16672 35284
rect 15427 35244 16672 35272
rect 15427 35241 15439 35244
rect 15381 35235 15439 35241
rect 16666 35232 16672 35244
rect 16724 35232 16730 35284
rect 16758 35232 16764 35284
rect 16816 35272 16822 35284
rect 16853 35275 16911 35281
rect 16853 35272 16865 35275
rect 16816 35244 16865 35272
rect 16816 35232 16822 35244
rect 16853 35241 16865 35244
rect 16899 35241 16911 35275
rect 16853 35235 16911 35241
rect 17954 35232 17960 35284
rect 18012 35272 18018 35284
rect 18506 35272 18512 35284
rect 18012 35244 18512 35272
rect 18012 35232 18018 35244
rect 18506 35232 18512 35244
rect 18564 35272 18570 35284
rect 18601 35275 18659 35281
rect 18601 35272 18613 35275
rect 18564 35244 18613 35272
rect 18564 35232 18570 35244
rect 18601 35241 18613 35244
rect 18647 35241 18659 35275
rect 18601 35235 18659 35241
rect 19610 35232 19616 35284
rect 19668 35272 19674 35284
rect 21913 35275 21971 35281
rect 21913 35272 21925 35275
rect 19668 35244 21925 35272
rect 19668 35232 19674 35244
rect 21913 35241 21925 35244
rect 21959 35272 21971 35275
rect 23382 35272 23388 35284
rect 21959 35244 22094 35272
rect 23343 35244 23388 35272
rect 21959 35241 21971 35244
rect 21913 35235 21971 35241
rect 17865 35207 17923 35213
rect 17865 35173 17877 35207
rect 17911 35204 17923 35207
rect 18138 35204 18144 35216
rect 17911 35176 18144 35204
rect 17911 35173 17923 35176
rect 17865 35167 17923 35173
rect 18138 35164 18144 35176
rect 18196 35164 18202 35216
rect 18874 35164 18880 35216
rect 18932 35204 18938 35216
rect 21266 35204 21272 35216
rect 18932 35176 19840 35204
rect 21227 35176 21272 35204
rect 18932 35164 18938 35176
rect 19812 35148 19840 35176
rect 21266 35164 21272 35176
rect 21324 35164 21330 35216
rect 19702 35136 19708 35148
rect 10888 35108 15608 35136
rect 1578 35068 1584 35080
rect 1539 35040 1584 35068
rect 1578 35028 1584 35040
rect 1636 35028 1642 35080
rect 10134 35028 10140 35080
rect 10192 35068 10198 35080
rect 10888 35077 10916 35108
rect 10873 35071 10931 35077
rect 10873 35068 10885 35071
rect 10192 35040 10885 35068
rect 10192 35028 10198 35040
rect 10873 35037 10885 35040
rect 10919 35037 10931 35071
rect 10873 35031 10931 35037
rect 12069 35071 12127 35077
rect 12069 35037 12081 35071
rect 12115 35037 12127 35071
rect 12250 35068 12256 35080
rect 12211 35040 12256 35068
rect 12069 35031 12127 35037
rect 12084 35000 12112 35031
rect 12250 35028 12256 35040
rect 12308 35028 12314 35080
rect 13357 35071 13415 35077
rect 13357 35037 13369 35071
rect 13403 35068 13415 35071
rect 15194 35068 15200 35080
rect 13403 35040 15200 35068
rect 13403 35037 13415 35040
rect 13357 35031 13415 35037
rect 15194 35028 15200 35040
rect 15252 35028 15258 35080
rect 15378 35068 15384 35080
rect 15291 35040 15384 35068
rect 15378 35028 15384 35040
rect 15436 35068 15442 35080
rect 15473 35071 15531 35077
rect 15473 35068 15485 35071
rect 15436 35040 15485 35068
rect 15436 35028 15442 35040
rect 15473 35037 15485 35040
rect 15519 35037 15531 35071
rect 15580 35068 15608 35108
rect 16500 35108 19708 35136
rect 16500 35068 16528 35108
rect 19702 35096 19708 35108
rect 19760 35096 19766 35148
rect 19794 35096 19800 35148
rect 19852 35136 19858 35148
rect 20346 35136 20352 35148
rect 19852 35108 20352 35136
rect 19852 35096 19858 35108
rect 20346 35096 20352 35108
rect 20404 35136 20410 35148
rect 20809 35139 20867 35145
rect 20809 35136 20821 35139
rect 20404 35108 20821 35136
rect 20404 35096 20410 35108
rect 20809 35105 20821 35108
rect 20855 35105 20867 35139
rect 20809 35099 20867 35105
rect 15580 35040 16528 35068
rect 15473 35031 15531 35037
rect 16758 35028 16764 35080
rect 16816 35068 16822 35080
rect 17438 35071 17496 35077
rect 17438 35068 17450 35071
rect 16816 35040 17450 35068
rect 16816 35028 16822 35040
rect 17438 35037 17450 35040
rect 17484 35037 17496 35071
rect 17438 35031 17496 35037
rect 17770 35028 17776 35080
rect 17828 35068 17834 35080
rect 17957 35071 18015 35077
rect 17957 35068 17969 35071
rect 17828 35040 17969 35068
rect 17828 35028 17834 35040
rect 17957 35037 17969 35040
rect 18003 35037 18015 35071
rect 17957 35031 18015 35037
rect 19058 35028 19064 35080
rect 19116 35068 19122 35080
rect 19245 35071 19303 35077
rect 19245 35068 19257 35071
rect 19116 35040 19257 35068
rect 19116 35028 19122 35040
rect 19245 35037 19257 35040
rect 19291 35037 19303 35071
rect 19245 35031 19303 35037
rect 19521 35071 19579 35077
rect 19521 35037 19533 35071
rect 19567 35068 19579 35071
rect 20438 35068 20444 35080
rect 19567 35040 20444 35068
rect 19567 35037 19579 35040
rect 19521 35031 19579 35037
rect 20438 35028 20444 35040
rect 20496 35028 20502 35080
rect 20533 35071 20591 35077
rect 20533 35037 20545 35071
rect 20579 35037 20591 35071
rect 20533 35031 20591 35037
rect 20717 35071 20775 35077
rect 20717 35037 20729 35071
rect 20763 35037 20775 35071
rect 20717 35031 20775 35037
rect 2746 34972 12112 35000
rect 1397 34935 1455 34941
rect 1397 34901 1409 34935
rect 1443 34932 1455 34935
rect 2746 34932 2774 34972
rect 13170 34960 13176 35012
rect 13228 35000 13234 35012
rect 14553 35003 14611 35009
rect 14553 35000 14565 35003
rect 13228 34972 14565 35000
rect 13228 34960 13234 34972
rect 14553 34969 14565 34972
rect 14599 34969 14611 35003
rect 14553 34963 14611 34969
rect 15654 34960 15660 35012
rect 15712 35009 15718 35012
rect 15712 35003 15776 35009
rect 15712 34969 15730 35003
rect 15764 34969 15776 35003
rect 15712 34963 15776 34969
rect 18509 35003 18567 35009
rect 18509 34969 18521 35003
rect 18555 35000 18567 35003
rect 20162 35000 20168 35012
rect 18555 34972 20168 35000
rect 18555 34969 18567 34972
rect 18509 34963 18567 34969
rect 15712 34960 15718 34963
rect 20162 34960 20168 34972
rect 20220 34960 20226 35012
rect 1443 34904 2774 34932
rect 11057 34935 11115 34941
rect 1443 34901 1455 34904
rect 1397 34895 1455 34901
rect 11057 34901 11069 34935
rect 11103 34932 11115 34935
rect 11238 34932 11244 34944
rect 11103 34904 11244 34932
rect 11103 34901 11115 34904
rect 11057 34895 11115 34901
rect 11238 34892 11244 34904
rect 11296 34892 11302 34944
rect 13449 34935 13507 34941
rect 13449 34901 13461 34935
rect 13495 34932 13507 34935
rect 14918 34932 14924 34944
rect 13495 34904 14924 34932
rect 13495 34901 13507 34904
rect 13449 34895 13507 34901
rect 14918 34892 14924 34904
rect 14976 34892 14982 34944
rect 17034 34892 17040 34944
rect 17092 34932 17098 34944
rect 17313 34935 17371 34941
rect 17313 34932 17325 34935
rect 17092 34904 17325 34932
rect 17092 34892 17098 34904
rect 17313 34901 17325 34904
rect 17359 34901 17371 34935
rect 17313 34895 17371 34901
rect 17402 34892 17408 34944
rect 17460 34932 17466 34944
rect 17497 34935 17555 34941
rect 17497 34932 17509 34935
rect 17460 34904 17509 34932
rect 17460 34892 17466 34904
rect 17497 34901 17509 34904
rect 17543 34901 17555 34935
rect 17497 34895 17555 34901
rect 19518 34892 19524 34944
rect 19576 34932 19582 34944
rect 20548 34932 20576 35031
rect 19576 34904 20576 34932
rect 20732 34932 20760 35031
rect 20898 35028 20904 35080
rect 20956 35068 20962 35080
rect 21085 35071 21143 35077
rect 20956 35040 21001 35068
rect 20956 35028 20962 35040
rect 21085 35037 21097 35071
rect 21131 35068 21143 35071
rect 21358 35068 21364 35080
rect 21131 35040 21364 35068
rect 21131 35037 21143 35040
rect 21085 35031 21143 35037
rect 21358 35028 21364 35040
rect 21416 35028 21422 35080
rect 22066 35068 22094 35244
rect 23382 35232 23388 35244
rect 23440 35232 23446 35284
rect 25130 35272 25136 35284
rect 25091 35244 25136 35272
rect 25130 35232 25136 35244
rect 25188 35232 25194 35284
rect 26605 35275 26663 35281
rect 26605 35241 26617 35275
rect 26651 35272 26663 35275
rect 26970 35272 26976 35284
rect 26651 35244 26976 35272
rect 26651 35241 26663 35244
rect 26605 35235 26663 35241
rect 26970 35232 26976 35244
rect 27028 35232 27034 35284
rect 28350 35272 28356 35284
rect 28000 35244 28356 35272
rect 24394 35164 24400 35216
rect 24452 35164 24458 35216
rect 25777 35207 25835 35213
rect 25777 35173 25789 35207
rect 25823 35204 25835 35207
rect 28000 35204 28028 35244
rect 28350 35232 28356 35244
rect 28408 35232 28414 35284
rect 28534 35232 28540 35284
rect 28592 35272 28598 35284
rect 29914 35272 29920 35284
rect 28592 35244 29684 35272
rect 29875 35244 29920 35272
rect 28592 35232 28598 35244
rect 25823 35176 28028 35204
rect 28077 35207 28135 35213
rect 25823 35173 25835 35176
rect 25777 35167 25835 35173
rect 28077 35173 28089 35207
rect 28123 35204 28135 35207
rect 29086 35204 29092 35216
rect 28123 35176 29092 35204
rect 28123 35173 28135 35176
rect 28077 35167 28135 35173
rect 29086 35164 29092 35176
rect 29144 35204 29150 35216
rect 29549 35207 29607 35213
rect 29549 35204 29561 35207
rect 29144 35176 29561 35204
rect 29144 35164 29150 35176
rect 29549 35173 29561 35176
rect 29595 35173 29607 35207
rect 29656 35204 29684 35244
rect 29914 35232 29920 35244
rect 29972 35232 29978 35284
rect 30101 35275 30159 35281
rect 30101 35241 30113 35275
rect 30147 35241 30159 35275
rect 30101 35235 30159 35241
rect 30116 35204 30144 35235
rect 29656 35176 30144 35204
rect 29549 35167 29607 35173
rect 24412 35136 24440 35164
rect 24673 35139 24731 35145
rect 24412 35108 24624 35136
rect 22649 35071 22707 35077
rect 22649 35068 22661 35071
rect 22066 35040 22661 35068
rect 22649 35037 22661 35040
rect 22695 35068 22707 35071
rect 23293 35071 23351 35077
rect 23293 35068 23305 35071
rect 22695 35040 23305 35068
rect 22695 35037 22707 35040
rect 22649 35031 22707 35037
rect 23293 35037 23305 35040
rect 23339 35037 23351 35071
rect 23293 35031 23351 35037
rect 23474 35028 23480 35080
rect 23532 35068 23538 35080
rect 24596 35077 24624 35108
rect 24673 35105 24685 35139
rect 24719 35136 24731 35139
rect 24854 35136 24860 35148
rect 24719 35108 24860 35136
rect 24719 35105 24731 35108
rect 24673 35099 24731 35105
rect 24854 35096 24860 35108
rect 24912 35096 24918 35148
rect 30098 35136 30104 35148
rect 27632 35108 30104 35136
rect 24397 35071 24455 35077
rect 24397 35068 24409 35071
rect 23532 35040 24409 35068
rect 23532 35028 23538 35040
rect 24397 35037 24409 35040
rect 24443 35037 24455 35071
rect 24397 35031 24455 35037
rect 24581 35071 24639 35077
rect 24581 35037 24593 35071
rect 24627 35037 24639 35071
rect 24581 35031 24639 35037
rect 24765 35071 24823 35077
rect 24765 35037 24777 35071
rect 24811 35037 24823 35071
rect 24946 35068 24952 35080
rect 24907 35040 24952 35068
rect 24765 35031 24823 35037
rect 21818 35000 21824 35012
rect 21779 34972 21824 35000
rect 21818 34960 21824 34972
rect 21876 34960 21882 35012
rect 24118 34960 24124 35012
rect 24176 35000 24182 35012
rect 24486 35000 24492 35012
rect 24176 34972 24492 35000
rect 24176 34960 24182 34972
rect 24486 34960 24492 34972
rect 24544 35000 24550 35012
rect 24780 35000 24808 35031
rect 24946 35028 24952 35040
rect 25004 35028 25010 35080
rect 25961 35071 26019 35077
rect 25961 35037 25973 35071
rect 26007 35037 26019 35071
rect 26418 35068 26424 35080
rect 26379 35040 26424 35068
rect 25961 35031 26019 35037
rect 24544 34972 24808 35000
rect 25976 35000 26004 35031
rect 26418 35028 26424 35040
rect 26476 35028 26482 35080
rect 27632 35077 27660 35108
rect 30098 35096 30104 35108
rect 30156 35096 30162 35148
rect 27617 35071 27675 35077
rect 27617 35037 27629 35071
rect 27663 35037 27675 35071
rect 28258 35068 28264 35080
rect 28219 35040 28264 35068
rect 27617 35031 27675 35037
rect 28258 35028 28264 35040
rect 28316 35028 28322 35080
rect 28718 35068 28724 35080
rect 28679 35040 28724 35068
rect 28718 35028 28724 35040
rect 28776 35028 28782 35080
rect 29454 35000 29460 35012
rect 25976 34972 29460 35000
rect 24544 34960 24550 34972
rect 29454 34960 29460 34972
rect 29512 34960 29518 35012
rect 22002 34932 22008 34944
rect 20732 34904 22008 34932
rect 19576 34892 19582 34904
rect 22002 34892 22008 34904
rect 22060 34892 22066 34944
rect 22370 34892 22376 34944
rect 22428 34932 22434 34944
rect 22741 34935 22799 34941
rect 22741 34932 22753 34935
rect 22428 34904 22753 34932
rect 22428 34892 22434 34904
rect 22741 34901 22753 34904
rect 22787 34901 22799 34935
rect 22741 34895 22799 34901
rect 27433 34935 27491 34941
rect 27433 34901 27445 34935
rect 27479 34932 27491 34935
rect 27982 34932 27988 34944
rect 27479 34904 27988 34932
rect 27479 34901 27491 34904
rect 27433 34895 27491 34901
rect 27982 34892 27988 34904
rect 28040 34892 28046 34944
rect 28902 34932 28908 34944
rect 28863 34904 28908 34932
rect 28902 34892 28908 34904
rect 28960 34892 28966 34944
rect 28994 34892 29000 34944
rect 29052 34932 29058 34944
rect 29917 34935 29975 34941
rect 29917 34932 29929 34935
rect 29052 34904 29929 34932
rect 29052 34892 29058 34904
rect 29917 34901 29929 34904
rect 29963 34901 29975 34935
rect 29917 34895 29975 34901
rect 1104 34842 30820 34864
rect 1104 34790 10880 34842
rect 10932 34790 10944 34842
rect 10996 34790 11008 34842
rect 11060 34790 11072 34842
rect 11124 34790 11136 34842
rect 11188 34790 20811 34842
rect 20863 34790 20875 34842
rect 20927 34790 20939 34842
rect 20991 34790 21003 34842
rect 21055 34790 21067 34842
rect 21119 34790 30820 34842
rect 1104 34768 30820 34790
rect 10686 34728 10692 34740
rect 10599 34700 10692 34728
rect 10686 34688 10692 34700
rect 10744 34728 10750 34740
rect 11330 34728 11336 34740
rect 10744 34700 11336 34728
rect 10744 34688 10750 34700
rect 11330 34688 11336 34700
rect 11388 34688 11394 34740
rect 14829 34731 14887 34737
rect 14829 34697 14841 34731
rect 14875 34728 14887 34731
rect 17218 34728 17224 34740
rect 14875 34700 16160 34728
rect 17179 34700 17224 34728
rect 14875 34697 14887 34700
rect 14829 34691 14887 34697
rect 13716 34663 13774 34669
rect 13716 34629 13728 34663
rect 13762 34660 13774 34663
rect 16025 34663 16083 34669
rect 16025 34660 16037 34663
rect 13762 34632 16037 34660
rect 13762 34629 13774 34632
rect 13716 34623 13774 34629
rect 16025 34629 16037 34632
rect 16071 34629 16083 34663
rect 16025 34623 16083 34629
rect 10042 34552 10048 34604
rect 10100 34592 10106 34604
rect 10505 34595 10563 34601
rect 10505 34592 10517 34595
rect 10100 34564 10517 34592
rect 10100 34552 10106 34564
rect 10505 34561 10517 34564
rect 10551 34561 10563 34595
rect 10505 34555 10563 34561
rect 11784 34595 11842 34601
rect 11784 34561 11796 34595
rect 11830 34592 11842 34595
rect 12158 34592 12164 34604
rect 11830 34564 12164 34592
rect 11830 34561 11842 34564
rect 11784 34555 11842 34561
rect 12158 34552 12164 34564
rect 12216 34552 12222 34604
rect 13449 34595 13507 34601
rect 13449 34561 13461 34595
rect 13495 34592 13507 34595
rect 13538 34592 13544 34604
rect 13495 34564 13544 34592
rect 13495 34561 13507 34564
rect 13449 34555 13507 34561
rect 13538 34552 13544 34564
rect 13596 34552 13602 34604
rect 14274 34552 14280 34604
rect 14332 34592 14338 34604
rect 14332 34564 14504 34592
rect 14332 34552 14338 34564
rect 11514 34524 11520 34536
rect 11475 34496 11520 34524
rect 11514 34484 11520 34496
rect 11572 34484 11578 34536
rect 14476 34524 14504 34564
rect 15010 34552 15016 34604
rect 15068 34592 15074 34604
rect 15289 34595 15347 34601
rect 15289 34592 15301 34595
rect 15068 34564 15301 34592
rect 15068 34552 15074 34564
rect 15289 34561 15301 34564
rect 15335 34561 15347 34595
rect 15289 34555 15347 34561
rect 15473 34595 15531 34601
rect 15473 34561 15485 34595
rect 15519 34561 15531 34595
rect 15473 34555 15531 34561
rect 15565 34595 15623 34601
rect 15565 34561 15577 34595
rect 15611 34592 15623 34595
rect 15841 34595 15899 34601
rect 15611 34564 15792 34592
rect 15611 34561 15623 34564
rect 15565 34555 15623 34561
rect 15488 34524 15516 34555
rect 14476 34496 15516 34524
rect 15657 34527 15715 34533
rect 15657 34493 15669 34527
rect 15703 34493 15715 34527
rect 15764 34524 15792 34564
rect 15841 34561 15853 34595
rect 15887 34592 15899 34595
rect 16132 34592 16160 34700
rect 17218 34688 17224 34700
rect 17276 34688 17282 34740
rect 17310 34688 17316 34740
rect 17368 34728 17374 34740
rect 17405 34731 17463 34737
rect 17405 34728 17417 34731
rect 17368 34700 17417 34728
rect 17368 34688 17374 34700
rect 17405 34697 17417 34700
rect 17451 34697 17463 34731
rect 17405 34691 17463 34697
rect 17926 34700 19820 34728
rect 17926 34660 17954 34700
rect 17880 34632 17954 34660
rect 17880 34601 17908 34632
rect 18782 34620 18788 34672
rect 18840 34620 18846 34672
rect 19242 34620 19248 34672
rect 19300 34660 19306 34672
rect 19300 34632 19472 34660
rect 19300 34620 19306 34632
rect 17346 34595 17404 34601
rect 17346 34592 17358 34595
rect 15887 34564 17358 34592
rect 15887 34561 15899 34564
rect 15841 34555 15899 34561
rect 17346 34561 17358 34564
rect 17392 34561 17404 34595
rect 17346 34555 17404 34561
rect 17865 34595 17923 34601
rect 17865 34561 17877 34595
rect 17911 34561 17923 34595
rect 17865 34555 17923 34561
rect 18325 34595 18383 34601
rect 18325 34561 18337 34595
rect 18371 34561 18383 34595
rect 18506 34592 18512 34604
rect 18467 34564 18512 34592
rect 18325 34555 18383 34561
rect 16206 34524 16212 34536
rect 15764 34496 16212 34524
rect 15657 34487 15715 34493
rect 15470 34416 15476 34468
rect 15528 34456 15534 34468
rect 15672 34456 15700 34487
rect 16206 34484 16212 34496
rect 16264 34484 16270 34536
rect 18340 34524 18368 34555
rect 18506 34552 18512 34564
rect 18564 34552 18570 34604
rect 18601 34595 18659 34601
rect 18601 34561 18613 34595
rect 18647 34594 18659 34595
rect 18647 34592 18724 34594
rect 18800 34592 18828 34620
rect 18647 34566 18828 34592
rect 18647 34561 18659 34566
rect 18696 34564 18828 34566
rect 18601 34555 18659 34561
rect 18874 34552 18880 34604
rect 18932 34592 18938 34604
rect 19061 34595 19119 34601
rect 18932 34564 18977 34592
rect 18932 34552 18938 34564
rect 19061 34561 19073 34595
rect 19107 34592 19119 34595
rect 19334 34592 19340 34604
rect 19107 34564 19340 34592
rect 19107 34561 19119 34564
rect 19061 34555 19119 34561
rect 19334 34552 19340 34564
rect 19392 34552 19398 34604
rect 19444 34602 19472 34632
rect 19610 34620 19616 34672
rect 19668 34660 19674 34672
rect 19792 34660 19820 34700
rect 20162 34688 20168 34740
rect 20220 34728 20226 34740
rect 20993 34731 21051 34737
rect 20993 34728 21005 34731
rect 20220 34700 21005 34728
rect 20220 34688 20226 34700
rect 20993 34697 21005 34700
rect 21039 34728 21051 34731
rect 21818 34728 21824 34740
rect 21039 34700 21824 34728
rect 21039 34697 21051 34700
rect 20993 34691 21051 34697
rect 21818 34688 21824 34700
rect 21876 34688 21882 34740
rect 22557 34731 22615 34737
rect 22557 34697 22569 34731
rect 22603 34728 22615 34731
rect 22646 34728 22652 34740
rect 22603 34700 22652 34728
rect 22603 34697 22615 34700
rect 22557 34691 22615 34697
rect 22646 34688 22652 34700
rect 22704 34688 22710 34740
rect 24670 34728 24676 34740
rect 24631 34700 24676 34728
rect 24670 34688 24676 34700
rect 24728 34688 24734 34740
rect 25317 34731 25375 34737
rect 25317 34697 25329 34731
rect 25363 34697 25375 34731
rect 25317 34691 25375 34697
rect 20257 34663 20315 34669
rect 19668 34632 19748 34660
rect 19792 34632 20199 34660
rect 19668 34620 19674 34632
rect 19518 34602 19524 34604
rect 19444 34574 19524 34602
rect 19518 34552 19524 34574
rect 19576 34592 19582 34604
rect 19720 34601 19748 34632
rect 19705 34595 19763 34601
rect 19576 34564 19621 34592
rect 19576 34552 19582 34564
rect 19705 34561 19717 34595
rect 19751 34561 19763 34595
rect 19705 34555 19763 34561
rect 19794 34552 19800 34604
rect 19852 34592 19858 34604
rect 20056 34595 20114 34601
rect 19852 34564 19897 34592
rect 19852 34552 19858 34564
rect 20056 34561 20068 34595
rect 20102 34561 20114 34595
rect 20171 34594 20199 34632
rect 20257 34629 20269 34663
rect 20303 34660 20315 34663
rect 20438 34660 20444 34672
rect 20303 34632 20444 34660
rect 20303 34629 20315 34632
rect 20257 34623 20315 34629
rect 20438 34620 20444 34632
rect 20496 34620 20502 34672
rect 20530 34620 20536 34672
rect 20588 34660 20594 34672
rect 20588 34632 23060 34660
rect 20588 34620 20594 34632
rect 20901 34595 20959 34601
rect 20171 34592 20208 34594
rect 20171 34566 20300 34592
rect 20180 34564 20300 34566
rect 20056 34555 20114 34561
rect 18693 34527 18751 34533
rect 18340 34496 18414 34524
rect 15528 34428 15700 34456
rect 15528 34416 15534 34428
rect 17862 34416 17868 34468
rect 17920 34456 17926 34468
rect 18386 34456 18414 34496
rect 18693 34493 18705 34527
rect 18739 34524 18751 34527
rect 19150 34524 19156 34536
rect 18739 34496 19156 34524
rect 18739 34493 18751 34496
rect 18693 34487 18751 34493
rect 19150 34484 19156 34496
rect 19208 34524 19214 34536
rect 19889 34527 19947 34533
rect 19208 34496 19748 34524
rect 19208 34484 19214 34496
rect 19242 34456 19248 34468
rect 17920 34428 18414 34456
rect 17920 34416 17926 34428
rect 12894 34388 12900 34400
rect 12855 34360 12900 34388
rect 12894 34348 12900 34360
rect 12952 34348 12958 34400
rect 17773 34391 17831 34397
rect 17773 34357 17785 34391
rect 17819 34388 17831 34391
rect 18138 34388 18144 34400
rect 17819 34360 18144 34388
rect 17819 34357 17831 34360
rect 17773 34351 17831 34357
rect 18138 34348 18144 34360
rect 18196 34348 18202 34400
rect 18386 34388 18414 34428
rect 18800 34428 19248 34456
rect 18800 34388 18828 34428
rect 19242 34416 19248 34428
rect 19300 34416 19306 34468
rect 19720 34456 19748 34496
rect 19889 34493 19901 34527
rect 19935 34493 19947 34527
rect 20071 34524 20099 34555
rect 20162 34524 20168 34536
rect 20071 34496 20168 34524
rect 19889 34487 19947 34493
rect 19904 34456 19932 34487
rect 20162 34484 20168 34496
rect 20220 34484 20226 34536
rect 20272 34524 20300 34564
rect 20901 34561 20913 34595
rect 20947 34592 20959 34595
rect 21174 34592 21180 34604
rect 20947 34564 21180 34592
rect 20947 34561 20959 34564
rect 20901 34555 20959 34561
rect 21174 34552 21180 34564
rect 21232 34552 21238 34604
rect 22370 34592 22376 34604
rect 22331 34564 22376 34592
rect 22370 34552 22376 34564
rect 22428 34552 22434 34604
rect 23032 34601 23060 34632
rect 23017 34595 23075 34601
rect 23017 34561 23029 34595
rect 23063 34561 23075 34595
rect 23842 34592 23848 34604
rect 23755 34564 23848 34592
rect 23017 34555 23075 34561
rect 23842 34552 23848 34564
rect 23900 34592 23906 34604
rect 24026 34592 24032 34604
rect 23900 34564 24032 34592
rect 23900 34552 23906 34564
rect 24026 34552 24032 34564
rect 24084 34552 24090 34604
rect 24486 34592 24492 34604
rect 24447 34564 24492 34592
rect 24486 34552 24492 34564
rect 24544 34552 24550 34604
rect 24854 34552 24860 34604
rect 24912 34592 24918 34604
rect 25133 34595 25191 34601
rect 25133 34592 25145 34595
rect 24912 34564 25145 34592
rect 24912 34552 24918 34564
rect 25133 34561 25145 34564
rect 25179 34561 25191 34595
rect 25332 34592 25360 34691
rect 26602 34688 26608 34740
rect 26660 34728 26666 34740
rect 28442 34728 28448 34740
rect 26660 34700 28304 34728
rect 28403 34700 28448 34728
rect 26660 34688 26666 34700
rect 28276 34660 28304 34700
rect 28442 34688 28448 34700
rect 28500 34688 28506 34740
rect 28994 34728 29000 34740
rect 28552 34700 29000 34728
rect 28552 34660 28580 34700
rect 28994 34688 29000 34700
rect 29052 34688 29058 34740
rect 29454 34688 29460 34740
rect 29512 34728 29518 34740
rect 29549 34731 29607 34737
rect 29549 34728 29561 34731
rect 29512 34700 29561 34728
rect 29512 34688 29518 34700
rect 29549 34697 29561 34700
rect 29595 34697 29607 34731
rect 29549 34691 29607 34697
rect 28276 34632 28580 34660
rect 28718 34620 28724 34672
rect 28776 34660 28782 34672
rect 29365 34663 29423 34669
rect 29365 34660 29377 34663
rect 28776 34632 29377 34660
rect 28776 34620 28782 34632
rect 29365 34629 29377 34632
rect 29411 34629 29423 34663
rect 29365 34623 29423 34629
rect 25777 34595 25835 34601
rect 25777 34592 25789 34595
rect 25332 34564 25789 34592
rect 25133 34555 25191 34561
rect 25777 34561 25789 34564
rect 25823 34561 25835 34595
rect 26970 34592 26976 34604
rect 26931 34564 26976 34592
rect 25777 34555 25835 34561
rect 26970 34552 26976 34564
rect 27028 34552 27034 34604
rect 27801 34595 27859 34601
rect 27801 34561 27813 34595
rect 27847 34592 27859 34595
rect 28166 34592 28172 34604
rect 27847 34564 28172 34592
rect 27847 34561 27859 34564
rect 27801 34555 27859 34561
rect 28166 34552 28172 34564
rect 28224 34552 28230 34604
rect 28261 34595 28319 34601
rect 28261 34561 28273 34595
rect 28307 34592 28319 34595
rect 28350 34592 28356 34604
rect 28307 34564 28356 34592
rect 28307 34561 28319 34564
rect 28261 34555 28319 34561
rect 28350 34552 28356 34564
rect 28408 34552 28414 34604
rect 28997 34595 29055 34601
rect 28997 34561 29009 34595
rect 29043 34592 29055 34595
rect 29086 34592 29092 34604
rect 29043 34564 29092 34592
rect 29043 34561 29055 34564
rect 28997 34555 29055 34561
rect 29086 34552 29092 34564
rect 29144 34552 29150 34604
rect 23109 34527 23167 34533
rect 23109 34524 23121 34527
rect 20272 34496 23121 34524
rect 23109 34493 23121 34496
rect 23155 34493 23167 34527
rect 29822 34524 29828 34536
rect 23109 34487 23167 34493
rect 27632 34496 29828 34524
rect 19720 34428 19932 34456
rect 24029 34459 24087 34465
rect 24029 34425 24041 34459
rect 24075 34456 24087 34459
rect 24302 34456 24308 34468
rect 24075 34428 24308 34456
rect 24075 34425 24087 34428
rect 24029 34419 24087 34425
rect 24302 34416 24308 34428
rect 24360 34456 24366 34468
rect 24670 34456 24676 34468
rect 24360 34428 24676 34456
rect 24360 34416 24366 34428
rect 24670 34416 24676 34428
rect 24728 34416 24734 34468
rect 27632 34465 27660 34496
rect 29822 34484 29828 34496
rect 29880 34484 29886 34536
rect 27617 34459 27675 34465
rect 27617 34425 27629 34459
rect 27663 34425 27675 34459
rect 27617 34419 27675 34425
rect 18386 34360 18828 34388
rect 19518 34348 19524 34400
rect 19576 34388 19582 34400
rect 21450 34388 21456 34400
rect 19576 34360 21456 34388
rect 19576 34348 19582 34360
rect 21450 34348 21456 34360
rect 21508 34348 21514 34400
rect 25222 34348 25228 34400
rect 25280 34388 25286 34400
rect 25961 34391 26019 34397
rect 25961 34388 25973 34391
rect 25280 34360 25973 34388
rect 25280 34348 25286 34360
rect 25961 34357 25973 34360
rect 26007 34357 26019 34391
rect 27154 34388 27160 34400
rect 27115 34360 27160 34388
rect 25961 34351 26019 34357
rect 27154 34348 27160 34360
rect 27212 34348 27218 34400
rect 29270 34348 29276 34400
rect 29328 34388 29334 34400
rect 29365 34391 29423 34397
rect 29365 34388 29377 34391
rect 29328 34360 29377 34388
rect 29328 34348 29334 34360
rect 29365 34357 29377 34360
rect 29411 34357 29423 34391
rect 29365 34351 29423 34357
rect 1104 34298 30820 34320
rect 1104 34246 5915 34298
rect 5967 34246 5979 34298
rect 6031 34246 6043 34298
rect 6095 34246 6107 34298
rect 6159 34246 6171 34298
rect 6223 34246 15846 34298
rect 15898 34246 15910 34298
rect 15962 34246 15974 34298
rect 16026 34246 16038 34298
rect 16090 34246 16102 34298
rect 16154 34246 25776 34298
rect 25828 34246 25840 34298
rect 25892 34246 25904 34298
rect 25956 34246 25968 34298
rect 26020 34246 26032 34298
rect 26084 34246 30820 34298
rect 1104 34224 30820 34246
rect 1394 34144 1400 34196
rect 1452 34184 1458 34196
rect 10965 34187 11023 34193
rect 1452 34156 10272 34184
rect 1452 34144 1458 34156
rect 10244 34048 10272 34156
rect 10965 34153 10977 34187
rect 11011 34184 11023 34187
rect 11514 34184 11520 34196
rect 11011 34156 11520 34184
rect 11011 34153 11023 34156
rect 10965 34147 11023 34153
rect 11514 34144 11520 34156
rect 11572 34144 11578 34196
rect 13170 34184 13176 34196
rect 13131 34156 13176 34184
rect 13170 34144 13176 34156
rect 13228 34144 13234 34196
rect 14829 34187 14887 34193
rect 14829 34153 14841 34187
rect 14875 34184 14887 34187
rect 17770 34184 17776 34196
rect 14875 34156 17776 34184
rect 14875 34153 14887 34156
rect 14829 34147 14887 34153
rect 17770 34144 17776 34156
rect 17828 34144 17834 34196
rect 23658 34184 23664 34196
rect 17880 34156 23664 34184
rect 11425 34119 11483 34125
rect 11425 34085 11437 34119
rect 11471 34116 11483 34119
rect 12250 34116 12256 34128
rect 11471 34088 12256 34116
rect 11471 34085 11483 34088
rect 11425 34079 11483 34085
rect 12250 34076 12256 34088
rect 12308 34076 12314 34128
rect 16666 34076 16672 34128
rect 16724 34116 16730 34128
rect 17880 34116 17908 34156
rect 23658 34144 23664 34156
rect 23716 34144 23722 34196
rect 24486 34144 24492 34196
rect 24544 34184 24550 34196
rect 24765 34187 24823 34193
rect 24765 34184 24777 34187
rect 24544 34156 24777 34184
rect 24544 34144 24550 34156
rect 24765 34153 24777 34156
rect 24811 34153 24823 34187
rect 26602 34184 26608 34196
rect 26563 34156 26608 34184
rect 24765 34147 24823 34153
rect 26602 34144 26608 34156
rect 26660 34144 26666 34196
rect 29270 34144 29276 34196
rect 29328 34184 29334 34196
rect 29914 34184 29920 34196
rect 29328 34156 29920 34184
rect 29328 34144 29334 34156
rect 29914 34144 29920 34156
rect 29972 34144 29978 34196
rect 30098 34184 30104 34196
rect 30059 34156 30104 34184
rect 30098 34144 30104 34156
rect 30156 34144 30162 34196
rect 16724 34088 17908 34116
rect 16724 34076 16730 34088
rect 19150 34076 19156 34128
rect 19208 34076 19214 34128
rect 20717 34119 20775 34125
rect 20717 34085 20729 34119
rect 20763 34085 20775 34119
rect 20717 34079 20775 34085
rect 12069 34051 12127 34057
rect 12069 34048 12081 34051
rect 10244 34020 12081 34048
rect 12069 34017 12081 34020
rect 12115 34017 12127 34051
rect 12069 34011 12127 34017
rect 12437 34051 12495 34057
rect 12437 34017 12449 34051
rect 12483 34048 12495 34051
rect 15378 34048 15384 34060
rect 12483 34020 15240 34048
rect 15339 34020 15384 34048
rect 12483 34017 12495 34020
rect 12437 34011 12495 34017
rect 10137 33983 10195 33989
rect 10137 33949 10149 33983
rect 10183 33980 10195 33983
rect 10226 33980 10232 33992
rect 10183 33952 10232 33980
rect 10183 33949 10195 33952
rect 10137 33943 10195 33949
rect 10226 33940 10232 33952
rect 10284 33940 10290 33992
rect 10321 33983 10379 33989
rect 10321 33949 10333 33983
rect 10367 33980 10379 33983
rect 10594 33980 10600 33992
rect 10367 33952 10600 33980
rect 10367 33949 10379 33952
rect 10321 33943 10379 33949
rect 10594 33940 10600 33952
rect 10652 33940 10658 33992
rect 10781 33983 10839 33989
rect 10781 33949 10793 33983
rect 10827 33980 10839 33983
rect 11238 33980 11244 33992
rect 10827 33952 11244 33980
rect 10827 33949 10839 33952
rect 10781 33943 10839 33949
rect 11238 33940 11244 33952
rect 11296 33940 11302 33992
rect 11609 33983 11667 33989
rect 11609 33949 11621 33983
rect 11655 33949 11667 33983
rect 12250 33980 12256 33992
rect 12211 33952 12256 33980
rect 11609 33943 11667 33949
rect 10042 33872 10048 33924
rect 10100 33912 10106 33924
rect 11624 33912 11652 33943
rect 12250 33940 12256 33952
rect 12308 33940 12314 33992
rect 14737 33983 14795 33989
rect 14737 33949 14749 33983
rect 14783 33980 14795 33983
rect 15102 33980 15108 33992
rect 14783 33952 15108 33980
rect 14783 33949 14795 33952
rect 14737 33943 14795 33949
rect 15102 33940 15108 33952
rect 15160 33940 15166 33992
rect 15212 33980 15240 34020
rect 15378 34008 15384 34020
rect 15436 34008 15442 34060
rect 17770 34008 17776 34060
rect 17828 34048 17834 34060
rect 18230 34048 18236 34060
rect 17828 34020 18092 34048
rect 18191 34020 18236 34048
rect 17828 34008 17834 34020
rect 17313 33983 17371 33989
rect 15212 33952 16804 33980
rect 10100 33884 11652 33912
rect 10100 33872 10106 33884
rect 12710 33872 12716 33924
rect 12768 33912 12774 33924
rect 13081 33915 13139 33921
rect 13081 33912 13093 33915
rect 12768 33884 13093 33912
rect 12768 33872 12774 33884
rect 13081 33881 13093 33884
rect 13127 33881 13139 33915
rect 13081 33875 13139 33881
rect 15648 33915 15706 33921
rect 15648 33881 15660 33915
rect 15694 33912 15706 33915
rect 15838 33912 15844 33924
rect 15694 33884 15844 33912
rect 15694 33881 15706 33884
rect 15648 33875 15706 33881
rect 15838 33872 15844 33884
rect 15896 33872 15902 33924
rect 16666 33912 16672 33924
rect 15948 33884 16672 33912
rect 10226 33844 10232 33856
rect 10187 33816 10232 33844
rect 10226 33804 10232 33816
rect 10284 33804 10290 33856
rect 11514 33804 11520 33856
rect 11572 33844 11578 33856
rect 15948 33844 15976 33884
rect 16666 33872 16672 33884
rect 16724 33872 16730 33924
rect 16776 33912 16804 33952
rect 17313 33949 17325 33983
rect 17359 33980 17371 33983
rect 17678 33980 17684 33992
rect 17359 33952 17684 33980
rect 17359 33949 17371 33952
rect 17313 33943 17371 33949
rect 17678 33940 17684 33952
rect 17736 33940 17742 33992
rect 17862 33940 17868 33992
rect 17920 33980 17926 33992
rect 17957 33983 18015 33989
rect 17957 33980 17969 33983
rect 17920 33952 17969 33980
rect 17920 33940 17926 33952
rect 17957 33949 17969 33952
rect 18003 33949 18015 33983
rect 18064 33980 18092 34020
rect 18230 34008 18236 34020
rect 18288 34008 18294 34060
rect 19168 34048 19196 34076
rect 19705 34051 19763 34057
rect 19705 34048 19717 34051
rect 19168 34020 19717 34048
rect 19705 34017 19717 34020
rect 19751 34017 19763 34051
rect 20732 34048 20760 34079
rect 29086 34076 29092 34128
rect 29144 34116 29150 34128
rect 29549 34119 29607 34125
rect 29549 34116 29561 34119
rect 29144 34088 29561 34116
rect 29144 34076 29150 34088
rect 29549 34085 29561 34088
rect 29595 34085 29607 34119
rect 29549 34079 29607 34085
rect 21177 34051 21235 34057
rect 21177 34048 21189 34051
rect 20732 34020 21189 34048
rect 19705 34011 19763 34017
rect 21177 34017 21189 34020
rect 21223 34017 21235 34051
rect 25222 34048 25228 34060
rect 25183 34020 25228 34048
rect 21177 34011 21235 34017
rect 25222 34008 25228 34020
rect 25280 34008 25286 34060
rect 26878 34008 26884 34060
rect 26936 34048 26942 34060
rect 27433 34051 27491 34057
rect 27433 34048 27445 34051
rect 26936 34020 27445 34048
rect 26936 34008 26942 34020
rect 27433 34017 27445 34020
rect 27479 34017 27491 34051
rect 27433 34011 27491 34017
rect 18141 33983 18199 33989
rect 18141 33980 18153 33983
rect 18064 33952 18153 33980
rect 17957 33943 18015 33949
rect 18141 33949 18153 33952
rect 18187 33949 18199 33983
rect 18141 33943 18199 33949
rect 18322 33940 18328 33992
rect 18380 33989 18386 33992
rect 18380 33983 18429 33989
rect 18380 33949 18383 33983
rect 18417 33949 18429 33983
rect 18380 33943 18429 33949
rect 18509 33983 18567 33989
rect 18509 33949 18521 33983
rect 18555 33980 18567 33983
rect 19153 33983 19211 33989
rect 19153 33980 19165 33983
rect 18555 33952 19165 33980
rect 18555 33949 18567 33952
rect 18509 33943 18567 33949
rect 19153 33949 19165 33952
rect 19199 33949 19211 33983
rect 19153 33943 19211 33949
rect 18380 33940 18386 33943
rect 19242 33940 19248 33992
rect 19300 33980 19306 33992
rect 19337 33983 19395 33989
rect 19337 33980 19349 33983
rect 19300 33952 19349 33980
rect 19300 33940 19306 33952
rect 19337 33949 19349 33952
rect 19383 33949 19395 33983
rect 19518 33980 19524 33992
rect 19479 33952 19524 33980
rect 19337 33943 19395 33949
rect 19518 33940 19524 33952
rect 19576 33940 19582 33992
rect 19613 33983 19671 33989
rect 19613 33949 19625 33983
rect 19659 33980 19671 33983
rect 19794 33980 19800 33992
rect 19659 33952 19800 33980
rect 19659 33949 19671 33952
rect 19613 33943 19671 33949
rect 19794 33940 19800 33952
rect 19852 33940 19858 33992
rect 19889 33983 19947 33989
rect 19889 33949 19901 33983
rect 19935 33980 19947 33983
rect 20438 33980 20444 33992
rect 19935 33952 20444 33980
rect 19935 33949 19947 33952
rect 19889 33943 19947 33949
rect 20438 33940 20444 33952
rect 20496 33940 20502 33992
rect 20533 33983 20591 33989
rect 20533 33949 20545 33983
rect 20579 33980 20591 33983
rect 21266 33980 21272 33992
rect 20579 33952 21272 33980
rect 20579 33949 20591 33952
rect 20533 33943 20591 33949
rect 21266 33940 21272 33952
rect 21324 33940 21330 33992
rect 22278 33940 22284 33992
rect 22336 33980 22342 33992
rect 23017 33983 23075 33989
rect 23017 33980 23029 33983
rect 22336 33952 23029 33980
rect 22336 33940 22342 33952
rect 23017 33949 23029 33952
rect 23063 33949 23075 33983
rect 23017 33943 23075 33949
rect 24581 33983 24639 33989
rect 24581 33949 24593 33983
rect 24627 33980 24639 33983
rect 24854 33980 24860 33992
rect 24627 33952 24860 33980
rect 24627 33949 24639 33952
rect 24581 33943 24639 33949
rect 24854 33940 24860 33952
rect 24912 33940 24918 33992
rect 27062 33980 27068 33992
rect 27023 33952 27068 33980
rect 27062 33940 27068 33952
rect 27120 33940 27126 33992
rect 27249 33983 27307 33989
rect 27249 33949 27261 33983
rect 27295 33949 27307 33983
rect 27249 33943 27307 33949
rect 27341 33983 27399 33989
rect 27341 33949 27353 33983
rect 27387 33949 27399 33983
rect 27341 33943 27399 33949
rect 27617 33983 27675 33989
rect 27617 33949 27629 33983
rect 27663 33980 27675 33983
rect 27663 33952 27936 33980
rect 27663 33949 27675 33952
rect 27617 33943 27675 33949
rect 21450 33921 21456 33924
rect 16776 33884 20208 33912
rect 16758 33844 16764 33856
rect 11572 33816 15976 33844
rect 16719 33816 16764 33844
rect 11572 33804 11578 33816
rect 16758 33804 16764 33816
rect 16816 33804 16822 33856
rect 17405 33847 17463 33853
rect 17405 33813 17417 33847
rect 17451 33844 17463 33847
rect 17586 33844 17592 33856
rect 17451 33816 17592 33844
rect 17451 33813 17463 33816
rect 17405 33807 17463 33813
rect 17586 33804 17592 33816
rect 17644 33804 17650 33856
rect 18506 33804 18512 33856
rect 18564 33844 18570 33856
rect 18693 33847 18751 33853
rect 18693 33844 18705 33847
rect 18564 33816 18705 33844
rect 18564 33804 18570 33816
rect 18693 33813 18705 33816
rect 18739 33813 18751 33847
rect 19242 33844 19248 33856
rect 19203 33816 19248 33844
rect 18693 33807 18751 33813
rect 19242 33804 19248 33816
rect 19300 33804 19306 33856
rect 19334 33804 19340 33856
rect 19392 33844 19398 33856
rect 19610 33844 19616 33856
rect 19392 33816 19616 33844
rect 19392 33804 19398 33816
rect 19610 33804 19616 33816
rect 19668 33804 19674 33856
rect 20070 33844 20076 33856
rect 20031 33816 20076 33844
rect 20070 33804 20076 33816
rect 20128 33804 20134 33856
rect 20180 33844 20208 33884
rect 21444 33875 21456 33921
rect 21508 33912 21514 33924
rect 24394 33912 24400 33924
rect 21508 33884 21544 33912
rect 22066 33884 24400 33912
rect 21450 33872 21456 33875
rect 21508 33872 21514 33884
rect 22066 33844 22094 33884
rect 24394 33872 24400 33884
rect 24452 33912 24458 33924
rect 24946 33912 24952 33924
rect 24452 33884 24952 33912
rect 24452 33872 24458 33884
rect 24946 33872 24952 33884
rect 25004 33872 25010 33924
rect 25492 33915 25550 33921
rect 25492 33881 25504 33915
rect 25538 33912 25550 33915
rect 26142 33912 26148 33924
rect 25538 33884 26148 33912
rect 25538 33881 25550 33884
rect 25492 33875 25550 33881
rect 26142 33872 26148 33884
rect 26200 33872 26206 33924
rect 26326 33872 26332 33924
rect 26384 33912 26390 33924
rect 27264 33912 27292 33943
rect 26384 33884 27292 33912
rect 27356 33912 27384 33943
rect 27430 33912 27436 33924
rect 27356 33884 27436 33912
rect 26384 33872 26390 33884
rect 27430 33872 27436 33884
rect 27488 33872 27494 33924
rect 22554 33844 22560 33856
rect 20180 33816 22094 33844
rect 22515 33816 22560 33844
rect 22554 33804 22560 33816
rect 22612 33804 22618 33856
rect 22738 33804 22744 33856
rect 22796 33844 22802 33856
rect 23201 33847 23259 33853
rect 23201 33844 23213 33847
rect 22796 33816 23213 33844
rect 22796 33804 22802 33816
rect 23201 33813 23213 33816
rect 23247 33813 23259 33847
rect 23201 33807 23259 33813
rect 27614 33804 27620 33856
rect 27672 33844 27678 33856
rect 27801 33847 27859 33853
rect 27801 33844 27813 33847
rect 27672 33816 27813 33844
rect 27672 33804 27678 33816
rect 27801 33813 27813 33816
rect 27847 33813 27859 33847
rect 27908 33844 27936 33952
rect 27982 33940 27988 33992
rect 28040 33980 28046 33992
rect 28721 33983 28779 33989
rect 28721 33980 28733 33983
rect 28040 33952 28733 33980
rect 28040 33940 28046 33952
rect 28721 33949 28733 33952
rect 28767 33949 28779 33983
rect 28721 33943 28779 33949
rect 28626 33872 28632 33924
rect 28684 33912 28690 33924
rect 29917 33915 29975 33921
rect 29917 33912 29929 33915
rect 28684 33884 29929 33912
rect 28684 33872 28690 33884
rect 29917 33881 29929 33884
rect 29963 33881 29975 33915
rect 29917 33875 29975 33881
rect 28718 33844 28724 33856
rect 27908 33816 28724 33844
rect 27801 33807 27859 33813
rect 28718 33804 28724 33816
rect 28776 33804 28782 33856
rect 28902 33844 28908 33856
rect 28863 33816 28908 33844
rect 28902 33804 28908 33816
rect 28960 33804 28966 33856
rect 1104 33754 30820 33776
rect 1104 33702 10880 33754
rect 10932 33702 10944 33754
rect 10996 33702 11008 33754
rect 11060 33702 11072 33754
rect 11124 33702 11136 33754
rect 11188 33702 20811 33754
rect 20863 33702 20875 33754
rect 20927 33702 20939 33754
rect 20991 33702 21003 33754
rect 21055 33702 21067 33754
rect 21119 33702 30820 33754
rect 1104 33680 30820 33702
rect 1394 33640 1400 33652
rect 1355 33612 1400 33640
rect 1394 33600 1400 33612
rect 1452 33600 1458 33652
rect 11422 33600 11428 33652
rect 11480 33640 11486 33652
rect 11793 33643 11851 33649
rect 11793 33640 11805 33643
rect 11480 33612 11805 33640
rect 11480 33600 11486 33612
rect 11793 33609 11805 33612
rect 11839 33609 11851 33643
rect 11793 33603 11851 33609
rect 11882 33600 11888 33652
rect 11940 33640 11946 33652
rect 12710 33640 12716 33652
rect 11940 33612 11985 33640
rect 12671 33612 12716 33640
rect 11940 33600 11946 33612
rect 12710 33600 12716 33612
rect 12768 33600 12774 33652
rect 13998 33640 14004 33652
rect 13188 33612 14004 33640
rect 11514 33572 11520 33584
rect 11475 33544 11520 33572
rect 11514 33532 11520 33544
rect 11572 33532 11578 33584
rect 1578 33504 1584 33516
rect 1539 33476 1584 33504
rect 1578 33464 1584 33476
rect 1636 33464 1642 33516
rect 10045 33507 10103 33513
rect 10045 33473 10057 33507
rect 10091 33504 10103 33507
rect 11333 33507 11391 33513
rect 11333 33504 11345 33507
rect 10091 33476 11345 33504
rect 10091 33473 10103 33476
rect 10045 33467 10103 33473
rect 11333 33473 11345 33476
rect 11379 33473 11391 33507
rect 11333 33467 11391 33473
rect 11701 33507 11759 33513
rect 11701 33473 11713 33507
rect 11747 33473 11759 33507
rect 12066 33504 12072 33516
rect 12027 33476 12072 33504
rect 11701 33467 11759 33473
rect 9950 33396 9956 33448
rect 10008 33436 10014 33448
rect 10137 33439 10195 33445
rect 10137 33436 10149 33439
rect 10008 33408 10149 33436
rect 10008 33396 10014 33408
rect 10137 33405 10149 33408
rect 10183 33405 10195 33439
rect 10137 33399 10195 33405
rect 10229 33439 10287 33445
rect 10229 33405 10241 33439
rect 10275 33405 10287 33439
rect 10229 33399 10287 33405
rect 10244 33368 10272 33399
rect 10318 33396 10324 33448
rect 10376 33436 10382 33448
rect 11716 33436 11744 33467
rect 12066 33464 12072 33476
rect 12124 33464 12130 33516
rect 12621 33507 12679 33513
rect 12621 33473 12633 33507
rect 12667 33473 12679 33507
rect 13188 33504 13216 33612
rect 13998 33600 14004 33612
rect 14056 33600 14062 33652
rect 14550 33600 14556 33652
rect 14608 33640 14614 33652
rect 17770 33640 17776 33652
rect 14608 33612 17776 33640
rect 14608 33600 14614 33612
rect 17770 33600 17776 33612
rect 17828 33640 17834 33652
rect 19337 33643 19395 33649
rect 19337 33640 19349 33643
rect 17828 33612 19349 33640
rect 17828 33600 17834 33612
rect 19337 33609 19349 33612
rect 19383 33609 19395 33643
rect 19337 33603 19395 33609
rect 19702 33600 19708 33652
rect 19760 33640 19766 33652
rect 20254 33640 20260 33652
rect 19760 33612 20260 33640
rect 19760 33600 19766 33612
rect 20254 33600 20260 33612
rect 20312 33600 20318 33652
rect 21269 33643 21327 33649
rect 21269 33609 21281 33643
rect 21315 33640 21327 33643
rect 21450 33640 21456 33652
rect 21315 33612 21456 33640
rect 21315 33609 21327 33612
rect 21269 33603 21327 33609
rect 21450 33600 21456 33612
rect 21508 33600 21514 33652
rect 22278 33640 22284 33652
rect 22239 33612 22284 33640
rect 22278 33600 22284 33612
rect 22336 33600 22342 33652
rect 26142 33640 26148 33652
rect 26103 33612 26148 33640
rect 26142 33600 26148 33612
rect 26200 33600 26206 33652
rect 27430 33640 27436 33652
rect 26243 33612 27436 33640
rect 15102 33572 15108 33584
rect 13372 33544 15108 33572
rect 13265 33507 13323 33513
rect 13265 33504 13277 33507
rect 13188 33476 13277 33504
rect 12621 33467 12679 33473
rect 13265 33473 13277 33476
rect 13311 33473 13323 33507
rect 13265 33467 13323 33473
rect 10376 33408 11744 33436
rect 12636 33436 12664 33467
rect 13372 33436 13400 33544
rect 15102 33532 15108 33544
rect 15160 33532 15166 33584
rect 15286 33532 15292 33584
rect 15344 33532 15350 33584
rect 16758 33572 16764 33584
rect 15580 33544 16764 33572
rect 13909 33507 13967 33513
rect 13909 33504 13921 33507
rect 12636 33408 13400 33436
rect 13464 33476 13921 33504
rect 10376 33396 10382 33408
rect 10686 33368 10692 33380
rect 10244 33340 10692 33368
rect 10686 33328 10692 33340
rect 10744 33328 10750 33380
rect 11333 33371 11391 33377
rect 11333 33337 11345 33371
rect 11379 33368 11391 33371
rect 13354 33368 13360 33380
rect 11379 33340 13360 33368
rect 11379 33337 11391 33340
rect 11333 33331 11391 33337
rect 13354 33328 13360 33340
rect 13412 33328 13418 33380
rect 13464 33377 13492 33476
rect 13909 33473 13921 33476
rect 13955 33473 13967 33507
rect 15010 33504 15016 33516
rect 14971 33476 15016 33504
rect 13909 33467 13967 33473
rect 15010 33464 15016 33476
rect 15068 33464 15074 33516
rect 15197 33507 15255 33513
rect 15197 33473 15209 33507
rect 15243 33504 15255 33507
rect 15304 33504 15332 33532
rect 15243 33476 15332 33504
rect 15381 33507 15439 33513
rect 15243 33473 15255 33476
rect 15197 33467 15255 33473
rect 15381 33473 15393 33507
rect 15427 33504 15439 33507
rect 15470 33504 15476 33516
rect 15427 33476 15476 33504
rect 15427 33473 15439 33476
rect 15381 33467 15439 33473
rect 15470 33464 15476 33476
rect 15528 33464 15534 33516
rect 15580 33513 15608 33544
rect 16758 33532 16764 33544
rect 16816 33532 16822 33584
rect 22186 33572 22192 33584
rect 21100 33544 22192 33572
rect 15565 33507 15623 33513
rect 15565 33473 15577 33507
rect 15611 33473 15623 33507
rect 15565 33467 15623 33473
rect 15749 33507 15807 33513
rect 15749 33473 15761 33507
rect 15795 33504 15807 33507
rect 15838 33504 15844 33516
rect 15795 33476 15844 33504
rect 15795 33473 15807 33476
rect 15749 33467 15807 33473
rect 15838 33464 15844 33476
rect 15896 33464 15902 33516
rect 16669 33507 16727 33513
rect 16669 33473 16681 33507
rect 16715 33473 16727 33507
rect 16850 33504 16856 33516
rect 16811 33476 16856 33504
rect 16669 33467 16727 33473
rect 13449 33371 13507 33377
rect 13449 33337 13461 33371
rect 13495 33337 13507 33371
rect 13449 33331 13507 33337
rect 14458 33328 14464 33380
rect 14516 33368 14522 33380
rect 15028 33368 15056 33464
rect 15286 33436 15292 33448
rect 15247 33408 15292 33436
rect 15286 33396 15292 33408
rect 15344 33396 15350 33448
rect 16684 33368 16712 33467
rect 16850 33464 16856 33476
rect 16908 33464 16914 33516
rect 17221 33507 17279 33513
rect 17221 33473 17233 33507
rect 17267 33504 17279 33507
rect 17770 33504 17776 33516
rect 17267 33476 17776 33504
rect 17267 33473 17279 33476
rect 17221 33467 17279 33473
rect 17770 33464 17776 33476
rect 17828 33464 17834 33516
rect 17954 33504 17960 33516
rect 17915 33476 17960 33504
rect 17954 33464 17960 33476
rect 18012 33464 18018 33516
rect 18233 33507 18291 33513
rect 18233 33473 18245 33507
rect 18279 33504 18291 33507
rect 18506 33504 18512 33516
rect 18279 33476 18512 33504
rect 18279 33473 18291 33476
rect 18233 33467 18291 33473
rect 18506 33464 18512 33476
rect 18564 33464 18570 33516
rect 19702 33464 19708 33516
rect 19760 33504 19766 33516
rect 20533 33507 20591 33513
rect 20533 33504 20545 33507
rect 19760 33476 20545 33504
rect 19760 33464 19766 33476
rect 20533 33473 20545 33476
rect 20579 33473 20591 33507
rect 20714 33504 20720 33516
rect 20675 33476 20720 33504
rect 20533 33467 20591 33473
rect 20714 33464 20720 33476
rect 20772 33464 20778 33516
rect 20806 33464 20812 33516
rect 20864 33504 20870 33516
rect 21100 33513 21128 33544
rect 22186 33532 22192 33544
rect 22244 33572 22250 33584
rect 22554 33572 22560 33584
rect 22244 33544 22560 33572
rect 22244 33532 22250 33544
rect 22554 33532 22560 33544
rect 22612 33532 22618 33584
rect 26243 33572 26271 33612
rect 27430 33600 27436 33612
rect 27488 33600 27494 33652
rect 27706 33640 27712 33652
rect 27632 33612 27712 33640
rect 25700 33544 26271 33572
rect 21085 33507 21143 33513
rect 20864 33476 20909 33504
rect 20864 33464 20870 33476
rect 21085 33473 21097 33507
rect 21131 33473 21143 33507
rect 21085 33467 21143 33473
rect 22094 33464 22100 33516
rect 22152 33504 22158 33516
rect 22738 33504 22744 33516
rect 22152 33476 22197 33504
rect 22699 33476 22744 33504
rect 22152 33464 22158 33476
rect 22738 33464 22744 33476
rect 22796 33464 22802 33516
rect 22830 33464 22836 33516
rect 22888 33504 22894 33516
rect 22997 33507 23055 33513
rect 22997 33504 23009 33507
rect 22888 33476 23009 33504
rect 22888 33464 22894 33476
rect 22997 33473 23009 33476
rect 23043 33473 23055 33507
rect 22997 33467 23055 33473
rect 23566 33464 23572 33516
rect 23624 33504 23630 33516
rect 24581 33507 24639 33513
rect 24581 33504 24593 33507
rect 23624 33476 24593 33504
rect 23624 33464 23630 33476
rect 24581 33473 24593 33476
rect 24627 33473 24639 33507
rect 24581 33467 24639 33473
rect 24670 33464 24676 33516
rect 24728 33504 24734 33516
rect 25409 33507 25467 33513
rect 25409 33504 25421 33507
rect 24728 33476 25421 33504
rect 24728 33464 24734 33476
rect 25409 33473 25421 33476
rect 25455 33473 25467 33507
rect 25409 33467 25467 33473
rect 25498 33464 25504 33516
rect 25556 33504 25562 33516
rect 25700 33513 25728 33544
rect 25593 33507 25651 33513
rect 25593 33504 25605 33507
rect 25556 33476 25605 33504
rect 25556 33464 25562 33476
rect 25593 33473 25605 33476
rect 25639 33473 25651 33507
rect 25593 33467 25651 33473
rect 25685 33507 25743 33513
rect 25685 33473 25697 33507
rect 25731 33473 25743 33507
rect 25685 33467 25743 33473
rect 25961 33507 26019 33513
rect 25961 33473 25973 33507
rect 26007 33504 26019 33507
rect 26602 33504 26608 33516
rect 26007 33476 26608 33504
rect 26007 33473 26019 33476
rect 25961 33467 26019 33473
rect 26602 33464 26608 33476
rect 26660 33464 26666 33516
rect 27249 33507 27307 33513
rect 27249 33504 27261 33507
rect 27172 33476 27261 33504
rect 16945 33439 17003 33445
rect 16945 33405 16957 33439
rect 16991 33405 17003 33439
rect 16945 33399 17003 33405
rect 17037 33439 17095 33445
rect 17037 33405 17049 33439
rect 17083 33436 17095 33439
rect 17678 33436 17684 33448
rect 17083 33408 17684 33436
rect 17083 33405 17095 33408
rect 17037 33399 17095 33405
rect 14516 33340 16712 33368
rect 16960 33368 16988 33399
rect 17678 33396 17684 33408
rect 17736 33396 17742 33448
rect 20901 33439 20959 33445
rect 20901 33405 20913 33439
rect 20947 33436 20959 33439
rect 22554 33436 22560 33448
rect 20947 33408 22560 33436
rect 20947 33405 20959 33408
rect 20901 33399 20959 33405
rect 22554 33396 22560 33408
rect 22612 33396 22618 33448
rect 25777 33439 25835 33445
rect 25777 33405 25789 33439
rect 25823 33436 25835 33439
rect 26878 33436 26884 33448
rect 25823 33408 26884 33436
rect 25823 33405 25835 33408
rect 25777 33399 25835 33405
rect 26878 33396 26884 33408
rect 26936 33396 26942 33448
rect 17862 33368 17868 33380
rect 16960 33340 17868 33368
rect 14516 33328 14522 33340
rect 9674 33300 9680 33312
rect 9635 33272 9680 33300
rect 9674 33260 9680 33272
rect 9732 33260 9738 33312
rect 12250 33260 12256 33312
rect 12308 33300 12314 33312
rect 12710 33300 12716 33312
rect 12308 33272 12716 33300
rect 12308 33260 12314 33272
rect 12710 33260 12716 33272
rect 12768 33260 12774 33312
rect 13262 33260 13268 33312
rect 13320 33300 13326 33312
rect 14093 33303 14151 33309
rect 14093 33300 14105 33303
rect 13320 33272 14105 33300
rect 13320 33260 13326 33272
rect 14093 33269 14105 33272
rect 14139 33269 14151 33303
rect 14093 33263 14151 33269
rect 15286 33260 15292 33312
rect 15344 33300 15350 33312
rect 16206 33300 16212 33312
rect 15344 33272 16212 33300
rect 15344 33260 15350 33272
rect 16206 33260 16212 33272
rect 16264 33300 16270 33312
rect 16960 33300 16988 33340
rect 17862 33328 17868 33340
rect 17920 33328 17926 33380
rect 17402 33300 17408 33312
rect 16264 33272 16988 33300
rect 17363 33272 17408 33300
rect 16264 33260 16270 33272
rect 17402 33260 17408 33272
rect 17460 33260 17466 33312
rect 24121 33303 24179 33309
rect 24121 33269 24133 33303
rect 24167 33300 24179 33303
rect 24394 33300 24400 33312
rect 24167 33272 24400 33300
rect 24167 33269 24179 33272
rect 24121 33263 24179 33269
rect 24394 33260 24400 33272
rect 24452 33260 24458 33312
rect 24765 33303 24823 33309
rect 24765 33269 24777 33303
rect 24811 33300 24823 33303
rect 24854 33300 24860 33312
rect 24811 33272 24860 33300
rect 24811 33269 24823 33272
rect 24765 33263 24823 33269
rect 24854 33260 24860 33272
rect 24912 33300 24918 33312
rect 25590 33300 25596 33312
rect 24912 33272 25596 33300
rect 24912 33260 24918 33272
rect 25590 33260 25596 33272
rect 25648 33260 25654 33312
rect 27172 33300 27200 33476
rect 27249 33473 27261 33476
rect 27295 33473 27307 33507
rect 27249 33467 27307 33473
rect 27516 33507 27574 33513
rect 27516 33473 27528 33507
rect 27562 33504 27574 33507
rect 27632 33504 27660 33612
rect 27706 33600 27712 33612
rect 27764 33600 27770 33652
rect 28626 33640 28632 33652
rect 28587 33612 28632 33640
rect 28626 33600 28632 33612
rect 28684 33600 28690 33652
rect 27562 33476 27660 33504
rect 27562 33473 27574 33476
rect 27516 33467 27574 33473
rect 27798 33464 27804 33516
rect 27856 33504 27862 33516
rect 29089 33507 29147 33513
rect 29089 33504 29101 33507
rect 27856 33476 29101 33504
rect 27856 33464 27862 33476
rect 29089 33473 29101 33476
rect 29135 33473 29147 33507
rect 29822 33504 29828 33516
rect 29783 33476 29828 33504
rect 29089 33467 29147 33473
rect 29822 33464 29828 33476
rect 29880 33464 29886 33516
rect 29273 33303 29331 33309
rect 29273 33300 29285 33303
rect 27172 33272 29285 33300
rect 29273 33269 29285 33272
rect 29319 33269 29331 33303
rect 30006 33300 30012 33312
rect 29967 33272 30012 33300
rect 29273 33263 29331 33269
rect 30006 33260 30012 33272
rect 30064 33260 30070 33312
rect 1104 33210 30820 33232
rect 1104 33158 5915 33210
rect 5967 33158 5979 33210
rect 6031 33158 6043 33210
rect 6095 33158 6107 33210
rect 6159 33158 6171 33210
rect 6223 33158 15846 33210
rect 15898 33158 15910 33210
rect 15962 33158 15974 33210
rect 16026 33158 16038 33210
rect 16090 33158 16102 33210
rect 16154 33158 25776 33210
rect 25828 33158 25840 33210
rect 25892 33158 25904 33210
rect 25956 33158 25968 33210
rect 26020 33158 26032 33210
rect 26084 33158 30820 33210
rect 1104 33136 30820 33158
rect 9950 33096 9956 33108
rect 9911 33068 9956 33096
rect 9950 33056 9956 33068
rect 10008 33056 10014 33108
rect 16298 33096 16304 33108
rect 11164 33068 16304 33096
rect 9401 33031 9459 33037
rect 9401 32997 9413 33031
rect 9447 33028 9459 33031
rect 10318 33028 10324 33040
rect 9447 33000 10324 33028
rect 9447 32997 9459 33000
rect 9401 32991 9459 32997
rect 10318 32988 10324 33000
rect 10376 32988 10382 33040
rect 11164 33037 11192 33068
rect 16298 33056 16304 33068
rect 16356 33056 16362 33108
rect 16666 33056 16672 33108
rect 16724 33096 16730 33108
rect 17126 33096 17132 33108
rect 16724 33068 17132 33096
rect 16724 33056 16730 33068
rect 17126 33056 17132 33068
rect 17184 33056 17190 33108
rect 17770 33096 17776 33108
rect 17731 33068 17776 33096
rect 17770 33056 17776 33068
rect 17828 33056 17834 33108
rect 22005 33099 22063 33105
rect 22005 33065 22017 33099
rect 22051 33065 22063 33099
rect 22005 33059 22063 33065
rect 26513 33099 26571 33105
rect 26513 33065 26525 33099
rect 26559 33096 26571 33099
rect 26970 33096 26976 33108
rect 26559 33068 26976 33096
rect 26559 33065 26571 33068
rect 26513 33059 26571 33065
rect 11149 33031 11207 33037
rect 11149 32997 11161 33031
rect 11195 32997 11207 33031
rect 11149 32991 11207 32997
rect 17954 32920 17960 32972
rect 18012 32960 18018 32972
rect 19242 32960 19248 32972
rect 18012 32932 19248 32960
rect 18012 32920 18018 32932
rect 19242 32920 19248 32932
rect 19300 32960 19306 32972
rect 19521 32963 19579 32969
rect 19521 32960 19533 32963
rect 19300 32932 19533 32960
rect 19300 32920 19306 32932
rect 19521 32929 19533 32932
rect 19567 32929 19579 32963
rect 22020 32960 22048 33059
rect 26970 33056 26976 33068
rect 27028 33056 27034 33108
rect 28258 33096 28264 33108
rect 27264 33068 28264 33096
rect 24762 32988 24768 33040
rect 24820 33028 24826 33040
rect 27264 33028 27292 33068
rect 28258 33056 28264 33068
rect 28316 33096 28322 33108
rect 28442 33096 28448 33108
rect 28316 33068 28448 33096
rect 28316 33056 28322 33068
rect 28442 33056 28448 33068
rect 28500 33056 28506 33108
rect 28629 33099 28687 33105
rect 28629 33065 28641 33099
rect 28675 33096 28687 33099
rect 28718 33096 28724 33108
rect 28675 33068 28724 33096
rect 28675 33065 28687 33068
rect 28629 33059 28687 33065
rect 28718 33056 28724 33068
rect 28776 33056 28782 33108
rect 24820 33000 27292 33028
rect 24820 32988 24826 33000
rect 22465 32963 22523 32969
rect 22465 32960 22477 32963
rect 22020 32932 22477 32960
rect 19521 32923 19579 32929
rect 22465 32929 22477 32932
rect 22511 32929 22523 32963
rect 22465 32923 22523 32929
rect 25041 32963 25099 32969
rect 25041 32929 25053 32963
rect 25087 32960 25099 32963
rect 25130 32960 25136 32972
rect 25087 32932 25136 32960
rect 25087 32929 25099 32932
rect 25041 32923 25099 32929
rect 25130 32920 25136 32932
rect 25188 32920 25194 32972
rect 25332 32969 25360 33000
rect 25317 32963 25375 32969
rect 25317 32929 25329 32963
rect 25363 32929 25375 32963
rect 25317 32923 25375 32929
rect 26234 32920 26240 32972
rect 26292 32960 26298 32972
rect 26510 32960 26516 32972
rect 26292 32932 26516 32960
rect 26292 32920 26298 32932
rect 26510 32920 26516 32932
rect 26568 32920 26574 32972
rect 27154 32920 27160 32972
rect 27212 32960 27218 32972
rect 27249 32963 27307 32969
rect 27249 32960 27261 32963
rect 27212 32932 27261 32960
rect 27212 32920 27218 32932
rect 27249 32929 27261 32932
rect 27295 32929 27307 32963
rect 27249 32923 27307 32929
rect 9309 32895 9367 32901
rect 9309 32861 9321 32895
rect 9355 32861 9367 32895
rect 9309 32855 9367 32861
rect 9493 32895 9551 32901
rect 9493 32861 9505 32895
rect 9539 32892 9551 32895
rect 9950 32892 9956 32904
rect 9539 32864 9956 32892
rect 9539 32861 9551 32864
rect 9493 32855 9551 32861
rect 9324 32824 9352 32855
rect 9950 32852 9956 32864
rect 10008 32852 10014 32904
rect 10137 32895 10195 32901
rect 10137 32861 10149 32895
rect 10183 32892 10195 32895
rect 10226 32892 10232 32904
rect 10183 32864 10232 32892
rect 10183 32861 10195 32864
rect 10137 32855 10195 32861
rect 10152 32824 10180 32855
rect 10226 32852 10232 32864
rect 10284 32852 10290 32904
rect 10410 32852 10416 32904
rect 10468 32892 10474 32904
rect 11238 32892 11244 32904
rect 10468 32864 11244 32892
rect 10468 32852 10474 32864
rect 11238 32852 11244 32864
rect 11296 32852 11302 32904
rect 11698 32892 11704 32904
rect 11611 32864 11704 32892
rect 11698 32852 11704 32864
rect 11756 32892 11762 32904
rect 12066 32892 12072 32904
rect 11756 32864 12072 32892
rect 11756 32852 11762 32864
rect 12066 32852 12072 32864
rect 12124 32852 12130 32904
rect 12161 32895 12219 32901
rect 12161 32861 12173 32895
rect 12207 32892 12219 32895
rect 13262 32892 13268 32904
rect 12207 32864 13268 32892
rect 12207 32861 12219 32864
rect 12161 32855 12219 32861
rect 13262 32852 13268 32864
rect 13320 32852 13326 32904
rect 14182 32892 14188 32904
rect 14143 32864 14188 32892
rect 14182 32852 14188 32864
rect 14240 32852 14246 32904
rect 16393 32895 16451 32901
rect 16393 32861 16405 32895
rect 16439 32892 16451 32895
rect 17972 32892 18000 32920
rect 16439 32864 18000 32892
rect 18233 32895 18291 32901
rect 16439 32861 16451 32864
rect 16393 32855 16451 32861
rect 18233 32861 18245 32895
rect 18279 32861 18291 32895
rect 18233 32855 18291 32861
rect 11330 32824 11336 32836
rect 9324 32796 10180 32824
rect 11291 32796 11336 32824
rect 11330 32784 11336 32796
rect 11388 32784 11394 32836
rect 12428 32827 12486 32833
rect 12428 32793 12440 32827
rect 12474 32824 12486 32827
rect 12986 32824 12992 32836
rect 12474 32796 12992 32824
rect 12474 32793 12486 32796
rect 12428 32787 12486 32793
rect 12986 32784 12992 32796
rect 13044 32784 13050 32836
rect 14452 32827 14510 32833
rect 14452 32793 14464 32827
rect 14498 32824 14510 32827
rect 15194 32824 15200 32836
rect 14498 32796 15200 32824
rect 14498 32793 14510 32796
rect 14452 32787 14510 32793
rect 15194 32784 15200 32796
rect 15252 32784 15258 32836
rect 16660 32827 16718 32833
rect 16660 32793 16672 32827
rect 16706 32824 16718 32827
rect 17402 32824 17408 32836
rect 16706 32796 17408 32824
rect 16706 32793 16718 32796
rect 16660 32787 16718 32793
rect 17402 32784 17408 32796
rect 17460 32784 17466 32836
rect 18248 32824 18276 32855
rect 19610 32852 19616 32904
rect 19668 32892 19674 32904
rect 19777 32895 19835 32901
rect 19777 32892 19789 32895
rect 19668 32864 19789 32892
rect 19668 32852 19674 32864
rect 19777 32861 19789 32864
rect 19823 32861 19835 32895
rect 19777 32855 19835 32861
rect 21821 32895 21879 32901
rect 21821 32861 21833 32895
rect 21867 32892 21879 32895
rect 23474 32892 23480 32904
rect 21867 32864 23480 32892
rect 21867 32861 21879 32864
rect 21821 32855 21879 32861
rect 23474 32852 23480 32864
rect 23532 32852 23538 32904
rect 24581 32895 24639 32901
rect 24581 32861 24593 32895
rect 24627 32892 24639 32895
rect 24854 32892 24860 32904
rect 24627 32864 24860 32892
rect 24627 32861 24639 32864
rect 24581 32855 24639 32861
rect 24854 32852 24860 32864
rect 24912 32852 24918 32904
rect 26142 32852 26148 32904
rect 26200 32892 26206 32904
rect 26329 32895 26387 32901
rect 26329 32892 26341 32895
rect 26200 32864 26341 32892
rect 26200 32852 26206 32864
rect 26329 32861 26341 32864
rect 26375 32861 26387 32895
rect 26329 32855 26387 32861
rect 28258 32852 28264 32904
rect 28316 32892 28322 32904
rect 29825 32895 29883 32901
rect 29825 32892 29837 32895
rect 28316 32864 29837 32892
rect 28316 32852 28322 32864
rect 29825 32861 29837 32864
rect 29871 32861 29883 32895
rect 29825 32855 29883 32861
rect 17512 32796 18276 32824
rect 10321 32759 10379 32765
rect 10321 32725 10333 32759
rect 10367 32756 10379 32759
rect 10594 32756 10600 32768
rect 10367 32728 10600 32756
rect 10367 32725 10379 32728
rect 10321 32719 10379 32725
rect 10594 32716 10600 32728
rect 10652 32716 10658 32768
rect 11422 32756 11428 32768
rect 11383 32728 11428 32756
rect 11422 32716 11428 32728
rect 11480 32716 11486 32768
rect 11517 32759 11575 32765
rect 11517 32725 11529 32759
rect 11563 32756 11575 32759
rect 11882 32756 11888 32768
rect 11563 32728 11888 32756
rect 11563 32725 11575 32728
rect 11517 32719 11575 32725
rect 11882 32716 11888 32728
rect 11940 32716 11946 32768
rect 12802 32716 12808 32768
rect 12860 32756 12866 32768
rect 13541 32759 13599 32765
rect 13541 32756 13553 32759
rect 12860 32728 13553 32756
rect 12860 32716 12866 32728
rect 13541 32725 13553 32728
rect 13587 32725 13599 32759
rect 13541 32719 13599 32725
rect 15010 32716 15016 32768
rect 15068 32756 15074 32768
rect 15565 32759 15623 32765
rect 15565 32756 15577 32759
rect 15068 32728 15577 32756
rect 15068 32716 15074 32728
rect 15565 32725 15577 32728
rect 15611 32725 15623 32759
rect 15565 32719 15623 32725
rect 16758 32716 16764 32768
rect 16816 32756 16822 32768
rect 17512 32756 17540 32796
rect 20714 32784 20720 32836
rect 20772 32824 20778 32836
rect 21358 32824 21364 32836
rect 20772 32796 21364 32824
rect 20772 32784 20778 32796
rect 21358 32784 21364 32796
rect 21416 32784 21422 32836
rect 22732 32827 22790 32833
rect 22732 32793 22744 32827
rect 22778 32824 22790 32827
rect 23106 32824 23112 32836
rect 22778 32796 23112 32824
rect 22778 32793 22790 32796
rect 22732 32787 22790 32793
rect 23106 32784 23112 32796
rect 23164 32784 23170 32836
rect 27516 32827 27574 32833
rect 27516 32793 27528 32827
rect 27562 32824 27574 32827
rect 27614 32824 27620 32836
rect 27562 32796 27620 32824
rect 27562 32793 27574 32796
rect 27516 32787 27574 32793
rect 27614 32784 27620 32796
rect 27672 32784 27678 32836
rect 16816 32728 17540 32756
rect 16816 32716 16822 32728
rect 17954 32716 17960 32768
rect 18012 32756 18018 32768
rect 18325 32759 18383 32765
rect 18325 32756 18337 32759
rect 18012 32728 18337 32756
rect 18012 32716 18018 32728
rect 18325 32725 18337 32728
rect 18371 32725 18383 32759
rect 18325 32719 18383 32725
rect 18874 32716 18880 32768
rect 18932 32756 18938 32768
rect 20901 32759 20959 32765
rect 20901 32756 20913 32759
rect 18932 32728 20913 32756
rect 18932 32716 18938 32728
rect 20901 32725 20913 32728
rect 20947 32725 20959 32759
rect 20901 32719 20959 32725
rect 23382 32716 23388 32768
rect 23440 32756 23446 32768
rect 23845 32759 23903 32765
rect 23845 32756 23857 32759
rect 23440 32728 23857 32756
rect 23440 32716 23446 32728
rect 23845 32725 23857 32728
rect 23891 32725 23903 32759
rect 23845 32719 23903 32725
rect 24397 32759 24455 32765
rect 24397 32725 24409 32759
rect 24443 32756 24455 32759
rect 25222 32756 25228 32768
rect 24443 32728 25228 32756
rect 24443 32725 24455 32728
rect 24397 32719 24455 32725
rect 25222 32716 25228 32728
rect 25280 32716 25286 32768
rect 30009 32759 30067 32765
rect 30009 32725 30021 32759
rect 30055 32756 30067 32759
rect 30098 32756 30104 32768
rect 30055 32728 30104 32756
rect 30055 32725 30067 32728
rect 30009 32719 30067 32725
rect 30098 32716 30104 32728
rect 30156 32716 30162 32768
rect 1104 32666 30820 32688
rect 1104 32614 10880 32666
rect 10932 32614 10944 32666
rect 10996 32614 11008 32666
rect 11060 32614 11072 32666
rect 11124 32614 11136 32666
rect 11188 32614 20811 32666
rect 20863 32614 20875 32666
rect 20927 32614 20939 32666
rect 20991 32614 21003 32666
rect 21055 32614 21067 32666
rect 21119 32614 30820 32666
rect 1104 32592 30820 32614
rect 11698 32552 11704 32564
rect 11659 32524 11704 32552
rect 11698 32512 11704 32524
rect 11756 32512 11762 32564
rect 12986 32552 12992 32564
rect 12947 32524 12992 32552
rect 12986 32512 12992 32524
rect 13044 32512 13050 32564
rect 15102 32512 15108 32564
rect 15160 32552 15166 32564
rect 17221 32555 17279 32561
rect 17221 32552 17233 32555
rect 15160 32524 17233 32552
rect 15160 32512 15166 32524
rect 17221 32521 17233 32524
rect 17267 32552 17279 32555
rect 20714 32552 20720 32564
rect 17267 32524 20720 32552
rect 17267 32521 17279 32524
rect 17221 32515 17279 32521
rect 20714 32512 20720 32524
rect 20772 32512 20778 32564
rect 21266 32552 21272 32564
rect 21227 32524 21272 32552
rect 21266 32512 21272 32524
rect 21324 32512 21330 32564
rect 22094 32552 22100 32564
rect 22066 32512 22100 32552
rect 22152 32512 22158 32564
rect 22830 32552 22836 32564
rect 22791 32524 22836 32552
rect 22830 32512 22836 32524
rect 22888 32512 22894 32564
rect 23474 32552 23480 32564
rect 23435 32524 23480 32552
rect 23474 32512 23480 32524
rect 23532 32512 23538 32564
rect 26421 32555 26479 32561
rect 26421 32521 26433 32555
rect 26467 32552 26479 32555
rect 27798 32552 27804 32564
rect 26467 32524 27804 32552
rect 26467 32521 26479 32524
rect 26421 32515 26479 32521
rect 27798 32512 27804 32524
rect 27856 32512 27862 32564
rect 28166 32512 28172 32564
rect 28224 32552 28230 32564
rect 29457 32555 29515 32561
rect 29457 32552 29469 32555
rect 28224 32524 29469 32552
rect 28224 32512 28230 32524
rect 29457 32521 29469 32524
rect 29503 32521 29515 32555
rect 29457 32515 29515 32521
rect 10229 32487 10287 32493
rect 10229 32453 10241 32487
rect 10275 32484 10287 32487
rect 13446 32484 13452 32496
rect 10275 32456 13452 32484
rect 10275 32453 10287 32456
rect 10229 32447 10287 32453
rect 13446 32444 13452 32456
rect 13504 32444 13510 32496
rect 13998 32444 14004 32496
rect 14056 32484 14062 32496
rect 22066 32484 22094 32512
rect 23198 32484 23204 32496
rect 14056 32456 23204 32484
rect 14056 32444 14062 32456
rect 11609 32419 11667 32425
rect 11609 32385 11621 32419
rect 11655 32416 11667 32419
rect 11790 32416 11796 32428
rect 11655 32388 11796 32416
rect 11655 32385 11667 32388
rect 11609 32379 11667 32385
rect 11790 32376 11796 32388
rect 11848 32376 11854 32428
rect 12253 32419 12311 32425
rect 12253 32385 12265 32419
rect 12299 32416 12311 32419
rect 12342 32416 12348 32428
rect 12299 32388 12348 32416
rect 12299 32385 12311 32388
rect 12253 32379 12311 32385
rect 12342 32376 12348 32388
rect 12400 32376 12406 32428
rect 12434 32376 12440 32428
rect 12492 32416 12498 32428
rect 12621 32419 12679 32425
rect 12492 32388 12537 32416
rect 12492 32376 12498 32388
rect 12621 32385 12633 32419
rect 12667 32385 12679 32419
rect 12802 32416 12808 32428
rect 12763 32388 12808 32416
rect 12621 32379 12679 32385
rect 10318 32348 10324 32360
rect 10279 32320 10324 32348
rect 10318 32308 10324 32320
rect 10376 32308 10382 32360
rect 10505 32351 10563 32357
rect 10505 32317 10517 32351
rect 10551 32348 10563 32351
rect 10686 32348 10692 32360
rect 10551 32320 10692 32348
rect 10551 32317 10563 32320
rect 10505 32311 10563 32317
rect 10686 32308 10692 32320
rect 10744 32308 10750 32360
rect 11514 32308 11520 32360
rect 11572 32348 11578 32360
rect 12529 32351 12587 32357
rect 12529 32348 12541 32351
rect 11572 32320 12541 32348
rect 11572 32308 11578 32320
rect 12529 32317 12541 32320
rect 12575 32317 12587 32351
rect 12636 32348 12664 32379
rect 12802 32376 12808 32388
rect 12860 32376 12866 32428
rect 13354 32376 13360 32428
rect 13412 32416 13418 32428
rect 13541 32419 13599 32425
rect 13541 32416 13553 32419
rect 13412 32388 13553 32416
rect 13412 32376 13418 32388
rect 13541 32385 13553 32388
rect 13587 32385 13599 32419
rect 14458 32416 14464 32428
rect 14419 32388 14464 32416
rect 13541 32379 13599 32385
rect 12636 32320 12747 32348
rect 12529 32311 12587 32317
rect 10704 32280 10732 32308
rect 12618 32280 12624 32292
rect 10704 32252 12624 32280
rect 12618 32240 12624 32252
rect 12676 32280 12682 32292
rect 12719 32280 12747 32320
rect 12676 32252 12747 32280
rect 13556 32280 13584 32379
rect 14458 32376 14464 32388
rect 14516 32376 14522 32428
rect 14645 32419 14703 32425
rect 14645 32385 14657 32419
rect 14691 32385 14703 32419
rect 15010 32416 15016 32428
rect 14971 32388 15016 32416
rect 14645 32379 14703 32385
rect 14274 32308 14280 32360
rect 14332 32348 14338 32360
rect 14660 32348 14688 32379
rect 15010 32376 15016 32388
rect 15068 32376 15074 32428
rect 15194 32416 15200 32428
rect 15155 32388 15200 32416
rect 15194 32376 15200 32388
rect 15252 32376 15258 32428
rect 15933 32419 15991 32425
rect 15933 32385 15945 32419
rect 15979 32416 15991 32419
rect 16206 32416 16212 32428
rect 15979 32388 16212 32416
rect 15979 32385 15991 32388
rect 15933 32379 15991 32385
rect 16206 32376 16212 32388
rect 16264 32376 16270 32428
rect 17126 32416 17132 32428
rect 17087 32388 17132 32416
rect 17126 32376 17132 32388
rect 17184 32376 17190 32428
rect 17770 32416 17776 32428
rect 17731 32388 17776 32416
rect 17770 32376 17776 32388
rect 17828 32376 17834 32428
rect 19242 32416 19248 32428
rect 19203 32388 19248 32416
rect 19242 32376 19248 32388
rect 19300 32376 19306 32428
rect 19512 32419 19570 32425
rect 19512 32385 19524 32419
rect 19558 32416 19570 32419
rect 20070 32416 20076 32428
rect 19558 32388 20076 32416
rect 19558 32385 19570 32388
rect 19512 32379 19570 32385
rect 20070 32376 20076 32388
rect 20128 32376 20134 32428
rect 21100 32425 21128 32456
rect 23198 32444 23204 32456
rect 23256 32484 23262 32496
rect 23256 32456 23336 32484
rect 23256 32444 23262 32456
rect 21085 32419 21143 32425
rect 21085 32385 21097 32419
rect 21131 32385 21143 32419
rect 22094 32416 22100 32428
rect 21085 32379 21143 32385
rect 21192 32388 22100 32416
rect 14332 32320 14688 32348
rect 14737 32351 14795 32357
rect 14332 32308 14338 32320
rect 14737 32317 14749 32351
rect 14783 32317 14795 32351
rect 14737 32311 14795 32317
rect 14829 32351 14887 32357
rect 14829 32317 14841 32351
rect 14875 32348 14887 32351
rect 15470 32348 15476 32360
rect 14875 32320 15476 32348
rect 14875 32317 14887 32320
rect 14829 32311 14887 32317
rect 14550 32280 14556 32292
rect 13556 32252 14556 32280
rect 12676 32240 12682 32252
rect 14550 32240 14556 32252
rect 14608 32240 14614 32292
rect 14752 32280 14780 32311
rect 15470 32308 15476 32320
rect 15528 32348 15534 32360
rect 16117 32351 16175 32357
rect 16117 32348 16129 32351
rect 15528 32320 16129 32348
rect 15528 32308 15534 32320
rect 16117 32317 16129 32320
rect 16163 32317 16175 32351
rect 21192 32348 21220 32388
rect 22094 32376 22100 32388
rect 22152 32416 22158 32428
rect 23308 32425 23336 32456
rect 26878 32444 26884 32496
rect 26936 32484 26942 32496
rect 27246 32484 27252 32496
rect 26936 32456 27252 32484
rect 26936 32444 26942 32456
rect 27246 32444 27252 32456
rect 27304 32484 27310 32496
rect 27706 32484 27712 32496
rect 27304 32456 27384 32484
rect 27667 32456 27712 32484
rect 27304 32444 27310 32456
rect 22281 32419 22339 32425
rect 22152 32388 22197 32416
rect 22152 32376 22158 32388
rect 22281 32385 22293 32419
rect 22327 32385 22339 32419
rect 22281 32379 22339 32385
rect 22649 32419 22707 32425
rect 22649 32385 22661 32419
rect 22695 32385 22707 32419
rect 22649 32379 22707 32385
rect 23293 32419 23351 32425
rect 23293 32385 23305 32419
rect 23339 32385 23351 32419
rect 23293 32379 23351 32385
rect 16117 32311 16175 32317
rect 20364 32320 21220 32348
rect 15286 32280 15292 32292
rect 14752 32252 15292 32280
rect 15286 32240 15292 32252
rect 15344 32240 15350 32292
rect 15654 32240 15660 32292
rect 15712 32280 15718 32292
rect 15712 32252 19288 32280
rect 15712 32240 15718 32252
rect 9582 32172 9588 32224
rect 9640 32212 9646 32224
rect 9861 32215 9919 32221
rect 9861 32212 9873 32215
rect 9640 32184 9873 32212
rect 9640 32172 9646 32184
rect 9861 32181 9873 32184
rect 9907 32181 9919 32215
rect 9861 32175 9919 32181
rect 13446 32172 13452 32224
rect 13504 32212 13510 32224
rect 13541 32215 13599 32221
rect 13541 32212 13553 32215
rect 13504 32184 13553 32212
rect 13504 32172 13510 32184
rect 13541 32181 13553 32184
rect 13587 32181 13599 32215
rect 13541 32175 13599 32181
rect 16850 32172 16856 32224
rect 16908 32212 16914 32224
rect 17865 32215 17923 32221
rect 17865 32212 17877 32215
rect 16908 32184 17877 32212
rect 16908 32172 16914 32184
rect 17865 32181 17877 32184
rect 17911 32181 17923 32215
rect 19260 32212 19288 32252
rect 19610 32212 19616 32224
rect 19260 32184 19616 32212
rect 17865 32175 17923 32181
rect 19610 32172 19616 32184
rect 19668 32212 19674 32224
rect 20364 32212 20392 32320
rect 21358 32308 21364 32360
rect 21416 32348 21422 32360
rect 22296 32348 22324 32379
rect 21416 32320 22324 32348
rect 22373 32351 22431 32357
rect 21416 32308 21422 32320
rect 22373 32317 22385 32351
rect 22419 32317 22431 32351
rect 22373 32311 22431 32317
rect 22465 32351 22523 32357
rect 22465 32317 22477 32351
rect 22511 32348 22523 32351
rect 22554 32348 22560 32360
rect 22511 32320 22560 32348
rect 22511 32317 22523 32320
rect 22465 32311 22523 32317
rect 20438 32240 20444 32292
rect 20496 32280 20502 32292
rect 20625 32283 20683 32289
rect 20625 32280 20637 32283
rect 20496 32252 20637 32280
rect 20496 32240 20502 32252
rect 20625 32249 20637 32252
rect 20671 32249 20683 32283
rect 22388 32280 22416 32311
rect 22554 32308 22560 32320
rect 22612 32308 22618 32360
rect 22664 32348 22692 32379
rect 23382 32376 23388 32428
rect 23440 32416 23446 32428
rect 24489 32419 24547 32425
rect 24489 32416 24501 32419
rect 23440 32388 24501 32416
rect 23440 32376 23446 32388
rect 24489 32385 24501 32388
rect 24535 32385 24547 32419
rect 25590 32416 25596 32428
rect 25503 32388 25596 32416
rect 24489 32379 24547 32385
rect 25590 32376 25596 32388
rect 25648 32416 25654 32428
rect 26142 32416 26148 32428
rect 25648 32388 26148 32416
rect 25648 32376 25654 32388
rect 26142 32376 26148 32388
rect 26200 32416 26206 32428
rect 26237 32419 26295 32425
rect 26237 32416 26249 32419
rect 26200 32388 26249 32416
rect 26200 32376 26206 32388
rect 26237 32385 26249 32388
rect 26283 32385 26295 32419
rect 26237 32379 26295 32385
rect 26418 32376 26424 32428
rect 26476 32416 26482 32428
rect 26973 32419 27031 32425
rect 26973 32416 26985 32419
rect 26476 32388 26985 32416
rect 26476 32376 26482 32388
rect 26973 32385 26985 32388
rect 27019 32416 27031 32419
rect 27062 32416 27068 32428
rect 27019 32388 27068 32416
rect 27019 32385 27031 32388
rect 26973 32379 27031 32385
rect 27062 32376 27068 32388
rect 27120 32376 27126 32428
rect 27154 32376 27160 32428
rect 27212 32416 27218 32428
rect 27356 32425 27384 32456
rect 27706 32444 27712 32456
rect 27764 32444 27770 32496
rect 28626 32484 28632 32496
rect 28368 32456 28632 32484
rect 27341 32419 27399 32425
rect 27212 32388 27257 32416
rect 27212 32376 27218 32388
rect 27341 32385 27353 32419
rect 27387 32385 27399 32419
rect 27341 32379 27399 32385
rect 27525 32419 27583 32425
rect 27525 32385 27537 32419
rect 27571 32416 27583 32419
rect 28368 32416 28396 32456
rect 28626 32444 28632 32456
rect 28684 32444 28690 32496
rect 28718 32444 28724 32496
rect 28776 32484 28782 32496
rect 29273 32487 29331 32493
rect 29273 32484 29285 32487
rect 28776 32456 29285 32484
rect 28776 32444 28782 32456
rect 29273 32453 29285 32456
rect 29319 32453 29331 32487
rect 29273 32447 29331 32453
rect 27571 32388 28396 32416
rect 27571 32385 27583 32388
rect 27525 32379 27583 32385
rect 28442 32376 28448 32428
rect 28500 32416 28506 32428
rect 28500 32388 28545 32416
rect 28500 32376 28506 32388
rect 29178 32376 29184 32428
rect 29236 32416 29242 32428
rect 30101 32419 30159 32425
rect 30101 32416 30113 32419
rect 29236 32388 30113 32416
rect 29236 32376 29242 32388
rect 30101 32385 30113 32388
rect 30147 32385 30159 32419
rect 30101 32379 30159 32385
rect 24394 32348 24400 32360
rect 22664 32320 24400 32348
rect 24394 32308 24400 32320
rect 24452 32308 24458 32360
rect 25498 32348 25504 32360
rect 24872 32320 25504 32348
rect 24872 32280 24900 32320
rect 25498 32308 25504 32320
rect 25556 32308 25562 32360
rect 27249 32351 27307 32357
rect 27249 32317 27261 32351
rect 27295 32348 27307 32351
rect 27430 32348 27436 32360
rect 27295 32320 27436 32348
rect 27295 32317 27307 32320
rect 27249 32311 27307 32317
rect 22388 32252 24900 32280
rect 24949 32283 25007 32289
rect 20625 32243 20683 32249
rect 24949 32249 24961 32283
rect 24995 32280 25007 32283
rect 26234 32280 26240 32292
rect 24995 32252 26240 32280
rect 24995 32249 25007 32252
rect 24949 32243 25007 32249
rect 26234 32240 26240 32252
rect 26292 32240 26298 32292
rect 26878 32240 26884 32292
rect 26936 32280 26942 32292
rect 27264 32280 27292 32311
rect 27430 32308 27436 32320
rect 27488 32308 27494 32360
rect 26936 32252 27292 32280
rect 28261 32283 28319 32289
rect 26936 32240 26942 32252
rect 28261 32249 28273 32283
rect 28307 32280 28319 32283
rect 28902 32280 28908 32292
rect 28307 32252 28908 32280
rect 28307 32249 28319 32252
rect 28261 32243 28319 32249
rect 28902 32240 28908 32252
rect 28960 32240 28966 32292
rect 24762 32212 24768 32224
rect 19668 32184 20392 32212
rect 24723 32184 24768 32212
rect 19668 32172 19674 32184
rect 24762 32172 24768 32184
rect 24820 32172 24826 32224
rect 25682 32172 25688 32224
rect 25740 32212 25746 32224
rect 25777 32215 25835 32221
rect 25777 32212 25789 32215
rect 25740 32184 25789 32212
rect 25740 32172 25746 32184
rect 25777 32181 25789 32184
rect 25823 32181 25835 32215
rect 25777 32175 25835 32181
rect 26786 32172 26792 32224
rect 26844 32212 26850 32224
rect 27154 32212 27160 32224
rect 26844 32184 27160 32212
rect 26844 32172 26850 32184
rect 27154 32172 27160 32184
rect 27212 32172 27218 32224
rect 29270 32212 29276 32224
rect 29231 32184 29276 32212
rect 29270 32172 29276 32184
rect 29328 32172 29334 32224
rect 29822 32172 29828 32224
rect 29880 32212 29886 32224
rect 29917 32215 29975 32221
rect 29917 32212 29929 32215
rect 29880 32184 29929 32212
rect 29880 32172 29886 32184
rect 29917 32181 29929 32184
rect 29963 32181 29975 32215
rect 29917 32175 29975 32181
rect 1104 32122 30820 32144
rect 1104 32070 5915 32122
rect 5967 32070 5979 32122
rect 6031 32070 6043 32122
rect 6095 32070 6107 32122
rect 6159 32070 6171 32122
rect 6223 32070 15846 32122
rect 15898 32070 15910 32122
rect 15962 32070 15974 32122
rect 16026 32070 16038 32122
rect 16090 32070 16102 32122
rect 16154 32070 25776 32122
rect 25828 32070 25840 32122
rect 25892 32070 25904 32122
rect 25956 32070 25968 32122
rect 26020 32070 26032 32122
rect 26084 32070 30820 32122
rect 1104 32048 30820 32070
rect 10137 32011 10195 32017
rect 10137 31977 10149 32011
rect 10183 32008 10195 32011
rect 10318 32008 10324 32020
rect 10183 31980 10324 32008
rect 10183 31977 10195 31980
rect 10137 31971 10195 31977
rect 10318 31968 10324 31980
rect 10376 31968 10382 32020
rect 11790 32008 11796 32020
rect 11751 31980 11796 32008
rect 11790 31968 11796 31980
rect 11848 31968 11854 32020
rect 12342 31968 12348 32020
rect 12400 32008 12406 32020
rect 15654 32008 15660 32020
rect 12400 31980 15660 32008
rect 12400 31968 12406 31980
rect 15654 31968 15660 31980
rect 15712 31968 15718 32020
rect 16298 31968 16304 32020
rect 16356 32008 16362 32020
rect 20993 32011 21051 32017
rect 20993 32008 21005 32011
rect 16356 31980 21005 32008
rect 16356 31968 16362 31980
rect 20993 31977 21005 31980
rect 21039 31977 21051 32011
rect 23106 32008 23112 32020
rect 23067 31980 23112 32008
rect 20993 31971 21051 31977
rect 23106 31968 23112 31980
rect 23164 31968 23170 32020
rect 24670 32008 24676 32020
rect 24631 31980 24676 32008
rect 24670 31968 24676 31980
rect 24728 31968 24734 32020
rect 24854 32008 24860 32020
rect 24815 31980 24860 32008
rect 24854 31968 24860 31980
rect 24912 31968 24918 32020
rect 26142 31968 26148 32020
rect 26200 32008 26206 32020
rect 26878 32008 26884 32020
rect 26200 31980 26884 32008
rect 26200 31968 26206 31980
rect 26878 31968 26884 31980
rect 26936 31968 26942 32020
rect 28169 32011 28227 32017
rect 26988 31980 28120 32008
rect 10226 31900 10232 31952
rect 10284 31940 10290 31952
rect 10505 31943 10563 31949
rect 10505 31940 10517 31943
rect 10284 31912 10517 31940
rect 10284 31900 10290 31912
rect 10505 31909 10517 31912
rect 10551 31909 10563 31943
rect 16666 31940 16672 31952
rect 10505 31903 10563 31909
rect 16592 31912 16672 31940
rect 10686 31832 10692 31884
rect 10744 31872 10750 31884
rect 11149 31875 11207 31881
rect 11149 31872 11161 31875
rect 10744 31844 11161 31872
rect 10744 31832 10750 31844
rect 11149 31841 11161 31844
rect 11195 31841 11207 31875
rect 11149 31835 11207 31841
rect 11882 31832 11888 31884
rect 11940 31872 11946 31884
rect 12253 31875 12311 31881
rect 12253 31872 12265 31875
rect 11940 31844 12265 31872
rect 11940 31832 11946 31844
rect 12253 31841 12265 31844
rect 12299 31841 12311 31875
rect 12253 31835 12311 31841
rect 12437 31875 12495 31881
rect 12437 31841 12449 31875
rect 12483 31872 12495 31875
rect 12618 31872 12624 31884
rect 12483 31844 12624 31872
rect 12483 31841 12495 31844
rect 12437 31835 12495 31841
rect 12618 31832 12624 31844
rect 12676 31832 12682 31884
rect 10321 31807 10379 31813
rect 10321 31773 10333 31807
rect 10367 31804 10379 31807
rect 10410 31804 10416 31816
rect 10367 31776 10416 31804
rect 10367 31773 10379 31776
rect 10321 31767 10379 31773
rect 10410 31764 10416 31776
rect 10468 31764 10474 31816
rect 10597 31807 10655 31813
rect 10597 31773 10609 31807
rect 10643 31804 10655 31807
rect 10778 31804 10784 31816
rect 10643 31776 10784 31804
rect 10643 31773 10655 31776
rect 10597 31767 10655 31773
rect 10778 31764 10784 31776
rect 10836 31764 10842 31816
rect 11057 31807 11115 31813
rect 11057 31773 11069 31807
rect 11103 31804 11115 31807
rect 11238 31804 11244 31816
rect 11103 31776 11244 31804
rect 11103 31773 11115 31776
rect 11057 31767 11115 31773
rect 11238 31764 11244 31776
rect 11296 31804 11302 31816
rect 11790 31804 11796 31816
rect 11296 31776 11796 31804
rect 11296 31764 11302 31776
rect 11790 31764 11796 31776
rect 11848 31764 11854 31816
rect 15010 31764 15016 31816
rect 15068 31804 15074 31816
rect 15749 31807 15807 31813
rect 15749 31804 15761 31807
rect 15068 31776 15761 31804
rect 15068 31764 15074 31776
rect 15749 31773 15761 31776
rect 15795 31773 15807 31807
rect 15749 31767 15807 31773
rect 15930 31764 15936 31816
rect 15988 31804 15994 31816
rect 16592 31813 16620 31912
rect 16666 31900 16672 31912
rect 16724 31900 16730 31952
rect 18230 31900 18236 31952
rect 18288 31940 18294 31952
rect 18601 31943 18659 31949
rect 18601 31940 18613 31943
rect 18288 31912 18613 31940
rect 18288 31900 18294 31912
rect 18601 31909 18613 31912
rect 18647 31909 18659 31943
rect 21450 31940 21456 31952
rect 18601 31903 18659 31909
rect 20916 31912 21456 31940
rect 16761 31875 16819 31881
rect 16761 31841 16773 31875
rect 16807 31872 16819 31875
rect 16807 31844 17908 31872
rect 16807 31841 16819 31844
rect 16761 31835 16819 31841
rect 16393 31807 16451 31813
rect 16393 31804 16405 31807
rect 15988 31776 16405 31804
rect 15988 31764 15994 31776
rect 16393 31773 16405 31776
rect 16439 31773 16451 31807
rect 16393 31767 16451 31773
rect 16577 31807 16635 31813
rect 16577 31773 16589 31807
rect 16623 31773 16635 31807
rect 16577 31767 16635 31773
rect 16669 31807 16727 31813
rect 16669 31773 16681 31807
rect 16715 31773 16727 31807
rect 16942 31804 16948 31816
rect 16903 31776 16948 31804
rect 16669 31767 16727 31773
rect 12161 31739 12219 31745
rect 12161 31705 12173 31739
rect 12207 31736 12219 31739
rect 12526 31736 12532 31748
rect 12207 31708 12532 31736
rect 12207 31705 12219 31708
rect 12161 31699 12219 31705
rect 12526 31696 12532 31708
rect 12584 31696 12590 31748
rect 16684 31736 16712 31767
rect 16942 31764 16948 31776
rect 17000 31764 17006 31816
rect 16758 31736 16764 31748
rect 16684 31708 16764 31736
rect 16758 31696 16764 31708
rect 16816 31696 16822 31748
rect 17880 31680 17908 31844
rect 18506 31832 18512 31884
rect 18564 31872 18570 31884
rect 19981 31875 20039 31881
rect 19981 31872 19993 31875
rect 18564 31844 19993 31872
rect 18564 31832 18570 31844
rect 19981 31841 19993 31844
rect 20027 31841 20039 31875
rect 19981 31835 20039 31841
rect 18322 31764 18328 31816
rect 18380 31804 18386 31816
rect 18417 31807 18475 31813
rect 18417 31804 18429 31807
rect 18380 31776 18429 31804
rect 18380 31764 18386 31776
rect 18417 31773 18429 31776
rect 18463 31773 18475 31807
rect 18417 31767 18475 31773
rect 19889 31807 19947 31813
rect 19889 31773 19901 31807
rect 19935 31804 19947 31807
rect 20916 31804 20944 31912
rect 21450 31900 21456 31912
rect 21508 31900 21514 31952
rect 22922 31900 22928 31952
rect 22980 31940 22986 31952
rect 23845 31943 23903 31949
rect 23845 31940 23857 31943
rect 22980 31912 23857 31940
rect 22980 31900 22986 31912
rect 23845 31909 23857 31912
rect 23891 31909 23903 31943
rect 23845 31903 23903 31909
rect 25961 31943 26019 31949
rect 25961 31909 25973 31943
rect 26007 31940 26019 31943
rect 26786 31940 26792 31952
rect 26007 31912 26792 31940
rect 26007 31909 26019 31912
rect 25961 31903 26019 31909
rect 26786 31900 26792 31912
rect 26844 31900 26850 31952
rect 20993 31875 21051 31881
rect 20993 31841 21005 31875
rect 21039 31872 21051 31875
rect 21085 31875 21143 31881
rect 21085 31872 21097 31875
rect 21039 31844 21097 31872
rect 21039 31841 21051 31844
rect 20993 31835 21051 31841
rect 21085 31841 21097 31844
rect 21131 31841 21143 31875
rect 21358 31872 21364 31884
rect 21319 31844 21364 31872
rect 21085 31835 21143 31841
rect 19935 31776 20944 31804
rect 21100 31804 21128 31835
rect 21358 31832 21364 31844
rect 21416 31872 21422 31884
rect 22002 31872 22008 31884
rect 21416 31844 22008 31872
rect 21416 31832 21422 31844
rect 22002 31832 22008 31844
rect 22060 31872 22066 31884
rect 22649 31875 22707 31881
rect 22060 31844 22600 31872
rect 22060 31832 22066 31844
rect 21266 31804 21272 31816
rect 21100 31776 21272 31804
rect 19935 31773 19947 31776
rect 19889 31767 19947 31773
rect 21266 31764 21272 31776
rect 21324 31764 21330 31816
rect 22094 31764 22100 31816
rect 22152 31804 22158 31816
rect 22572 31813 22600 31844
rect 22649 31841 22661 31875
rect 22695 31872 22707 31875
rect 26326 31872 26332 31884
rect 22695 31844 26332 31872
rect 22695 31841 22707 31844
rect 22649 31835 22707 31841
rect 26326 31832 26332 31844
rect 26384 31832 26390 31884
rect 26697 31875 26755 31881
rect 26697 31841 26709 31875
rect 26743 31872 26755 31875
rect 26878 31872 26884 31884
rect 26743 31844 26884 31872
rect 26743 31841 26755 31844
rect 26697 31835 26755 31841
rect 26878 31832 26884 31844
rect 26936 31832 26942 31884
rect 22373 31807 22431 31813
rect 22373 31804 22385 31807
rect 22152 31776 22385 31804
rect 22152 31764 22158 31776
rect 22373 31773 22385 31776
rect 22419 31773 22431 31807
rect 22373 31767 22431 31773
rect 22557 31807 22615 31813
rect 22557 31773 22569 31807
rect 22603 31773 22615 31807
rect 22557 31767 22615 31773
rect 22741 31807 22799 31813
rect 22741 31773 22753 31807
rect 22787 31804 22799 31807
rect 22925 31807 22983 31813
rect 22787 31776 22821 31804
rect 22787 31773 22799 31776
rect 22741 31767 22799 31773
rect 22925 31773 22937 31807
rect 22971 31804 22983 31807
rect 23382 31804 23388 31816
rect 22971 31776 23388 31804
rect 22971 31773 22983 31776
rect 22925 31767 22983 31773
rect 18598 31696 18604 31748
rect 18656 31736 18662 31748
rect 19242 31736 19248 31748
rect 18656 31708 19248 31736
rect 18656 31696 18662 31708
rect 19242 31696 19248 31708
rect 19300 31696 19306 31748
rect 10502 31628 10508 31680
rect 10560 31668 10566 31680
rect 15378 31668 15384 31680
rect 10560 31640 15384 31668
rect 10560 31628 10566 31640
rect 15378 31628 15384 31640
rect 15436 31628 15442 31680
rect 15841 31671 15899 31677
rect 15841 31637 15853 31671
rect 15887 31668 15899 31671
rect 16942 31668 16948 31680
rect 15887 31640 16948 31668
rect 15887 31637 15899 31640
rect 15841 31631 15899 31637
rect 16942 31628 16948 31640
rect 17000 31628 17006 31680
rect 17129 31671 17187 31677
rect 17129 31637 17141 31671
rect 17175 31668 17187 31671
rect 17402 31668 17408 31680
rect 17175 31640 17408 31668
rect 17175 31637 17187 31640
rect 17129 31631 17187 31637
rect 17402 31628 17408 31640
rect 17460 31628 17466 31680
rect 17862 31628 17868 31680
rect 17920 31628 17926 31680
rect 22554 31628 22560 31680
rect 22612 31668 22618 31680
rect 22756 31668 22784 31767
rect 23382 31764 23388 31776
rect 23440 31764 23446 31816
rect 23658 31804 23664 31816
rect 23619 31776 23664 31804
rect 23658 31764 23664 31776
rect 23716 31764 23722 31816
rect 24394 31804 24400 31816
rect 24355 31776 24400 31804
rect 24394 31764 24400 31776
rect 24452 31764 24458 31816
rect 25682 31764 25688 31816
rect 25740 31804 25746 31816
rect 25777 31807 25835 31813
rect 25777 31804 25789 31807
rect 25740 31776 25789 31804
rect 25740 31764 25746 31776
rect 25777 31773 25789 31776
rect 25823 31773 25835 31807
rect 26418 31804 26424 31816
rect 26379 31776 26424 31804
rect 25777 31767 25835 31773
rect 26418 31764 26424 31776
rect 26476 31764 26482 31816
rect 26605 31807 26663 31813
rect 26605 31773 26617 31807
rect 26651 31804 26663 31807
rect 26651 31776 26685 31804
rect 26651 31773 26663 31776
rect 26605 31767 26663 31773
rect 26510 31696 26516 31748
rect 26568 31736 26574 31748
rect 26620 31736 26648 31767
rect 26786 31764 26792 31816
rect 26844 31804 26850 31816
rect 26988 31813 27016 31980
rect 28092 31940 28120 31980
rect 28169 31977 28181 32011
rect 28215 32008 28227 32011
rect 28258 32008 28264 32020
rect 28215 31980 28264 32008
rect 28215 31977 28227 31980
rect 28169 31971 28227 31977
rect 28258 31968 28264 31980
rect 28316 31968 28322 32020
rect 28718 31940 28724 31952
rect 28092 31912 28724 31940
rect 28718 31900 28724 31912
rect 28776 31900 28782 31952
rect 28813 31943 28871 31949
rect 28813 31909 28825 31943
rect 28859 31909 28871 31943
rect 28813 31903 28871 31909
rect 28828 31872 28856 31903
rect 28828 31844 29868 31872
rect 26973 31807 27031 31813
rect 26844 31776 26937 31804
rect 26844 31764 26850 31776
rect 26568 31708 26648 31736
rect 26896 31736 26924 31776
rect 26973 31773 26985 31807
rect 27019 31773 27031 31807
rect 27246 31804 27252 31816
rect 26973 31767 27031 31773
rect 27080 31776 27252 31804
rect 27080 31736 27108 31776
rect 27246 31764 27252 31776
rect 27304 31764 27310 31816
rect 28353 31807 28411 31813
rect 28353 31773 28365 31807
rect 28399 31804 28411 31807
rect 28994 31804 29000 31816
rect 28399 31776 28856 31804
rect 28955 31776 29000 31804
rect 28399 31773 28411 31776
rect 28353 31767 28411 31773
rect 26896 31708 27108 31736
rect 28828 31736 28856 31776
rect 28994 31764 29000 31776
rect 29052 31764 29058 31816
rect 29840 31813 29868 31844
rect 29825 31807 29883 31813
rect 29825 31773 29837 31807
rect 29871 31773 29883 31807
rect 29825 31767 29883 31773
rect 30098 31736 30104 31748
rect 28828 31708 30104 31736
rect 26568 31696 26574 31708
rect 30098 31696 30104 31708
rect 30156 31696 30162 31748
rect 22612 31640 22784 31668
rect 27157 31671 27215 31677
rect 22612 31628 22618 31640
rect 27157 31637 27169 31671
rect 27203 31668 27215 31671
rect 27430 31668 27436 31680
rect 27203 31640 27436 31668
rect 27203 31637 27215 31640
rect 27157 31631 27215 31637
rect 27430 31628 27436 31640
rect 27488 31628 27494 31680
rect 30006 31668 30012 31680
rect 29967 31640 30012 31668
rect 30006 31628 30012 31640
rect 30064 31628 30070 31680
rect 1104 31578 30820 31600
rect 1104 31526 10880 31578
rect 10932 31526 10944 31578
rect 10996 31526 11008 31578
rect 11060 31526 11072 31578
rect 11124 31526 11136 31578
rect 11188 31526 20811 31578
rect 20863 31526 20875 31578
rect 20927 31526 20939 31578
rect 20991 31526 21003 31578
rect 21055 31526 21067 31578
rect 21119 31526 30820 31578
rect 1104 31504 30820 31526
rect 10410 31424 10416 31476
rect 10468 31464 10474 31476
rect 10686 31464 10692 31476
rect 10468 31436 10692 31464
rect 10468 31424 10474 31436
rect 10686 31424 10692 31436
rect 10744 31424 10750 31476
rect 10965 31467 11023 31473
rect 10965 31433 10977 31467
rect 11011 31464 11023 31467
rect 11330 31464 11336 31476
rect 11011 31436 11336 31464
rect 11011 31433 11023 31436
rect 10965 31427 11023 31433
rect 11330 31424 11336 31436
rect 11388 31424 11394 31476
rect 12802 31464 12808 31476
rect 12763 31436 12808 31464
rect 12802 31424 12808 31436
rect 12860 31424 12866 31476
rect 15565 31467 15623 31473
rect 15565 31433 15577 31467
rect 15611 31464 15623 31467
rect 15930 31464 15936 31476
rect 15611 31436 15936 31464
rect 15611 31433 15623 31436
rect 15565 31427 15623 31433
rect 15930 31424 15936 31436
rect 15988 31424 15994 31476
rect 23198 31464 23204 31476
rect 23159 31436 23204 31464
rect 23198 31424 23204 31436
rect 23256 31424 23262 31476
rect 26142 31424 26148 31476
rect 26200 31464 26206 31476
rect 28537 31467 28595 31473
rect 26200 31436 27568 31464
rect 26200 31424 26206 31436
rect 12434 31396 12440 31408
rect 2746 31368 12440 31396
rect 1673 31331 1731 31337
rect 1673 31297 1685 31331
rect 1719 31328 1731 31331
rect 2746 31328 2774 31368
rect 12434 31356 12440 31368
rect 12492 31396 12498 31408
rect 12492 31368 13032 31396
rect 12492 31356 12498 31368
rect 1719 31300 2774 31328
rect 7929 31331 7987 31337
rect 1719 31297 1731 31300
rect 1673 31291 1731 31297
rect 7929 31297 7941 31331
rect 7975 31328 7987 31331
rect 8202 31328 8208 31340
rect 7975 31300 8208 31328
rect 7975 31297 7987 31300
rect 7929 31291 7987 31297
rect 8202 31288 8208 31300
rect 8260 31288 8266 31340
rect 8846 31337 8852 31340
rect 8840 31291 8852 31337
rect 8904 31328 8910 31340
rect 8904 31300 8940 31328
rect 8846 31288 8852 31291
rect 8904 31288 8910 31300
rect 10410 31288 10416 31340
rect 10468 31328 10474 31340
rect 10597 31331 10655 31337
rect 10597 31328 10609 31331
rect 10468 31300 10609 31328
rect 10468 31288 10474 31300
rect 10597 31297 10609 31300
rect 10643 31297 10655 31331
rect 10597 31291 10655 31297
rect 11514 31288 11520 31340
rect 11572 31328 11578 31340
rect 11609 31331 11667 31337
rect 11609 31328 11621 31331
rect 11572 31300 11621 31328
rect 11572 31288 11578 31300
rect 11609 31297 11621 31300
rect 11655 31328 11667 31331
rect 11698 31328 11704 31340
rect 11655 31300 11704 31328
rect 11655 31297 11667 31300
rect 11609 31291 11667 31297
rect 11698 31288 11704 31300
rect 11756 31288 11762 31340
rect 11790 31288 11796 31340
rect 11848 31328 11854 31340
rect 12894 31328 12900 31340
rect 11848 31300 12900 31328
rect 11848 31288 11854 31300
rect 12894 31288 12900 31300
rect 12952 31288 12958 31340
rect 1394 31260 1400 31272
rect 1355 31232 1400 31260
rect 1394 31220 1400 31232
rect 1452 31220 1458 31272
rect 8573 31263 8631 31269
rect 8573 31260 8585 31263
rect 8128 31232 8585 31260
rect 8128 31201 8156 31232
rect 8573 31229 8585 31232
rect 8619 31229 8631 31263
rect 8573 31223 8631 31229
rect 10689 31263 10747 31269
rect 10689 31229 10701 31263
rect 10735 31260 10747 31263
rect 10778 31260 10784 31272
rect 10735 31232 10784 31260
rect 10735 31229 10747 31232
rect 10689 31223 10747 31229
rect 8113 31195 8171 31201
rect 8113 31161 8125 31195
rect 8159 31161 8171 31195
rect 9950 31192 9956 31204
rect 9863 31164 9956 31192
rect 8113 31155 8171 31161
rect 9950 31152 9956 31164
rect 10008 31192 10014 31204
rect 10502 31192 10508 31204
rect 10008 31164 10508 31192
rect 10008 31152 10014 31164
rect 10502 31152 10508 31164
rect 10560 31192 10566 31204
rect 10704 31192 10732 31223
rect 10778 31220 10784 31232
rect 10836 31220 10842 31272
rect 11882 31220 11888 31272
rect 11940 31220 11946 31272
rect 12805 31263 12863 31269
rect 12805 31229 12817 31263
rect 12851 31260 12863 31263
rect 13004 31260 13032 31368
rect 13446 31356 13452 31408
rect 13504 31396 13510 31408
rect 15381 31399 15439 31405
rect 15381 31396 15393 31399
rect 13504 31368 15393 31396
rect 13504 31356 13510 31368
rect 15381 31365 15393 31368
rect 15427 31365 15439 31399
rect 15381 31359 15439 31365
rect 17678 31356 17684 31408
rect 17736 31396 17742 31408
rect 17736 31368 18092 31396
rect 17736 31356 17742 31368
rect 15197 31331 15255 31337
rect 15197 31297 15209 31331
rect 15243 31328 15255 31331
rect 15286 31328 15292 31340
rect 15243 31300 15292 31328
rect 15243 31297 15255 31300
rect 15197 31291 15255 31297
rect 15286 31288 15292 31300
rect 15344 31288 15350 31340
rect 17773 31331 17831 31337
rect 17773 31297 17785 31331
rect 17819 31297 17831 31331
rect 17954 31328 17960 31340
rect 17915 31300 17960 31328
rect 17773 31291 17831 31297
rect 13078 31260 13084 31272
rect 12851 31232 13084 31260
rect 12851 31229 12863 31232
rect 12805 31223 12863 31229
rect 13078 31220 13084 31232
rect 13136 31220 13142 31272
rect 17788 31260 17816 31291
rect 17954 31288 17960 31300
rect 18012 31288 18018 31340
rect 18064 31337 18092 31368
rect 18230 31356 18236 31408
rect 18288 31396 18294 31408
rect 18969 31399 19027 31405
rect 18969 31396 18981 31399
rect 18288 31368 18981 31396
rect 18288 31356 18294 31368
rect 18969 31365 18981 31368
rect 19015 31365 19027 31399
rect 18969 31359 19027 31365
rect 19245 31399 19303 31405
rect 19245 31365 19257 31399
rect 19291 31396 19303 31399
rect 20162 31396 20168 31408
rect 19291 31368 20168 31396
rect 19291 31365 19303 31368
rect 19245 31359 19303 31365
rect 20162 31356 20168 31368
rect 20220 31356 20226 31408
rect 20714 31356 20720 31408
rect 20772 31396 20778 31408
rect 21085 31399 21143 31405
rect 21085 31396 21097 31399
rect 20772 31368 21097 31396
rect 20772 31356 20778 31368
rect 21085 31365 21097 31368
rect 21131 31365 21143 31399
rect 21085 31359 21143 31365
rect 21726 31356 21732 31408
rect 21784 31396 21790 31408
rect 21910 31396 21916 31408
rect 21784 31368 21916 31396
rect 21784 31356 21790 31368
rect 21910 31356 21916 31368
rect 21968 31356 21974 31408
rect 26694 31396 26700 31408
rect 22112 31368 26700 31396
rect 18049 31331 18107 31337
rect 18049 31297 18061 31331
rect 18095 31297 18107 31331
rect 18049 31291 18107 31297
rect 18325 31331 18383 31337
rect 18325 31297 18337 31331
rect 18371 31328 18383 31331
rect 18414 31328 18420 31340
rect 18371 31300 18420 31328
rect 18371 31297 18383 31300
rect 18325 31291 18383 31297
rect 18414 31288 18420 31300
rect 18472 31288 18478 31340
rect 19058 31288 19064 31340
rect 19116 31328 19122 31340
rect 19153 31331 19211 31337
rect 19153 31328 19165 31331
rect 19116 31300 19165 31328
rect 19116 31288 19122 31300
rect 19153 31297 19165 31300
rect 19199 31297 19211 31331
rect 19153 31291 19211 31297
rect 19334 31288 19340 31340
rect 19392 31337 19398 31340
rect 19392 31328 19400 31337
rect 19392 31300 19437 31328
rect 19392 31291 19400 31300
rect 19392 31288 19398 31291
rect 19702 31288 19708 31340
rect 19760 31328 19766 31340
rect 20349 31331 20407 31337
rect 20349 31328 20361 31331
rect 19760 31300 20361 31328
rect 19760 31288 19766 31300
rect 20349 31297 20361 31300
rect 20395 31297 20407 31331
rect 20349 31291 20407 31297
rect 21821 31331 21879 31337
rect 21821 31297 21833 31331
rect 21867 31297 21879 31331
rect 22002 31328 22008 31340
rect 21963 31300 22008 31328
rect 21821 31291 21879 31297
rect 18138 31260 18144 31272
rect 17788 31232 17908 31260
rect 18051 31232 18144 31260
rect 10560 31164 10732 31192
rect 10560 31152 10566 31164
rect 11422 31152 11428 31204
rect 11480 31192 11486 31204
rect 11900 31192 11928 31220
rect 12345 31195 12403 31201
rect 12345 31192 12357 31195
rect 11480 31164 12357 31192
rect 11480 31152 11486 31164
rect 12345 31161 12357 31164
rect 12391 31161 12403 31195
rect 17880 31192 17908 31232
rect 18138 31220 18144 31232
rect 18196 31260 18202 31272
rect 18506 31260 18512 31272
rect 18196 31232 18512 31260
rect 18196 31220 18202 31232
rect 18506 31220 18512 31232
rect 18564 31220 18570 31272
rect 21836 31260 21864 31291
rect 22002 31288 22008 31300
rect 22060 31288 22066 31340
rect 22112 31337 22140 31368
rect 26694 31356 26700 31368
rect 26752 31396 26758 31408
rect 27062 31396 27068 31408
rect 26752 31368 27068 31396
rect 26752 31356 26758 31368
rect 27062 31356 27068 31368
rect 27120 31356 27126 31408
rect 27430 31405 27436 31408
rect 27424 31396 27436 31405
rect 27391 31368 27436 31396
rect 27424 31359 27436 31368
rect 27430 31356 27436 31359
rect 27488 31356 27494 31408
rect 27540 31396 27568 31436
rect 28537 31433 28549 31467
rect 28583 31464 28595 31467
rect 28718 31464 28724 31476
rect 28583 31436 28724 31464
rect 28583 31433 28595 31436
rect 28537 31427 28595 31433
rect 28718 31424 28724 31436
rect 28776 31424 28782 31476
rect 28994 31424 29000 31476
rect 29052 31464 29058 31476
rect 29549 31467 29607 31473
rect 29549 31464 29561 31467
rect 29052 31436 29561 31464
rect 29052 31424 29058 31436
rect 29549 31433 29561 31436
rect 29595 31433 29607 31467
rect 29549 31427 29607 31433
rect 29365 31399 29423 31405
rect 29365 31396 29377 31399
rect 27540 31368 29377 31396
rect 29365 31365 29377 31368
rect 29411 31365 29423 31399
rect 29365 31359 29423 31365
rect 22097 31331 22155 31337
rect 22097 31297 22109 31331
rect 22143 31297 22155 31331
rect 22097 31291 22155 31297
rect 22373 31331 22431 31337
rect 22373 31297 22385 31331
rect 22419 31328 22431 31331
rect 22830 31328 22836 31340
rect 22419 31300 22836 31328
rect 22419 31297 22431 31300
rect 22373 31291 22431 31297
rect 22830 31288 22836 31300
rect 22888 31288 22894 31340
rect 23017 31331 23075 31337
rect 23017 31297 23029 31331
rect 23063 31328 23075 31331
rect 23566 31328 23572 31340
rect 23063 31300 23572 31328
rect 23063 31297 23075 31300
rect 23017 31291 23075 31297
rect 23566 31288 23572 31300
rect 23624 31288 23630 31340
rect 27154 31328 27160 31340
rect 27115 31300 27160 31328
rect 27154 31288 27160 31300
rect 27212 31288 27218 31340
rect 21910 31260 21916 31272
rect 21836 31232 21916 31260
rect 21910 31220 21916 31232
rect 21968 31220 21974 31272
rect 22189 31263 22247 31269
rect 22189 31229 22201 31263
rect 22235 31260 22247 31263
rect 22554 31260 22560 31272
rect 22235 31232 22560 31260
rect 22235 31229 22247 31232
rect 22189 31223 22247 31229
rect 22554 31220 22560 31232
rect 22612 31220 22618 31272
rect 23937 31263 23995 31269
rect 23937 31229 23949 31263
rect 23983 31260 23995 31263
rect 24026 31260 24032 31272
rect 23983 31232 24032 31260
rect 23983 31229 23995 31232
rect 23937 31223 23995 31229
rect 24026 31220 24032 31232
rect 24084 31220 24090 31272
rect 24210 31260 24216 31272
rect 24171 31232 24216 31260
rect 24210 31220 24216 31232
rect 24268 31220 24274 31272
rect 24854 31220 24860 31272
rect 24912 31260 24918 31272
rect 25409 31263 25467 31269
rect 25409 31260 25421 31263
rect 24912 31232 25421 31260
rect 24912 31220 24918 31232
rect 25409 31229 25421 31232
rect 25455 31229 25467 31263
rect 25682 31260 25688 31272
rect 25643 31232 25688 31260
rect 25409 31223 25467 31229
rect 25682 31220 25688 31232
rect 25740 31260 25746 31272
rect 26050 31260 26056 31272
rect 25740 31232 26056 31260
rect 25740 31220 25746 31232
rect 26050 31220 26056 31232
rect 26108 31220 26114 31272
rect 18969 31195 19027 31201
rect 18969 31192 18981 31195
rect 17880 31164 18981 31192
rect 12345 31155 12403 31161
rect 18969 31161 18981 31164
rect 19015 31161 19027 31195
rect 18969 31155 19027 31161
rect 28626 31152 28632 31204
rect 28684 31192 28690 31204
rect 28902 31192 28908 31204
rect 28684 31164 28908 31192
rect 28684 31152 28690 31164
rect 28902 31152 28908 31164
rect 28960 31192 28966 31204
rect 28997 31195 29055 31201
rect 28997 31192 29009 31195
rect 28960 31164 29009 31192
rect 28960 31152 28966 31164
rect 28997 31161 29009 31164
rect 29043 31161 29055 31195
rect 28997 31155 29055 31161
rect 10594 31124 10600 31136
rect 10555 31096 10600 31124
rect 10594 31084 10600 31096
rect 10652 31084 10658 31136
rect 11609 31127 11667 31133
rect 11609 31093 11621 31127
rect 11655 31124 11667 31127
rect 11882 31124 11888 31136
rect 11655 31096 11888 31124
rect 11655 31093 11667 31096
rect 11609 31087 11667 31093
rect 11882 31084 11888 31096
rect 11940 31084 11946 31136
rect 16758 31084 16764 31136
rect 16816 31124 16822 31136
rect 17954 31124 17960 31136
rect 16816 31096 17960 31124
rect 16816 31084 16822 31096
rect 17954 31084 17960 31096
rect 18012 31084 18018 31136
rect 18509 31127 18567 31133
rect 18509 31093 18521 31127
rect 18555 31124 18567 31127
rect 18598 31124 18604 31136
rect 18555 31096 18604 31124
rect 18555 31093 18567 31096
rect 18509 31087 18567 31093
rect 18598 31084 18604 31096
rect 18656 31084 18662 31136
rect 20346 31084 20352 31136
rect 20404 31124 20410 31136
rect 20533 31127 20591 31133
rect 20533 31124 20545 31127
rect 20404 31096 20545 31124
rect 20404 31084 20410 31096
rect 20533 31093 20545 31096
rect 20579 31093 20591 31127
rect 21174 31124 21180 31136
rect 21135 31096 21180 31124
rect 20533 31087 20591 31093
rect 21174 31084 21180 31096
rect 21232 31084 21238 31136
rect 21358 31084 21364 31136
rect 21416 31124 21422 31136
rect 22557 31127 22615 31133
rect 22557 31124 22569 31127
rect 21416 31096 22569 31124
rect 21416 31084 21422 31096
rect 22557 31093 22569 31096
rect 22603 31093 22615 31127
rect 22557 31087 22615 31093
rect 23014 31084 23020 31136
rect 23072 31124 23078 31136
rect 29086 31124 29092 31136
rect 23072 31096 29092 31124
rect 23072 31084 23078 31096
rect 29086 31084 29092 31096
rect 29144 31124 29150 31136
rect 29365 31127 29423 31133
rect 29365 31124 29377 31127
rect 29144 31096 29377 31124
rect 29144 31084 29150 31096
rect 29365 31093 29377 31096
rect 29411 31124 29423 31127
rect 29914 31124 29920 31136
rect 29411 31096 29920 31124
rect 29411 31093 29423 31096
rect 29365 31087 29423 31093
rect 29914 31084 29920 31096
rect 29972 31084 29978 31136
rect 1104 31034 30820 31056
rect 1104 30982 5915 31034
rect 5967 30982 5979 31034
rect 6031 30982 6043 31034
rect 6095 30982 6107 31034
rect 6159 30982 6171 31034
rect 6223 30982 15846 31034
rect 15898 30982 15910 31034
rect 15962 30982 15974 31034
rect 16026 30982 16038 31034
rect 16090 30982 16102 31034
rect 16154 30982 25776 31034
rect 25828 30982 25840 31034
rect 25892 30982 25904 31034
rect 25956 30982 25968 31034
rect 26020 30982 26032 31034
rect 26084 30982 30820 31034
rect 1104 30960 30820 30982
rect 10594 30880 10600 30932
rect 10652 30920 10658 30932
rect 10689 30923 10747 30929
rect 10689 30920 10701 30923
rect 10652 30892 10701 30920
rect 10652 30880 10658 30892
rect 10689 30889 10701 30892
rect 10735 30889 10747 30923
rect 18233 30923 18291 30929
rect 18233 30920 18245 30923
rect 10689 30883 10747 30889
rect 17135 30892 18245 30920
rect 11974 30812 11980 30864
rect 12032 30852 12038 30864
rect 12342 30852 12348 30864
rect 12032 30824 12348 30852
rect 12032 30812 12038 30824
rect 12342 30812 12348 30824
rect 12400 30812 12406 30864
rect 11701 30787 11759 30793
rect 11701 30753 11713 30787
rect 11747 30784 11759 30787
rect 12710 30784 12716 30796
rect 11747 30756 12716 30784
rect 11747 30753 11759 30756
rect 11701 30747 11759 30753
rect 12710 30744 12716 30756
rect 12768 30744 12774 30796
rect 13998 30744 14004 30796
rect 14056 30784 14062 30796
rect 14093 30787 14151 30793
rect 14093 30784 14105 30787
rect 14056 30756 14105 30784
rect 14056 30744 14062 30756
rect 14093 30753 14105 30756
rect 14139 30753 14151 30787
rect 17135 30784 17163 30892
rect 18233 30889 18245 30892
rect 18279 30889 18291 30923
rect 18233 30883 18291 30889
rect 23658 30880 23664 30932
rect 23716 30920 23722 30932
rect 23753 30923 23811 30929
rect 23753 30920 23765 30923
rect 23716 30892 23765 30920
rect 23716 30880 23722 30892
rect 23753 30889 23765 30892
rect 23799 30920 23811 30923
rect 25961 30923 26019 30929
rect 23799 30892 25636 30920
rect 23799 30889 23811 30892
rect 23753 30883 23811 30889
rect 17954 30852 17960 30864
rect 17420 30824 17960 30852
rect 17420 30793 17448 30824
rect 17954 30812 17960 30824
rect 18012 30812 18018 30864
rect 21729 30855 21787 30861
rect 21729 30821 21741 30855
rect 21775 30852 21787 30855
rect 22830 30852 22836 30864
rect 21775 30824 22836 30852
rect 21775 30821 21787 30824
rect 21729 30815 21787 30821
rect 22830 30812 22836 30824
rect 22888 30812 22894 30864
rect 14093 30747 14151 30753
rect 17052 30756 17163 30784
rect 17313 30787 17371 30793
rect 9861 30719 9919 30725
rect 9861 30685 9873 30719
rect 9907 30716 9919 30719
rect 11422 30716 11428 30728
rect 9907 30688 11284 30716
rect 11383 30688 11428 30716
rect 9907 30685 9919 30688
rect 9861 30679 9919 30685
rect 10042 30608 10048 30660
rect 10100 30648 10106 30660
rect 10505 30651 10563 30657
rect 10505 30648 10517 30651
rect 10100 30620 10517 30648
rect 10100 30608 10106 30620
rect 10505 30617 10517 30620
rect 10551 30617 10563 30651
rect 11256 30648 11284 30688
rect 11422 30676 11428 30688
rect 11480 30676 11486 30728
rect 11517 30719 11575 30725
rect 11517 30685 11529 30719
rect 11563 30716 11575 30719
rect 11974 30716 11980 30728
rect 11563 30688 11980 30716
rect 11563 30685 11575 30688
rect 11517 30679 11575 30685
rect 11974 30676 11980 30688
rect 12032 30676 12038 30728
rect 12250 30716 12256 30728
rect 12211 30688 12256 30716
rect 12250 30676 12256 30688
rect 12308 30676 12314 30728
rect 13078 30716 13084 30728
rect 13039 30688 13084 30716
rect 13078 30676 13084 30688
rect 13136 30676 13142 30728
rect 14366 30716 14372 30728
rect 14327 30688 14372 30716
rect 14366 30676 14372 30688
rect 14424 30676 14430 30728
rect 17052 30725 17080 30756
rect 17313 30753 17325 30787
rect 17359 30753 17371 30787
rect 17313 30747 17371 30753
rect 17405 30787 17463 30793
rect 17405 30753 17417 30787
rect 17451 30753 17463 30787
rect 17405 30747 17463 30753
rect 17037 30719 17095 30725
rect 17037 30685 17049 30719
rect 17083 30685 17095 30719
rect 17209 30713 17267 30719
rect 17209 30710 17221 30713
rect 17037 30679 17095 30685
rect 17144 30682 17221 30710
rect 11701 30651 11759 30657
rect 11701 30648 11713 30651
rect 11256 30620 11713 30648
rect 10505 30611 10563 30617
rect 11701 30617 11713 30620
rect 11747 30648 11759 30651
rect 12066 30648 12072 30660
rect 11747 30620 12072 30648
rect 11747 30617 11759 30620
rect 11701 30611 11759 30617
rect 12066 30608 12072 30620
rect 12124 30608 12130 30660
rect 12434 30608 12440 30660
rect 12492 30648 12498 30660
rect 12897 30651 12955 30657
rect 12492 30620 12537 30648
rect 12492 30608 12498 30620
rect 12897 30617 12909 30651
rect 12943 30648 12955 30651
rect 16206 30648 16212 30660
rect 12943 30620 14228 30648
rect 12943 30617 12955 30620
rect 12897 30611 12955 30617
rect 9490 30540 9496 30592
rect 9548 30580 9554 30592
rect 9766 30580 9772 30592
rect 9548 30552 9772 30580
rect 9548 30540 9554 30552
rect 9766 30540 9772 30552
rect 9824 30540 9830 30592
rect 9953 30583 10011 30589
rect 9953 30549 9965 30583
rect 9999 30580 10011 30583
rect 10226 30580 10232 30592
rect 9999 30552 10232 30580
rect 9999 30549 10011 30552
rect 9953 30543 10011 30549
rect 10226 30540 10232 30552
rect 10284 30540 10290 30592
rect 10410 30540 10416 30592
rect 10468 30580 10474 30592
rect 10705 30583 10763 30589
rect 10705 30580 10717 30583
rect 10468 30552 10717 30580
rect 10468 30540 10474 30552
rect 10705 30549 10717 30552
rect 10751 30549 10763 30583
rect 10705 30543 10763 30549
rect 10873 30583 10931 30589
rect 10873 30549 10885 30583
rect 10919 30580 10931 30583
rect 11790 30580 11796 30592
rect 10919 30552 11796 30580
rect 10919 30549 10931 30552
rect 10873 30543 10931 30549
rect 11790 30540 11796 30552
rect 11848 30540 11854 30592
rect 12986 30540 12992 30592
rect 13044 30580 13050 30592
rect 13265 30583 13323 30589
rect 13265 30580 13277 30583
rect 13044 30552 13277 30580
rect 13044 30540 13050 30552
rect 13265 30549 13277 30552
rect 13311 30549 13323 30583
rect 14200 30580 14228 30620
rect 15120 30620 16212 30648
rect 15120 30580 15148 30620
rect 16206 30608 16212 30620
rect 16264 30608 16270 30660
rect 16850 30608 16856 30660
rect 16908 30648 16914 30660
rect 17144 30648 17172 30682
rect 17209 30679 17221 30682
rect 17255 30679 17267 30713
rect 17209 30673 17267 30679
rect 16908 30620 17172 30648
rect 16908 30608 16914 30620
rect 17328 30592 17356 30747
rect 17678 30744 17684 30796
rect 17736 30744 17742 30796
rect 18138 30744 18144 30796
rect 18196 30784 18202 30796
rect 19245 30787 19303 30793
rect 19245 30784 19257 30787
rect 18196 30756 19257 30784
rect 18196 30744 18202 30756
rect 19245 30753 19257 30756
rect 19291 30753 19303 30787
rect 20346 30784 20352 30796
rect 20307 30756 20352 30784
rect 19245 30747 19303 30753
rect 20346 30744 20352 30756
rect 20404 30744 20410 30796
rect 22002 30744 22008 30796
rect 22060 30784 22066 30796
rect 22465 30787 22523 30793
rect 22060 30756 22416 30784
rect 22060 30744 22066 30756
rect 17589 30719 17647 30725
rect 17589 30716 17601 30719
rect 17512 30688 17601 30716
rect 17512 30660 17540 30688
rect 17589 30685 17601 30688
rect 17635 30685 17647 30719
rect 17589 30679 17647 30685
rect 17494 30608 17500 30660
rect 17552 30608 17558 30660
rect 17696 30648 17724 30744
rect 18637 30719 18695 30725
rect 18637 30685 18649 30719
rect 18683 30716 18695 30719
rect 19334 30716 19340 30728
rect 18683 30688 19340 30716
rect 18683 30685 18695 30688
rect 18637 30679 18695 30685
rect 19334 30676 19340 30688
rect 19392 30716 19398 30728
rect 19618 30719 19676 30725
rect 19618 30716 19630 30719
rect 19392 30688 19630 30716
rect 19392 30676 19398 30688
rect 19618 30685 19630 30688
rect 19664 30685 19676 30719
rect 19618 30679 19676 30685
rect 20616 30719 20674 30725
rect 20616 30685 20628 30719
rect 20662 30716 20674 30719
rect 21358 30716 21364 30728
rect 20662 30688 21364 30716
rect 20662 30685 20674 30688
rect 20616 30679 20674 30685
rect 21358 30676 21364 30688
rect 21416 30676 21422 30728
rect 21450 30676 21456 30728
rect 21508 30716 21514 30728
rect 21910 30716 21916 30728
rect 21508 30688 21916 30716
rect 21508 30676 21514 30688
rect 21910 30676 21916 30688
rect 21968 30716 21974 30728
rect 22388 30725 22416 30756
rect 22465 30753 22477 30787
rect 22511 30784 22523 30787
rect 22511 30756 24716 30784
rect 22511 30753 22523 30756
rect 22465 30747 22523 30753
rect 22189 30719 22247 30725
rect 22189 30716 22201 30719
rect 21968 30688 22201 30716
rect 21968 30676 21974 30688
rect 22189 30685 22201 30688
rect 22235 30685 22247 30719
rect 22189 30679 22247 30685
rect 22373 30719 22431 30725
rect 22373 30685 22385 30719
rect 22419 30685 22431 30719
rect 22373 30679 22431 30685
rect 22554 30676 22560 30728
rect 22612 30716 22618 30728
rect 22741 30719 22799 30725
rect 22612 30688 22657 30716
rect 22612 30676 22618 30688
rect 22741 30685 22753 30719
rect 22787 30685 22799 30719
rect 23566 30716 23572 30728
rect 23527 30688 23572 30716
rect 22741 30679 22799 30685
rect 17604 30620 17724 30648
rect 14200 30552 15148 30580
rect 13265 30543 13323 30549
rect 15194 30540 15200 30592
rect 15252 30580 15258 30592
rect 15473 30583 15531 30589
rect 15473 30580 15485 30583
rect 15252 30552 15485 30580
rect 15252 30540 15258 30552
rect 15473 30549 15485 30552
rect 15519 30549 15531 30583
rect 15473 30543 15531 30549
rect 17310 30540 17316 30592
rect 17368 30580 17374 30592
rect 17604 30580 17632 30620
rect 17954 30608 17960 30660
rect 18012 30648 18018 30660
rect 18230 30648 18236 30660
rect 18012 30620 18236 30648
rect 18012 30608 18018 30620
rect 18230 30608 18236 30620
rect 18288 30608 18294 30660
rect 18414 30648 18420 30660
rect 18375 30620 18420 30648
rect 18414 30608 18420 30620
rect 18472 30608 18478 30660
rect 18509 30651 18567 30657
rect 18509 30617 18521 30651
rect 18555 30648 18567 30651
rect 18874 30648 18880 30660
rect 18555 30620 18880 30648
rect 18555 30617 18567 30620
rect 18509 30611 18567 30617
rect 18874 30608 18880 30620
rect 18932 30608 18938 30660
rect 19245 30651 19303 30657
rect 19245 30617 19257 30651
rect 19291 30617 19303 30651
rect 19245 30611 19303 30617
rect 19429 30651 19487 30657
rect 19429 30617 19441 30651
rect 19475 30617 19487 30651
rect 19429 30611 19487 30617
rect 19521 30651 19579 30657
rect 19521 30617 19533 30651
rect 19567 30648 19579 30651
rect 20438 30648 20444 30660
rect 19567 30620 20444 30648
rect 19567 30617 19579 30620
rect 19521 30611 19579 30617
rect 17770 30580 17776 30592
rect 17368 30552 17632 30580
rect 17731 30552 17776 30580
rect 17368 30540 17374 30552
rect 17770 30540 17776 30552
rect 17828 30540 17834 30592
rect 18248 30580 18276 30608
rect 19260 30580 19288 30611
rect 18248 30552 19288 30580
rect 19444 30580 19472 30611
rect 20438 30608 20444 30620
rect 20496 30608 20502 30660
rect 22756 30648 22784 30679
rect 23566 30676 23572 30688
rect 23624 30676 23630 30728
rect 24578 30716 24584 30728
rect 24539 30688 24584 30716
rect 24578 30676 24584 30688
rect 24636 30676 24642 30728
rect 24688 30716 24716 30756
rect 25608 30716 25636 30892
rect 25961 30889 25973 30923
rect 26007 30920 26019 30923
rect 26142 30920 26148 30932
rect 26007 30892 26148 30920
rect 26007 30889 26019 30892
rect 25961 30883 26019 30889
rect 26142 30880 26148 30892
rect 26200 30880 26206 30932
rect 29914 30920 29920 30932
rect 29875 30892 29920 30920
rect 29914 30880 29920 30892
rect 29972 30880 29978 30932
rect 30098 30920 30104 30932
rect 30059 30892 30104 30920
rect 30098 30880 30104 30892
rect 30156 30880 30162 30932
rect 26421 30719 26479 30725
rect 26421 30716 26433 30719
rect 24688 30688 25544 30716
rect 25608 30688 26433 30716
rect 23474 30648 23480 30660
rect 22756 30620 23480 30648
rect 23474 30608 23480 30620
rect 23532 30608 23538 30660
rect 24848 30651 24906 30657
rect 24848 30617 24860 30651
rect 24894 30648 24906 30651
rect 25130 30648 25136 30660
rect 24894 30620 25136 30648
rect 24894 30617 24906 30620
rect 24848 30611 24906 30617
rect 25130 30608 25136 30620
rect 25188 30608 25194 30660
rect 25516 30648 25544 30688
rect 26421 30685 26433 30688
rect 26467 30685 26479 30719
rect 26421 30679 26479 30685
rect 27065 30719 27123 30725
rect 27065 30685 27077 30719
rect 27111 30716 27123 30719
rect 28350 30716 28356 30728
rect 27111 30688 28356 30716
rect 27111 30685 27123 30688
rect 27065 30679 27123 30685
rect 28350 30676 28356 30688
rect 28408 30676 28414 30728
rect 28626 30676 28632 30728
rect 28684 30716 28690 30728
rect 29549 30719 29607 30725
rect 29549 30716 29561 30719
rect 28684 30688 29561 30716
rect 28684 30676 28690 30688
rect 29549 30685 29561 30688
rect 29595 30685 29607 30719
rect 29549 30679 29607 30685
rect 26510 30648 26516 30660
rect 25516 30620 26516 30648
rect 26510 30608 26516 30620
rect 26568 30608 26574 30660
rect 27332 30651 27390 30657
rect 27332 30617 27344 30651
rect 27378 30648 27390 30651
rect 27706 30648 27712 30660
rect 27378 30620 27712 30648
rect 27378 30617 27390 30620
rect 27332 30611 27390 30617
rect 27706 30608 27712 30620
rect 27764 30608 27770 30660
rect 19886 30580 19892 30592
rect 19444 30552 19892 30580
rect 19886 30540 19892 30552
rect 19944 30540 19950 30592
rect 22370 30540 22376 30592
rect 22428 30580 22434 30592
rect 22925 30583 22983 30589
rect 22925 30580 22937 30583
rect 22428 30552 22937 30580
rect 22428 30540 22434 30552
rect 22925 30549 22937 30552
rect 22971 30549 22983 30583
rect 22925 30543 22983 30549
rect 26605 30583 26663 30589
rect 26605 30549 26617 30583
rect 26651 30580 26663 30583
rect 28166 30580 28172 30592
rect 26651 30552 28172 30580
rect 26651 30549 26663 30552
rect 26605 30543 26663 30549
rect 28166 30540 28172 30552
rect 28224 30540 28230 30592
rect 28442 30580 28448 30592
rect 28355 30552 28448 30580
rect 28442 30540 28448 30552
rect 28500 30580 28506 30592
rect 29917 30583 29975 30589
rect 29917 30580 29929 30583
rect 28500 30552 29929 30580
rect 28500 30540 28506 30552
rect 29917 30549 29929 30552
rect 29963 30549 29975 30583
rect 29917 30543 29975 30549
rect 1104 30490 30820 30512
rect 1104 30438 10880 30490
rect 10932 30438 10944 30490
rect 10996 30438 11008 30490
rect 11060 30438 11072 30490
rect 11124 30438 11136 30490
rect 11188 30438 20811 30490
rect 20863 30438 20875 30490
rect 20927 30438 20939 30490
rect 20991 30438 21003 30490
rect 21055 30438 21067 30490
rect 21119 30438 30820 30490
rect 1104 30416 30820 30438
rect 8846 30336 8852 30388
rect 8904 30376 8910 30388
rect 8941 30379 8999 30385
rect 8941 30376 8953 30379
rect 8904 30348 8953 30376
rect 8904 30336 8910 30348
rect 8941 30345 8953 30348
rect 8987 30345 8999 30379
rect 8941 30339 8999 30345
rect 10318 30336 10324 30388
rect 10376 30376 10382 30388
rect 11238 30376 11244 30388
rect 10376 30348 11244 30376
rect 10376 30336 10382 30348
rect 11238 30336 11244 30348
rect 11296 30376 11302 30388
rect 12710 30376 12716 30388
rect 11296 30348 11744 30376
rect 12671 30348 12716 30376
rect 11296 30336 11302 30348
rect 9766 30268 9772 30320
rect 9824 30308 9830 30320
rect 9861 30311 9919 30317
rect 9861 30308 9873 30311
rect 9824 30280 9873 30308
rect 9824 30268 9830 30280
rect 9861 30277 9873 30280
rect 9907 30308 9919 30311
rect 9907 30280 11652 30308
rect 9907 30277 9919 30280
rect 9861 30271 9919 30277
rect 8846 30240 8852 30252
rect 8807 30212 8852 30240
rect 8846 30200 8852 30212
rect 8904 30200 8910 30252
rect 9033 30243 9091 30249
rect 9033 30209 9045 30243
rect 9079 30240 9091 30243
rect 9306 30240 9312 30252
rect 9079 30212 9312 30240
rect 9079 30209 9091 30212
rect 9033 30203 9091 30209
rect 9306 30200 9312 30212
rect 9364 30200 9370 30252
rect 10137 30243 10195 30249
rect 10137 30209 10149 30243
rect 10183 30240 10195 30243
rect 10226 30240 10232 30252
rect 10183 30212 10232 30240
rect 10183 30209 10195 30212
rect 10137 30203 10195 30209
rect 10226 30200 10232 30212
rect 10284 30200 10290 30252
rect 10318 30200 10324 30252
rect 10376 30240 10382 30252
rect 10376 30212 10421 30240
rect 10376 30200 10382 30212
rect 10502 30200 10508 30252
rect 10560 30240 10566 30252
rect 10597 30243 10655 30249
rect 10597 30240 10609 30243
rect 10560 30212 10609 30240
rect 10560 30200 10566 30212
rect 10597 30209 10609 30212
rect 10643 30209 10655 30243
rect 10597 30203 10655 30209
rect 11517 30243 11575 30249
rect 11517 30209 11529 30243
rect 11563 30209 11575 30243
rect 11517 30203 11575 30209
rect 10413 30175 10471 30181
rect 10413 30141 10425 30175
rect 10459 30172 10471 30175
rect 10459 30144 10640 30172
rect 10459 30141 10471 30144
rect 10413 30135 10471 30141
rect 10612 30116 10640 30144
rect 10594 30064 10600 30116
rect 10652 30064 10658 30116
rect 11532 30104 11560 30203
rect 11624 30172 11652 30280
rect 11716 30249 11744 30348
rect 12710 30336 12716 30348
rect 12768 30336 12774 30388
rect 12802 30336 12808 30388
rect 12860 30376 12866 30388
rect 25130 30376 25136 30388
rect 12860 30348 19334 30376
rect 25091 30348 25136 30376
rect 12860 30336 12866 30348
rect 12158 30268 12164 30320
rect 12216 30308 12222 30320
rect 12253 30311 12311 30317
rect 12253 30308 12265 30311
rect 12216 30280 12265 30308
rect 12216 30268 12222 30280
rect 12253 30277 12265 30280
rect 12299 30277 12311 30311
rect 12253 30271 12311 30277
rect 12618 30268 12624 30320
rect 12676 30308 12682 30320
rect 13081 30311 13139 30317
rect 13081 30308 13093 30311
rect 12676 30280 13093 30308
rect 12676 30268 12682 30280
rect 13081 30277 13093 30280
rect 13127 30277 13139 30311
rect 13081 30271 13139 30277
rect 16850 30268 16856 30320
rect 16908 30268 16914 30320
rect 16942 30268 16948 30320
rect 17000 30308 17006 30320
rect 17000 30280 17172 30308
rect 17000 30268 17006 30280
rect 11701 30243 11759 30249
rect 11701 30209 11713 30243
rect 11747 30209 11759 30243
rect 11882 30240 11888 30252
rect 11843 30212 11888 30240
rect 11701 30203 11759 30209
rect 11882 30200 11888 30212
rect 11940 30200 11946 30252
rect 12066 30240 12072 30252
rect 12027 30212 12072 30240
rect 12066 30200 12072 30212
rect 12124 30200 12130 30252
rect 14182 30200 14188 30252
rect 14240 30240 14246 30252
rect 14734 30249 14740 30252
rect 14461 30243 14519 30249
rect 14461 30240 14473 30243
rect 14240 30212 14473 30240
rect 14240 30200 14246 30212
rect 14461 30209 14473 30212
rect 14507 30209 14519 30243
rect 14461 30203 14519 30209
rect 14728 30203 14740 30249
rect 14792 30240 14798 30252
rect 16868 30240 16896 30268
rect 17037 30243 17095 30249
rect 17037 30240 17049 30243
rect 14792 30212 14828 30240
rect 16868 30212 17049 30240
rect 14734 30200 14740 30203
rect 14792 30200 14798 30212
rect 17037 30209 17049 30212
rect 17083 30209 17095 30243
rect 17144 30238 17172 30280
rect 18138 30268 18144 30320
rect 18196 30308 18202 30320
rect 18969 30311 19027 30317
rect 18969 30308 18981 30311
rect 18196 30280 18981 30308
rect 18196 30268 18202 30280
rect 18969 30277 18981 30280
rect 19015 30277 19027 30311
rect 19306 30308 19334 30348
rect 25130 30336 25136 30348
rect 25188 30336 25194 30388
rect 28350 30376 28356 30388
rect 28311 30348 28356 30376
rect 28350 30336 28356 30348
rect 28408 30336 28414 30388
rect 19306 30280 20852 30308
rect 18969 30271 19027 30277
rect 17221 30243 17279 30249
rect 17221 30238 17233 30243
rect 17144 30210 17233 30238
rect 17037 30203 17095 30209
rect 17221 30209 17233 30210
rect 17267 30209 17279 30243
rect 17221 30203 17279 30209
rect 17310 30200 17316 30252
rect 17368 30240 17374 30252
rect 17586 30240 17592 30252
rect 17368 30212 17413 30240
rect 17547 30212 17592 30240
rect 17368 30200 17374 30212
rect 17586 30200 17592 30212
rect 17644 30200 17650 30252
rect 18230 30240 18236 30252
rect 18191 30212 18236 30240
rect 18230 30200 18236 30212
rect 18288 30200 18294 30252
rect 18417 30243 18475 30249
rect 18417 30209 18429 30243
rect 18463 30240 18475 30243
rect 18690 30240 18696 30252
rect 18463 30212 18696 30240
rect 18463 30209 18475 30212
rect 18417 30203 18475 30209
rect 18690 30200 18696 30212
rect 18748 30200 18754 30252
rect 18782 30200 18788 30252
rect 18840 30240 18846 30252
rect 19429 30243 19487 30249
rect 18840 30212 18885 30240
rect 18840 30200 18846 30212
rect 19429 30209 19441 30243
rect 19475 30240 19487 30243
rect 19518 30240 19524 30252
rect 19475 30212 19524 30240
rect 19475 30209 19487 30212
rect 19429 30203 19487 30209
rect 19518 30200 19524 30212
rect 19576 30240 19582 30252
rect 19794 30240 19800 30252
rect 19576 30212 19800 30240
rect 19576 30200 19582 30212
rect 19794 30200 19800 30212
rect 19852 30200 19858 30252
rect 20714 30240 20720 30252
rect 20675 30212 20720 30240
rect 20714 30200 20720 30212
rect 20772 30200 20778 30252
rect 20824 30240 20852 30280
rect 21358 30268 21364 30320
rect 21416 30308 21422 30320
rect 21726 30308 21732 30320
rect 21416 30280 21732 30308
rect 21416 30268 21422 30280
rect 21726 30268 21732 30280
rect 21784 30268 21790 30320
rect 22370 30317 22376 30320
rect 22364 30308 22376 30317
rect 22331 30280 22376 30308
rect 22364 30271 22376 30280
rect 22370 30268 22376 30271
rect 22428 30268 22434 30320
rect 23750 30268 23756 30320
rect 23808 30308 23814 30320
rect 23808 30280 24624 30308
rect 23808 30268 23814 30280
rect 24118 30240 24124 30252
rect 20824 30212 24124 30240
rect 24118 30200 24124 30212
rect 24176 30200 24182 30252
rect 24210 30200 24216 30252
rect 24268 30240 24274 30252
rect 24596 30249 24624 30280
rect 25682 30268 25688 30320
rect 25740 30308 25746 30320
rect 27706 30308 27712 30320
rect 25740 30280 27292 30308
rect 27667 30280 27712 30308
rect 25740 30268 25746 30280
rect 24397 30243 24455 30249
rect 24397 30240 24409 30243
rect 24268 30212 24409 30240
rect 24268 30200 24274 30212
rect 24397 30209 24409 30212
rect 24443 30209 24455 30243
rect 24397 30203 24455 30209
rect 24581 30243 24639 30249
rect 24581 30209 24593 30243
rect 24627 30209 24639 30243
rect 24581 30203 24639 30209
rect 24673 30243 24731 30249
rect 24673 30209 24685 30243
rect 24719 30240 24731 30243
rect 24854 30240 24860 30252
rect 24719 30212 24860 30240
rect 24719 30209 24731 30212
rect 24673 30203 24731 30209
rect 11793 30175 11851 30181
rect 11793 30172 11805 30175
rect 11624 30144 11805 30172
rect 11793 30141 11805 30144
rect 11839 30141 11851 30175
rect 11793 30135 11851 30141
rect 13173 30175 13231 30181
rect 13173 30141 13185 30175
rect 13219 30172 13231 30175
rect 13262 30172 13268 30184
rect 13219 30144 13268 30172
rect 13219 30141 13231 30144
rect 13173 30135 13231 30141
rect 13262 30132 13268 30144
rect 13320 30132 13326 30184
rect 13357 30175 13415 30181
rect 13357 30141 13369 30175
rect 13403 30172 13415 30175
rect 13630 30172 13636 30184
rect 13403 30144 13636 30172
rect 13403 30141 13415 30144
rect 13357 30135 13415 30141
rect 13630 30132 13636 30144
rect 13688 30132 13694 30184
rect 16758 30132 16764 30184
rect 16816 30172 16822 30184
rect 17405 30175 17463 30181
rect 17405 30172 17417 30175
rect 16816 30144 17417 30172
rect 16816 30132 16822 30144
rect 17405 30141 17417 30144
rect 17451 30172 17463 30175
rect 18509 30175 18567 30181
rect 18509 30172 18521 30175
rect 17451 30144 18521 30172
rect 17451 30141 17463 30144
rect 17405 30135 17463 30141
rect 18509 30141 18521 30144
rect 18555 30141 18567 30175
rect 18509 30135 18567 30141
rect 18601 30175 18659 30181
rect 18601 30141 18613 30175
rect 18647 30141 18659 30175
rect 18601 30135 18659 30141
rect 12710 30104 12716 30116
rect 11532 30076 12716 30104
rect 12710 30064 12716 30076
rect 12768 30064 12774 30116
rect 18616 30104 18644 30135
rect 19242 30132 19248 30184
rect 19300 30172 19306 30184
rect 20162 30172 20168 30184
rect 19300 30144 20168 30172
rect 19300 30132 19306 30144
rect 20162 30132 20168 30144
rect 20220 30132 20226 30184
rect 20254 30132 20260 30184
rect 20312 30172 20318 30184
rect 22097 30175 22155 30181
rect 22097 30172 22109 30175
rect 20312 30144 22109 30172
rect 20312 30132 20318 30144
rect 22097 30141 22109 30144
rect 22143 30141 22155 30175
rect 22097 30135 22155 30141
rect 18524 30076 18644 30104
rect 18524 30048 18552 30076
rect 19426 30064 19432 30116
rect 19484 30104 19490 30116
rect 19613 30107 19671 30113
rect 19613 30104 19625 30107
rect 19484 30076 19625 30104
rect 19484 30064 19490 30076
rect 19613 30073 19625 30076
rect 19659 30104 19671 30107
rect 20438 30104 20444 30116
rect 19659 30076 20444 30104
rect 19659 30073 19671 30076
rect 19613 30067 19671 30073
rect 20438 30064 20444 30076
rect 20496 30064 20502 30116
rect 24412 30104 24440 30203
rect 24854 30200 24860 30212
rect 24912 30200 24918 30252
rect 24949 30243 25007 30249
rect 24949 30209 24961 30243
rect 24995 30240 25007 30243
rect 26142 30240 26148 30252
rect 24995 30212 26148 30240
rect 24995 30209 25007 30212
rect 24949 30203 25007 30209
rect 26142 30200 26148 30212
rect 26200 30200 26206 30252
rect 26418 30200 26424 30252
rect 26476 30240 26482 30252
rect 26973 30243 27031 30249
rect 26973 30240 26985 30243
rect 26476 30212 26985 30240
rect 26476 30200 26482 30212
rect 26973 30209 26985 30212
rect 27019 30209 27031 30243
rect 26973 30203 27031 30209
rect 27062 30200 27068 30252
rect 27120 30240 27126 30252
rect 27264 30249 27292 30280
rect 27706 30268 27712 30280
rect 27764 30268 27770 30320
rect 28442 30308 28448 30320
rect 28000 30280 28448 30308
rect 27157 30243 27215 30249
rect 27157 30240 27169 30243
rect 27120 30212 27169 30240
rect 27120 30200 27126 30212
rect 27157 30209 27169 30212
rect 27203 30209 27215 30243
rect 27157 30203 27215 30209
rect 27249 30243 27307 30249
rect 27249 30209 27261 30243
rect 27295 30209 27307 30243
rect 27249 30203 27307 30209
rect 27525 30243 27583 30249
rect 27525 30209 27537 30243
rect 27571 30240 27583 30243
rect 28000 30240 28028 30280
rect 28442 30268 28448 30280
rect 28500 30268 28506 30320
rect 28166 30240 28172 30252
rect 27571 30212 28028 30240
rect 28127 30212 28172 30240
rect 27571 30209 27583 30212
rect 27525 30203 27583 30209
rect 28166 30200 28172 30212
rect 28224 30200 28230 30252
rect 28994 30200 29000 30252
rect 29052 30240 29058 30252
rect 29365 30243 29423 30249
rect 29365 30240 29377 30243
rect 29052 30212 29377 30240
rect 29052 30200 29058 30212
rect 29365 30209 29377 30212
rect 29411 30209 29423 30243
rect 29365 30203 29423 30209
rect 29825 30243 29883 30249
rect 29825 30209 29837 30243
rect 29871 30209 29883 30243
rect 29825 30203 29883 30209
rect 24762 30172 24768 30184
rect 24723 30144 24768 30172
rect 24762 30132 24768 30144
rect 24820 30172 24826 30184
rect 25593 30175 25651 30181
rect 25593 30172 25605 30175
rect 24820 30144 25605 30172
rect 24820 30132 24826 30144
rect 25593 30141 25605 30144
rect 25639 30141 25651 30175
rect 25593 30135 25651 30141
rect 25869 30175 25927 30181
rect 25869 30141 25881 30175
rect 25915 30172 25927 30175
rect 26786 30172 26792 30184
rect 25915 30144 26792 30172
rect 25915 30141 25927 30144
rect 25869 30135 25927 30141
rect 26786 30132 26792 30144
rect 26844 30172 26850 30184
rect 27341 30175 27399 30181
rect 27341 30172 27353 30175
rect 26844 30144 27353 30172
rect 26844 30132 26850 30144
rect 27341 30141 27353 30144
rect 27387 30141 27399 30175
rect 29840 30172 29868 30203
rect 27341 30135 27399 30141
rect 29196 30144 29868 30172
rect 26418 30104 26424 30116
rect 24412 30076 26424 30104
rect 26418 30064 26424 30076
rect 26476 30064 26482 30116
rect 29196 30113 29224 30144
rect 29181 30107 29239 30113
rect 29181 30073 29193 30107
rect 29227 30073 29239 30107
rect 29181 30067 29239 30073
rect 10229 30039 10287 30045
rect 10229 30005 10241 30039
rect 10275 30036 10287 30039
rect 11974 30036 11980 30048
rect 10275 30008 11980 30036
rect 10275 30005 10287 30008
rect 10229 29999 10287 30005
rect 11974 29996 11980 30008
rect 12032 29996 12038 30048
rect 13538 29996 13544 30048
rect 13596 30036 13602 30048
rect 15194 30036 15200 30048
rect 13596 30008 15200 30036
rect 13596 29996 13602 30008
rect 15194 29996 15200 30008
rect 15252 29996 15258 30048
rect 15470 29996 15476 30048
rect 15528 30036 15534 30048
rect 15841 30039 15899 30045
rect 15841 30036 15853 30039
rect 15528 30008 15853 30036
rect 15528 29996 15534 30008
rect 15841 30005 15853 30008
rect 15887 30005 15899 30039
rect 15841 29999 15899 30005
rect 16942 29996 16948 30048
rect 17000 30036 17006 30048
rect 17773 30039 17831 30045
rect 17773 30036 17785 30039
rect 17000 30008 17785 30036
rect 17000 29996 17006 30008
rect 17773 30005 17785 30008
rect 17819 30005 17831 30039
rect 17773 29999 17831 30005
rect 17862 29996 17868 30048
rect 17920 30036 17926 30048
rect 18506 30036 18512 30048
rect 17920 30008 18512 30036
rect 17920 29996 17926 30008
rect 18506 29996 18512 30008
rect 18564 29996 18570 30048
rect 20070 29996 20076 30048
rect 20128 30036 20134 30048
rect 20901 30039 20959 30045
rect 20901 30036 20913 30039
rect 20128 30008 20913 30036
rect 20128 29996 20134 30008
rect 20901 30005 20913 30008
rect 20947 30005 20959 30039
rect 23474 30036 23480 30048
rect 23435 30008 23480 30036
rect 20901 29999 20959 30005
rect 23474 29996 23480 30008
rect 23532 29996 23538 30048
rect 23842 29996 23848 30048
rect 23900 30036 23906 30048
rect 28074 30036 28080 30048
rect 23900 30008 28080 30036
rect 23900 29996 23906 30008
rect 28074 29996 28080 30008
rect 28132 29996 28138 30048
rect 30006 30036 30012 30048
rect 29967 30008 30012 30036
rect 30006 29996 30012 30008
rect 30064 29996 30070 30048
rect 1104 29946 30820 29968
rect 1104 29894 5915 29946
rect 5967 29894 5979 29946
rect 6031 29894 6043 29946
rect 6095 29894 6107 29946
rect 6159 29894 6171 29946
rect 6223 29894 15846 29946
rect 15898 29894 15910 29946
rect 15962 29894 15974 29946
rect 16026 29894 16038 29946
rect 16090 29894 16102 29946
rect 16154 29894 25776 29946
rect 25828 29894 25840 29946
rect 25892 29894 25904 29946
rect 25956 29894 25968 29946
rect 26020 29894 26032 29946
rect 26084 29894 30820 29946
rect 1104 29872 30820 29894
rect 8846 29792 8852 29844
rect 8904 29832 8910 29844
rect 9401 29835 9459 29841
rect 9401 29832 9413 29835
rect 8904 29804 9413 29832
rect 8904 29792 8910 29804
rect 9401 29801 9413 29804
rect 9447 29801 9459 29835
rect 11514 29832 11520 29844
rect 9401 29795 9459 29801
rect 11164 29804 11520 29832
rect 9953 29699 10011 29705
rect 9953 29665 9965 29699
rect 9999 29696 10011 29699
rect 10226 29696 10232 29708
rect 9999 29668 10232 29696
rect 9999 29665 10011 29668
rect 9953 29659 10011 29665
rect 10226 29656 10232 29668
rect 10284 29696 10290 29708
rect 10686 29696 10692 29708
rect 10284 29668 10692 29696
rect 10284 29656 10290 29668
rect 10686 29656 10692 29668
rect 10744 29656 10750 29708
rect 8205 29631 8263 29637
rect 8205 29597 8217 29631
rect 8251 29597 8263 29631
rect 8205 29591 8263 29597
rect 8389 29631 8447 29637
rect 8389 29597 8401 29631
rect 8435 29628 8447 29631
rect 9306 29628 9312 29640
rect 8435 29600 9312 29628
rect 8435 29597 8447 29600
rect 8389 29591 8447 29597
rect 8220 29560 8248 29591
rect 9306 29588 9312 29600
rect 9364 29588 9370 29640
rect 9582 29588 9588 29640
rect 9640 29628 9646 29640
rect 10042 29628 10048 29640
rect 9640 29600 9682 29628
rect 10003 29600 10048 29628
rect 9640 29588 9646 29600
rect 10042 29588 10048 29600
rect 10100 29588 10106 29640
rect 10505 29631 10563 29637
rect 10505 29597 10517 29631
rect 10551 29628 10563 29631
rect 10594 29628 10600 29640
rect 10551 29600 10600 29628
rect 10551 29597 10563 29600
rect 10505 29591 10563 29597
rect 10594 29588 10600 29600
rect 10652 29588 10658 29640
rect 11164 29637 11192 29804
rect 11514 29792 11520 29804
rect 11572 29792 11578 29844
rect 13541 29835 13599 29841
rect 13541 29801 13553 29835
rect 13587 29832 13599 29835
rect 14366 29832 14372 29844
rect 13587 29804 14372 29832
rect 13587 29801 13599 29804
rect 13541 29795 13599 29801
rect 14366 29792 14372 29804
rect 14424 29792 14430 29844
rect 14734 29792 14740 29844
rect 14792 29832 14798 29844
rect 14921 29835 14979 29841
rect 14921 29832 14933 29835
rect 14792 29804 14933 29832
rect 14792 29792 14798 29804
rect 14921 29801 14933 29804
rect 14967 29801 14979 29835
rect 14921 29795 14979 29801
rect 15289 29835 15347 29841
rect 15289 29801 15301 29835
rect 15335 29832 15347 29835
rect 15378 29832 15384 29844
rect 15335 29804 15384 29832
rect 15335 29801 15347 29804
rect 15289 29795 15347 29801
rect 15378 29792 15384 29804
rect 15436 29792 15442 29844
rect 16482 29792 16488 29844
rect 16540 29832 16546 29844
rect 18782 29832 18788 29844
rect 16540 29804 18788 29832
rect 16540 29792 16546 29804
rect 18782 29792 18788 29804
rect 18840 29792 18846 29844
rect 19702 29832 19708 29844
rect 19663 29804 19708 29832
rect 19702 29792 19708 29804
rect 19760 29792 19766 29844
rect 21683 29835 21741 29841
rect 21683 29801 21695 29835
rect 21729 29832 21741 29835
rect 22554 29832 22560 29844
rect 21729 29804 22560 29832
rect 21729 29801 21741 29804
rect 21683 29795 21741 29801
rect 22554 29792 22560 29804
rect 22612 29792 22618 29844
rect 23109 29835 23167 29841
rect 23109 29801 23121 29835
rect 23155 29832 23167 29835
rect 24578 29832 24584 29844
rect 23155 29804 24584 29832
rect 23155 29801 23167 29804
rect 23109 29795 23167 29801
rect 24578 29792 24584 29804
rect 24636 29792 24642 29844
rect 27338 29832 27344 29844
rect 24780 29804 25268 29832
rect 24780 29776 24808 29804
rect 11422 29724 11428 29776
rect 11480 29724 11486 29776
rect 11885 29767 11943 29773
rect 11885 29733 11897 29767
rect 11931 29764 11943 29767
rect 12802 29764 12808 29776
rect 11931 29736 12808 29764
rect 11931 29733 11943 29736
rect 11885 29727 11943 29733
rect 12802 29724 12808 29736
rect 12860 29724 12866 29776
rect 16656 29736 18276 29764
rect 11440 29696 11468 29724
rect 15381 29699 15439 29705
rect 11440 29668 11744 29696
rect 11149 29631 11207 29637
rect 11149 29597 11161 29631
rect 11195 29597 11207 29631
rect 11330 29628 11336 29640
rect 11291 29600 11336 29628
rect 11149 29591 11207 29597
rect 11330 29588 11336 29600
rect 11388 29588 11394 29640
rect 11716 29637 11744 29668
rect 13188 29668 14136 29696
rect 13188 29640 13216 29668
rect 11422 29631 11480 29637
rect 11422 29597 11434 29631
rect 11468 29597 11480 29631
rect 11422 29591 11480 29597
rect 11517 29631 11575 29637
rect 11517 29597 11529 29631
rect 11563 29597 11575 29631
rect 11517 29591 11575 29597
rect 11701 29631 11759 29637
rect 11701 29597 11713 29631
rect 11747 29628 11759 29631
rect 12066 29628 12072 29640
rect 11747 29600 12072 29628
rect 11747 29597 11759 29600
rect 11701 29591 11759 29597
rect 9858 29560 9864 29572
rect 8220 29532 9864 29560
rect 9858 29520 9864 29532
rect 9916 29520 9922 29572
rect 11440 29504 11468 29591
rect 11532 29560 11560 29591
rect 12066 29588 12072 29600
rect 12124 29588 12130 29640
rect 12897 29631 12955 29637
rect 12897 29597 12909 29631
rect 12943 29597 12955 29631
rect 12897 29591 12955 29597
rect 11974 29560 11980 29572
rect 11532 29532 11980 29560
rect 11974 29520 11980 29532
rect 12032 29520 12038 29572
rect 8297 29495 8355 29501
rect 8297 29461 8309 29495
rect 8343 29492 8355 29495
rect 8386 29492 8392 29504
rect 8343 29464 8392 29492
rect 8343 29461 8355 29464
rect 8297 29455 8355 29461
rect 8386 29452 8392 29464
rect 8444 29452 8450 29504
rect 9585 29495 9643 29501
rect 9585 29461 9597 29495
rect 9631 29492 9643 29495
rect 9766 29492 9772 29504
rect 9631 29464 9772 29492
rect 9631 29461 9643 29464
rect 9585 29455 9643 29461
rect 9766 29452 9772 29464
rect 9824 29452 9830 29504
rect 10597 29495 10655 29501
rect 10597 29461 10609 29495
rect 10643 29492 10655 29495
rect 10778 29492 10784 29504
rect 10643 29464 10784 29492
rect 10643 29461 10655 29464
rect 10597 29455 10655 29461
rect 10778 29452 10784 29464
rect 10836 29452 10842 29504
rect 11422 29452 11428 29504
rect 11480 29452 11486 29504
rect 12912 29492 12940 29591
rect 12986 29588 12992 29640
rect 13044 29628 13050 29640
rect 13044 29600 13089 29628
rect 13044 29588 13050 29600
rect 13170 29588 13176 29640
rect 13228 29628 13234 29640
rect 14108 29637 14136 29668
rect 15381 29665 15393 29699
rect 15427 29696 15439 29699
rect 15470 29696 15476 29708
rect 15427 29668 15476 29696
rect 15427 29665 15439 29668
rect 15381 29659 15439 29665
rect 15470 29656 15476 29668
rect 15528 29656 15534 29708
rect 13403 29631 13461 29637
rect 13228 29600 13321 29628
rect 13228 29588 13234 29600
rect 13403 29597 13415 29631
rect 13449 29628 13461 29631
rect 14093 29631 14151 29637
rect 13449 29600 13860 29628
rect 13449 29597 13461 29600
rect 13403 29591 13461 29597
rect 13265 29563 13323 29569
rect 13265 29529 13277 29563
rect 13311 29560 13323 29563
rect 13538 29560 13544 29572
rect 13311 29532 13544 29560
rect 13311 29529 13323 29532
rect 13265 29523 13323 29529
rect 13538 29520 13544 29532
rect 13596 29520 13602 29572
rect 13832 29560 13860 29600
rect 14093 29597 14105 29631
rect 14139 29597 14151 29631
rect 14093 29591 14151 29597
rect 15105 29631 15163 29637
rect 15105 29597 15117 29631
rect 15151 29628 15163 29631
rect 15562 29628 15568 29640
rect 15151 29600 15568 29628
rect 15151 29597 15163 29600
rect 15105 29591 15163 29597
rect 15562 29588 15568 29600
rect 15620 29588 15626 29640
rect 15654 29588 15660 29640
rect 15712 29628 15718 29640
rect 15841 29631 15899 29637
rect 15841 29628 15853 29631
rect 15712 29600 15853 29628
rect 15712 29588 15718 29600
rect 15841 29597 15853 29600
rect 15887 29597 15899 29631
rect 16022 29628 16028 29640
rect 15983 29600 16028 29628
rect 15841 29591 15899 29597
rect 16022 29588 16028 29600
rect 16080 29588 16086 29640
rect 16114 29588 16120 29640
rect 16172 29628 16178 29640
rect 16656 29639 16684 29736
rect 16853 29699 16911 29705
rect 16853 29665 16865 29699
rect 16899 29696 16911 29699
rect 17862 29696 17868 29708
rect 16899 29668 17868 29696
rect 16899 29665 16911 29668
rect 16853 29659 16911 29665
rect 17862 29656 17868 29668
rect 17920 29656 17926 29708
rect 16485 29631 16543 29637
rect 16485 29628 16497 29631
rect 16172 29600 16497 29628
rect 16172 29588 16178 29600
rect 16485 29597 16497 29600
rect 16531 29597 16543 29631
rect 16485 29591 16543 29597
rect 16641 29633 16699 29639
rect 16641 29599 16653 29633
rect 16687 29599 16699 29633
rect 16641 29593 16699 29599
rect 16758 29588 16764 29640
rect 16816 29628 16822 29640
rect 17037 29631 17095 29637
rect 16816 29600 16861 29628
rect 16816 29588 16822 29600
rect 17037 29597 17049 29631
rect 17083 29597 17095 29631
rect 17221 29631 17279 29637
rect 17221 29628 17233 29631
rect 17037 29591 17095 29597
rect 17135 29600 17233 29628
rect 14185 29563 14243 29569
rect 14185 29560 14197 29563
rect 13832 29532 14197 29560
rect 14185 29529 14197 29532
rect 14231 29529 14243 29563
rect 14185 29523 14243 29529
rect 14918 29520 14924 29572
rect 14976 29560 14982 29572
rect 17052 29560 17080 29591
rect 14976 29532 17080 29560
rect 14976 29520 14982 29532
rect 14090 29492 14096 29504
rect 12912 29464 14096 29492
rect 14090 29452 14096 29464
rect 14148 29452 14154 29504
rect 15194 29452 15200 29504
rect 15252 29492 15258 29504
rect 15933 29495 15991 29501
rect 15933 29492 15945 29495
rect 15252 29464 15945 29492
rect 15252 29452 15258 29464
rect 15933 29461 15945 29464
rect 15979 29461 15991 29495
rect 15933 29455 15991 29461
rect 16850 29452 16856 29504
rect 16908 29492 16914 29504
rect 17135 29492 17163 29600
rect 17221 29597 17233 29600
rect 17267 29597 17279 29631
rect 17221 29591 17279 29597
rect 17957 29631 18015 29637
rect 17957 29597 17969 29631
rect 18003 29628 18015 29631
rect 18138 29628 18144 29640
rect 18003 29600 18144 29628
rect 18003 29597 18015 29600
rect 17957 29591 18015 29597
rect 18138 29588 18144 29600
rect 18196 29588 18202 29640
rect 18049 29563 18107 29569
rect 18049 29560 18061 29563
rect 17236 29532 18061 29560
rect 17236 29504 17264 29532
rect 18049 29529 18061 29532
rect 18095 29529 18107 29563
rect 18049 29523 18107 29529
rect 16908 29464 17163 29492
rect 16908 29452 16914 29464
rect 17218 29452 17224 29504
rect 17276 29452 17282 29504
rect 18248 29492 18276 29736
rect 19150 29724 19156 29776
rect 19208 29764 19214 29776
rect 24762 29764 24768 29776
rect 19208 29736 24768 29764
rect 19208 29724 19214 29736
rect 24762 29724 24768 29736
rect 24820 29724 24826 29776
rect 24854 29724 24860 29776
rect 24912 29764 24918 29776
rect 24912 29736 25176 29764
rect 24912 29724 24918 29736
rect 23842 29696 23848 29708
rect 23803 29668 23848 29696
rect 23842 29656 23848 29668
rect 23900 29656 23906 29708
rect 24946 29656 24952 29708
rect 25004 29656 25010 29708
rect 25148 29705 25176 29736
rect 25240 29705 25268 29804
rect 25424 29804 27344 29832
rect 25133 29699 25191 29705
rect 25133 29665 25145 29699
rect 25179 29665 25191 29699
rect 25133 29659 25191 29665
rect 25225 29699 25283 29705
rect 25225 29665 25237 29699
rect 25271 29665 25283 29699
rect 25225 29659 25283 29665
rect 19426 29588 19432 29640
rect 19484 29628 19490 29640
rect 19521 29631 19579 29637
rect 19521 29628 19533 29631
rect 19484 29600 19533 29628
rect 19484 29588 19490 29600
rect 19521 29597 19533 29600
rect 19567 29597 19579 29631
rect 19521 29591 19579 29597
rect 20165 29631 20223 29637
rect 20165 29597 20177 29631
rect 20211 29628 20223 29631
rect 20346 29628 20352 29640
rect 20211 29600 20352 29628
rect 20211 29597 20223 29600
rect 20165 29591 20223 29597
rect 20346 29588 20352 29600
rect 20404 29588 20410 29640
rect 20809 29631 20867 29637
rect 20809 29597 20821 29631
rect 20855 29628 20867 29631
rect 21266 29628 21272 29640
rect 20855 29600 21272 29628
rect 20855 29597 20867 29600
rect 20809 29591 20867 29597
rect 21266 29588 21272 29600
rect 21324 29588 21330 29640
rect 21453 29631 21511 29637
rect 21453 29597 21465 29631
rect 21499 29597 21511 29631
rect 22922 29628 22928 29640
rect 22883 29600 22928 29628
rect 21453 29591 21511 29597
rect 21358 29560 21364 29572
rect 19444 29532 21364 29560
rect 19444 29492 19472 29532
rect 21358 29520 21364 29532
rect 21416 29520 21422 29572
rect 18248 29464 19472 29492
rect 19518 29452 19524 29504
rect 19576 29492 19582 29504
rect 20349 29495 20407 29501
rect 20349 29492 20361 29495
rect 19576 29464 20361 29492
rect 19576 29452 19582 29464
rect 20349 29461 20361 29464
rect 20395 29492 20407 29495
rect 20714 29492 20720 29504
rect 20395 29464 20720 29492
rect 20395 29461 20407 29464
rect 20349 29455 20407 29461
rect 20714 29452 20720 29464
rect 20772 29452 20778 29504
rect 20901 29495 20959 29501
rect 20901 29461 20913 29495
rect 20947 29492 20959 29495
rect 21468 29492 21496 29591
rect 22922 29588 22928 29600
rect 22980 29588 22986 29640
rect 24670 29588 24676 29640
rect 24728 29628 24734 29640
rect 24857 29631 24915 29637
rect 24857 29628 24869 29631
rect 24728 29600 24869 29628
rect 24728 29588 24734 29600
rect 24857 29597 24869 29600
rect 24903 29597 24915 29631
rect 24964 29628 24992 29656
rect 25424 29637 25452 29804
rect 27338 29792 27344 29804
rect 27396 29792 27402 29844
rect 28813 29835 28871 29841
rect 28813 29801 28825 29835
rect 28859 29801 28871 29835
rect 28994 29832 29000 29844
rect 28955 29804 29000 29832
rect 28813 29795 28871 29801
rect 28828 29764 28856 29795
rect 28994 29792 29000 29804
rect 29052 29792 29058 29844
rect 30009 29835 30067 29841
rect 30009 29801 30021 29835
rect 30055 29832 30067 29835
rect 30098 29832 30104 29844
rect 30055 29804 30104 29832
rect 30055 29801 30067 29804
rect 30009 29795 30067 29801
rect 30098 29792 30104 29804
rect 30156 29792 30162 29844
rect 29086 29764 29092 29776
rect 28828 29736 29092 29764
rect 29086 29724 29092 29736
rect 29144 29724 29150 29776
rect 25041 29631 25099 29637
rect 25041 29628 25053 29631
rect 24964 29600 25053 29628
rect 24857 29591 24915 29597
rect 25041 29597 25053 29600
rect 25087 29597 25099 29631
rect 25041 29591 25099 29597
rect 25409 29631 25467 29637
rect 25409 29597 25421 29631
rect 25455 29597 25467 29631
rect 25409 29591 25467 29597
rect 26053 29631 26111 29637
rect 26053 29597 26065 29631
rect 26099 29628 26111 29631
rect 27154 29628 27160 29640
rect 26099 29600 27160 29628
rect 26099 29597 26111 29600
rect 26053 29591 26111 29597
rect 23661 29563 23719 29569
rect 23661 29529 23673 29563
rect 23707 29560 23719 29563
rect 24946 29560 24952 29572
rect 23707 29532 24952 29560
rect 23707 29529 23719 29532
rect 23661 29523 23719 29529
rect 24946 29520 24952 29532
rect 25004 29520 25010 29572
rect 25056 29504 25084 29591
rect 27154 29588 27160 29600
rect 27212 29588 27218 29640
rect 28445 29631 28503 29637
rect 28445 29597 28457 29631
rect 28491 29628 28503 29631
rect 28626 29628 28632 29640
rect 28491 29600 28632 29628
rect 28491 29597 28503 29600
rect 28445 29591 28503 29597
rect 28626 29588 28632 29600
rect 28684 29588 28690 29640
rect 29822 29628 29828 29640
rect 29783 29600 29828 29628
rect 29822 29588 29828 29600
rect 29880 29588 29886 29640
rect 25498 29520 25504 29572
rect 25556 29560 25562 29572
rect 26298 29563 26356 29569
rect 26298 29560 26310 29563
rect 25556 29532 26310 29560
rect 25556 29520 25562 29532
rect 26298 29529 26310 29532
rect 26344 29529 26356 29563
rect 26298 29523 26356 29529
rect 27338 29520 27344 29572
rect 27396 29560 27402 29572
rect 28813 29563 28871 29569
rect 28813 29560 28825 29563
rect 27396 29532 28825 29560
rect 27396 29520 27402 29532
rect 28813 29529 28825 29532
rect 28859 29529 28871 29563
rect 28813 29523 28871 29529
rect 21726 29492 21732 29504
rect 20947 29464 21732 29492
rect 20947 29461 20959 29464
rect 20901 29455 20959 29461
rect 21726 29452 21732 29464
rect 21784 29452 21790 29504
rect 22738 29452 22744 29504
rect 22796 29492 22802 29504
rect 23750 29492 23756 29504
rect 22796 29464 23756 29492
rect 22796 29452 22802 29464
rect 23750 29452 23756 29464
rect 23808 29452 23814 29504
rect 25038 29452 25044 29504
rect 25096 29452 25102 29504
rect 25593 29495 25651 29501
rect 25593 29461 25605 29495
rect 25639 29492 25651 29495
rect 26418 29492 26424 29504
rect 25639 29464 26424 29492
rect 25639 29461 25651 29464
rect 25593 29455 25651 29461
rect 26418 29452 26424 29464
rect 26476 29452 26482 29504
rect 27430 29492 27436 29504
rect 27391 29464 27436 29492
rect 27430 29452 27436 29464
rect 27488 29452 27494 29504
rect 1104 29402 30820 29424
rect 1104 29350 10880 29402
rect 10932 29350 10944 29402
rect 10996 29350 11008 29402
rect 11060 29350 11072 29402
rect 11124 29350 11136 29402
rect 11188 29350 20811 29402
rect 20863 29350 20875 29402
rect 20927 29350 20939 29402
rect 20991 29350 21003 29402
rect 21055 29350 21067 29402
rect 21119 29350 30820 29402
rect 1104 29328 30820 29350
rect 9766 29248 9772 29300
rect 9824 29288 9830 29300
rect 10321 29291 10379 29297
rect 10321 29288 10333 29291
rect 9824 29260 10333 29288
rect 9824 29248 9830 29260
rect 10321 29257 10333 29260
rect 10367 29257 10379 29291
rect 10321 29251 10379 29257
rect 11238 29248 11244 29300
rect 11296 29288 11302 29300
rect 12250 29288 12256 29300
rect 11296 29260 12256 29288
rect 11296 29248 11302 29260
rect 12250 29248 12256 29260
rect 12308 29248 12314 29300
rect 12713 29291 12771 29297
rect 12713 29257 12725 29291
rect 12759 29288 12771 29291
rect 13170 29288 13176 29300
rect 12759 29260 13176 29288
rect 12759 29257 12771 29260
rect 12713 29251 12771 29257
rect 13170 29248 13176 29260
rect 13228 29248 13234 29300
rect 16114 29288 16120 29300
rect 16075 29260 16120 29288
rect 16114 29248 16120 29260
rect 16172 29248 16178 29300
rect 16758 29248 16764 29300
rect 16816 29288 16822 29300
rect 16899 29291 16957 29297
rect 16899 29288 16911 29291
rect 16816 29260 16911 29288
rect 16816 29248 16822 29260
rect 16899 29257 16911 29260
rect 16945 29257 16957 29291
rect 16899 29251 16957 29257
rect 18969 29291 19027 29297
rect 18969 29257 18981 29291
rect 19015 29257 19027 29291
rect 20254 29288 20260 29300
rect 20215 29260 20260 29288
rect 18969 29251 19027 29257
rect 7834 29220 7840 29232
rect 7668 29192 7840 29220
rect 1397 29155 1455 29161
rect 1397 29121 1409 29155
rect 1443 29152 1455 29155
rect 2314 29152 2320 29164
rect 1443 29124 2320 29152
rect 1443 29121 1455 29124
rect 1397 29115 1455 29121
rect 2314 29112 2320 29124
rect 2372 29112 2378 29164
rect 7668 29161 7696 29192
rect 7834 29180 7840 29192
rect 7892 29220 7898 29232
rect 10134 29220 10140 29232
rect 7892 29192 10140 29220
rect 7892 29180 7898 29192
rect 10134 29180 10140 29192
rect 10192 29180 10198 29232
rect 12434 29180 12440 29232
rect 12492 29220 12498 29232
rect 14001 29223 14059 29229
rect 14001 29220 14013 29223
rect 12492 29192 14013 29220
rect 12492 29180 12498 29192
rect 14001 29189 14013 29192
rect 14047 29189 14059 29223
rect 14182 29220 14188 29232
rect 14143 29192 14188 29220
rect 14001 29183 14059 29189
rect 14182 29180 14188 29192
rect 14240 29180 14246 29232
rect 15197 29223 15255 29229
rect 15197 29189 15209 29223
rect 15243 29220 15255 29223
rect 18230 29220 18236 29232
rect 15243 29192 18236 29220
rect 15243 29189 15255 29192
rect 15197 29183 15255 29189
rect 18230 29180 18236 29192
rect 18288 29180 18294 29232
rect 18984 29220 19012 29251
rect 20254 29248 20260 29260
rect 20312 29248 20318 29300
rect 25498 29288 25504 29300
rect 25459 29260 25504 29288
rect 25498 29248 25504 29260
rect 25556 29248 25562 29300
rect 26145 29291 26203 29297
rect 26145 29257 26157 29291
rect 26191 29257 26203 29291
rect 27154 29288 27160 29300
rect 27115 29260 27160 29288
rect 26145 29251 26203 29257
rect 18984 29192 22048 29220
rect 7653 29155 7711 29161
rect 7653 29121 7665 29155
rect 7699 29121 7711 29155
rect 7653 29115 7711 29121
rect 8386 29112 8392 29164
rect 8444 29152 8450 29164
rect 8553 29155 8611 29161
rect 8553 29152 8565 29155
rect 8444 29124 8565 29152
rect 8444 29112 8450 29124
rect 8553 29121 8565 29124
rect 8599 29121 8611 29155
rect 8553 29115 8611 29121
rect 9674 29112 9680 29164
rect 9732 29152 9738 29164
rect 10262 29155 10320 29161
rect 10262 29152 10274 29155
rect 9732 29124 10274 29152
rect 9732 29112 9738 29124
rect 10262 29121 10274 29124
rect 10308 29121 10320 29155
rect 10686 29152 10692 29164
rect 10647 29124 10692 29152
rect 10262 29115 10320 29121
rect 10686 29112 10692 29124
rect 10744 29112 10750 29164
rect 10778 29112 10784 29164
rect 10836 29152 10842 29164
rect 11514 29152 11520 29164
rect 10836 29124 10881 29152
rect 11475 29124 11520 29152
rect 10836 29112 10842 29124
rect 11514 29112 11520 29124
rect 11572 29112 11578 29164
rect 11682 29155 11740 29161
rect 11682 29152 11694 29155
rect 11624 29124 11694 29152
rect 8294 29084 8300 29096
rect 8255 29056 8300 29084
rect 8294 29044 8300 29056
rect 8352 29044 8358 29096
rect 9306 29044 9312 29096
rect 9364 29084 9370 29096
rect 11146 29084 11152 29096
rect 9364 29056 11152 29084
rect 9364 29044 9370 29056
rect 11146 29044 11152 29056
rect 11204 29044 11210 29096
rect 11330 29044 11336 29096
rect 11388 29084 11394 29096
rect 11624 29084 11652 29124
rect 11682 29121 11694 29124
rect 11728 29121 11740 29155
rect 11682 29115 11740 29121
rect 11790 29112 11796 29164
rect 11848 29152 11854 29164
rect 12066 29152 12072 29164
rect 11848 29124 11893 29152
rect 12027 29124 12072 29152
rect 11848 29112 11854 29124
rect 12066 29112 12072 29124
rect 12124 29112 12130 29164
rect 12618 29112 12624 29164
rect 12676 29152 12682 29164
rect 13081 29155 13139 29161
rect 13081 29152 13093 29155
rect 12676 29124 13093 29152
rect 12676 29112 12682 29124
rect 13081 29121 13093 29124
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 14829 29155 14887 29161
rect 14829 29121 14841 29155
rect 14875 29121 14887 29155
rect 14829 29115 14887 29121
rect 11882 29084 11888 29096
rect 11388 29056 11652 29084
rect 11843 29056 11888 29084
rect 11388 29044 11394 29056
rect 11882 29044 11888 29056
rect 11940 29044 11946 29096
rect 13173 29087 13231 29093
rect 13173 29053 13185 29087
rect 13219 29084 13231 29087
rect 13262 29084 13268 29096
rect 13219 29056 13268 29084
rect 13219 29053 13231 29056
rect 13173 29047 13231 29053
rect 13262 29044 13268 29056
rect 13320 29044 13326 29096
rect 13357 29087 13415 29093
rect 13357 29053 13369 29087
rect 13403 29084 13415 29087
rect 13630 29084 13636 29096
rect 13403 29056 13636 29084
rect 13403 29053 13415 29056
rect 13357 29047 13415 29053
rect 13630 29044 13636 29056
rect 13688 29044 13694 29096
rect 1578 29016 1584 29028
rect 1539 28988 1584 29016
rect 1578 28976 1584 28988
rect 1636 28976 1642 29028
rect 9858 28976 9864 29028
rect 9916 29016 9922 29028
rect 10137 29019 10195 29025
rect 10137 29016 10149 29019
rect 9916 28988 10149 29016
rect 9916 28976 9922 28988
rect 10137 28985 10149 28988
rect 10183 28985 10195 29019
rect 10137 28979 10195 28985
rect 11790 28976 11796 29028
rect 11848 29016 11854 29028
rect 11974 29016 11980 29028
rect 11848 28988 11980 29016
rect 11848 28976 11854 28988
rect 11974 28976 11980 28988
rect 12032 28976 12038 29028
rect 12253 29019 12311 29025
rect 12253 28985 12265 29019
rect 12299 29016 12311 29019
rect 12802 29016 12808 29028
rect 12299 28988 12808 29016
rect 12299 28985 12311 28988
rect 12253 28979 12311 28985
rect 12802 28976 12808 28988
rect 12860 28976 12866 29028
rect 14844 29016 14872 29115
rect 14918 29112 14924 29164
rect 14976 29152 14982 29164
rect 15013 29155 15071 29161
rect 15013 29152 15025 29155
rect 14976 29124 15025 29152
rect 14976 29112 14982 29124
rect 15013 29121 15025 29124
rect 15059 29121 15071 29155
rect 15013 29115 15071 29121
rect 15470 29112 15476 29164
rect 15528 29152 15534 29164
rect 15657 29155 15715 29161
rect 15657 29152 15669 29155
rect 15528 29124 15669 29152
rect 15528 29112 15534 29124
rect 15657 29121 15669 29124
rect 15703 29121 15715 29155
rect 15657 29115 15715 29121
rect 16850 29112 16856 29164
rect 16908 29152 16914 29164
rect 17218 29152 17224 29164
rect 16908 29124 17224 29152
rect 16908 29112 16914 29124
rect 17218 29112 17224 29124
rect 17276 29112 17282 29164
rect 18046 29112 18052 29164
rect 18104 29152 18110 29164
rect 18141 29155 18199 29161
rect 18141 29152 18153 29155
rect 18104 29124 18153 29152
rect 18104 29112 18110 29124
rect 18141 29121 18153 29124
rect 18187 29121 18199 29155
rect 18141 29115 18199 29121
rect 18325 29155 18383 29161
rect 18325 29121 18337 29155
rect 18371 29121 18383 29155
rect 18325 29115 18383 29121
rect 18785 29155 18843 29161
rect 18785 29121 18797 29155
rect 18831 29121 18843 29155
rect 19426 29152 19432 29164
rect 19387 29124 19432 29152
rect 18785 29115 18843 29121
rect 16669 29087 16727 29093
rect 16669 29053 16681 29087
rect 16715 29084 16727 29087
rect 16758 29084 16764 29096
rect 16715 29056 16764 29084
rect 16715 29053 16727 29056
rect 16669 29047 16727 29053
rect 16758 29044 16764 29056
rect 16816 29044 16822 29096
rect 18340 29084 18368 29115
rect 18064 29056 18368 29084
rect 18800 29084 18828 29115
rect 19426 29112 19432 29124
rect 19484 29112 19490 29164
rect 20070 29152 20076 29164
rect 20031 29124 20076 29152
rect 20070 29112 20076 29124
rect 20128 29112 20134 29164
rect 20809 29155 20867 29161
rect 20809 29121 20821 29155
rect 20855 29152 20867 29155
rect 21174 29152 21180 29164
rect 20855 29124 21180 29152
rect 20855 29121 20867 29124
rect 20809 29115 20867 29121
rect 21174 29112 21180 29124
rect 21232 29112 21238 29164
rect 22020 29161 22048 29192
rect 23658 29180 23664 29232
rect 23716 29220 23722 29232
rect 24486 29220 24492 29232
rect 23716 29192 24492 29220
rect 23716 29180 23722 29192
rect 24486 29180 24492 29192
rect 24544 29220 24550 29232
rect 24544 29192 26004 29220
rect 24544 29180 24550 29192
rect 22005 29155 22063 29161
rect 22005 29121 22017 29155
rect 22051 29121 22063 29155
rect 22005 29115 22063 29121
rect 22094 29112 22100 29164
rect 22152 29152 22158 29164
rect 22261 29155 22319 29161
rect 22261 29152 22273 29155
rect 22152 29124 22273 29152
rect 22152 29112 22158 29124
rect 22261 29121 22273 29124
rect 22307 29121 22319 29155
rect 23845 29155 23903 29161
rect 23845 29152 23857 29155
rect 22261 29115 22319 29121
rect 23400 29124 23857 29152
rect 18800 29056 19656 29084
rect 14844 28988 15424 29016
rect 15396 28960 15424 28988
rect 16482 28976 16488 29028
rect 16540 29016 16546 29028
rect 18064 29016 18092 29056
rect 16540 28988 18092 29016
rect 18141 29019 18199 29025
rect 16540 28976 16546 28988
rect 18141 28985 18153 29019
rect 18187 29016 18199 29019
rect 19150 29016 19156 29028
rect 18187 28988 19156 29016
rect 18187 28985 18199 28988
rect 18141 28979 18199 28985
rect 19150 28976 19156 28988
rect 19208 28976 19214 29028
rect 19628 29025 19656 29056
rect 23400 29028 23428 29124
rect 23845 29121 23857 29124
rect 23891 29121 23903 29155
rect 23845 29115 23903 29121
rect 24210 29112 24216 29164
rect 24268 29152 24274 29164
rect 24670 29152 24676 29164
rect 24268 29124 24676 29152
rect 24268 29112 24274 29124
rect 24670 29112 24676 29124
rect 24728 29152 24734 29164
rect 25976 29161 26004 29192
rect 24765 29155 24823 29161
rect 24765 29152 24777 29155
rect 24728 29124 24777 29152
rect 24728 29112 24734 29124
rect 24765 29121 24777 29124
rect 24811 29121 24823 29155
rect 24765 29115 24823 29121
rect 24949 29155 25007 29161
rect 24949 29121 24961 29155
rect 24995 29152 25007 29155
rect 25317 29155 25375 29161
rect 24995 29124 25268 29152
rect 24995 29121 25007 29124
rect 24949 29115 25007 29121
rect 24854 29044 24860 29096
rect 24912 29084 24918 29096
rect 25041 29087 25099 29093
rect 25041 29084 25053 29087
rect 24912 29056 25053 29084
rect 24912 29044 24918 29056
rect 25041 29053 25053 29056
rect 25087 29053 25099 29087
rect 25041 29047 25099 29053
rect 25133 29087 25191 29093
rect 25133 29053 25145 29087
rect 25179 29053 25191 29087
rect 25133 29047 25191 29053
rect 19613 29019 19671 29025
rect 19613 28985 19625 29019
rect 19659 28985 19671 29019
rect 19613 28979 19671 28985
rect 20993 29019 21051 29025
rect 20993 28985 21005 29019
rect 21039 29016 21051 29019
rect 21174 29016 21180 29028
rect 21039 28988 21180 29016
rect 21039 28985 21051 28988
rect 20993 28979 21051 28985
rect 21174 28976 21180 28988
rect 21232 28976 21238 29028
rect 23382 29016 23388 29028
rect 23343 28988 23388 29016
rect 23382 28976 23388 28988
rect 23440 28976 23446 29028
rect 24305 29019 24363 29025
rect 23768 28988 24072 29016
rect 7837 28951 7895 28957
rect 7837 28917 7849 28951
rect 7883 28948 7895 28951
rect 7926 28948 7932 28960
rect 7883 28920 7932 28948
rect 7883 28917 7895 28920
rect 7837 28911 7895 28917
rect 7926 28908 7932 28920
rect 7984 28908 7990 28960
rect 9677 28951 9735 28957
rect 9677 28917 9689 28951
rect 9723 28948 9735 28951
rect 10594 28948 10600 28960
rect 9723 28920 10600 28948
rect 9723 28917 9735 28920
rect 9677 28911 9735 28917
rect 10594 28908 10600 28920
rect 10652 28908 10658 28960
rect 15378 28908 15384 28960
rect 15436 28948 15442 28960
rect 15749 28951 15807 28957
rect 15749 28948 15761 28951
rect 15436 28920 15761 28948
rect 15436 28908 15442 28920
rect 15749 28917 15761 28920
rect 15795 28917 15807 28951
rect 15749 28911 15807 28917
rect 16666 28908 16672 28960
rect 16724 28948 16730 28960
rect 19978 28948 19984 28960
rect 16724 28920 19984 28948
rect 16724 28908 16730 28920
rect 19978 28908 19984 28920
rect 20036 28908 20042 28960
rect 22278 28908 22284 28960
rect 22336 28948 22342 28960
rect 23768 28948 23796 28988
rect 22336 28920 23796 28948
rect 22336 28908 22342 28920
rect 23842 28908 23848 28960
rect 23900 28948 23906 28960
rect 23937 28951 23995 28957
rect 23937 28948 23949 28951
rect 23900 28920 23949 28948
rect 23900 28908 23906 28920
rect 23937 28917 23949 28920
rect 23983 28917 23995 28951
rect 24044 28948 24072 28988
rect 24305 28985 24317 29019
rect 24351 29016 24363 29019
rect 24578 29016 24584 29028
rect 24351 28988 24584 29016
rect 24351 28985 24363 28988
rect 24305 28979 24363 28985
rect 24578 28976 24584 28988
rect 24636 28976 24642 29028
rect 24762 28976 24768 29028
rect 24820 29016 24826 29028
rect 25148 29016 25176 29047
rect 24820 28988 25176 29016
rect 24820 28976 24826 28988
rect 25240 28948 25268 29124
rect 25317 29121 25329 29155
rect 25363 29121 25375 29155
rect 25317 29115 25375 29121
rect 25961 29155 26019 29161
rect 25961 29121 25973 29155
rect 26007 29121 26019 29155
rect 26160 29152 26188 29251
rect 27154 29248 27160 29260
rect 27212 29248 27218 29300
rect 27430 29248 27436 29300
rect 27488 29288 27494 29300
rect 28997 29291 29055 29297
rect 28997 29288 29009 29291
rect 27488 29260 29009 29288
rect 27488 29248 27494 29260
rect 28997 29257 29009 29260
rect 29043 29257 29055 29291
rect 29178 29288 29184 29300
rect 29139 29260 29184 29288
rect 28997 29251 29055 29257
rect 29178 29248 29184 29260
rect 29236 29248 29242 29300
rect 26973 29155 27031 29161
rect 26973 29152 26985 29155
rect 26160 29124 26985 29152
rect 25961 29115 26019 29121
rect 26973 29121 26985 29124
rect 27019 29121 27031 29155
rect 26973 29115 27031 29121
rect 25332 29084 25360 29115
rect 27062 29112 27068 29164
rect 27120 29152 27126 29164
rect 27617 29155 27675 29161
rect 27617 29152 27629 29155
rect 27120 29124 27629 29152
rect 27120 29112 27126 29124
rect 27617 29121 27629 29124
rect 27663 29121 27675 29155
rect 28626 29152 28632 29164
rect 28587 29124 28632 29152
rect 27617 29115 27675 29121
rect 28626 29112 28632 29124
rect 28684 29112 28690 29164
rect 29825 29155 29883 29161
rect 29825 29121 29837 29155
rect 29871 29121 29883 29155
rect 29825 29115 29883 29121
rect 27430 29084 27436 29096
rect 25332 29056 27436 29084
rect 27430 29044 27436 29056
rect 27488 29044 27494 29096
rect 27522 29044 27528 29096
rect 27580 29084 27586 29096
rect 29840 29084 29868 29115
rect 27580 29056 29868 29084
rect 27580 29044 27586 29056
rect 26510 28976 26516 29028
rect 26568 29016 26574 29028
rect 27801 29019 27859 29025
rect 27801 29016 27813 29019
rect 26568 28988 27813 29016
rect 26568 28976 26574 28988
rect 27801 28985 27813 28988
rect 27847 28985 27859 29019
rect 30006 29016 30012 29028
rect 29967 28988 30012 29016
rect 27801 28979 27859 28985
rect 30006 28976 30012 28988
rect 30064 28976 30070 29028
rect 24044 28920 25268 28948
rect 28997 28951 29055 28957
rect 23937 28911 23995 28917
rect 28997 28917 29009 28951
rect 29043 28948 29055 28951
rect 29086 28948 29092 28960
rect 29043 28920 29092 28948
rect 29043 28917 29055 28920
rect 28997 28911 29055 28917
rect 29086 28908 29092 28920
rect 29144 28908 29150 28960
rect 1104 28858 30820 28880
rect 1104 28806 5915 28858
rect 5967 28806 5979 28858
rect 6031 28806 6043 28858
rect 6095 28806 6107 28858
rect 6159 28806 6171 28858
rect 6223 28806 15846 28858
rect 15898 28806 15910 28858
rect 15962 28806 15974 28858
rect 16026 28806 16038 28858
rect 16090 28806 16102 28858
rect 16154 28806 25776 28858
rect 25828 28806 25840 28858
rect 25892 28806 25904 28858
rect 25956 28806 25968 28858
rect 26020 28806 26032 28858
rect 26084 28806 30820 28858
rect 1104 28784 30820 28806
rect 8113 28747 8171 28753
rect 8113 28713 8125 28747
rect 8159 28744 8171 28747
rect 8294 28744 8300 28756
rect 8159 28716 8300 28744
rect 8159 28713 8171 28716
rect 8113 28707 8171 28713
rect 8294 28704 8300 28716
rect 8352 28704 8358 28756
rect 10318 28704 10324 28756
rect 10376 28744 10382 28756
rect 10689 28747 10747 28753
rect 10689 28744 10701 28747
rect 10376 28716 10701 28744
rect 10376 28704 10382 28716
rect 10689 28713 10701 28716
rect 10735 28713 10747 28747
rect 10689 28707 10747 28713
rect 10873 28747 10931 28753
rect 10873 28713 10885 28747
rect 10919 28744 10931 28747
rect 11422 28744 11428 28756
rect 10919 28716 11428 28744
rect 10919 28713 10931 28716
rect 10873 28707 10931 28713
rect 11422 28704 11428 28716
rect 11480 28704 11486 28756
rect 12250 28704 12256 28756
rect 12308 28744 12314 28756
rect 12897 28747 12955 28753
rect 12897 28744 12909 28747
rect 12308 28716 12909 28744
rect 12308 28704 12314 28716
rect 12897 28713 12909 28716
rect 12943 28713 12955 28747
rect 22922 28744 22928 28756
rect 12897 28707 12955 28713
rect 16868 28716 20208 28744
rect 22883 28716 22928 28744
rect 9953 28679 10011 28685
rect 9953 28645 9965 28679
rect 9999 28676 10011 28679
rect 11514 28676 11520 28688
rect 9999 28648 11520 28676
rect 9999 28645 10011 28648
rect 9953 28639 10011 28645
rect 11514 28636 11520 28648
rect 11572 28636 11578 28688
rect 14090 28636 14096 28688
rect 14148 28676 14154 28688
rect 15013 28679 15071 28685
rect 15013 28676 15025 28679
rect 14148 28648 15025 28676
rect 14148 28636 14154 28648
rect 15013 28645 15025 28648
rect 15059 28645 15071 28679
rect 15013 28639 15071 28645
rect 8202 28568 8208 28620
rect 8260 28608 8266 28620
rect 16868 28608 16896 28716
rect 18233 28679 18291 28685
rect 18233 28645 18245 28679
rect 18279 28676 18291 28679
rect 18414 28676 18420 28688
rect 18279 28648 18420 28676
rect 18279 28645 18291 28648
rect 18233 28639 18291 28645
rect 18414 28636 18420 28648
rect 18472 28636 18478 28688
rect 20180 28676 20208 28716
rect 22922 28704 22928 28716
rect 22980 28704 22986 28756
rect 24854 28744 24860 28756
rect 24815 28716 24860 28744
rect 24854 28704 24860 28716
rect 24912 28704 24918 28756
rect 27338 28744 27344 28756
rect 27299 28716 27344 28744
rect 27338 28704 27344 28716
rect 27396 28704 27402 28756
rect 23845 28679 23903 28685
rect 23845 28676 23857 28679
rect 20180 28648 23857 28676
rect 23845 28645 23857 28648
rect 23891 28645 23903 28679
rect 23845 28639 23903 28645
rect 8260 28580 16896 28608
rect 8260 28568 8266 28580
rect 18874 28568 18880 28620
rect 18932 28608 18938 28620
rect 18932 28580 19196 28608
rect 18932 28568 18938 28580
rect 19168 28552 19196 28580
rect 21266 28568 21272 28620
rect 21324 28608 21330 28620
rect 21726 28608 21732 28620
rect 21324 28580 21588 28608
rect 21687 28580 21732 28608
rect 21324 28568 21330 28580
rect 7926 28540 7932 28552
rect 7887 28512 7932 28540
rect 7926 28500 7932 28512
rect 7984 28500 7990 28552
rect 9858 28540 9864 28552
rect 9819 28512 9864 28540
rect 9858 28500 9864 28512
rect 9916 28500 9922 28552
rect 11790 28500 11796 28552
rect 11848 28540 11854 28552
rect 12069 28543 12127 28549
rect 12069 28540 12081 28543
rect 11848 28512 12081 28540
rect 11848 28500 11854 28512
rect 12069 28509 12081 28512
rect 12115 28509 12127 28543
rect 12069 28503 12127 28509
rect 12158 28500 12164 28552
rect 12216 28540 12222 28552
rect 12805 28543 12863 28549
rect 12805 28540 12817 28543
rect 12216 28512 12817 28540
rect 12216 28500 12222 28512
rect 12805 28509 12817 28512
rect 12851 28509 12863 28543
rect 12805 28503 12863 28509
rect 13906 28500 13912 28552
rect 13964 28540 13970 28552
rect 14185 28543 14243 28549
rect 14185 28540 14197 28543
rect 13964 28512 14197 28540
rect 13964 28500 13970 28512
rect 14185 28509 14197 28512
rect 14231 28509 14243 28543
rect 14185 28503 14243 28509
rect 10505 28475 10563 28481
rect 10505 28441 10517 28475
rect 10551 28472 10563 28475
rect 10594 28472 10600 28484
rect 10551 28444 10600 28472
rect 10551 28441 10563 28444
rect 10505 28435 10563 28441
rect 10594 28432 10600 28444
rect 10652 28432 10658 28484
rect 11425 28475 11483 28481
rect 11425 28441 11437 28475
rect 11471 28472 11483 28475
rect 12434 28472 12440 28484
rect 11471 28444 12440 28472
rect 11471 28441 11483 28444
rect 11425 28435 11483 28441
rect 12434 28432 12440 28444
rect 12492 28432 12498 28484
rect 14200 28472 14228 28503
rect 14734 28500 14740 28552
rect 14792 28540 14798 28552
rect 14829 28543 14887 28549
rect 14829 28540 14841 28543
rect 14792 28512 14841 28540
rect 14792 28500 14798 28512
rect 14829 28509 14841 28512
rect 14875 28540 14887 28543
rect 15562 28540 15568 28552
rect 14875 28512 15424 28540
rect 15523 28512 15568 28540
rect 14875 28509 14887 28512
rect 14829 28503 14887 28509
rect 15102 28472 15108 28484
rect 14200 28444 15108 28472
rect 15102 28432 15108 28444
rect 15160 28432 15166 28484
rect 15396 28472 15424 28512
rect 15562 28500 15568 28512
rect 15620 28500 15626 28552
rect 15841 28543 15899 28549
rect 15841 28509 15853 28543
rect 15887 28540 15899 28543
rect 16666 28540 16672 28552
rect 15887 28512 16672 28540
rect 15887 28509 15899 28512
rect 15841 28503 15899 28509
rect 16666 28500 16672 28512
rect 16724 28500 16730 28552
rect 16850 28540 16856 28552
rect 16811 28512 16856 28540
rect 16850 28500 16856 28512
rect 16908 28500 16914 28552
rect 17052 28512 18192 28540
rect 17052 28472 17080 28512
rect 15396 28444 17080 28472
rect 17120 28475 17178 28481
rect 17120 28441 17132 28475
rect 17166 28472 17178 28475
rect 17862 28472 17868 28484
rect 17166 28444 17868 28472
rect 17166 28441 17178 28444
rect 17120 28435 17178 28441
rect 17862 28432 17868 28444
rect 17920 28432 17926 28484
rect 18164 28472 18192 28512
rect 18230 28500 18236 28552
rect 18288 28540 18294 28552
rect 19058 28540 19064 28552
rect 18288 28512 19064 28540
rect 18288 28500 18294 28512
rect 19058 28500 19064 28512
rect 19116 28500 19122 28552
rect 19150 28500 19156 28552
rect 19208 28500 19214 28552
rect 19245 28543 19303 28549
rect 19245 28509 19257 28543
rect 19291 28540 19303 28543
rect 19334 28540 19340 28552
rect 19291 28512 19340 28540
rect 19291 28509 19303 28512
rect 19245 28503 19303 28509
rect 19334 28500 19340 28512
rect 19392 28500 19398 28552
rect 21361 28543 21419 28549
rect 21361 28509 21373 28543
rect 21407 28540 21419 28543
rect 21450 28540 21456 28552
rect 21407 28512 21456 28540
rect 21407 28509 21419 28512
rect 21361 28503 21419 28509
rect 21450 28500 21456 28512
rect 21508 28500 21514 28552
rect 21560 28549 21588 28580
rect 21726 28568 21732 28580
rect 21784 28568 21790 28620
rect 23382 28608 23388 28620
rect 22066 28580 23388 28608
rect 21545 28543 21603 28549
rect 21545 28509 21557 28543
rect 21591 28509 21603 28543
rect 21545 28503 21603 28509
rect 21634 28500 21640 28552
rect 21692 28540 21698 28552
rect 21913 28543 21971 28549
rect 21692 28512 21737 28540
rect 21692 28500 21698 28512
rect 21913 28509 21925 28543
rect 21959 28540 21971 28543
rect 22066 28540 22094 28580
rect 23382 28568 23388 28580
rect 23440 28568 23446 28620
rect 21959 28512 22094 28540
rect 21959 28509 21971 28512
rect 21913 28503 21971 28509
rect 22186 28500 22192 28552
rect 22244 28540 22250 28552
rect 22741 28543 22799 28549
rect 22741 28540 22753 28543
rect 22244 28512 22753 28540
rect 22244 28500 22250 28512
rect 22741 28509 22753 28512
rect 22787 28509 22799 28543
rect 23658 28540 23664 28552
rect 23619 28512 23664 28540
rect 22741 28503 22799 28509
rect 23658 28500 23664 28512
rect 23716 28500 23722 28552
rect 24762 28540 24768 28552
rect 24723 28512 24768 28540
rect 24762 28500 24768 28512
rect 24820 28500 24826 28552
rect 25961 28543 26019 28549
rect 25961 28509 25973 28543
rect 26007 28540 26019 28543
rect 26510 28540 26516 28552
rect 26007 28512 26516 28540
rect 26007 28509 26019 28512
rect 25961 28503 26019 28509
rect 26510 28500 26516 28512
rect 26568 28500 26574 28552
rect 29822 28540 29828 28552
rect 29783 28512 29828 28540
rect 29822 28500 29828 28512
rect 29880 28500 29886 28552
rect 18164 28444 19196 28472
rect 10042 28364 10048 28416
rect 10100 28404 10106 28416
rect 10686 28404 10692 28416
rect 10744 28413 10750 28416
rect 10744 28407 10763 28413
rect 10100 28376 10692 28404
rect 10100 28364 10106 28376
rect 10686 28364 10692 28376
rect 10751 28373 10763 28407
rect 11514 28404 11520 28416
rect 11475 28376 11520 28404
rect 10744 28367 10763 28373
rect 10744 28364 10750 28367
rect 11514 28364 11520 28376
rect 11572 28364 11578 28416
rect 11698 28364 11704 28416
rect 11756 28404 11762 28416
rect 12250 28404 12256 28416
rect 11756 28376 12256 28404
rect 11756 28364 11762 28376
rect 12250 28364 12256 28376
rect 12308 28364 12314 28416
rect 14277 28407 14335 28413
rect 14277 28373 14289 28407
rect 14323 28404 14335 28407
rect 14826 28404 14832 28416
rect 14323 28376 14832 28404
rect 14323 28373 14335 28376
rect 14277 28367 14335 28373
rect 14826 28364 14832 28376
rect 14884 28364 14890 28416
rect 17310 28364 17316 28416
rect 17368 28404 17374 28416
rect 18782 28404 18788 28416
rect 17368 28376 18788 28404
rect 17368 28364 17374 28376
rect 18782 28364 18788 28376
rect 18840 28364 18846 28416
rect 19168 28404 19196 28444
rect 19509 28432 19515 28484
rect 19567 28472 19573 28484
rect 26228 28475 26286 28481
rect 19567 28444 19612 28472
rect 19567 28432 19573 28444
rect 26228 28441 26240 28475
rect 26274 28472 26286 28475
rect 26418 28472 26424 28484
rect 26274 28444 26424 28472
rect 26274 28441 26286 28444
rect 26228 28435 26286 28441
rect 26418 28432 26424 28444
rect 26476 28432 26482 28484
rect 19334 28404 19340 28416
rect 19168 28376 19340 28404
rect 19334 28364 19340 28376
rect 19392 28364 19398 28416
rect 19886 28364 19892 28416
rect 19944 28404 19950 28416
rect 20625 28407 20683 28413
rect 20625 28404 20637 28407
rect 19944 28376 20637 28404
rect 19944 28364 19950 28376
rect 20625 28373 20637 28376
rect 20671 28373 20683 28407
rect 20625 28367 20683 28373
rect 22094 28364 22100 28416
rect 22152 28404 22158 28416
rect 23201 28407 23259 28413
rect 22152 28376 22197 28404
rect 22152 28364 22158 28376
rect 23201 28373 23213 28407
rect 23247 28404 23259 28407
rect 23842 28404 23848 28416
rect 23247 28376 23848 28404
rect 23247 28373 23259 28376
rect 23201 28367 23259 28373
rect 23842 28364 23848 28376
rect 23900 28364 23906 28416
rect 24118 28364 24124 28416
rect 24176 28404 24182 28416
rect 25038 28404 25044 28416
rect 24176 28376 25044 28404
rect 24176 28364 24182 28376
rect 25038 28364 25044 28376
rect 25096 28364 25102 28416
rect 30006 28404 30012 28416
rect 29967 28376 30012 28404
rect 30006 28364 30012 28376
rect 30064 28364 30070 28416
rect 1104 28314 30820 28336
rect 1104 28262 10880 28314
rect 10932 28262 10944 28314
rect 10996 28262 11008 28314
rect 11060 28262 11072 28314
rect 11124 28262 11136 28314
rect 11188 28262 20811 28314
rect 20863 28262 20875 28314
rect 20927 28262 20939 28314
rect 20991 28262 21003 28314
rect 21055 28262 21067 28314
rect 21119 28262 30820 28314
rect 1104 28240 30820 28262
rect 9950 28160 9956 28212
rect 10008 28200 10014 28212
rect 16666 28200 16672 28212
rect 10008 28172 16672 28200
rect 10008 28160 10014 28172
rect 16666 28160 16672 28172
rect 16724 28160 16730 28212
rect 17310 28160 17316 28212
rect 17368 28200 17374 28212
rect 17862 28200 17868 28212
rect 17368 28172 17448 28200
rect 17823 28172 17868 28200
rect 17368 28160 17374 28172
rect 11793 28135 11851 28141
rect 11793 28101 11805 28135
rect 11839 28132 11851 28135
rect 11882 28132 11888 28144
rect 11839 28104 11888 28132
rect 11839 28101 11851 28104
rect 11793 28095 11851 28101
rect 11882 28092 11888 28104
rect 11940 28092 11946 28144
rect 14544 28135 14602 28141
rect 12452 28104 14228 28132
rect 7834 28024 7840 28076
rect 7892 28064 7898 28076
rect 7929 28067 7987 28073
rect 7929 28064 7941 28067
rect 7892 28036 7941 28064
rect 7892 28024 7898 28036
rect 7929 28033 7941 28036
rect 7975 28033 7987 28067
rect 7929 28027 7987 28033
rect 9493 28067 9551 28073
rect 9493 28033 9505 28067
rect 9539 28064 9551 28067
rect 10502 28064 10508 28076
rect 9539 28036 10508 28064
rect 9539 28033 9551 28036
rect 9493 28027 9551 28033
rect 10502 28024 10508 28036
rect 10560 28024 10566 28076
rect 12452 28073 12480 28104
rect 14200 28076 14228 28104
rect 14544 28101 14556 28135
rect 14590 28132 14602 28135
rect 15194 28132 15200 28144
rect 14590 28104 15200 28132
rect 14590 28101 14602 28104
rect 14544 28095 14602 28101
rect 15194 28092 15200 28104
rect 15252 28092 15258 28144
rect 15746 28092 15752 28144
rect 15804 28132 15810 28144
rect 17420 28132 17448 28172
rect 17862 28160 17868 28172
rect 17920 28160 17926 28212
rect 19242 28160 19248 28212
rect 19300 28200 19306 28212
rect 19429 28203 19487 28209
rect 19300 28172 19380 28200
rect 19300 28160 19306 28172
rect 15804 28104 17356 28132
rect 15804 28092 15810 28104
rect 12437 28067 12495 28073
rect 12437 28033 12449 28067
rect 12483 28033 12495 28067
rect 12437 28027 12495 28033
rect 12704 28067 12762 28073
rect 12704 28033 12716 28067
rect 12750 28064 12762 28067
rect 13262 28064 13268 28076
rect 12750 28036 13268 28064
rect 12750 28033 12762 28036
rect 12704 28027 12762 28033
rect 13262 28024 13268 28036
rect 13320 28024 13326 28076
rect 14182 28024 14188 28076
rect 14240 28064 14246 28076
rect 17328 28073 17356 28104
rect 17420 28104 18828 28132
rect 17420 28073 17448 28104
rect 14277 28067 14335 28073
rect 14277 28064 14289 28067
rect 14240 28036 14289 28064
rect 14240 28024 14246 28036
rect 14277 28033 14289 28036
rect 14323 28033 14335 28067
rect 14277 28027 14335 28033
rect 17129 28067 17187 28073
rect 17129 28033 17141 28067
rect 17175 28033 17187 28067
rect 17129 28027 17187 28033
rect 17313 28067 17371 28073
rect 17313 28033 17325 28067
rect 17359 28033 17371 28067
rect 17313 28027 17371 28033
rect 17405 28067 17463 28073
rect 17405 28033 17417 28067
rect 17451 28033 17463 28067
rect 17405 28027 17463 28033
rect 17497 28067 17555 28073
rect 17497 28033 17509 28067
rect 17543 28064 17555 28067
rect 17586 28064 17592 28076
rect 17543 28036 17592 28064
rect 17543 28033 17555 28036
rect 17497 28027 17555 28033
rect 9585 27999 9643 28005
rect 9585 27965 9597 27999
rect 9631 27996 9643 27999
rect 10134 27996 10140 28008
rect 9631 27968 10140 27996
rect 9631 27965 9643 27968
rect 9585 27959 9643 27965
rect 10134 27956 10140 27968
rect 10192 27956 10198 28008
rect 10413 27999 10471 28005
rect 10413 27965 10425 27999
rect 10459 27996 10471 27999
rect 10594 27996 10600 28008
rect 10459 27968 10600 27996
rect 10459 27965 10471 27968
rect 10413 27959 10471 27965
rect 10594 27956 10600 27968
rect 10652 27956 10658 28008
rect 17144 27996 17172 28027
rect 17586 28024 17592 28036
rect 17644 28024 17650 28076
rect 17681 28067 17739 28073
rect 17681 28033 17693 28067
rect 17727 28064 17739 28067
rect 18414 28064 18420 28076
rect 17727 28036 18420 28064
rect 17727 28033 17739 28036
rect 17681 28027 17739 28033
rect 18414 28024 18420 28036
rect 18472 28024 18478 28076
rect 18693 28067 18751 28073
rect 18693 28033 18705 28067
rect 18739 28033 18751 28067
rect 18693 28027 18751 28033
rect 17604 27996 17632 28024
rect 17862 27996 17868 28008
rect 17144 27968 17356 27996
rect 17604 27968 17868 27996
rect 17328 27940 17356 27968
rect 17862 27956 17868 27968
rect 17920 27956 17926 28008
rect 17310 27888 17316 27940
rect 17368 27928 17374 27940
rect 18708 27928 18736 28027
rect 18800 27996 18828 28104
rect 18966 28092 18972 28144
rect 19024 28092 19030 28144
rect 19352 28132 19380 28172
rect 19429 28169 19441 28203
rect 19475 28200 19487 28203
rect 19518 28200 19524 28212
rect 19475 28172 19524 28200
rect 19475 28169 19487 28172
rect 19429 28163 19487 28169
rect 19518 28160 19524 28172
rect 19576 28160 19582 28212
rect 21634 28160 21640 28212
rect 21692 28200 21698 28212
rect 24118 28200 24124 28212
rect 21692 28172 24124 28200
rect 21692 28160 21698 28172
rect 24118 28160 24124 28172
rect 24176 28160 24182 28212
rect 24946 28200 24952 28212
rect 24228 28172 24952 28200
rect 20257 28135 20315 28141
rect 19352 28104 20208 28132
rect 18865 28067 18923 28073
rect 18865 28033 18877 28067
rect 18911 28064 18923 28067
rect 18984 28064 19012 28092
rect 18911 28036 19012 28064
rect 18911 28033 18923 28036
rect 18865 28027 18923 28033
rect 19058 28024 19064 28076
rect 19116 28064 19122 28076
rect 19245 28068 19303 28073
rect 19245 28067 19472 28068
rect 19116 28036 19161 28064
rect 19116 28024 19122 28036
rect 19245 28033 19257 28067
rect 19291 28064 19472 28067
rect 19886 28064 19892 28076
rect 19291 28040 19892 28064
rect 19291 28033 19303 28040
rect 19444 28036 19892 28040
rect 19245 28027 19303 28033
rect 19886 28024 19892 28036
rect 19944 28024 19950 28076
rect 20180 28064 20208 28104
rect 20257 28101 20269 28135
rect 20303 28132 20315 28135
rect 20806 28132 20812 28144
rect 20303 28104 20812 28132
rect 20303 28101 20315 28104
rect 20257 28095 20315 28101
rect 20806 28092 20812 28104
rect 20864 28092 20870 28144
rect 21266 28092 21272 28144
rect 21324 28132 21330 28144
rect 21324 28104 22048 28132
rect 21324 28092 21330 28104
rect 20180 28036 20484 28064
rect 18969 27999 19027 28005
rect 18969 27996 18981 27999
rect 18800 27968 18981 27996
rect 18969 27965 18981 27968
rect 19015 27965 19027 27999
rect 20346 27996 20352 28008
rect 20307 27968 20352 27996
rect 18969 27959 19027 27965
rect 20346 27956 20352 27968
rect 20404 27956 20410 28008
rect 20456 28005 20484 28036
rect 20714 28024 20720 28076
rect 20772 28064 20778 28076
rect 21085 28067 21143 28073
rect 21085 28064 21097 28067
rect 20772 28036 21097 28064
rect 20772 28024 20778 28036
rect 21085 28033 21097 28036
rect 21131 28033 21143 28067
rect 21085 28027 21143 28033
rect 21450 28024 21456 28076
rect 21508 28064 21514 28076
rect 22020 28073 22048 28104
rect 21821 28067 21879 28073
rect 21821 28064 21833 28067
rect 21508 28036 21833 28064
rect 21508 28024 21514 28036
rect 21821 28033 21833 28036
rect 21867 28033 21879 28067
rect 21821 28027 21879 28033
rect 22005 28067 22063 28073
rect 22005 28033 22017 28067
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 22091 28067 22149 28073
rect 22091 28033 22103 28067
rect 22137 28064 22149 28067
rect 22278 28064 22284 28076
rect 22137 28036 22284 28064
rect 22137 28033 22149 28036
rect 22091 28027 22149 28033
rect 22278 28024 22284 28036
rect 22336 28024 22342 28076
rect 22373 28067 22431 28073
rect 22373 28033 22385 28067
rect 22419 28064 22431 28067
rect 22554 28064 22560 28076
rect 22419 28036 22560 28064
rect 22419 28033 22431 28036
rect 22373 28027 22431 28033
rect 22554 28024 22560 28036
rect 22612 28024 22618 28076
rect 23109 28067 23167 28073
rect 23109 28033 23121 28067
rect 23155 28064 23167 28067
rect 23474 28064 23480 28076
rect 23155 28036 23480 28064
rect 23155 28033 23167 28036
rect 23109 28027 23167 28033
rect 23474 28024 23480 28036
rect 23532 28024 23538 28076
rect 24228 28073 24256 28172
rect 24946 28160 24952 28172
rect 25004 28160 25010 28212
rect 25777 28203 25835 28209
rect 25777 28169 25789 28203
rect 25823 28200 25835 28203
rect 27062 28200 27068 28212
rect 25823 28172 27068 28200
rect 25823 28169 25835 28172
rect 25777 28163 25835 28169
rect 27062 28160 27068 28172
rect 27120 28160 27126 28212
rect 24486 28092 24492 28144
rect 24544 28132 24550 28144
rect 24544 28104 25636 28132
rect 24544 28092 24550 28104
rect 24213 28067 24271 28073
rect 24213 28033 24225 28067
rect 24259 28033 24271 28067
rect 24213 28027 24271 28033
rect 24673 28067 24731 28073
rect 24673 28033 24685 28067
rect 24719 28033 24731 28067
rect 24854 28064 24860 28076
rect 24815 28036 24860 28064
rect 24673 28027 24731 28033
rect 20441 27999 20499 28005
rect 20441 27965 20453 27999
rect 20487 27965 20499 27999
rect 20441 27959 20499 27965
rect 21726 27956 21732 28008
rect 21784 27996 21790 28008
rect 21910 27996 21916 28008
rect 21784 27968 21916 27996
rect 21784 27956 21790 27968
rect 21910 27956 21916 27968
rect 21968 27996 21974 28008
rect 22189 27999 22247 28005
rect 22189 27996 22201 27999
rect 21968 27968 22201 27996
rect 21968 27956 21974 27968
rect 22189 27965 22201 27968
rect 22235 27965 22247 27999
rect 22189 27959 22247 27965
rect 23566 27956 23572 28008
rect 23624 27996 23630 28008
rect 24688 27996 24716 28027
rect 24854 28024 24860 28036
rect 24912 28024 24918 28076
rect 25608 28073 25636 28104
rect 25593 28067 25651 28073
rect 25593 28033 25605 28067
rect 25639 28033 25651 28067
rect 25593 28027 25651 28033
rect 29825 28067 29883 28073
rect 29825 28033 29837 28067
rect 29871 28033 29883 28067
rect 29825 28027 29883 28033
rect 23624 27968 24716 27996
rect 24765 27999 24823 28005
rect 23624 27956 23630 27968
rect 24765 27965 24777 27999
rect 24811 27996 24823 27999
rect 29840 27996 29868 28027
rect 24811 27968 29868 27996
rect 24811 27965 24823 27968
rect 24765 27959 24823 27965
rect 17368 27900 18736 27928
rect 17368 27888 17374 27900
rect 19334 27888 19340 27940
rect 19392 27928 19398 27940
rect 19889 27931 19947 27937
rect 19889 27928 19901 27931
rect 19392 27900 19901 27928
rect 19392 27888 19398 27900
rect 19889 27897 19901 27900
rect 19935 27897 19947 27931
rect 19889 27891 19947 27897
rect 22278 27888 22284 27940
rect 22336 27928 22342 27940
rect 22557 27931 22615 27937
rect 22557 27928 22569 27931
rect 22336 27900 22569 27928
rect 22336 27888 22342 27900
rect 22557 27897 22569 27900
rect 22603 27897 22615 27931
rect 24029 27931 24087 27937
rect 24029 27928 24041 27931
rect 22557 27891 22615 27897
rect 23216 27900 24041 27928
rect 8018 27820 8024 27872
rect 8076 27860 8082 27872
rect 8113 27863 8171 27869
rect 8113 27860 8125 27863
rect 8076 27832 8125 27860
rect 8076 27820 8082 27832
rect 8113 27829 8125 27832
rect 8159 27829 8171 27863
rect 8113 27823 8171 27829
rect 9766 27820 9772 27872
rect 9824 27860 9830 27872
rect 11790 27860 11796 27872
rect 9824 27832 11796 27860
rect 9824 27820 9830 27832
rect 11790 27820 11796 27832
rect 11848 27860 11854 27872
rect 11885 27863 11943 27869
rect 11885 27860 11897 27863
rect 11848 27832 11897 27860
rect 11848 27820 11854 27832
rect 11885 27829 11897 27832
rect 11931 27829 11943 27863
rect 11885 27823 11943 27829
rect 13817 27863 13875 27869
rect 13817 27829 13829 27863
rect 13863 27860 13875 27863
rect 14274 27860 14280 27872
rect 13863 27832 14280 27860
rect 13863 27829 13875 27832
rect 13817 27823 13875 27829
rect 14274 27820 14280 27832
rect 14332 27820 14338 27872
rect 15286 27820 15292 27872
rect 15344 27860 15350 27872
rect 15657 27863 15715 27869
rect 15657 27860 15669 27863
rect 15344 27832 15669 27860
rect 15344 27820 15350 27832
rect 15657 27829 15669 27832
rect 15703 27829 15715 27863
rect 15657 27823 15715 27829
rect 19058 27820 19064 27872
rect 19116 27860 19122 27872
rect 19794 27860 19800 27872
rect 19116 27832 19800 27860
rect 19116 27820 19122 27832
rect 19794 27820 19800 27832
rect 19852 27820 19858 27872
rect 21269 27863 21327 27869
rect 21269 27829 21281 27863
rect 21315 27860 21327 27863
rect 22462 27860 22468 27872
rect 21315 27832 22468 27860
rect 21315 27829 21327 27832
rect 21269 27823 21327 27829
rect 22462 27820 22468 27832
rect 22520 27820 22526 27872
rect 22646 27820 22652 27872
rect 22704 27860 22710 27872
rect 22922 27860 22928 27872
rect 22704 27832 22928 27860
rect 22704 27820 22710 27832
rect 22922 27820 22928 27832
rect 22980 27860 22986 27872
rect 23216 27869 23244 27900
rect 24029 27897 24041 27900
rect 24075 27897 24087 27931
rect 24029 27891 24087 27897
rect 23201 27863 23259 27869
rect 23201 27860 23213 27863
rect 22980 27832 23213 27860
rect 22980 27820 22986 27832
rect 23201 27829 23213 27832
rect 23247 27829 23259 27863
rect 23201 27823 23259 27829
rect 23569 27863 23627 27869
rect 23569 27829 23581 27863
rect 23615 27860 23627 27863
rect 23934 27860 23940 27872
rect 23615 27832 23940 27860
rect 23615 27829 23627 27832
rect 23569 27823 23627 27829
rect 23934 27820 23940 27832
rect 23992 27820 23998 27872
rect 30006 27860 30012 27872
rect 29967 27832 30012 27860
rect 30006 27820 30012 27832
rect 30064 27820 30070 27872
rect 1104 27770 30820 27792
rect 1104 27718 5915 27770
rect 5967 27718 5979 27770
rect 6031 27718 6043 27770
rect 6095 27718 6107 27770
rect 6159 27718 6171 27770
rect 6223 27718 15846 27770
rect 15898 27718 15910 27770
rect 15962 27718 15974 27770
rect 16026 27718 16038 27770
rect 16090 27718 16102 27770
rect 16154 27718 25776 27770
rect 25828 27718 25840 27770
rect 25892 27718 25904 27770
rect 25956 27718 25968 27770
rect 26020 27718 26032 27770
rect 26084 27718 30820 27770
rect 1104 27696 30820 27718
rect 12066 27616 12072 27668
rect 12124 27656 12130 27668
rect 14734 27656 14740 27668
rect 12124 27628 14740 27656
rect 12124 27616 12130 27628
rect 14734 27616 14740 27628
rect 14792 27616 14798 27668
rect 15562 27616 15568 27668
rect 15620 27656 15626 27668
rect 16485 27659 16543 27665
rect 16485 27656 16497 27659
rect 15620 27628 16497 27656
rect 15620 27616 15626 27628
rect 16485 27625 16497 27628
rect 16531 27625 16543 27659
rect 16485 27619 16543 27625
rect 16666 27616 16672 27668
rect 16724 27656 16730 27668
rect 18414 27656 18420 27668
rect 16724 27628 18420 27656
rect 16724 27616 16730 27628
rect 18414 27616 18420 27628
rect 18472 27656 18478 27668
rect 20346 27656 20352 27668
rect 18472 27628 19196 27656
rect 18472 27616 18478 27628
rect 9950 27548 9956 27600
rect 10008 27588 10014 27600
rect 11422 27588 11428 27600
rect 10008 27560 11428 27588
rect 10008 27548 10014 27560
rect 11422 27548 11428 27560
rect 11480 27548 11486 27600
rect 11609 27591 11667 27597
rect 11609 27557 11621 27591
rect 11655 27588 11667 27591
rect 11882 27588 11888 27600
rect 11655 27560 11888 27588
rect 11655 27557 11667 27560
rect 11609 27551 11667 27557
rect 9769 27523 9827 27529
rect 9769 27489 9781 27523
rect 9815 27520 9827 27523
rect 10042 27520 10048 27532
rect 9815 27492 10048 27520
rect 9815 27489 9827 27492
rect 9769 27483 9827 27489
rect 10042 27480 10048 27492
rect 10100 27480 10106 27532
rect 10229 27523 10287 27529
rect 10229 27489 10241 27523
rect 10275 27520 10287 27523
rect 11238 27520 11244 27532
rect 10275 27492 11244 27520
rect 10275 27489 10287 27492
rect 10229 27483 10287 27489
rect 11238 27480 11244 27492
rect 11296 27480 11302 27532
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27412 1458 27464
rect 8018 27452 8024 27464
rect 7979 27424 8024 27452
rect 8018 27412 8024 27424
rect 8076 27412 8082 27464
rect 10134 27412 10140 27464
rect 10192 27452 10198 27464
rect 10413 27455 10471 27461
rect 10413 27452 10425 27455
rect 10192 27424 10425 27452
rect 10192 27412 10198 27424
rect 10413 27421 10425 27424
rect 10459 27421 10471 27455
rect 10413 27415 10471 27421
rect 10781 27455 10839 27461
rect 10781 27421 10793 27455
rect 10827 27452 10839 27455
rect 11624 27452 11652 27551
rect 11882 27548 11888 27560
rect 11940 27548 11946 27600
rect 14274 27548 14280 27600
rect 14332 27588 14338 27600
rect 15059 27591 15117 27597
rect 15059 27588 15071 27591
rect 14332 27560 15071 27588
rect 14332 27548 14338 27560
rect 15059 27557 15071 27560
rect 15105 27557 15117 27591
rect 15059 27551 15117 27557
rect 15194 27548 15200 27600
rect 15252 27588 15258 27600
rect 15654 27588 15660 27600
rect 15252 27560 15660 27588
rect 15252 27548 15258 27560
rect 15654 27548 15660 27560
rect 15712 27548 15718 27600
rect 17678 27548 17684 27600
rect 17736 27588 17742 27600
rect 19168 27588 19196 27628
rect 19306 27628 20352 27656
rect 19306 27588 19334 27628
rect 20346 27616 20352 27628
rect 20404 27616 20410 27668
rect 21450 27656 21456 27668
rect 21192 27628 21456 27656
rect 17736 27560 18368 27588
rect 19168 27560 19334 27588
rect 17736 27548 17742 27560
rect 12250 27480 12256 27532
rect 12308 27520 12314 27532
rect 14366 27520 14372 27532
rect 12308 27492 14372 27520
rect 12308 27480 12314 27492
rect 14366 27480 14372 27492
rect 14424 27480 14430 27532
rect 14461 27523 14519 27529
rect 14461 27489 14473 27523
rect 14507 27520 14519 27523
rect 15286 27520 15292 27532
rect 14507 27492 15148 27520
rect 15247 27492 15292 27520
rect 14507 27489 14519 27492
rect 14461 27483 14519 27489
rect 10827 27424 11652 27452
rect 12069 27455 12127 27461
rect 10827 27421 10839 27424
rect 10781 27415 10839 27421
rect 12069 27421 12081 27455
rect 12115 27452 12127 27455
rect 12437 27455 12495 27461
rect 12115 27424 12388 27452
rect 12115 27421 12127 27424
rect 12069 27415 12127 27421
rect 9582 27384 9588 27396
rect 9543 27356 9588 27384
rect 9582 27344 9588 27356
rect 9640 27344 9646 27396
rect 9858 27344 9864 27396
rect 9916 27384 9922 27396
rect 10226 27384 10232 27396
rect 9916 27356 10232 27384
rect 9916 27344 9922 27356
rect 10226 27344 10232 27356
rect 10284 27384 10290 27396
rect 11241 27387 11299 27393
rect 11241 27384 11253 27387
rect 10284 27356 11253 27384
rect 10284 27344 10290 27356
rect 11241 27353 11253 27356
rect 11287 27353 11299 27387
rect 11422 27384 11428 27396
rect 11383 27356 11428 27384
rect 11241 27347 11299 27353
rect 11422 27344 11428 27356
rect 11480 27344 11486 27396
rect 12253 27387 12311 27393
rect 12253 27384 12265 27387
rect 12084 27356 12265 27384
rect 12084 27328 12112 27356
rect 12253 27353 12265 27356
rect 12299 27353 12311 27387
rect 12360 27384 12388 27424
rect 12437 27421 12449 27455
rect 12483 27452 12495 27455
rect 12897 27455 12955 27461
rect 12897 27452 12909 27455
rect 12483 27424 12909 27452
rect 12483 27421 12495 27424
rect 12437 27415 12495 27421
rect 12897 27421 12909 27424
rect 12943 27421 12955 27455
rect 12897 27415 12955 27421
rect 12986 27412 12992 27464
rect 13044 27452 13050 27464
rect 14734 27452 14740 27464
rect 13044 27424 14740 27452
rect 13044 27412 13050 27424
rect 14734 27412 14740 27424
rect 14792 27412 14798 27464
rect 12618 27384 12624 27396
rect 12360 27356 12624 27384
rect 12253 27347 12311 27353
rect 12618 27344 12624 27356
rect 12676 27344 12682 27396
rect 14277 27387 14335 27393
rect 14277 27353 14289 27387
rect 14323 27353 14335 27387
rect 14277 27347 14335 27353
rect 1578 27316 1584 27328
rect 1539 27288 1584 27316
rect 1578 27276 1584 27288
rect 1636 27276 1642 27328
rect 7742 27276 7748 27328
rect 7800 27316 7806 27328
rect 8205 27319 8263 27325
rect 8205 27316 8217 27319
rect 7800 27288 8217 27316
rect 7800 27276 7806 27288
rect 8205 27285 8217 27288
rect 8251 27285 8263 27319
rect 10502 27316 10508 27328
rect 10463 27288 10508 27316
rect 8205 27279 8263 27285
rect 10502 27276 10508 27288
rect 10560 27276 10566 27328
rect 10597 27319 10655 27325
rect 10597 27285 10609 27319
rect 10643 27316 10655 27319
rect 10686 27316 10692 27328
rect 10643 27288 10692 27316
rect 10643 27285 10655 27288
rect 10597 27279 10655 27285
rect 10686 27276 10692 27288
rect 10744 27276 10750 27328
rect 12066 27276 12072 27328
rect 12124 27276 12130 27328
rect 13078 27316 13084 27328
rect 13039 27288 13084 27316
rect 13078 27276 13084 27288
rect 13136 27276 13142 27328
rect 14292 27316 14320 27347
rect 14458 27344 14464 27396
rect 14516 27384 14522 27396
rect 14921 27387 14979 27393
rect 14921 27384 14933 27387
rect 14516 27356 14933 27384
rect 14516 27344 14522 27356
rect 14921 27353 14933 27356
rect 14967 27353 14979 27387
rect 15120 27384 15148 27492
rect 15286 27480 15292 27492
rect 15344 27520 15350 27532
rect 17788 27529 17816 27560
rect 17773 27523 17831 27529
rect 15344 27492 16344 27520
rect 15344 27480 15350 27492
rect 16114 27452 16120 27464
rect 16075 27424 16120 27452
rect 16114 27412 16120 27424
rect 16172 27412 16178 27464
rect 16316 27461 16344 27492
rect 17773 27489 17785 27523
rect 17819 27489 17831 27523
rect 17773 27483 17831 27489
rect 17862 27480 17868 27532
rect 17920 27520 17926 27532
rect 18230 27520 18236 27532
rect 17920 27492 17965 27520
rect 18191 27492 18236 27520
rect 17920 27480 17926 27492
rect 18230 27480 18236 27492
rect 18288 27480 18294 27532
rect 18340 27520 18368 27560
rect 20070 27520 20076 27532
rect 18340 27492 20076 27520
rect 20070 27480 20076 27492
rect 20128 27480 20134 27532
rect 20165 27523 20223 27529
rect 20165 27489 20177 27523
rect 20211 27520 20223 27523
rect 20530 27520 20536 27532
rect 20211 27492 20536 27520
rect 20211 27489 20223 27492
rect 20165 27483 20223 27489
rect 20530 27480 20536 27492
rect 20588 27520 20594 27532
rect 21192 27520 21220 27628
rect 21450 27616 21456 27628
rect 21508 27616 21514 27668
rect 22554 27656 22560 27668
rect 22515 27628 22560 27656
rect 22554 27616 22560 27628
rect 22612 27616 22618 27668
rect 23201 27591 23259 27597
rect 23201 27557 23213 27591
rect 23247 27557 23259 27591
rect 23201 27551 23259 27557
rect 26329 27591 26387 27597
rect 26329 27557 26341 27591
rect 26375 27588 26387 27591
rect 27522 27588 27528 27600
rect 26375 27560 27528 27588
rect 26375 27557 26387 27560
rect 26329 27551 26387 27557
rect 23216 27520 23244 27551
rect 27522 27548 27528 27560
rect 27580 27548 27586 27600
rect 20588 27492 21220 27520
rect 22664 27492 23244 27520
rect 20588 27480 20594 27492
rect 16301 27455 16359 27461
rect 16301 27421 16313 27455
rect 16347 27421 16359 27455
rect 16301 27415 16359 27421
rect 17310 27412 17316 27464
rect 17368 27452 17374 27464
rect 17405 27455 17463 27461
rect 17405 27452 17417 27455
rect 17368 27424 17417 27452
rect 17368 27412 17374 27424
rect 17405 27421 17417 27424
rect 17451 27452 17463 27455
rect 17497 27455 17555 27461
rect 17497 27452 17509 27455
rect 17451 27424 17509 27452
rect 17451 27421 17463 27424
rect 17405 27415 17463 27421
rect 17497 27421 17509 27424
rect 17543 27421 17555 27455
rect 17678 27452 17684 27464
rect 17639 27424 17684 27452
rect 17497 27415 17555 27421
rect 17678 27412 17684 27424
rect 17736 27412 17742 27464
rect 18049 27455 18107 27461
rect 18049 27421 18061 27455
rect 18095 27452 18107 27455
rect 18322 27452 18328 27464
rect 18095 27424 18328 27452
rect 18095 27421 18107 27424
rect 18049 27415 18107 27421
rect 18322 27412 18328 27424
rect 18380 27412 18386 27464
rect 19245 27455 19303 27461
rect 19245 27421 19257 27455
rect 19291 27452 19303 27455
rect 19426 27452 19432 27464
rect 19291 27424 19432 27452
rect 19291 27421 19303 27424
rect 19245 27415 19303 27421
rect 19426 27412 19432 27424
rect 19484 27412 19490 27464
rect 19886 27452 19892 27464
rect 19847 27424 19892 27452
rect 19886 27412 19892 27424
rect 19944 27412 19950 27464
rect 21177 27455 21235 27461
rect 21177 27421 21189 27455
rect 21223 27452 21235 27455
rect 22664 27452 22692 27492
rect 24854 27480 24860 27532
rect 24912 27520 24918 27532
rect 25777 27523 25835 27529
rect 24912 27492 25268 27520
rect 24912 27480 24918 27492
rect 21223 27424 22692 27452
rect 23017 27455 23075 27461
rect 21223 27421 21235 27424
rect 21177 27415 21235 27421
rect 23017 27421 23029 27455
rect 23063 27421 23075 27455
rect 23842 27452 23848 27464
rect 23803 27424 23848 27452
rect 23017 27415 23075 27421
rect 19702 27384 19708 27396
rect 15120 27356 19708 27384
rect 14921 27347 14979 27353
rect 19702 27344 19708 27356
rect 19760 27344 19766 27396
rect 20622 27344 20628 27396
rect 20680 27384 20686 27396
rect 21266 27384 21272 27396
rect 20680 27356 21272 27384
rect 20680 27344 20686 27356
rect 21266 27344 21272 27356
rect 21324 27344 21330 27396
rect 21444 27387 21502 27393
rect 21444 27353 21456 27387
rect 21490 27384 21502 27387
rect 22278 27384 22284 27396
rect 21490 27356 22284 27384
rect 21490 27353 21502 27356
rect 21444 27347 21502 27353
rect 22278 27344 22284 27356
rect 22336 27344 22342 27396
rect 23032 27384 23060 27415
rect 23842 27412 23848 27424
rect 23900 27412 23906 27464
rect 23934 27412 23940 27464
rect 23992 27452 23998 27464
rect 24581 27455 24639 27461
rect 24581 27452 24593 27455
rect 23992 27424 24593 27452
rect 23992 27412 23998 27424
rect 24581 27421 24593 27424
rect 24627 27421 24639 27455
rect 25038 27452 25044 27464
rect 24999 27424 25044 27452
rect 24581 27415 24639 27421
rect 25038 27412 25044 27424
rect 25096 27412 25102 27464
rect 25240 27461 25268 27492
rect 25777 27489 25789 27523
rect 25823 27520 25835 27523
rect 29822 27520 29828 27532
rect 25823 27492 29828 27520
rect 25823 27489 25835 27492
rect 25777 27483 25835 27489
rect 29822 27480 29828 27492
rect 29880 27480 29886 27532
rect 25225 27455 25283 27461
rect 25225 27421 25237 27455
rect 25271 27421 25283 27455
rect 25225 27415 25283 27421
rect 25240 27384 25268 27415
rect 25682 27412 25688 27464
rect 25740 27452 25746 27464
rect 25869 27455 25927 27461
rect 25740 27424 25785 27452
rect 25740 27412 25746 27424
rect 25869 27421 25881 27455
rect 25915 27421 25927 27455
rect 26326 27452 26332 27464
rect 26287 27424 26332 27452
rect 25869 27415 25927 27421
rect 25314 27384 25320 27396
rect 22480 27356 23060 27384
rect 25227 27356 25320 27384
rect 15562 27316 15568 27328
rect 14292 27288 15568 27316
rect 15562 27276 15568 27288
rect 15620 27276 15626 27328
rect 15746 27276 15752 27328
rect 15804 27316 15810 27328
rect 16206 27316 16212 27328
rect 15804 27288 16212 27316
rect 15804 27276 15810 27288
rect 16206 27276 16212 27288
rect 16264 27276 16270 27328
rect 17405 27319 17463 27325
rect 17405 27285 17417 27319
rect 17451 27316 17463 27319
rect 19058 27316 19064 27328
rect 17451 27288 19064 27316
rect 17451 27285 17463 27288
rect 17405 27279 17463 27285
rect 19058 27276 19064 27288
rect 19116 27276 19122 27328
rect 19429 27319 19487 27325
rect 19429 27285 19441 27319
rect 19475 27316 19487 27319
rect 22480 27316 22508 27356
rect 25314 27344 25320 27356
rect 25372 27384 25378 27396
rect 25884 27384 25912 27415
rect 26326 27412 26332 27424
rect 26384 27412 26390 27464
rect 26513 27455 26571 27461
rect 26513 27421 26525 27455
rect 26559 27421 26571 27455
rect 26513 27415 26571 27421
rect 26528 27384 26556 27415
rect 25372 27356 26556 27384
rect 25372 27344 25378 27356
rect 19475 27288 22508 27316
rect 23661 27319 23719 27325
rect 19475 27285 19487 27288
rect 19429 27279 19487 27285
rect 23661 27285 23673 27319
rect 23707 27316 23719 27319
rect 23934 27316 23940 27328
rect 23707 27288 23940 27316
rect 23707 27285 23719 27288
rect 23661 27279 23719 27285
rect 23934 27276 23940 27288
rect 23992 27276 23998 27328
rect 24394 27316 24400 27328
rect 24355 27288 24400 27316
rect 24394 27276 24400 27288
rect 24452 27276 24458 27328
rect 25130 27316 25136 27328
rect 25091 27288 25136 27316
rect 25130 27276 25136 27288
rect 25188 27276 25194 27328
rect 1104 27226 30820 27248
rect 1104 27174 10880 27226
rect 10932 27174 10944 27226
rect 10996 27174 11008 27226
rect 11060 27174 11072 27226
rect 11124 27174 11136 27226
rect 11188 27174 20811 27226
rect 20863 27174 20875 27226
rect 20927 27174 20939 27226
rect 20991 27174 21003 27226
rect 21055 27174 21067 27226
rect 21119 27174 30820 27226
rect 1104 27152 30820 27174
rect 10502 27072 10508 27124
rect 10560 27112 10566 27124
rect 11793 27115 11851 27121
rect 11793 27112 11805 27115
rect 10560 27084 11805 27112
rect 10560 27072 10566 27084
rect 11793 27081 11805 27084
rect 11839 27081 11851 27115
rect 11793 27075 11851 27081
rect 11885 27115 11943 27121
rect 11885 27081 11897 27115
rect 11931 27081 11943 27115
rect 12986 27112 12992 27124
rect 11885 27075 11943 27081
rect 12406 27084 12992 27112
rect 11900 27044 11928 27075
rect 10704 27016 11928 27044
rect 12069 27047 12127 27053
rect 10704 26988 10732 27016
rect 12069 27013 12081 27047
rect 12115 27044 12127 27047
rect 12406 27044 12434 27084
rect 12986 27072 12992 27084
rect 13044 27072 13050 27124
rect 13262 27112 13268 27124
rect 13223 27084 13268 27112
rect 13262 27072 13268 27084
rect 13320 27072 13326 27124
rect 13817 27115 13875 27121
rect 13817 27081 13829 27115
rect 13863 27112 13875 27115
rect 15010 27112 15016 27124
rect 13863 27084 14596 27112
rect 14923 27084 15016 27112
rect 13863 27081 13875 27084
rect 13817 27075 13875 27081
rect 14458 27044 14464 27056
rect 12115 27016 12434 27044
rect 12544 27016 14464 27044
rect 12115 27013 12127 27016
rect 12069 27007 12127 27013
rect 9306 26976 9312 26988
rect 9267 26948 9312 26976
rect 9306 26936 9312 26948
rect 9364 26936 9370 26988
rect 9401 26979 9459 26985
rect 9401 26945 9413 26979
rect 9447 26976 9459 26979
rect 9950 26976 9956 26988
rect 9447 26948 9956 26976
rect 9447 26945 9459 26948
rect 9401 26939 9459 26945
rect 9950 26936 9956 26948
rect 10008 26936 10014 26988
rect 10042 26936 10048 26988
rect 10100 26976 10106 26988
rect 10321 26979 10379 26985
rect 10321 26976 10333 26979
rect 10100 26948 10333 26976
rect 10100 26936 10106 26948
rect 10321 26945 10333 26948
rect 10367 26945 10379 26979
rect 10321 26939 10379 26945
rect 10413 26979 10471 26985
rect 10413 26945 10425 26979
rect 10459 26976 10471 26979
rect 10686 26976 10692 26988
rect 10459 26948 10692 26976
rect 10459 26945 10471 26948
rect 10413 26939 10471 26945
rect 10686 26936 10692 26948
rect 10744 26936 10750 26988
rect 10778 26936 10784 26988
rect 10836 26976 10842 26988
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 10836 26948 11713 26976
rect 10836 26936 10842 26948
rect 11701 26945 11713 26948
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 12434 26936 12440 26988
rect 12492 26976 12498 26988
rect 12544 26985 12572 27016
rect 14458 27004 14464 27016
rect 14516 27004 14522 27056
rect 12529 26979 12587 26985
rect 12529 26976 12541 26979
rect 12492 26948 12541 26976
rect 12492 26936 12498 26948
rect 12529 26945 12541 26948
rect 12575 26945 12587 26979
rect 12529 26939 12587 26945
rect 12802 26936 12808 26988
rect 12860 26976 12866 26988
rect 13173 26979 13231 26985
rect 13173 26976 13185 26979
rect 12860 26948 13185 26976
rect 12860 26936 12866 26948
rect 13173 26945 13185 26948
rect 13219 26945 13231 26979
rect 13173 26939 13231 26945
rect 13262 26936 13268 26988
rect 13320 26976 13326 26988
rect 13357 26979 13415 26985
rect 13357 26976 13369 26979
rect 13320 26948 13369 26976
rect 13320 26936 13326 26948
rect 13357 26945 13369 26948
rect 13403 26945 13415 26979
rect 13357 26939 13415 26945
rect 14093 26979 14151 26985
rect 14093 26945 14105 26979
rect 14139 26945 14151 26979
rect 14274 26976 14280 26988
rect 14235 26948 14280 26976
rect 14093 26939 14151 26945
rect 8846 26868 8852 26920
rect 8904 26908 8910 26920
rect 9493 26911 9551 26917
rect 9493 26908 9505 26911
rect 8904 26880 9505 26908
rect 8904 26868 8910 26880
rect 9493 26877 9505 26880
rect 9539 26877 9551 26911
rect 10502 26908 10508 26920
rect 10463 26880 10508 26908
rect 9493 26871 9551 26877
rect 10502 26868 10508 26880
rect 10560 26868 10566 26920
rect 10597 26911 10655 26917
rect 10597 26877 10609 26911
rect 10643 26908 10655 26911
rect 13078 26908 13084 26920
rect 10643 26880 13084 26908
rect 10643 26877 10655 26880
rect 10597 26871 10655 26877
rect 1670 26800 1676 26852
rect 1728 26840 1734 26852
rect 10612 26840 10640 26871
rect 13078 26868 13084 26880
rect 13136 26868 13142 26920
rect 1728 26812 10640 26840
rect 11517 26843 11575 26849
rect 1728 26800 1734 26812
rect 11517 26809 11529 26843
rect 11563 26840 11575 26843
rect 12618 26840 12624 26852
rect 11563 26812 12434 26840
rect 12531 26812 12624 26840
rect 11563 26809 11575 26812
rect 11517 26803 11575 26809
rect 8938 26772 8944 26784
rect 8899 26744 8944 26772
rect 8938 26732 8944 26744
rect 8996 26732 9002 26784
rect 10137 26775 10195 26781
rect 10137 26741 10149 26775
rect 10183 26772 10195 26775
rect 10226 26772 10232 26784
rect 10183 26744 10232 26772
rect 10183 26741 10195 26744
rect 10137 26735 10195 26741
rect 10226 26732 10232 26744
rect 10284 26732 10290 26784
rect 12406 26772 12434 26812
rect 12618 26800 12624 26812
rect 12676 26840 12682 26852
rect 13817 26843 13875 26849
rect 13817 26840 13829 26843
rect 12676 26812 13829 26840
rect 12676 26800 12682 26812
rect 13817 26809 13829 26812
rect 13863 26809 13875 26843
rect 13817 26803 13875 26809
rect 13722 26772 13728 26784
rect 12406 26744 13728 26772
rect 13722 26732 13728 26744
rect 13780 26732 13786 26784
rect 13906 26772 13912 26784
rect 13867 26744 13912 26772
rect 13906 26732 13912 26744
rect 13964 26732 13970 26784
rect 14108 26772 14136 26939
rect 14274 26936 14280 26948
rect 14332 26936 14338 26988
rect 14369 26979 14427 26985
rect 14369 26945 14381 26979
rect 14415 26976 14427 26979
rect 14568 26976 14596 27084
rect 15010 27072 15016 27084
rect 15068 27112 15074 27124
rect 16114 27112 16120 27124
rect 15068 27084 16120 27112
rect 15068 27072 15074 27084
rect 16114 27072 16120 27084
rect 16172 27072 16178 27124
rect 17678 27072 17684 27124
rect 17736 27112 17742 27124
rect 18785 27115 18843 27121
rect 18785 27112 18797 27115
rect 17736 27084 18797 27112
rect 17736 27072 17742 27084
rect 18785 27081 18797 27084
rect 18831 27081 18843 27115
rect 19150 27112 19156 27124
rect 19111 27084 19156 27112
rect 18785 27075 18843 27081
rect 19150 27072 19156 27084
rect 19208 27072 19214 27124
rect 21910 27112 21916 27124
rect 20916 27084 21916 27112
rect 20916 27056 20944 27084
rect 21910 27072 21916 27084
rect 21968 27072 21974 27124
rect 22094 27072 22100 27124
rect 22152 27112 22158 27124
rect 22370 27112 22376 27124
rect 22152 27084 22376 27112
rect 22152 27072 22158 27084
rect 22370 27072 22376 27084
rect 22428 27072 22434 27124
rect 23566 27112 23572 27124
rect 23527 27084 23572 27112
rect 23566 27072 23572 27084
rect 23624 27072 23630 27124
rect 23934 27112 23940 27124
rect 23895 27084 23940 27112
rect 23934 27072 23940 27084
rect 23992 27072 23998 27124
rect 25317 27115 25375 27121
rect 25317 27081 25329 27115
rect 25363 27112 25375 27115
rect 26145 27115 26203 27121
rect 26145 27112 26157 27115
rect 25363 27084 26157 27112
rect 25363 27081 25375 27084
rect 25317 27075 25375 27081
rect 26145 27081 26157 27084
rect 26191 27081 26203 27115
rect 26145 27075 26203 27081
rect 15749 27047 15807 27053
rect 15749 27013 15761 27047
rect 15795 27044 15807 27047
rect 17212 27047 17270 27053
rect 15795 27016 17172 27044
rect 15795 27013 15807 27016
rect 15749 27007 15807 27013
rect 14415 26948 14596 26976
rect 14921 26979 14979 26985
rect 14415 26945 14427 26948
rect 14369 26939 14427 26945
rect 14921 26945 14933 26979
rect 14967 26945 14979 26979
rect 14921 26939 14979 26945
rect 14292 26908 14320 26936
rect 14936 26908 14964 26939
rect 16850 26936 16856 26988
rect 16908 26976 16914 26988
rect 16945 26979 17003 26985
rect 16945 26976 16957 26979
rect 16908 26948 16957 26976
rect 16908 26936 16914 26948
rect 16945 26945 16957 26948
rect 16991 26945 17003 26979
rect 17144 26976 17172 27016
rect 17212 27013 17224 27047
rect 17258 27044 17270 27047
rect 18230 27044 18236 27056
rect 17258 27016 18236 27044
rect 17258 27013 17270 27016
rect 17212 27007 17270 27013
rect 18230 27004 18236 27016
rect 18288 27004 18294 27056
rect 19886 27044 19892 27056
rect 18432 27016 19892 27044
rect 18432 26976 18460 27016
rect 19886 27004 19892 27016
rect 19944 27004 19950 27056
rect 20898 27004 20904 27056
rect 20956 27004 20962 27056
rect 23750 27044 23756 27056
rect 21008 27016 23756 27044
rect 17144 26948 18460 26976
rect 16945 26939 17003 26945
rect 18874 26936 18880 26988
rect 18932 26976 18938 26988
rect 20530 26976 20536 26988
rect 18932 26948 19380 26976
rect 20491 26948 20536 26976
rect 18932 26936 18938 26948
rect 14292 26880 14964 26908
rect 18230 26868 18236 26920
rect 18288 26908 18294 26920
rect 18690 26908 18696 26920
rect 18288 26880 18696 26908
rect 18288 26868 18294 26880
rect 18690 26868 18696 26880
rect 18748 26868 18754 26920
rect 19352 26917 19380 26948
rect 20530 26936 20536 26948
rect 20588 26936 20594 26988
rect 20622 26936 20628 26988
rect 20680 26976 20686 26988
rect 20717 26979 20775 26985
rect 20717 26976 20729 26979
rect 20680 26948 20729 26976
rect 20680 26936 20686 26948
rect 20717 26945 20729 26948
rect 20763 26945 20775 26979
rect 20717 26939 20775 26945
rect 20809 26979 20867 26985
rect 20809 26945 20821 26979
rect 20855 26976 20867 26979
rect 21008 26976 21036 27016
rect 23750 27004 23756 27016
rect 23808 27004 23814 27056
rect 25130 27004 25136 27056
rect 25188 27044 25194 27056
rect 25188 27016 29868 27044
rect 25188 27004 25194 27016
rect 20855 26948 21036 26976
rect 21085 26979 21143 26985
rect 20855 26945 20867 26948
rect 20809 26939 20867 26945
rect 21085 26945 21097 26979
rect 21131 26945 21143 26979
rect 21085 26939 21143 26945
rect 19245 26911 19303 26917
rect 19245 26877 19257 26911
rect 19291 26877 19303 26911
rect 19245 26871 19303 26877
rect 19337 26911 19395 26917
rect 19337 26877 19349 26911
rect 19383 26877 19395 26911
rect 20898 26908 20904 26920
rect 20859 26880 20904 26908
rect 19337 26871 19395 26877
rect 14185 26843 14243 26849
rect 14185 26809 14197 26843
rect 14231 26840 14243 26843
rect 15194 26840 15200 26852
rect 14231 26812 15200 26840
rect 14231 26809 14243 26812
rect 14185 26803 14243 26809
rect 15194 26800 15200 26812
rect 15252 26800 15258 26852
rect 18322 26840 18328 26852
rect 18283 26812 18328 26840
rect 18322 26800 18328 26812
rect 18380 26800 18386 26852
rect 18874 26800 18880 26852
rect 18932 26840 18938 26852
rect 19260 26840 19288 26871
rect 20898 26868 20904 26880
rect 20956 26868 20962 26920
rect 21100 26908 21128 26939
rect 21174 26936 21180 26988
rect 21232 26976 21238 26988
rect 22281 26979 22339 26985
rect 22281 26976 22293 26979
rect 21232 26948 22293 26976
rect 21232 26936 21238 26948
rect 22281 26945 22293 26948
rect 22327 26945 22339 26979
rect 22281 26939 22339 26945
rect 22462 26936 22468 26988
rect 22520 26976 22526 26988
rect 22925 26979 22983 26985
rect 22925 26976 22937 26979
rect 22520 26948 22937 26976
rect 22520 26936 22526 26948
rect 22925 26945 22937 26948
rect 22971 26945 22983 26979
rect 22925 26939 22983 26945
rect 24029 26979 24087 26985
rect 24029 26945 24041 26979
rect 24075 26976 24087 26979
rect 24302 26976 24308 26988
rect 24075 26948 24308 26976
rect 24075 26945 24087 26948
rect 24029 26939 24087 26945
rect 24302 26936 24308 26948
rect 24360 26936 24366 26988
rect 26234 26936 26240 26988
rect 26292 26976 26298 26988
rect 29840 26985 29868 27016
rect 26329 26979 26387 26985
rect 26329 26976 26341 26979
rect 26292 26948 26341 26976
rect 26292 26936 26298 26948
rect 26329 26945 26341 26948
rect 26375 26945 26387 26979
rect 26329 26939 26387 26945
rect 29825 26979 29883 26985
rect 29825 26945 29837 26979
rect 29871 26945 29883 26979
rect 29825 26939 29883 26945
rect 21910 26908 21916 26920
rect 21100 26880 21916 26908
rect 21910 26868 21916 26880
rect 21968 26868 21974 26920
rect 24213 26911 24271 26917
rect 24213 26877 24225 26911
rect 24259 26877 24271 26911
rect 25406 26908 25412 26920
rect 25367 26880 25412 26908
rect 24213 26871 24271 26877
rect 18932 26812 19288 26840
rect 18932 26800 18938 26812
rect 20530 26800 20536 26852
rect 20588 26840 20594 26852
rect 23109 26843 23167 26849
rect 23109 26840 23121 26843
rect 20588 26812 23121 26840
rect 20588 26800 20594 26812
rect 23109 26809 23121 26812
rect 23155 26809 23167 26843
rect 24228 26840 24256 26871
rect 25406 26868 25412 26880
rect 25464 26868 25470 26920
rect 25498 26868 25504 26920
rect 25556 26908 25562 26920
rect 25556 26880 25601 26908
rect 25556 26868 25562 26880
rect 24670 26840 24676 26852
rect 24228 26812 24676 26840
rect 23109 26803 23167 26809
rect 24670 26800 24676 26812
rect 24728 26840 24734 26852
rect 25516 26840 25544 26868
rect 30006 26840 30012 26852
rect 24728 26812 25544 26840
rect 29967 26812 30012 26840
rect 24728 26800 24734 26812
rect 30006 26800 30012 26812
rect 30064 26800 30070 26852
rect 14642 26772 14648 26784
rect 14108 26744 14648 26772
rect 14642 26732 14648 26744
rect 14700 26772 14706 26784
rect 15286 26772 15292 26784
rect 14700 26744 15292 26772
rect 14700 26732 14706 26744
rect 15286 26732 15292 26744
rect 15344 26732 15350 26784
rect 15470 26732 15476 26784
rect 15528 26772 15534 26784
rect 16025 26775 16083 26781
rect 16025 26772 16037 26775
rect 15528 26744 16037 26772
rect 15528 26732 15534 26744
rect 16025 26741 16037 26744
rect 16071 26772 16083 26775
rect 16298 26772 16304 26784
rect 16071 26744 16304 26772
rect 16071 26741 16083 26744
rect 16025 26735 16083 26741
rect 16298 26732 16304 26744
rect 16356 26732 16362 26784
rect 21266 26772 21272 26784
rect 21227 26744 21272 26772
rect 21266 26732 21272 26744
rect 21324 26732 21330 26784
rect 24949 26775 25007 26781
rect 24949 26741 24961 26775
rect 24995 26772 25007 26775
rect 25682 26772 25688 26784
rect 24995 26744 25688 26772
rect 24995 26741 25007 26744
rect 24949 26735 25007 26741
rect 25682 26732 25688 26744
rect 25740 26732 25746 26784
rect 1104 26682 30820 26704
rect 1104 26630 5915 26682
rect 5967 26630 5979 26682
rect 6031 26630 6043 26682
rect 6095 26630 6107 26682
rect 6159 26630 6171 26682
rect 6223 26630 15846 26682
rect 15898 26630 15910 26682
rect 15962 26630 15974 26682
rect 16026 26630 16038 26682
rect 16090 26630 16102 26682
rect 16154 26630 25776 26682
rect 25828 26630 25840 26682
rect 25892 26630 25904 26682
rect 25956 26630 25968 26682
rect 26020 26630 26032 26682
rect 26084 26630 30820 26682
rect 1104 26608 30820 26630
rect 9582 26528 9588 26580
rect 9640 26568 9646 26580
rect 10873 26571 10931 26577
rect 10873 26568 10885 26571
rect 9640 26540 10885 26568
rect 9640 26528 9646 26540
rect 10873 26537 10885 26540
rect 10919 26568 10931 26571
rect 11330 26568 11336 26580
rect 10919 26540 11336 26568
rect 10919 26537 10931 26540
rect 10873 26531 10931 26537
rect 11330 26528 11336 26540
rect 11388 26528 11394 26580
rect 12802 26568 12808 26580
rect 12763 26540 12808 26568
rect 12802 26528 12808 26540
rect 12860 26528 12866 26580
rect 14553 26571 14611 26577
rect 13004 26540 14504 26568
rect 9674 26460 9680 26512
rect 9732 26500 9738 26512
rect 13004 26500 13032 26540
rect 9732 26472 13032 26500
rect 13081 26503 13139 26509
rect 9732 26460 9738 26472
rect 13081 26469 13093 26503
rect 13127 26500 13139 26503
rect 13906 26500 13912 26512
rect 13127 26472 13912 26500
rect 13127 26469 13139 26472
rect 13081 26463 13139 26469
rect 13906 26460 13912 26472
rect 13964 26460 13970 26512
rect 14476 26500 14504 26540
rect 14553 26537 14565 26571
rect 14599 26568 14611 26571
rect 15194 26568 15200 26580
rect 14599 26540 15200 26568
rect 14599 26537 14611 26540
rect 14553 26531 14611 26537
rect 15194 26528 15200 26540
rect 15252 26528 15258 26580
rect 16850 26528 16856 26580
rect 16908 26568 16914 26580
rect 17310 26568 17316 26580
rect 16908 26540 17316 26568
rect 16908 26528 16914 26540
rect 17310 26528 17316 26540
rect 17368 26568 17374 26580
rect 19981 26571 20039 26577
rect 19981 26568 19993 26571
rect 17368 26540 19993 26568
rect 17368 26528 17374 26540
rect 19981 26537 19993 26540
rect 20027 26537 20039 26571
rect 19981 26531 20039 26537
rect 20070 26528 20076 26580
rect 20128 26568 20134 26580
rect 21910 26568 21916 26580
rect 20128 26540 21496 26568
rect 21871 26540 21916 26568
rect 20128 26528 20134 26540
rect 15289 26503 15347 26509
rect 14476 26472 15240 26500
rect 8938 26392 8944 26444
rect 8996 26432 9002 26444
rect 10689 26435 10747 26441
rect 10689 26432 10701 26435
rect 8996 26404 10701 26432
rect 8996 26392 9002 26404
rect 10689 26401 10701 26404
rect 10735 26401 10747 26435
rect 10689 26395 10747 26401
rect 13265 26435 13323 26441
rect 13265 26401 13277 26435
rect 13311 26432 13323 26435
rect 13814 26432 13820 26444
rect 13311 26404 13820 26432
rect 13311 26401 13323 26404
rect 13265 26395 13323 26401
rect 13814 26392 13820 26404
rect 13872 26392 13878 26444
rect 14185 26435 14243 26441
rect 14185 26401 14197 26435
rect 14231 26432 14243 26435
rect 14274 26432 14280 26444
rect 14231 26404 14280 26432
rect 14231 26401 14243 26404
rect 14185 26395 14243 26401
rect 14274 26392 14280 26404
rect 14332 26392 14338 26444
rect 15010 26432 15016 26444
rect 14384 26404 15016 26432
rect 9030 26364 9036 26376
rect 8991 26336 9036 26364
rect 9030 26324 9036 26336
rect 9088 26324 9094 26376
rect 9122 26324 9128 26376
rect 9180 26364 9186 26376
rect 9309 26367 9367 26373
rect 9309 26364 9321 26367
rect 9180 26336 9321 26364
rect 9180 26324 9186 26336
rect 9309 26333 9321 26336
rect 9355 26364 9367 26367
rect 10321 26367 10379 26373
rect 10321 26364 10333 26367
rect 9355 26336 10333 26364
rect 9355 26333 9367 26336
rect 9309 26327 9367 26333
rect 10321 26333 10333 26336
rect 10367 26333 10379 26367
rect 10321 26327 10379 26333
rect 11238 26324 11244 26376
rect 11296 26364 11302 26376
rect 12158 26364 12164 26376
rect 11296 26336 12164 26364
rect 11296 26324 11302 26336
rect 12158 26324 12164 26336
rect 12216 26324 12222 26376
rect 12986 26364 12992 26376
rect 12947 26336 12992 26364
rect 12986 26324 12992 26336
rect 13044 26324 13050 26376
rect 13170 26364 13176 26376
rect 13131 26336 13176 26364
rect 13170 26324 13176 26336
rect 13228 26324 13234 26376
rect 14384 26373 14412 26404
rect 15010 26392 15016 26404
rect 15068 26392 15074 26444
rect 15212 26432 15240 26472
rect 15289 26469 15301 26503
rect 15335 26500 15347 26503
rect 16022 26500 16028 26512
rect 15335 26472 16028 26500
rect 15335 26469 15347 26472
rect 15289 26463 15347 26469
rect 16022 26460 16028 26472
rect 16080 26460 16086 26512
rect 21468 26500 21496 26540
rect 21910 26528 21916 26540
rect 21968 26528 21974 26580
rect 22646 26568 22652 26580
rect 22607 26540 22652 26568
rect 22646 26528 22652 26540
rect 22704 26528 22710 26580
rect 24857 26571 24915 26577
rect 24857 26537 24869 26571
rect 24903 26568 24915 26571
rect 26326 26568 26332 26580
rect 24903 26540 26332 26568
rect 24903 26537 24915 26540
rect 24857 26531 24915 26537
rect 26326 26528 26332 26540
rect 26384 26528 26390 26580
rect 26237 26503 26295 26509
rect 26237 26500 26249 26503
rect 21468 26472 26249 26500
rect 26237 26469 26249 26472
rect 26283 26469 26295 26503
rect 26237 26463 26295 26469
rect 18874 26432 18880 26444
rect 15212 26404 18880 26432
rect 13449 26367 13507 26373
rect 13449 26333 13461 26367
rect 13495 26364 13507 26367
rect 14369 26367 14427 26373
rect 14369 26364 14381 26367
rect 13495 26336 14381 26364
rect 13495 26333 13507 26336
rect 13449 26327 13507 26333
rect 14369 26333 14381 26336
rect 14415 26333 14427 26367
rect 14369 26327 14427 26333
rect 14642 26324 14648 26376
rect 14700 26364 14706 26376
rect 15470 26364 15476 26376
rect 14700 26336 14745 26364
rect 15431 26336 15476 26364
rect 14700 26324 14706 26336
rect 15470 26324 15476 26336
rect 15528 26324 15534 26376
rect 15948 26373 15976 26404
rect 18874 26392 18880 26404
rect 18932 26392 18938 26444
rect 20530 26432 20536 26444
rect 20491 26404 20536 26432
rect 20530 26392 20536 26404
rect 20588 26392 20594 26444
rect 22925 26435 22983 26441
rect 22925 26401 22937 26435
rect 22971 26432 22983 26435
rect 23658 26432 23664 26444
rect 22971 26404 23664 26432
rect 22971 26401 22983 26404
rect 22925 26395 22983 26401
rect 23658 26392 23664 26404
rect 23716 26392 23722 26444
rect 25498 26432 25504 26444
rect 25459 26404 25504 26432
rect 25498 26392 25504 26404
rect 25556 26392 25562 26444
rect 15933 26367 15991 26373
rect 15933 26333 15945 26367
rect 15979 26333 15991 26367
rect 15933 26327 15991 26333
rect 16761 26367 16819 26373
rect 16761 26333 16773 26367
rect 16807 26364 16819 26367
rect 17954 26364 17960 26376
rect 16807 26336 17960 26364
rect 16807 26333 16819 26336
rect 16761 26327 16819 26333
rect 17954 26324 17960 26336
rect 18012 26324 18018 26376
rect 18414 26324 18420 26376
rect 18472 26364 18478 26376
rect 18509 26367 18567 26373
rect 18509 26364 18521 26367
rect 18472 26336 18521 26364
rect 18472 26324 18478 26336
rect 18509 26333 18521 26336
rect 18555 26364 18567 26367
rect 19150 26364 19156 26376
rect 18555 26336 19156 26364
rect 18555 26333 18567 26336
rect 18509 26327 18567 26333
rect 19150 26324 19156 26336
rect 19208 26324 19214 26376
rect 19889 26367 19947 26373
rect 19889 26333 19901 26367
rect 19935 26364 19947 26367
rect 21174 26364 21180 26376
rect 19935 26336 21180 26364
rect 19935 26333 19947 26336
rect 19889 26327 19947 26333
rect 21174 26324 21180 26336
rect 21232 26324 21238 26376
rect 22465 26367 22523 26373
rect 22465 26333 22477 26367
rect 22511 26364 22523 26367
rect 22554 26364 22560 26376
rect 22511 26336 22560 26364
rect 22511 26333 22523 26336
rect 22465 26327 22523 26333
rect 22554 26324 22560 26336
rect 22612 26324 22618 26376
rect 23566 26364 23572 26376
rect 23527 26336 23572 26364
rect 23566 26324 23572 26336
rect 23624 26324 23630 26376
rect 25222 26364 25228 26376
rect 25183 26336 25228 26364
rect 25222 26324 25228 26336
rect 25280 26324 25286 26376
rect 26053 26367 26111 26373
rect 26053 26333 26065 26367
rect 26099 26364 26111 26367
rect 26786 26364 26792 26376
rect 26099 26336 26792 26364
rect 26099 26333 26111 26336
rect 26053 26327 26111 26333
rect 26786 26324 26792 26336
rect 26844 26324 26850 26376
rect 29822 26364 29828 26376
rect 29783 26336 29828 26364
rect 29822 26324 29828 26336
rect 29880 26324 29886 26376
rect 12253 26299 12311 26305
rect 10428 26268 10732 26296
rect 2222 26188 2228 26240
rect 2280 26228 2286 26240
rect 10428 26228 10456 26268
rect 2280 26200 10456 26228
rect 2280 26188 2286 26200
rect 10502 26188 10508 26240
rect 10560 26228 10566 26240
rect 10704 26228 10732 26268
rect 12253 26265 12265 26299
rect 12299 26296 12311 26299
rect 13354 26296 13360 26308
rect 12299 26268 13360 26296
rect 12299 26265 12311 26268
rect 12253 26259 12311 26265
rect 13354 26256 13360 26268
rect 13412 26256 13418 26308
rect 13722 26256 13728 26308
rect 13780 26296 13786 26308
rect 15194 26296 15200 26308
rect 13780 26268 15200 26296
rect 13780 26256 13786 26268
rect 15194 26256 15200 26268
rect 15252 26256 15258 26308
rect 16025 26299 16083 26305
rect 16025 26265 16037 26299
rect 16071 26296 16083 26299
rect 16482 26296 16488 26308
rect 16071 26268 16488 26296
rect 16071 26265 16083 26268
rect 16025 26259 16083 26265
rect 16482 26256 16488 26268
rect 16540 26256 16546 26308
rect 16666 26256 16672 26308
rect 16724 26296 16730 26308
rect 17497 26299 17555 26305
rect 17497 26296 17509 26299
rect 16724 26268 17509 26296
rect 16724 26256 16730 26268
rect 17497 26265 17509 26268
rect 17543 26265 17555 26299
rect 17497 26259 17555 26265
rect 18601 26299 18659 26305
rect 18601 26265 18613 26299
rect 18647 26296 18659 26299
rect 19518 26296 19524 26308
rect 18647 26268 19524 26296
rect 18647 26265 18659 26268
rect 18601 26259 18659 26265
rect 19518 26256 19524 26268
rect 19576 26296 19582 26308
rect 20254 26296 20260 26308
rect 19576 26268 20260 26296
rect 19576 26256 19582 26268
rect 20254 26256 20260 26268
rect 20312 26256 20318 26308
rect 20800 26299 20858 26305
rect 20800 26265 20812 26299
rect 20846 26296 20858 26299
rect 21266 26296 21272 26308
rect 20846 26268 21272 26296
rect 20846 26265 20858 26268
rect 20800 26259 20858 26265
rect 21266 26256 21272 26268
rect 21324 26256 21330 26308
rect 24486 26256 24492 26308
rect 24544 26296 24550 26308
rect 25317 26299 25375 26305
rect 25317 26296 25329 26299
rect 24544 26268 25329 26296
rect 24544 26256 24550 26268
rect 25317 26265 25329 26268
rect 25363 26265 25375 26299
rect 25317 26259 25375 26265
rect 15930 26228 15936 26240
rect 10560 26200 10605 26228
rect 10704 26200 15936 26228
rect 10560 26188 10566 26200
rect 15930 26188 15936 26200
rect 15988 26188 15994 26240
rect 23385 26231 23443 26237
rect 23385 26197 23397 26231
rect 23431 26228 23443 26231
rect 23474 26228 23480 26240
rect 23431 26200 23480 26228
rect 23431 26197 23443 26200
rect 23385 26191 23443 26197
rect 23474 26188 23480 26200
rect 23532 26188 23538 26240
rect 30006 26228 30012 26240
rect 29967 26200 30012 26228
rect 30006 26188 30012 26200
rect 30064 26188 30070 26240
rect 1104 26138 30820 26160
rect 1104 26086 10880 26138
rect 10932 26086 10944 26138
rect 10996 26086 11008 26138
rect 11060 26086 11072 26138
rect 11124 26086 11136 26138
rect 11188 26086 20811 26138
rect 20863 26086 20875 26138
rect 20927 26086 20939 26138
rect 20991 26086 21003 26138
rect 21055 26086 21067 26138
rect 21119 26086 30820 26138
rect 1104 26064 30820 26086
rect 1394 25984 1400 26036
rect 1452 26024 1458 26036
rect 1673 26027 1731 26033
rect 1673 26024 1685 26027
rect 1452 25996 1685 26024
rect 1452 25984 1458 25996
rect 1673 25993 1685 25996
rect 1719 25993 1731 26027
rect 2314 26024 2320 26036
rect 2275 25996 2320 26024
rect 1673 25987 1731 25993
rect 2314 25984 2320 25996
rect 2372 25984 2378 26036
rect 11517 26027 11575 26033
rect 11517 25993 11529 26027
rect 11563 26024 11575 26027
rect 11563 25996 12434 26024
rect 11563 25993 11575 25996
rect 11517 25987 11575 25993
rect 5258 25956 5264 25968
rect 1596 25928 5264 25956
rect 1596 25897 1624 25928
rect 5258 25916 5264 25928
rect 5316 25916 5322 25968
rect 9769 25959 9827 25965
rect 9769 25956 9781 25959
rect 5368 25928 9781 25956
rect 1581 25891 1639 25897
rect 1581 25857 1593 25891
rect 1627 25857 1639 25891
rect 1762 25888 1768 25900
rect 1723 25860 1768 25888
rect 1581 25851 1639 25857
rect 1762 25848 1768 25860
rect 1820 25848 1826 25900
rect 2222 25888 2228 25900
rect 2183 25860 2228 25888
rect 2222 25848 2228 25860
rect 2280 25848 2286 25900
rect 2409 25891 2467 25897
rect 2409 25857 2421 25891
rect 2455 25888 2467 25891
rect 5368 25888 5396 25928
rect 9769 25925 9781 25928
rect 9815 25925 9827 25959
rect 10781 25959 10839 25965
rect 10781 25956 10793 25959
rect 9769 25919 9827 25925
rect 9876 25928 10793 25956
rect 9122 25888 9128 25900
rect 2455 25860 5396 25888
rect 9083 25860 9128 25888
rect 2455 25857 2467 25860
rect 2409 25851 2467 25857
rect 1780 25820 1808 25848
rect 2424 25820 2452 25851
rect 9122 25848 9128 25860
rect 9180 25848 9186 25900
rect 9214 25848 9220 25900
rect 9272 25888 9278 25900
rect 9309 25891 9367 25897
rect 9309 25888 9321 25891
rect 9272 25860 9321 25888
rect 9272 25848 9278 25860
rect 9309 25857 9321 25860
rect 9355 25888 9367 25891
rect 9876 25888 9904 25928
rect 10781 25925 10793 25928
rect 10827 25956 10839 25959
rect 12406 25956 12434 25996
rect 13814 25984 13820 26036
rect 13872 26024 13878 26036
rect 14185 26027 14243 26033
rect 14185 26024 14197 26027
rect 13872 25996 14197 26024
rect 13872 25984 13878 25996
rect 14185 25993 14197 25996
rect 14231 25993 14243 26027
rect 14185 25987 14243 25993
rect 15930 25984 15936 26036
rect 15988 26024 15994 26036
rect 17037 26027 17095 26033
rect 17037 26024 17049 26027
rect 15988 25996 17049 26024
rect 15988 25984 15994 25996
rect 17037 25993 17049 25996
rect 17083 25993 17095 26027
rect 17037 25987 17095 25993
rect 18046 25984 18052 26036
rect 18104 26024 18110 26036
rect 20441 26027 20499 26033
rect 18104 25996 20208 26024
rect 18104 25984 18110 25996
rect 12986 25956 12992 25968
rect 10827 25928 12112 25956
rect 12406 25928 12992 25956
rect 10827 25925 10839 25928
rect 10781 25919 10839 25925
rect 9355 25860 9904 25888
rect 10597 25891 10655 25897
rect 9355 25857 9367 25860
rect 9309 25851 9367 25857
rect 10597 25857 10609 25891
rect 10643 25857 10655 25891
rect 11885 25891 11943 25897
rect 11885 25888 11897 25891
rect 10597 25851 10655 25857
rect 11164 25860 11897 25888
rect 1780 25792 2452 25820
rect 9033 25823 9091 25829
rect 9033 25789 9045 25823
rect 9079 25789 9091 25823
rect 9140 25820 9168 25848
rect 10612 25820 10640 25851
rect 11164 25832 11192 25860
rect 11885 25857 11897 25860
rect 11931 25857 11943 25891
rect 11885 25851 11943 25857
rect 11146 25820 11152 25832
rect 9140 25792 11152 25820
rect 9033 25783 9091 25789
rect 9048 25752 9076 25783
rect 11146 25780 11152 25792
rect 11204 25780 11210 25832
rect 11974 25820 11980 25832
rect 11935 25792 11980 25820
rect 11974 25780 11980 25792
rect 12032 25780 12038 25832
rect 12084 25829 12112 25928
rect 12986 25916 12992 25928
rect 13044 25956 13050 25968
rect 14461 25959 14519 25965
rect 14461 25956 14473 25959
rect 13044 25928 14473 25956
rect 13044 25916 13050 25928
rect 14461 25925 14473 25928
rect 14507 25925 14519 25959
rect 14461 25919 14519 25925
rect 15562 25916 15568 25968
rect 15620 25956 15626 25968
rect 18877 25959 18935 25965
rect 15620 25928 18184 25956
rect 15620 25916 15626 25928
rect 13078 25848 13084 25900
rect 13136 25888 13142 25900
rect 13265 25891 13323 25897
rect 13265 25888 13277 25891
rect 13136 25860 13277 25888
rect 13136 25848 13142 25860
rect 13265 25857 13277 25860
rect 13311 25857 13323 25891
rect 13265 25851 13323 25857
rect 13354 25848 13360 25900
rect 13412 25888 13418 25900
rect 13449 25891 13507 25897
rect 13449 25888 13461 25891
rect 13412 25860 13461 25888
rect 13412 25848 13418 25860
rect 13449 25857 13461 25860
rect 13495 25857 13507 25891
rect 13449 25851 13507 25857
rect 13541 25891 13599 25897
rect 13541 25857 13553 25891
rect 13587 25857 13599 25891
rect 13722 25888 13728 25900
rect 13683 25860 13728 25888
rect 13541 25851 13599 25857
rect 12069 25823 12127 25829
rect 12069 25789 12081 25823
rect 12115 25789 12127 25823
rect 12069 25783 12127 25789
rect 12710 25780 12716 25832
rect 12768 25820 12774 25832
rect 13556 25820 13584 25851
rect 13722 25848 13728 25860
rect 13780 25848 13786 25900
rect 13814 25848 13820 25900
rect 13872 25888 13878 25900
rect 14185 25891 14243 25897
rect 14185 25888 14197 25891
rect 13872 25860 14197 25888
rect 13872 25848 13878 25860
rect 14185 25857 14197 25860
rect 14231 25888 14243 25891
rect 14550 25888 14556 25900
rect 14231 25860 14556 25888
rect 14231 25857 14243 25860
rect 14185 25851 14243 25857
rect 14550 25848 14556 25860
rect 14608 25848 14614 25900
rect 14918 25848 14924 25900
rect 14976 25888 14982 25900
rect 15749 25891 15807 25897
rect 15749 25888 15761 25891
rect 14976 25860 15761 25888
rect 14976 25848 14982 25860
rect 15749 25857 15761 25860
rect 15795 25857 15807 25891
rect 15749 25851 15807 25857
rect 17221 25891 17279 25897
rect 17221 25857 17233 25891
rect 17267 25857 17279 25891
rect 17221 25851 17279 25857
rect 17313 25891 17371 25897
rect 17313 25857 17325 25891
rect 17359 25888 17371 25891
rect 17494 25888 17500 25900
rect 17359 25860 17500 25888
rect 17359 25857 17371 25860
rect 17313 25851 17371 25857
rect 12768 25792 13584 25820
rect 12768 25780 12774 25792
rect 13280 25764 13308 25792
rect 15654 25780 15660 25832
rect 15712 25820 15718 25832
rect 15841 25823 15899 25829
rect 15841 25820 15853 25823
rect 15712 25792 15853 25820
rect 15712 25780 15718 25792
rect 15841 25789 15853 25792
rect 15887 25789 15899 25823
rect 15841 25783 15899 25789
rect 15933 25823 15991 25829
rect 15933 25789 15945 25823
rect 15979 25789 15991 25823
rect 15933 25783 15991 25789
rect 10594 25752 10600 25764
rect 9048 25724 10600 25752
rect 10594 25712 10600 25724
rect 10652 25712 10658 25764
rect 10965 25755 11023 25761
rect 10965 25721 10977 25755
rect 11011 25752 11023 25755
rect 12434 25752 12440 25764
rect 11011 25724 12440 25752
rect 11011 25721 11023 25724
rect 10965 25715 11023 25721
rect 12434 25712 12440 25724
rect 12492 25752 12498 25764
rect 12894 25752 12900 25764
rect 12492 25724 12900 25752
rect 12492 25712 12498 25724
rect 12894 25712 12900 25724
rect 12952 25712 12958 25764
rect 13262 25712 13268 25764
rect 13320 25712 13326 25764
rect 13357 25755 13415 25761
rect 13357 25721 13369 25755
rect 13403 25752 13415 25755
rect 13906 25752 13912 25764
rect 13403 25724 13912 25752
rect 13403 25721 13415 25724
rect 13357 25715 13415 25721
rect 13906 25712 13912 25724
rect 13964 25752 13970 25764
rect 14277 25755 14335 25761
rect 14277 25752 14289 25755
rect 13964 25724 14289 25752
rect 13964 25712 13970 25724
rect 14277 25721 14289 25724
rect 14323 25721 14335 25755
rect 14277 25715 14335 25721
rect 15102 25712 15108 25764
rect 15160 25752 15166 25764
rect 15470 25752 15476 25764
rect 15160 25724 15476 25752
rect 15160 25712 15166 25724
rect 15470 25712 15476 25724
rect 15528 25752 15534 25764
rect 15948 25752 15976 25783
rect 16390 25780 16396 25832
rect 16448 25820 16454 25832
rect 16850 25820 16856 25832
rect 16448 25792 16856 25820
rect 16448 25780 16454 25792
rect 16850 25780 16856 25792
rect 16908 25780 16914 25832
rect 15528 25724 15976 25752
rect 17236 25752 17264 25851
rect 17494 25848 17500 25860
rect 17552 25848 17558 25900
rect 17589 25891 17647 25897
rect 17589 25857 17601 25891
rect 17635 25888 17647 25891
rect 17862 25888 17868 25900
rect 17635 25860 17868 25888
rect 17635 25857 17647 25860
rect 17589 25851 17647 25857
rect 17862 25848 17868 25860
rect 17920 25848 17926 25900
rect 18046 25888 18052 25900
rect 18007 25860 18052 25888
rect 18046 25848 18052 25860
rect 18104 25848 18110 25900
rect 18156 25888 18184 25928
rect 18877 25925 18889 25959
rect 18923 25956 18935 25959
rect 18966 25956 18972 25968
rect 18923 25928 18972 25956
rect 18923 25925 18935 25928
rect 18877 25919 18935 25925
rect 18966 25916 18972 25928
rect 19024 25916 19030 25968
rect 18156 25860 19092 25888
rect 18322 25780 18328 25832
rect 18380 25820 18386 25832
rect 18969 25823 19027 25829
rect 18969 25820 18981 25823
rect 18380 25792 18981 25820
rect 18380 25780 18386 25792
rect 18969 25789 18981 25792
rect 19015 25789 19027 25823
rect 19064 25820 19092 25860
rect 19150 25848 19156 25900
rect 19208 25888 19214 25900
rect 20070 25888 20076 25900
rect 19208 25860 19253 25888
rect 20031 25860 20076 25888
rect 19208 25848 19214 25860
rect 20070 25848 20076 25860
rect 20128 25848 20134 25900
rect 20180 25888 20208 25996
rect 20441 25993 20453 26027
rect 20487 26024 20499 26027
rect 20622 26024 20628 26036
rect 20487 25996 20628 26024
rect 20487 25993 20499 25996
rect 20441 25987 20499 25993
rect 20622 25984 20628 25996
rect 20680 25984 20686 26036
rect 20714 25984 20720 26036
rect 20772 26024 20778 26036
rect 20993 26027 21051 26033
rect 20993 26024 21005 26027
rect 20772 25996 21005 26024
rect 20772 25984 20778 25996
rect 20993 25993 21005 25996
rect 21039 25993 21051 26027
rect 20993 25987 21051 25993
rect 23385 26027 23443 26033
rect 23385 25993 23397 26027
rect 23431 26024 23443 26027
rect 23566 26024 23572 26036
rect 23431 25996 23572 26024
rect 23431 25993 23443 25996
rect 23385 25987 23443 25993
rect 23566 25984 23572 25996
rect 23624 25984 23630 26036
rect 24305 26027 24363 26033
rect 24305 25993 24317 26027
rect 24351 26024 24363 26027
rect 24394 26024 24400 26036
rect 24351 25996 24400 26024
rect 24351 25993 24363 25996
rect 24305 25987 24363 25993
rect 24394 25984 24400 25996
rect 24452 25984 24458 26036
rect 25225 26027 25283 26033
rect 25225 25993 25237 26027
rect 25271 26024 25283 26027
rect 29822 26024 29828 26036
rect 25271 25996 29828 26024
rect 25271 25993 25283 25996
rect 25225 25987 25283 25993
rect 29822 25984 29828 25996
rect 29880 25984 29886 26036
rect 20254 25916 20260 25968
rect 20312 25956 20318 25968
rect 26694 25956 26700 25968
rect 20312 25928 21128 25956
rect 20312 25916 20318 25928
rect 21100 25897 21128 25928
rect 23032 25928 26700 25956
rect 20901 25891 20959 25897
rect 20901 25888 20913 25891
rect 20180 25860 20913 25888
rect 20901 25857 20913 25860
rect 20947 25857 20959 25891
rect 20901 25851 20959 25857
rect 21085 25891 21143 25897
rect 21085 25857 21097 25891
rect 21131 25857 21143 25891
rect 21085 25851 21143 25857
rect 21910 25848 21916 25900
rect 21968 25888 21974 25900
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21968 25860 22017 25888
rect 21968 25848 21974 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 22830 25848 22836 25900
rect 22888 25888 22894 25900
rect 22925 25891 22983 25897
rect 22925 25888 22937 25891
rect 22888 25860 22937 25888
rect 22888 25848 22894 25860
rect 22925 25857 22937 25860
rect 22971 25857 22983 25891
rect 22925 25851 22983 25857
rect 23032 25820 23060 25928
rect 26694 25916 26700 25928
rect 26752 25956 26758 25968
rect 27433 25959 27491 25965
rect 27433 25956 27445 25959
rect 26752 25928 27445 25956
rect 26752 25916 26758 25928
rect 27433 25925 27445 25928
rect 27479 25925 27491 25959
rect 27433 25919 27491 25925
rect 23106 25848 23112 25900
rect 23164 25888 23170 25900
rect 25133 25891 25191 25897
rect 25133 25888 25145 25891
rect 23164 25860 25145 25888
rect 23164 25848 23170 25860
rect 25133 25857 25145 25860
rect 25179 25857 25191 25891
rect 25314 25888 25320 25900
rect 25275 25860 25320 25888
rect 25133 25851 25191 25857
rect 25314 25848 25320 25860
rect 25372 25848 25378 25900
rect 29825 25891 29883 25897
rect 29825 25857 29837 25891
rect 29871 25857 29883 25891
rect 29825 25851 29883 25857
rect 24394 25820 24400 25832
rect 19064 25792 23060 25820
rect 24355 25792 24400 25820
rect 18969 25783 19027 25789
rect 24394 25780 24400 25792
rect 24452 25780 24458 25832
rect 24581 25823 24639 25829
rect 24581 25789 24593 25823
rect 24627 25820 24639 25823
rect 24670 25820 24676 25832
rect 24627 25792 24676 25820
rect 24627 25789 24639 25792
rect 24581 25783 24639 25789
rect 24670 25780 24676 25792
rect 24728 25780 24734 25832
rect 26326 25780 26332 25832
rect 26384 25820 26390 25832
rect 29840 25820 29868 25851
rect 26384 25792 29868 25820
rect 26384 25780 26390 25792
rect 17586 25752 17592 25764
rect 17236 25724 17592 25752
rect 15528 25712 15534 25724
rect 17586 25712 17592 25724
rect 17644 25712 17650 25764
rect 17678 25712 17684 25764
rect 17736 25752 17742 25764
rect 18233 25755 18291 25761
rect 18233 25752 18245 25755
rect 17736 25724 18245 25752
rect 17736 25712 17742 25724
rect 18233 25721 18245 25724
rect 18279 25752 18291 25755
rect 18279 25724 20576 25752
rect 18279 25721 18291 25724
rect 18233 25715 18291 25721
rect 1302 25644 1308 25696
rect 1360 25684 1366 25696
rect 9490 25684 9496 25696
rect 1360 25656 9496 25684
rect 1360 25644 1366 25656
rect 9490 25644 9496 25656
rect 9548 25644 9554 25696
rect 13081 25687 13139 25693
rect 13081 25653 13093 25687
rect 13127 25684 13139 25687
rect 13998 25684 14004 25696
rect 13127 25656 14004 25684
rect 13127 25653 13139 25656
rect 13081 25647 13139 25653
rect 13998 25644 14004 25656
rect 14056 25644 14062 25696
rect 15381 25687 15439 25693
rect 15381 25653 15393 25687
rect 15427 25684 15439 25687
rect 16390 25684 16396 25696
rect 15427 25656 16396 25684
rect 15427 25653 15439 25656
rect 15381 25647 15439 25653
rect 16390 25644 16396 25656
rect 16448 25644 16454 25696
rect 17494 25684 17500 25696
rect 17455 25656 17500 25684
rect 17494 25644 17500 25656
rect 17552 25644 17558 25696
rect 18874 25684 18880 25696
rect 18835 25656 18880 25684
rect 18874 25644 18880 25656
rect 18932 25644 18938 25696
rect 19337 25687 19395 25693
rect 19337 25653 19349 25687
rect 19383 25684 19395 25687
rect 20346 25684 20352 25696
rect 19383 25656 20352 25684
rect 19383 25653 19395 25656
rect 19337 25647 19395 25653
rect 20346 25644 20352 25656
rect 20404 25644 20410 25696
rect 20548 25684 20576 25724
rect 20622 25712 20628 25764
rect 20680 25752 20686 25764
rect 22186 25752 22192 25764
rect 20680 25724 22192 25752
rect 20680 25712 20686 25724
rect 22186 25712 22192 25724
rect 22244 25712 22250 25764
rect 22646 25752 22652 25764
rect 22296 25724 22652 25752
rect 21450 25684 21456 25696
rect 20548 25656 21456 25684
rect 21450 25644 21456 25656
rect 21508 25644 21514 25696
rect 22296 25693 22324 25724
rect 22646 25712 22652 25724
rect 22704 25752 22710 25764
rect 23937 25755 23995 25761
rect 22704 25724 23060 25752
rect 22704 25712 22710 25724
rect 22281 25687 22339 25693
rect 22281 25653 22293 25687
rect 22327 25653 22339 25687
rect 22462 25684 22468 25696
rect 22423 25656 22468 25684
rect 22281 25647 22339 25653
rect 22462 25644 22468 25656
rect 22520 25644 22526 25696
rect 23032 25693 23060 25724
rect 23937 25721 23949 25755
rect 23983 25752 23995 25755
rect 25038 25752 25044 25764
rect 23983 25724 25044 25752
rect 23983 25721 23995 25724
rect 23937 25715 23995 25721
rect 25038 25712 25044 25724
rect 25096 25712 25102 25764
rect 27614 25752 27620 25764
rect 27575 25724 27620 25752
rect 27614 25712 27620 25724
rect 27672 25712 27678 25764
rect 23017 25687 23075 25693
rect 23017 25653 23029 25687
rect 23063 25653 23075 25687
rect 30006 25684 30012 25696
rect 29967 25656 30012 25684
rect 23017 25647 23075 25653
rect 30006 25644 30012 25656
rect 30064 25644 30070 25696
rect 1104 25594 30820 25616
rect 1104 25542 5915 25594
rect 5967 25542 5979 25594
rect 6031 25542 6043 25594
rect 6095 25542 6107 25594
rect 6159 25542 6171 25594
rect 6223 25542 15846 25594
rect 15898 25542 15910 25594
rect 15962 25542 15974 25594
rect 16026 25542 16038 25594
rect 16090 25542 16102 25594
rect 16154 25542 25776 25594
rect 25828 25542 25840 25594
rect 25892 25542 25904 25594
rect 25956 25542 25968 25594
rect 26020 25542 26032 25594
rect 26084 25542 30820 25594
rect 1104 25520 30820 25542
rect 9030 25440 9036 25492
rect 9088 25480 9094 25492
rect 9309 25483 9367 25489
rect 9309 25480 9321 25483
rect 9088 25452 9321 25480
rect 9088 25440 9094 25452
rect 9309 25449 9321 25452
rect 9355 25449 9367 25483
rect 9309 25443 9367 25449
rect 10781 25483 10839 25489
rect 10781 25449 10793 25483
rect 10827 25480 10839 25483
rect 13078 25480 13084 25492
rect 10827 25452 13084 25480
rect 10827 25449 10839 25452
rect 10781 25443 10839 25449
rect 13078 25440 13084 25452
rect 13136 25440 13142 25492
rect 13449 25483 13507 25489
rect 13449 25449 13461 25483
rect 13495 25480 13507 25483
rect 13722 25480 13728 25492
rect 13495 25452 13728 25480
rect 13495 25449 13507 25452
rect 13449 25443 13507 25449
rect 13722 25440 13728 25452
rect 13780 25440 13786 25492
rect 18693 25483 18751 25489
rect 18693 25449 18705 25483
rect 18739 25480 18751 25483
rect 19058 25480 19064 25492
rect 18739 25452 19064 25480
rect 18739 25449 18751 25452
rect 18693 25443 18751 25449
rect 19058 25440 19064 25452
rect 19116 25480 19122 25492
rect 19245 25483 19303 25489
rect 19245 25480 19257 25483
rect 19116 25452 19257 25480
rect 19116 25440 19122 25452
rect 19245 25449 19257 25452
rect 19291 25449 19303 25483
rect 19245 25443 19303 25449
rect 20441 25483 20499 25489
rect 20441 25449 20453 25483
rect 20487 25480 20499 25483
rect 20714 25480 20720 25492
rect 20487 25452 20720 25480
rect 20487 25449 20499 25452
rect 20441 25443 20499 25449
rect 20714 25440 20720 25452
rect 20772 25440 20778 25492
rect 23106 25480 23112 25492
rect 23067 25452 23112 25480
rect 23106 25440 23112 25452
rect 23164 25440 23170 25492
rect 5258 25372 5264 25424
rect 5316 25412 5322 25424
rect 13219 25415 13277 25421
rect 5316 25384 12434 25412
rect 5316 25372 5322 25384
rect 10686 25304 10692 25356
rect 10744 25344 10750 25356
rect 11333 25347 11391 25353
rect 11333 25344 11345 25347
rect 10744 25316 11345 25344
rect 10744 25304 10750 25316
rect 11333 25313 11345 25316
rect 11379 25344 11391 25347
rect 11379 25316 12204 25344
rect 11379 25313 11391 25316
rect 11333 25307 11391 25313
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 11146 25276 11152 25288
rect 11107 25248 11152 25276
rect 11146 25236 11152 25248
rect 11204 25236 11210 25288
rect 8846 25168 8852 25220
rect 8904 25208 8910 25220
rect 8941 25211 8999 25217
rect 8941 25208 8953 25211
rect 8904 25180 8953 25208
rect 8904 25168 8910 25180
rect 8941 25177 8953 25180
rect 8987 25177 8999 25211
rect 8941 25171 8999 25177
rect 9125 25211 9183 25217
rect 9125 25177 9137 25211
rect 9171 25208 9183 25211
rect 9306 25208 9312 25220
rect 9171 25180 9312 25208
rect 9171 25177 9183 25180
rect 9125 25171 9183 25177
rect 9306 25168 9312 25180
rect 9364 25168 9370 25220
rect 10042 25168 10048 25220
rect 10100 25208 10106 25220
rect 10137 25211 10195 25217
rect 10137 25208 10149 25211
rect 10100 25180 10149 25208
rect 10100 25168 10106 25180
rect 10137 25177 10149 25180
rect 10183 25177 10195 25211
rect 10137 25171 10195 25177
rect 10594 25168 10600 25220
rect 10652 25208 10658 25220
rect 11974 25208 11980 25220
rect 10652 25180 11980 25208
rect 10652 25168 10658 25180
rect 11974 25168 11980 25180
rect 12032 25168 12038 25220
rect 12176 25217 12204 25316
rect 12161 25211 12219 25217
rect 12161 25177 12173 25211
rect 12207 25177 12219 25211
rect 12406 25208 12434 25384
rect 13219 25381 13231 25415
rect 13265 25412 13277 25415
rect 13906 25412 13912 25424
rect 13265 25384 13912 25412
rect 13265 25381 13277 25384
rect 13219 25375 13277 25381
rect 13906 25372 13912 25384
rect 13964 25372 13970 25424
rect 16850 25372 16856 25424
rect 16908 25412 16914 25424
rect 18322 25412 18328 25424
rect 16908 25384 18328 25412
rect 16908 25372 16914 25384
rect 18322 25372 18328 25384
rect 18380 25372 18386 25424
rect 19150 25372 19156 25424
rect 19208 25412 19214 25424
rect 19208 25384 21404 25412
rect 19208 25372 19214 25384
rect 13357 25347 13415 25353
rect 13357 25313 13369 25347
rect 13403 25344 13415 25347
rect 13814 25344 13820 25356
rect 13403 25316 13820 25344
rect 13403 25313 13415 25316
rect 13357 25307 13415 25313
rect 13814 25304 13820 25316
rect 13872 25304 13878 25356
rect 16390 25344 16396 25356
rect 16351 25316 16396 25344
rect 16390 25304 16396 25316
rect 16448 25304 16454 25356
rect 16485 25347 16543 25353
rect 16485 25313 16497 25347
rect 16531 25344 16543 25347
rect 16666 25344 16672 25356
rect 16531 25316 16672 25344
rect 16531 25313 16543 25316
rect 16485 25307 16543 25313
rect 13078 25276 13084 25288
rect 13039 25248 13084 25276
rect 13078 25236 13084 25248
rect 13136 25236 13142 25288
rect 13541 25279 13599 25285
rect 13541 25245 13553 25279
rect 13587 25276 13599 25279
rect 13906 25276 13912 25288
rect 13587 25248 13912 25276
rect 13587 25245 13599 25248
rect 13541 25239 13599 25245
rect 13906 25236 13912 25248
rect 13964 25236 13970 25288
rect 14093 25279 14151 25285
rect 14093 25245 14105 25279
rect 14139 25276 14151 25279
rect 14182 25276 14188 25288
rect 14139 25248 14188 25276
rect 14139 25245 14151 25248
rect 14093 25239 14151 25245
rect 14182 25236 14188 25248
rect 14240 25236 14246 25288
rect 14734 25236 14740 25288
rect 14792 25276 14798 25288
rect 16500 25276 16528 25307
rect 16666 25304 16672 25316
rect 16724 25304 16730 25356
rect 17589 25347 17647 25353
rect 17589 25313 17601 25347
rect 17635 25344 17647 25347
rect 17770 25344 17776 25356
rect 17635 25316 17776 25344
rect 17635 25313 17647 25316
rect 17589 25307 17647 25313
rect 17770 25304 17776 25316
rect 17828 25304 17834 25356
rect 14792 25248 16528 25276
rect 17313 25279 17371 25285
rect 14792 25236 14798 25248
rect 17313 25245 17325 25279
rect 17359 25245 17371 25279
rect 17313 25239 17371 25245
rect 12406 25180 13952 25208
rect 12161 25171 12219 25177
rect 1578 25140 1584 25152
rect 1539 25112 1584 25140
rect 1578 25100 1584 25112
rect 1636 25100 1642 25152
rect 9950 25100 9956 25152
rect 10008 25140 10014 25152
rect 10229 25143 10287 25149
rect 10229 25140 10241 25143
rect 10008 25112 10241 25140
rect 10008 25100 10014 25112
rect 10229 25109 10241 25112
rect 10275 25109 10287 25143
rect 10229 25103 10287 25109
rect 10318 25100 10324 25152
rect 10376 25140 10382 25152
rect 11241 25143 11299 25149
rect 11241 25140 11253 25143
rect 10376 25112 11253 25140
rect 10376 25100 10382 25112
rect 11241 25109 11253 25112
rect 11287 25109 11299 25143
rect 11241 25103 11299 25109
rect 12345 25143 12403 25149
rect 12345 25109 12357 25143
rect 12391 25140 12403 25143
rect 13078 25140 13084 25152
rect 12391 25112 13084 25140
rect 12391 25109 12403 25112
rect 12345 25103 12403 25109
rect 13078 25100 13084 25112
rect 13136 25100 13142 25152
rect 13924 25140 13952 25180
rect 13998 25168 14004 25220
rect 14056 25208 14062 25220
rect 14338 25211 14396 25217
rect 14338 25208 14350 25211
rect 14056 25180 14350 25208
rect 14056 25168 14062 25180
rect 14338 25177 14350 25180
rect 14384 25177 14396 25211
rect 17129 25211 17187 25217
rect 17129 25208 17141 25211
rect 14338 25171 14396 25177
rect 14476 25180 17141 25208
rect 14476 25140 14504 25180
rect 17129 25177 17141 25180
rect 17175 25177 17187 25211
rect 17328 25208 17356 25239
rect 17402 25236 17408 25288
rect 17460 25276 17466 25288
rect 17681 25279 17739 25285
rect 17460 25248 17505 25276
rect 17460 25236 17466 25248
rect 17681 25245 17693 25279
rect 17727 25276 17739 25279
rect 17862 25276 17868 25288
rect 17727 25248 17868 25276
rect 17727 25245 17739 25248
rect 17681 25239 17739 25245
rect 17862 25236 17868 25248
rect 17920 25236 17926 25288
rect 18340 25285 18368 25372
rect 18874 25304 18880 25356
rect 18932 25344 18938 25356
rect 19337 25347 19395 25353
rect 19337 25344 19349 25347
rect 18932 25316 19349 25344
rect 18932 25304 18938 25316
rect 19337 25313 19349 25316
rect 19383 25313 19395 25347
rect 19337 25307 19395 25313
rect 18325 25279 18383 25285
rect 18325 25245 18337 25279
rect 18371 25245 18383 25279
rect 18325 25239 18383 25245
rect 18966 25236 18972 25288
rect 19024 25276 19030 25288
rect 19245 25279 19303 25285
rect 19245 25276 19257 25279
rect 19024 25248 19257 25276
rect 19024 25236 19030 25248
rect 19245 25245 19257 25248
rect 19291 25245 19303 25279
rect 19518 25276 19524 25288
rect 19479 25248 19524 25276
rect 19245 25239 19303 25245
rect 19518 25236 19524 25248
rect 19576 25236 19582 25288
rect 17586 25208 17592 25220
rect 17328 25180 17592 25208
rect 17129 25171 17187 25177
rect 17586 25168 17592 25180
rect 17644 25168 17650 25220
rect 18509 25211 18567 25217
rect 18509 25177 18521 25211
rect 18555 25177 18567 25211
rect 18509 25171 18567 25177
rect 15470 25140 15476 25152
rect 13924 25112 14504 25140
rect 15431 25112 15476 25140
rect 15470 25100 15476 25112
rect 15528 25100 15534 25152
rect 15746 25100 15752 25152
rect 15804 25140 15810 25152
rect 15933 25143 15991 25149
rect 15933 25140 15945 25143
rect 15804 25112 15945 25140
rect 15804 25100 15810 25112
rect 15933 25109 15945 25112
rect 15979 25109 15991 25143
rect 16298 25140 16304 25152
rect 16259 25112 16304 25140
rect 15933 25103 15991 25109
rect 16298 25100 16304 25112
rect 16356 25100 16362 25152
rect 16574 25100 16580 25152
rect 16632 25140 16638 25152
rect 18524 25140 18552 25171
rect 19426 25168 19432 25220
rect 19484 25208 19490 25220
rect 20070 25208 20076 25220
rect 19484 25180 20076 25208
rect 19484 25168 19490 25180
rect 20070 25168 20076 25180
rect 20128 25208 20134 25220
rect 21376 25217 21404 25384
rect 21450 25372 21456 25424
rect 21508 25412 21514 25424
rect 25130 25412 25136 25424
rect 21508 25384 25136 25412
rect 21508 25372 21514 25384
rect 25130 25372 25136 25384
rect 25188 25372 25194 25424
rect 27522 25372 27528 25424
rect 27580 25412 27586 25424
rect 29917 25415 29975 25421
rect 29917 25412 29929 25415
rect 27580 25384 29929 25412
rect 27580 25372 27586 25384
rect 29917 25381 29929 25384
rect 29963 25381 29975 25415
rect 29917 25375 29975 25381
rect 21542 25304 21548 25356
rect 21600 25304 21606 25356
rect 22097 25347 22155 25353
rect 22097 25313 22109 25347
rect 22143 25344 22155 25347
rect 23290 25344 23296 25356
rect 22143 25316 23296 25344
rect 22143 25313 22155 25316
rect 22097 25307 22155 25313
rect 23290 25304 23296 25316
rect 23348 25344 23354 25356
rect 23661 25347 23719 25353
rect 23661 25344 23673 25347
rect 23348 25316 23673 25344
rect 23348 25304 23354 25316
rect 23661 25313 23673 25316
rect 23707 25344 23719 25347
rect 24670 25344 24676 25356
rect 23707 25316 24676 25344
rect 23707 25313 23719 25316
rect 23661 25307 23719 25313
rect 24670 25304 24676 25316
rect 24728 25304 24734 25356
rect 21560 25276 21588 25304
rect 22005 25279 22063 25285
rect 22005 25276 22017 25279
rect 21468 25248 22017 25276
rect 20257 25211 20315 25217
rect 20257 25208 20269 25211
rect 20128 25180 20269 25208
rect 20128 25168 20134 25180
rect 20257 25177 20269 25180
rect 20303 25208 20315 25211
rect 21177 25211 21235 25217
rect 21177 25208 21189 25211
rect 20303 25180 21189 25208
rect 20303 25177 20315 25180
rect 20257 25171 20315 25177
rect 21177 25177 21189 25180
rect 21223 25177 21235 25211
rect 21177 25171 21235 25177
rect 21361 25211 21419 25217
rect 21361 25177 21373 25211
rect 21407 25177 21419 25211
rect 21361 25171 21419 25177
rect 19334 25140 19340 25152
rect 16632 25112 19340 25140
rect 16632 25100 16638 25112
rect 19334 25100 19340 25112
rect 19392 25100 19398 25152
rect 19702 25140 19708 25152
rect 19663 25112 19708 25140
rect 19702 25100 19708 25112
rect 19760 25100 19766 25152
rect 20346 25100 20352 25152
rect 20404 25140 20410 25152
rect 20441 25143 20499 25149
rect 20441 25140 20453 25143
rect 20404 25112 20453 25140
rect 20404 25100 20410 25112
rect 20441 25109 20453 25112
rect 20487 25109 20499 25143
rect 20441 25103 20499 25109
rect 20625 25143 20683 25149
rect 20625 25109 20637 25143
rect 20671 25140 20683 25143
rect 21468 25140 21496 25248
rect 22005 25245 22017 25248
rect 22051 25245 22063 25279
rect 23474 25276 23480 25288
rect 23435 25248 23480 25276
rect 22005 25239 22063 25245
rect 23474 25236 23480 25248
rect 23532 25236 23538 25288
rect 23750 25236 23756 25288
rect 23808 25276 23814 25288
rect 24397 25279 24455 25285
rect 24397 25276 24409 25279
rect 23808 25248 24409 25276
rect 23808 25236 23814 25248
rect 24397 25245 24409 25248
rect 24443 25245 24455 25279
rect 24397 25239 24455 25245
rect 24581 25279 24639 25285
rect 24581 25245 24593 25279
rect 24627 25276 24639 25279
rect 25314 25276 25320 25288
rect 24627 25248 25320 25276
rect 24627 25245 24639 25248
rect 24581 25239 24639 25245
rect 21545 25211 21603 25217
rect 21545 25177 21557 25211
rect 21591 25208 21603 25211
rect 21634 25208 21640 25220
rect 21591 25180 21640 25208
rect 21591 25177 21603 25180
rect 21545 25171 21603 25177
rect 21634 25168 21640 25180
rect 21692 25168 21698 25220
rect 23106 25168 23112 25220
rect 23164 25208 23170 25220
rect 24596 25208 24624 25239
rect 25314 25236 25320 25248
rect 25372 25236 25378 25288
rect 28902 25236 28908 25288
rect 28960 25276 28966 25288
rect 28997 25279 29055 25285
rect 28997 25276 29009 25279
rect 28960 25248 29009 25276
rect 28960 25236 28966 25248
rect 28997 25245 29009 25248
rect 29043 25245 29055 25279
rect 28997 25239 29055 25245
rect 30101 25279 30159 25285
rect 30101 25245 30113 25279
rect 30147 25245 30159 25279
rect 30101 25239 30159 25245
rect 23164 25180 24624 25208
rect 23164 25168 23170 25180
rect 25682 25168 25688 25220
rect 25740 25208 25746 25220
rect 26053 25211 26111 25217
rect 26053 25208 26065 25211
rect 25740 25180 26065 25208
rect 25740 25168 25746 25180
rect 26053 25177 26065 25180
rect 26099 25177 26111 25211
rect 26234 25208 26240 25220
rect 26195 25180 26240 25208
rect 26053 25171 26111 25177
rect 26234 25168 26240 25180
rect 26292 25168 26298 25220
rect 26786 25208 26792 25220
rect 26699 25180 26792 25208
rect 26786 25168 26792 25180
rect 26844 25208 26850 25220
rect 27614 25208 27620 25220
rect 26844 25180 27620 25208
rect 26844 25168 26850 25180
rect 27614 25168 27620 25180
rect 27672 25168 27678 25220
rect 28626 25168 28632 25220
rect 28684 25208 28690 25220
rect 30116 25208 30144 25239
rect 28684 25180 30144 25208
rect 28684 25168 28690 25180
rect 20671 25112 21496 25140
rect 20671 25109 20683 25112
rect 20625 25103 20683 25109
rect 23566 25100 23572 25152
rect 23624 25140 23630 25152
rect 24489 25143 24547 25149
rect 23624 25112 23669 25140
rect 23624 25100 23630 25112
rect 24489 25109 24501 25143
rect 24535 25140 24547 25143
rect 25958 25140 25964 25152
rect 24535 25112 25964 25140
rect 24535 25109 24547 25112
rect 24489 25103 24547 25109
rect 25958 25100 25964 25112
rect 26016 25100 26022 25152
rect 26878 25140 26884 25152
rect 26839 25112 26884 25140
rect 26878 25100 26884 25112
rect 26936 25100 26942 25152
rect 28810 25140 28816 25152
rect 28771 25112 28816 25140
rect 28810 25100 28816 25112
rect 28868 25100 28874 25152
rect 1104 25050 30820 25072
rect 1104 24998 10880 25050
rect 10932 24998 10944 25050
rect 10996 24998 11008 25050
rect 11060 24998 11072 25050
rect 11124 24998 11136 25050
rect 11188 24998 20811 25050
rect 20863 24998 20875 25050
rect 20927 24998 20939 25050
rect 20991 24998 21003 25050
rect 21055 24998 21067 25050
rect 21119 24998 30820 25050
rect 1104 24976 30820 24998
rect 1394 24896 1400 24948
rect 1452 24936 1458 24948
rect 1673 24939 1731 24945
rect 1673 24936 1685 24939
rect 1452 24908 1685 24936
rect 1452 24896 1458 24908
rect 1673 24905 1685 24908
rect 1719 24905 1731 24939
rect 9214 24936 9220 24948
rect 1673 24899 1731 24905
rect 8680 24908 9220 24936
rect 8680 24812 8708 24908
rect 9214 24896 9220 24908
rect 9272 24896 9278 24948
rect 11974 24896 11980 24948
rect 12032 24936 12038 24948
rect 12345 24939 12403 24945
rect 12345 24936 12357 24939
rect 12032 24908 12357 24936
rect 12032 24896 12038 24908
rect 12345 24905 12357 24908
rect 12391 24905 12403 24939
rect 12345 24899 12403 24905
rect 13262 24896 13268 24948
rect 13320 24936 13326 24948
rect 16850 24936 16856 24948
rect 13320 24908 16856 24936
rect 13320 24896 13326 24908
rect 16850 24896 16856 24908
rect 16908 24896 16914 24948
rect 18046 24896 18052 24948
rect 18104 24936 18110 24948
rect 18874 24936 18880 24948
rect 18104 24908 18880 24936
rect 18104 24896 18110 24908
rect 18874 24896 18880 24908
rect 18932 24896 18938 24948
rect 19426 24936 19432 24948
rect 18984 24908 19288 24936
rect 19387 24908 19432 24936
rect 8846 24828 8852 24880
rect 8904 24868 8910 24880
rect 8941 24871 8999 24877
rect 8941 24868 8953 24871
rect 8904 24840 8953 24868
rect 8904 24828 8910 24840
rect 8941 24837 8953 24840
rect 8987 24868 8999 24871
rect 9030 24868 9036 24880
rect 8987 24840 9036 24868
rect 8987 24837 8999 24840
rect 8941 24831 8999 24837
rect 9030 24828 9036 24840
rect 9088 24828 9094 24880
rect 9306 24828 9312 24880
rect 9364 24868 9370 24880
rect 9364 24840 9904 24868
rect 9364 24828 9370 24840
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24760 1642 24812
rect 1762 24760 1768 24812
rect 1820 24800 1826 24812
rect 2314 24800 2320 24812
rect 1820 24772 2320 24800
rect 1820 24760 1826 24772
rect 2314 24760 2320 24772
rect 2372 24760 2378 24812
rect 8297 24803 8355 24809
rect 8297 24769 8309 24803
rect 8343 24800 8355 24803
rect 8662 24800 8668 24812
rect 8343 24772 8668 24800
rect 8343 24769 8355 24772
rect 8297 24763 8355 24769
rect 8662 24760 8668 24772
rect 8720 24760 8726 24812
rect 9122 24800 9128 24812
rect 9083 24772 9128 24800
rect 9122 24760 9128 24772
rect 9180 24760 9186 24812
rect 9766 24800 9772 24812
rect 9727 24772 9772 24800
rect 9766 24760 9772 24772
rect 9824 24760 9830 24812
rect 9876 24800 9904 24840
rect 10042 24828 10048 24880
rect 10100 24868 10106 24880
rect 10781 24871 10839 24877
rect 10781 24868 10793 24871
rect 10100 24840 10793 24868
rect 10100 24828 10106 24840
rect 10781 24837 10793 24840
rect 10827 24837 10839 24871
rect 10781 24831 10839 24837
rect 9953 24803 10011 24809
rect 9953 24800 9965 24803
rect 9876 24772 9965 24800
rect 9953 24769 9965 24772
rect 9999 24800 10011 24803
rect 10410 24800 10416 24812
rect 9999 24772 10416 24800
rect 9999 24769 10011 24772
rect 9953 24763 10011 24769
rect 10410 24760 10416 24772
rect 10468 24760 10474 24812
rect 10594 24800 10600 24812
rect 10555 24772 10600 24800
rect 10594 24760 10600 24772
rect 10652 24760 10658 24812
rect 10796 24800 10824 24831
rect 11238 24828 11244 24880
rect 11296 24868 11302 24880
rect 11517 24871 11575 24877
rect 11517 24868 11529 24871
rect 11296 24840 11529 24868
rect 11296 24828 11302 24840
rect 11517 24837 11529 24840
rect 11563 24837 11575 24871
rect 11517 24831 11575 24837
rect 11882 24828 11888 24880
rect 11940 24868 11946 24880
rect 13722 24868 13728 24880
rect 11940 24840 13728 24868
rect 11940 24828 11946 24840
rect 13722 24828 13728 24840
rect 13780 24828 13786 24880
rect 14553 24871 14611 24877
rect 14553 24837 14565 24871
rect 14599 24868 14611 24871
rect 14918 24868 14924 24880
rect 14599 24840 14924 24868
rect 14599 24837 14611 24840
rect 14553 24831 14611 24837
rect 14918 24828 14924 24840
rect 14976 24828 14982 24880
rect 15028 24840 15332 24868
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 10796 24798 11468 24800
rect 11624 24798 11713 24800
rect 10796 24772 11713 24798
rect 11440 24770 11652 24772
rect 11701 24769 11713 24772
rect 11747 24769 11759 24803
rect 12529 24803 12587 24809
rect 12529 24800 12541 24803
rect 11701 24763 11759 24769
rect 12406 24772 12541 24800
rect 9309 24735 9367 24741
rect 9309 24701 9321 24735
rect 9355 24732 9367 24735
rect 12406 24732 12434 24772
rect 12529 24769 12541 24772
rect 12575 24769 12587 24803
rect 12529 24763 12587 24769
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 9355 24704 12434 24732
rect 9355 24701 9367 24704
rect 9309 24695 9367 24701
rect 8389 24667 8447 24673
rect 8389 24633 8401 24667
rect 8435 24664 8447 24667
rect 10042 24664 10048 24676
rect 8435 24636 10048 24664
rect 8435 24633 8447 24636
rect 8389 24627 8447 24633
rect 10042 24624 10048 24636
rect 10100 24624 10106 24676
rect 13004 24664 13032 24763
rect 13078 24760 13084 24812
rect 13136 24800 13142 24812
rect 13633 24803 13691 24809
rect 13633 24800 13645 24803
rect 13136 24772 13645 24800
rect 13136 24760 13142 24772
rect 13633 24769 13645 24772
rect 13679 24800 13691 24803
rect 14458 24800 14464 24812
rect 13679 24772 14320 24800
rect 14419 24772 14464 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 10888 24636 13032 24664
rect 13081 24667 13139 24673
rect 10134 24596 10140 24608
rect 10095 24568 10140 24596
rect 10134 24556 10140 24568
rect 10192 24556 10198 24608
rect 10778 24556 10784 24608
rect 10836 24596 10842 24608
rect 10888 24605 10916 24636
rect 13081 24633 13093 24667
rect 13127 24664 13139 24667
rect 13170 24664 13176 24676
rect 13127 24636 13176 24664
rect 13127 24633 13139 24636
rect 13081 24627 13139 24633
rect 13170 24624 13176 24636
rect 13228 24624 13234 24676
rect 10873 24599 10931 24605
rect 10873 24596 10885 24599
rect 10836 24568 10885 24596
rect 10836 24556 10842 24568
rect 10873 24565 10885 24568
rect 10919 24565 10931 24599
rect 11790 24596 11796 24608
rect 11751 24568 11796 24596
rect 10873 24559 10931 24565
rect 11790 24556 11796 24568
rect 11848 24556 11854 24608
rect 12158 24556 12164 24608
rect 12216 24596 12222 24608
rect 13446 24596 13452 24608
rect 12216 24568 13452 24596
rect 12216 24556 12222 24568
rect 13446 24556 13452 24568
rect 13504 24556 13510 24608
rect 14292 24596 14320 24772
rect 14458 24760 14464 24772
rect 14516 24760 14522 24812
rect 14645 24803 14703 24809
rect 14645 24769 14657 24803
rect 14691 24800 14703 24803
rect 15028 24800 15056 24840
rect 14691 24772 15056 24800
rect 15197 24803 15255 24809
rect 14691 24769 14703 24772
rect 14645 24763 14703 24769
rect 15197 24769 15209 24803
rect 15243 24769 15255 24803
rect 15304 24800 15332 24840
rect 17494 24828 17500 24880
rect 17552 24868 17558 24880
rect 18984 24868 19012 24908
rect 17552 24840 19012 24868
rect 19260 24868 19288 24908
rect 19426 24896 19432 24908
rect 19484 24896 19490 24948
rect 25222 24936 25228 24948
rect 22066 24908 25228 24936
rect 22066 24868 22094 24908
rect 25222 24896 25228 24908
rect 25280 24896 25286 24948
rect 19260 24840 22094 24868
rect 17552 24828 17558 24840
rect 25314 24828 25320 24880
rect 25372 24868 25378 24880
rect 25372 24840 25728 24868
rect 25372 24828 25378 24840
rect 15841 24803 15899 24809
rect 15304 24772 15424 24800
rect 15197 24763 15255 24769
rect 14826 24624 14832 24676
rect 14884 24664 14890 24676
rect 15212 24664 15240 24763
rect 15396 24673 15424 24772
rect 15841 24769 15853 24803
rect 15887 24800 15899 24803
rect 16761 24803 16819 24809
rect 16761 24800 16773 24803
rect 15887 24772 16773 24800
rect 15887 24769 15899 24772
rect 15841 24763 15899 24769
rect 16761 24769 16773 24772
rect 16807 24769 16819 24803
rect 18230 24800 18236 24812
rect 18191 24772 18236 24800
rect 16761 24763 16819 24769
rect 14884 24636 15240 24664
rect 15381 24667 15439 24673
rect 14884 24624 14890 24636
rect 15381 24633 15393 24667
rect 15427 24664 15439 24667
rect 15562 24664 15568 24676
rect 15427 24636 15568 24664
rect 15427 24633 15439 24636
rect 15381 24627 15439 24633
rect 15562 24624 15568 24636
rect 15620 24624 15626 24676
rect 15856 24596 15884 24763
rect 18230 24760 18236 24772
rect 18288 24760 18294 24812
rect 18966 24760 18972 24812
rect 19024 24800 19030 24812
rect 19061 24803 19119 24809
rect 19061 24800 19073 24803
rect 19024 24772 19073 24800
rect 19024 24760 19030 24772
rect 19061 24769 19073 24772
rect 19107 24769 19119 24803
rect 19061 24763 19119 24769
rect 19150 24760 19156 24812
rect 19208 24800 19214 24812
rect 19208 24772 19253 24800
rect 19208 24760 19214 24772
rect 19702 24760 19708 24812
rect 19760 24800 19766 24812
rect 20438 24800 20444 24812
rect 19760 24772 20444 24800
rect 19760 24760 19766 24772
rect 20438 24760 20444 24772
rect 20496 24760 20502 24812
rect 22646 24800 22652 24812
rect 22607 24772 22652 24800
rect 22646 24760 22652 24772
rect 22704 24760 22710 24812
rect 23658 24800 23664 24812
rect 23619 24772 23664 24800
rect 23658 24760 23664 24772
rect 23716 24760 23722 24812
rect 24670 24800 24676 24812
rect 24631 24772 24676 24800
rect 24670 24760 24676 24772
rect 24728 24760 24734 24812
rect 25700 24809 25728 24840
rect 25501 24803 25559 24809
rect 25501 24769 25513 24803
rect 25547 24769 25559 24803
rect 25501 24763 25559 24769
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24769 25743 24803
rect 28350 24800 28356 24812
rect 28311 24772 28356 24800
rect 25685 24763 25743 24769
rect 17037 24735 17095 24741
rect 17037 24701 17049 24735
rect 17083 24732 17095 24735
rect 17586 24732 17592 24744
rect 17083 24704 17592 24732
rect 17083 24701 17095 24704
rect 17037 24695 17095 24701
rect 17586 24692 17592 24704
rect 17644 24692 17650 24744
rect 18046 24692 18052 24744
rect 18104 24732 18110 24744
rect 18509 24735 18567 24741
rect 18509 24732 18521 24735
rect 18104 24704 18521 24732
rect 18104 24692 18110 24704
rect 18509 24701 18521 24704
rect 18555 24732 18567 24735
rect 19610 24732 19616 24744
rect 18555 24704 19616 24732
rect 18555 24701 18567 24704
rect 18509 24695 18567 24701
rect 19610 24692 19616 24704
rect 19668 24692 19674 24744
rect 20714 24732 20720 24744
rect 20675 24704 20720 24732
rect 20714 24692 20720 24704
rect 20772 24692 20778 24744
rect 22370 24692 22376 24744
rect 22428 24732 22434 24744
rect 22741 24735 22799 24741
rect 22741 24732 22753 24735
rect 22428 24704 22753 24732
rect 22428 24692 22434 24704
rect 22741 24701 22753 24704
rect 22787 24701 22799 24735
rect 22741 24695 22799 24701
rect 22925 24735 22983 24741
rect 22925 24701 22937 24735
rect 22971 24732 22983 24735
rect 23290 24732 23296 24744
rect 22971 24704 23296 24732
rect 22971 24701 22983 24704
rect 22925 24695 22983 24701
rect 23290 24692 23296 24704
rect 23348 24692 23354 24744
rect 23382 24692 23388 24744
rect 23440 24732 23446 24744
rect 24765 24735 24823 24741
rect 24765 24732 24777 24735
rect 23440 24704 24777 24732
rect 23440 24692 23446 24704
rect 24765 24701 24777 24704
rect 24811 24701 24823 24735
rect 24765 24695 24823 24701
rect 24854 24692 24860 24744
rect 24912 24732 24918 24744
rect 24912 24704 24957 24732
rect 24912 24692 24918 24704
rect 15930 24624 15936 24676
rect 15988 24664 15994 24676
rect 16025 24667 16083 24673
rect 16025 24664 16037 24667
rect 15988 24636 16037 24664
rect 15988 24624 15994 24636
rect 16025 24633 16037 24636
rect 16071 24633 16083 24667
rect 16025 24627 16083 24633
rect 14292 24568 15884 24596
rect 16040 24596 16068 24627
rect 16482 24624 16488 24676
rect 16540 24664 16546 24676
rect 19150 24664 19156 24676
rect 16540 24636 19156 24664
rect 16540 24624 16546 24636
rect 19150 24624 19156 24636
rect 19208 24624 19214 24676
rect 19426 24624 19432 24676
rect 19484 24664 19490 24676
rect 24210 24664 24216 24676
rect 19484 24636 24216 24664
rect 19484 24624 19490 24636
rect 24210 24624 24216 24636
rect 24268 24624 24274 24676
rect 24305 24667 24363 24673
rect 24305 24633 24317 24667
rect 24351 24664 24363 24667
rect 25516 24664 25544 24763
rect 28350 24760 28356 24772
rect 28408 24760 28414 24812
rect 28534 24760 28540 24812
rect 28592 24800 28598 24812
rect 28997 24803 29055 24809
rect 28997 24800 29009 24803
rect 28592 24772 29009 24800
rect 28592 24760 28598 24772
rect 28997 24769 29009 24772
rect 29043 24769 29055 24803
rect 28997 24763 29055 24769
rect 29825 24803 29883 24809
rect 29825 24769 29837 24803
rect 29871 24769 29883 24803
rect 29825 24763 29883 24769
rect 25593 24735 25651 24741
rect 25593 24701 25605 24735
rect 25639 24701 25651 24735
rect 25593 24695 25651 24701
rect 24351 24636 25544 24664
rect 25608 24664 25636 24695
rect 25958 24692 25964 24744
rect 26016 24732 26022 24744
rect 29840 24732 29868 24763
rect 26016 24704 29868 24732
rect 26016 24692 26022 24704
rect 29822 24664 29828 24676
rect 25608 24636 29828 24664
rect 24351 24633 24363 24636
rect 24305 24627 24363 24633
rect 29822 24624 29828 24636
rect 29880 24624 29886 24676
rect 30006 24664 30012 24676
rect 29967 24636 30012 24664
rect 30006 24624 30012 24636
rect 30064 24624 30070 24676
rect 17494 24596 17500 24608
rect 16040 24568 17500 24596
rect 17494 24556 17500 24568
rect 17552 24556 17558 24608
rect 19058 24596 19064 24608
rect 19019 24568 19064 24596
rect 19058 24556 19064 24568
rect 19116 24556 19122 24608
rect 22281 24599 22339 24605
rect 22281 24565 22293 24599
rect 22327 24596 22339 24599
rect 22922 24596 22928 24608
rect 22327 24568 22928 24596
rect 22327 24565 22339 24568
rect 22281 24559 22339 24565
rect 22922 24556 22928 24568
rect 22980 24556 22986 24608
rect 23474 24596 23480 24608
rect 23435 24568 23480 24596
rect 23474 24556 23480 24568
rect 23532 24556 23538 24608
rect 25038 24556 25044 24608
rect 25096 24596 25102 24608
rect 28169 24599 28227 24605
rect 28169 24596 28181 24599
rect 25096 24568 28181 24596
rect 25096 24556 25102 24568
rect 28169 24565 28181 24568
rect 28215 24565 28227 24599
rect 28169 24559 28227 24565
rect 28718 24556 28724 24608
rect 28776 24596 28782 24608
rect 28813 24599 28871 24605
rect 28813 24596 28825 24599
rect 28776 24568 28825 24596
rect 28776 24556 28782 24568
rect 28813 24565 28825 24568
rect 28859 24565 28871 24599
rect 28813 24559 28871 24565
rect 1104 24506 30820 24528
rect 1104 24454 5915 24506
rect 5967 24454 5979 24506
rect 6031 24454 6043 24506
rect 6095 24454 6107 24506
rect 6159 24454 6171 24506
rect 6223 24454 15846 24506
rect 15898 24454 15910 24506
rect 15962 24454 15974 24506
rect 16026 24454 16038 24506
rect 16090 24454 16102 24506
rect 16154 24454 25776 24506
rect 25828 24454 25840 24506
rect 25892 24454 25904 24506
rect 25956 24454 25968 24506
rect 26020 24454 26032 24506
rect 26084 24454 30820 24506
rect 1104 24432 30820 24454
rect 8294 24352 8300 24404
rect 8352 24392 8358 24404
rect 9122 24392 9128 24404
rect 8352 24364 9128 24392
rect 8352 24352 8358 24364
rect 9122 24352 9128 24364
rect 9180 24392 9186 24404
rect 9582 24392 9588 24404
rect 9180 24364 9588 24392
rect 9180 24352 9186 24364
rect 9582 24352 9588 24364
rect 9640 24392 9646 24404
rect 10505 24395 10563 24401
rect 10505 24392 10517 24395
rect 9640 24364 10517 24392
rect 9640 24352 9646 24364
rect 10505 24361 10517 24364
rect 10551 24361 10563 24395
rect 10505 24355 10563 24361
rect 11517 24395 11575 24401
rect 11517 24361 11529 24395
rect 11563 24392 11575 24395
rect 12158 24392 12164 24404
rect 11563 24364 12164 24392
rect 11563 24361 11575 24364
rect 11517 24355 11575 24361
rect 12158 24352 12164 24364
rect 12216 24352 12222 24404
rect 12345 24395 12403 24401
rect 12345 24361 12357 24395
rect 12391 24392 12403 24395
rect 13170 24392 13176 24404
rect 12391 24364 13176 24392
rect 12391 24361 12403 24364
rect 12345 24355 12403 24361
rect 13170 24352 13176 24364
rect 13228 24352 13234 24404
rect 15654 24352 15660 24404
rect 15712 24392 15718 24404
rect 16025 24395 16083 24401
rect 16025 24392 16037 24395
rect 15712 24364 16037 24392
rect 15712 24352 15718 24364
rect 16025 24361 16037 24364
rect 16071 24361 16083 24395
rect 16025 24355 16083 24361
rect 16298 24352 16304 24404
rect 16356 24392 16362 24404
rect 22278 24392 22284 24404
rect 16356 24364 22284 24392
rect 16356 24352 16362 24364
rect 22278 24352 22284 24364
rect 22336 24352 22342 24404
rect 22465 24395 22523 24401
rect 22465 24361 22477 24395
rect 22511 24392 22523 24395
rect 22646 24392 22652 24404
rect 22511 24364 22652 24392
rect 22511 24361 22523 24364
rect 22465 24355 22523 24361
rect 22646 24352 22652 24364
rect 22704 24352 22710 24404
rect 23109 24395 23167 24401
rect 23109 24361 23121 24395
rect 23155 24392 23167 24395
rect 23750 24392 23756 24404
rect 23155 24364 23756 24392
rect 23155 24361 23167 24364
rect 23109 24355 23167 24361
rect 23750 24352 23756 24364
rect 23808 24352 23814 24404
rect 24397 24395 24455 24401
rect 24397 24361 24409 24395
rect 24443 24392 24455 24395
rect 24670 24392 24676 24404
rect 24443 24364 24676 24392
rect 24443 24361 24455 24364
rect 24397 24355 24455 24361
rect 24670 24352 24676 24364
rect 24728 24352 24734 24404
rect 26234 24392 26240 24404
rect 25056 24364 26240 24392
rect 1578 24284 1584 24336
rect 1636 24324 1642 24336
rect 12529 24327 12587 24333
rect 1636 24296 11652 24324
rect 1636 24284 1642 24296
rect 11330 24256 11336 24268
rect 8956 24228 11336 24256
rect 8956 24200 8984 24228
rect 11330 24216 11336 24228
rect 11388 24216 11394 24268
rect 8938 24188 8944 24200
rect 8851 24160 8944 24188
rect 8938 24148 8944 24160
rect 8996 24148 9002 24200
rect 9030 24148 9036 24200
rect 9088 24188 9094 24200
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 9088 24160 9137 24188
rect 9088 24148 9094 24160
rect 9125 24157 9137 24160
rect 9171 24157 9183 24191
rect 9125 24151 9183 24157
rect 9214 24148 9220 24200
rect 9272 24188 9278 24200
rect 9355 24191 9413 24197
rect 9272 24160 9317 24188
rect 9272 24148 9278 24160
rect 9355 24157 9367 24191
rect 9401 24188 9413 24191
rect 9493 24191 9551 24197
rect 9401 24157 9435 24188
rect 9355 24151 9435 24157
rect 9493 24157 9505 24191
rect 9539 24157 9551 24191
rect 9493 24151 9551 24157
rect 8846 24080 8852 24132
rect 8904 24120 8910 24132
rect 9407 24120 9435 24151
rect 8904 24092 9435 24120
rect 9508 24120 9536 24151
rect 9766 24148 9772 24200
rect 9824 24188 9830 24200
rect 10505 24191 10563 24197
rect 10505 24188 10517 24191
rect 9824 24160 10517 24188
rect 9824 24148 9830 24160
rect 10505 24157 10517 24160
rect 10551 24157 10563 24191
rect 10686 24188 10692 24200
rect 10647 24160 10692 24188
rect 10505 24151 10563 24157
rect 10686 24148 10692 24160
rect 10744 24148 10750 24200
rect 11238 24148 11244 24200
rect 11296 24188 11302 24200
rect 11425 24191 11483 24197
rect 11425 24188 11437 24191
rect 11296 24160 11437 24188
rect 11296 24148 11302 24160
rect 11425 24157 11437 24160
rect 11471 24157 11483 24191
rect 11425 24151 11483 24157
rect 9858 24120 9864 24132
rect 9508 24092 9864 24120
rect 8904 24080 8910 24092
rect 9858 24080 9864 24092
rect 9916 24080 9922 24132
rect 11624 24120 11652 24296
rect 12529 24293 12541 24327
rect 12575 24293 12587 24327
rect 12529 24287 12587 24293
rect 11701 24259 11759 24265
rect 11701 24225 11713 24259
rect 11747 24256 11759 24259
rect 11882 24256 11888 24268
rect 11747 24228 11888 24256
rect 11747 24225 11759 24228
rect 11701 24219 11759 24225
rect 11882 24216 11888 24228
rect 11940 24216 11946 24268
rect 11974 24148 11980 24200
rect 12032 24188 12038 24200
rect 12161 24191 12219 24197
rect 12161 24188 12173 24191
rect 12032 24160 12173 24188
rect 12032 24148 12038 24160
rect 12161 24157 12173 24160
rect 12207 24157 12219 24191
rect 12161 24151 12219 24157
rect 12345 24191 12403 24197
rect 12345 24157 12357 24191
rect 12391 24188 12403 24191
rect 12434 24188 12440 24200
rect 12391 24160 12440 24188
rect 12391 24157 12403 24160
rect 12345 24151 12403 24157
rect 12434 24148 12440 24160
rect 12492 24148 12498 24200
rect 12544 24188 12572 24287
rect 17218 24284 17224 24336
rect 17276 24324 17282 24336
rect 17276 24296 17356 24324
rect 17276 24284 17282 24296
rect 13906 24216 13912 24268
rect 13964 24256 13970 24268
rect 14918 24256 14924 24268
rect 13964 24228 14924 24256
rect 13964 24216 13970 24228
rect 14918 24216 14924 24228
rect 14976 24256 14982 24268
rect 15105 24259 15163 24265
rect 15105 24256 15117 24259
rect 14976 24228 15117 24256
rect 14976 24216 14982 24228
rect 15105 24225 15117 24228
rect 15151 24225 15163 24259
rect 15105 24219 15163 24225
rect 12710 24188 12716 24200
rect 12544 24160 12716 24188
rect 12710 24148 12716 24160
rect 12768 24148 12774 24200
rect 12989 24191 13047 24197
rect 12989 24157 13001 24191
rect 13035 24188 13047 24191
rect 13078 24188 13084 24200
rect 13035 24160 13084 24188
rect 13035 24157 13047 24160
rect 12989 24151 13047 24157
rect 13078 24148 13084 24160
rect 13136 24148 13142 24200
rect 15013 24191 15071 24197
rect 15013 24157 15025 24191
rect 15059 24188 15071 24191
rect 15470 24188 15476 24200
rect 15059 24160 15476 24188
rect 15059 24157 15071 24160
rect 15013 24151 15071 24157
rect 15470 24148 15476 24160
rect 15528 24148 15534 24200
rect 16206 24188 16212 24200
rect 16167 24160 16212 24188
rect 16206 24148 16212 24160
rect 16264 24148 16270 24200
rect 17218 24188 17224 24200
rect 17179 24160 17224 24188
rect 17218 24148 17224 24160
rect 17276 24148 17282 24200
rect 17328 24197 17356 24296
rect 17402 24284 17408 24336
rect 17460 24324 17466 24336
rect 19613 24327 19671 24333
rect 19613 24324 19625 24327
rect 17460 24296 19625 24324
rect 17460 24284 17466 24296
rect 19613 24293 19625 24296
rect 19659 24293 19671 24327
rect 19613 24287 19671 24293
rect 19794 24284 19800 24336
rect 19852 24324 19858 24336
rect 25056 24324 25084 24364
rect 26234 24352 26240 24364
rect 26292 24392 26298 24404
rect 26602 24392 26608 24404
rect 26292 24364 26608 24392
rect 26292 24352 26298 24364
rect 26602 24352 26608 24364
rect 26660 24352 26666 24404
rect 19852 24296 25084 24324
rect 19852 24284 19858 24296
rect 17497 24259 17555 24265
rect 17497 24225 17509 24259
rect 17543 24256 17555 24259
rect 17543 24228 22094 24256
rect 17543 24225 17555 24228
rect 17497 24219 17555 24225
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24157 17371 24191
rect 17313 24151 17371 24157
rect 17589 24191 17647 24197
rect 17589 24157 17601 24191
rect 17635 24188 17647 24191
rect 17862 24188 17868 24200
rect 17635 24160 17868 24188
rect 17635 24157 17647 24160
rect 17589 24151 17647 24157
rect 17862 24148 17868 24160
rect 17920 24148 17926 24200
rect 19518 24188 19524 24200
rect 19479 24160 19524 24188
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 20438 24148 20444 24200
rect 20496 24188 20502 24200
rect 20809 24191 20867 24197
rect 20809 24188 20821 24191
rect 20496 24160 20821 24188
rect 20496 24148 20502 24160
rect 20809 24157 20821 24160
rect 20855 24157 20867 24191
rect 20809 24151 20867 24157
rect 20993 24191 21051 24197
rect 20993 24157 21005 24191
rect 21039 24188 21051 24191
rect 21266 24188 21272 24200
rect 21039 24160 21272 24188
rect 21039 24157 21051 24160
rect 20993 24151 21051 24157
rect 21266 24148 21272 24160
rect 21324 24188 21330 24200
rect 21818 24188 21824 24200
rect 21324 24160 21824 24188
rect 21324 24148 21330 24160
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 17037 24123 17095 24129
rect 17037 24120 17049 24123
rect 11624 24092 17049 24120
rect 17037 24089 17049 24092
rect 17083 24089 17095 24123
rect 17037 24083 17095 24089
rect 18230 24080 18236 24132
rect 18288 24120 18294 24132
rect 18325 24123 18383 24129
rect 18325 24120 18337 24123
rect 18288 24092 18337 24120
rect 18288 24080 18294 24092
rect 18325 24089 18337 24092
rect 18371 24120 18383 24123
rect 19886 24120 19892 24132
rect 18371 24092 19892 24120
rect 18371 24089 18383 24092
rect 18325 24083 18383 24089
rect 19886 24080 19892 24092
rect 19944 24120 19950 24132
rect 20070 24120 20076 24132
rect 19944 24092 20076 24120
rect 19944 24080 19950 24092
rect 20070 24080 20076 24092
rect 20128 24080 20134 24132
rect 21177 24123 21235 24129
rect 21177 24089 21189 24123
rect 21223 24089 21235 24123
rect 22066 24120 22094 24228
rect 22278 24216 22284 24268
rect 22336 24256 22342 24268
rect 23198 24256 23204 24268
rect 22336 24228 23204 24256
rect 22336 24216 22342 24228
rect 23198 24216 23204 24228
rect 23256 24216 23262 24268
rect 23290 24216 23296 24268
rect 23348 24256 23354 24268
rect 23661 24259 23719 24265
rect 23661 24256 23673 24259
rect 23348 24228 23673 24256
rect 23348 24216 23354 24228
rect 23661 24225 23673 24228
rect 23707 24225 23719 24259
rect 23661 24219 23719 24225
rect 22462 24148 22468 24200
rect 22520 24188 22526 24200
rect 22649 24191 22707 24197
rect 22649 24188 22661 24191
rect 22520 24160 22661 24188
rect 22520 24148 22526 24160
rect 22649 24157 22661 24160
rect 22695 24157 22707 24191
rect 23474 24188 23480 24200
rect 23435 24160 23480 24188
rect 22649 24151 22707 24157
rect 23474 24148 23480 24160
rect 23532 24148 23538 24200
rect 24578 24188 24584 24200
rect 24539 24160 24584 24188
rect 24578 24148 24584 24160
rect 24636 24148 24642 24200
rect 25056 24197 25084 24296
rect 25130 24284 25136 24336
rect 25188 24324 25194 24336
rect 28810 24324 28816 24336
rect 25188 24296 25452 24324
rect 25188 24284 25194 24296
rect 25314 24256 25320 24268
rect 25275 24228 25320 24256
rect 25314 24216 25320 24228
rect 25372 24216 25378 24268
rect 25424 24265 25452 24296
rect 26804 24296 28816 24324
rect 25409 24259 25467 24265
rect 25409 24225 25421 24259
rect 25455 24225 25467 24259
rect 25409 24219 25467 24225
rect 25041 24191 25099 24197
rect 25041 24157 25053 24191
rect 25087 24157 25099 24191
rect 25041 24151 25099 24157
rect 25130 24148 25136 24200
rect 25188 24188 25194 24200
rect 25225 24191 25283 24197
rect 25225 24188 25237 24191
rect 25188 24160 25237 24188
rect 25188 24148 25194 24160
rect 25225 24157 25237 24160
rect 25271 24157 25283 24191
rect 25225 24151 25283 24157
rect 25590 24148 25596 24200
rect 25648 24188 25654 24200
rect 26602 24188 26608 24200
rect 25648 24160 25693 24188
rect 26563 24160 26608 24188
rect 25648 24148 25654 24160
rect 26602 24148 26608 24160
rect 26660 24148 26666 24200
rect 26804 24197 26832 24296
rect 28810 24284 28816 24296
rect 28868 24284 28874 24336
rect 26973 24259 27031 24265
rect 26973 24225 26985 24259
rect 27019 24256 27031 24259
rect 28074 24256 28080 24268
rect 27019 24228 28080 24256
rect 27019 24225 27031 24228
rect 26973 24219 27031 24225
rect 28074 24216 28080 24228
rect 28132 24216 28138 24268
rect 26789 24191 26847 24197
rect 26789 24157 26801 24191
rect 26835 24157 26847 24191
rect 26789 24151 26847 24157
rect 26878 24148 26884 24200
rect 26936 24188 26942 24200
rect 27154 24188 27160 24200
rect 26936 24160 26981 24188
rect 27115 24160 27160 24188
rect 26936 24148 26942 24160
rect 27154 24148 27160 24160
rect 27212 24148 27218 24200
rect 27798 24188 27804 24200
rect 27759 24160 27804 24188
rect 27798 24148 27804 24160
rect 27856 24148 27862 24200
rect 28258 24148 28264 24200
rect 28316 24188 28322 24200
rect 28997 24191 29055 24197
rect 28997 24188 29009 24191
rect 28316 24160 29009 24188
rect 28316 24148 28322 24160
rect 28997 24157 29009 24160
rect 29043 24157 29055 24191
rect 29822 24188 29828 24200
rect 29783 24160 29828 24188
rect 28997 24151 29055 24157
rect 29822 24148 29828 24160
rect 29880 24148 29886 24200
rect 22066 24092 25912 24120
rect 21177 24083 21235 24089
rect 7558 24012 7564 24064
rect 7616 24052 7622 24064
rect 9677 24055 9735 24061
rect 9677 24052 9689 24055
rect 7616 24024 9689 24052
rect 7616 24012 7622 24024
rect 9677 24021 9689 24024
rect 9723 24021 9735 24055
rect 9677 24015 9735 24021
rect 10873 24055 10931 24061
rect 10873 24021 10885 24055
rect 10919 24052 10931 24055
rect 11330 24052 11336 24064
rect 10919 24024 11336 24052
rect 10919 24021 10931 24024
rect 10873 24015 10931 24021
rect 11330 24012 11336 24024
rect 11388 24012 11394 24064
rect 11698 24052 11704 24064
rect 11659 24024 11704 24052
rect 11698 24012 11704 24024
rect 11756 24012 11762 24064
rect 13173 24055 13231 24061
rect 13173 24021 13185 24055
rect 13219 24052 13231 24055
rect 15286 24052 15292 24064
rect 13219 24024 15292 24052
rect 13219 24021 13231 24024
rect 13173 24015 13231 24021
rect 15286 24012 15292 24024
rect 15344 24012 15350 24064
rect 16850 24012 16856 24064
rect 16908 24052 16914 24064
rect 18417 24055 18475 24061
rect 18417 24052 18429 24055
rect 16908 24024 18429 24052
rect 16908 24012 16914 24024
rect 18417 24021 18429 24024
rect 18463 24052 18475 24055
rect 19426 24052 19432 24064
rect 18463 24024 19432 24052
rect 18463 24021 18475 24024
rect 18417 24015 18475 24021
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 21192 24052 21220 24083
rect 22278 24052 22284 24064
rect 21192 24024 22284 24052
rect 22278 24012 22284 24024
rect 22336 24012 22342 24064
rect 23474 24012 23480 24064
rect 23532 24052 23538 24064
rect 23569 24055 23627 24061
rect 23569 24052 23581 24055
rect 23532 24024 23581 24052
rect 23532 24012 23538 24024
rect 23569 24021 23581 24024
rect 23615 24021 23627 24055
rect 25774 24052 25780 24064
rect 25735 24024 25780 24052
rect 23569 24015 23627 24021
rect 25774 24012 25780 24024
rect 25832 24012 25838 24064
rect 25884 24052 25912 24092
rect 27062 24052 27068 24064
rect 25884 24024 27068 24052
rect 27062 24012 27068 24024
rect 27120 24012 27126 24064
rect 27338 24052 27344 24064
rect 27299 24024 27344 24052
rect 27338 24012 27344 24024
rect 27396 24012 27402 24064
rect 27430 24012 27436 24064
rect 27488 24052 27494 24064
rect 27893 24055 27951 24061
rect 27893 24052 27905 24055
rect 27488 24024 27905 24052
rect 27488 24012 27494 24024
rect 27893 24021 27905 24024
rect 27939 24021 27951 24055
rect 27893 24015 27951 24021
rect 28166 24012 28172 24064
rect 28224 24052 28230 24064
rect 28813 24055 28871 24061
rect 28813 24052 28825 24055
rect 28224 24024 28825 24052
rect 28224 24012 28230 24024
rect 28813 24021 28825 24024
rect 28859 24021 28871 24055
rect 30006 24052 30012 24064
rect 29967 24024 30012 24052
rect 28813 24015 28871 24021
rect 30006 24012 30012 24024
rect 30064 24012 30070 24064
rect 1104 23962 30820 23984
rect 1104 23910 10880 23962
rect 10932 23910 10944 23962
rect 10996 23910 11008 23962
rect 11060 23910 11072 23962
rect 11124 23910 11136 23962
rect 11188 23910 20811 23962
rect 20863 23910 20875 23962
rect 20927 23910 20939 23962
rect 20991 23910 21003 23962
rect 21055 23910 21067 23962
rect 21119 23910 30820 23962
rect 1104 23888 30820 23910
rect 8665 23851 8723 23857
rect 8665 23817 8677 23851
rect 8711 23848 8723 23851
rect 9030 23848 9036 23860
rect 8711 23820 9036 23848
rect 8711 23817 8723 23820
rect 8665 23811 8723 23817
rect 9030 23808 9036 23820
rect 9088 23808 9094 23860
rect 12989 23851 13047 23857
rect 12989 23848 13001 23851
rect 9140 23820 13001 23848
rect 7300 23752 8524 23780
rect 7300 23656 7328 23752
rect 7558 23721 7564 23724
rect 7552 23712 7564 23721
rect 7519 23684 7564 23712
rect 7552 23675 7564 23684
rect 7558 23672 7564 23675
rect 7616 23672 7622 23724
rect 8496 23712 8524 23752
rect 8846 23740 8852 23792
rect 8904 23780 8910 23792
rect 9140 23780 9168 23820
rect 12989 23817 13001 23820
rect 13035 23817 13047 23851
rect 12989 23811 13047 23817
rect 14274 23808 14280 23860
rect 14332 23848 14338 23860
rect 14458 23848 14464 23860
rect 14332 23820 14464 23848
rect 14332 23808 14338 23820
rect 14458 23808 14464 23820
rect 14516 23808 14522 23860
rect 14918 23808 14924 23860
rect 14976 23848 14982 23860
rect 24305 23851 24363 23857
rect 14976 23820 20300 23848
rect 14976 23808 14982 23820
rect 11422 23780 11428 23792
rect 8904 23752 9168 23780
rect 9223 23752 11428 23780
rect 8904 23740 8910 23752
rect 9125 23715 9183 23721
rect 9125 23712 9137 23715
rect 8496 23684 9137 23712
rect 9125 23681 9137 23684
rect 9171 23712 9183 23715
rect 9223 23712 9251 23752
rect 11422 23740 11428 23752
rect 11480 23740 11486 23792
rect 11517 23783 11575 23789
rect 11517 23749 11529 23783
rect 11563 23780 11575 23783
rect 11698 23780 11704 23792
rect 11563 23752 11704 23780
rect 11563 23749 11575 23752
rect 11517 23743 11575 23749
rect 11698 23740 11704 23752
rect 11756 23780 11762 23792
rect 11756 23752 12940 23780
rect 11756 23740 11762 23752
rect 9171 23684 9251 23712
rect 9392 23715 9450 23721
rect 9171 23681 9183 23684
rect 9125 23675 9183 23681
rect 9392 23681 9404 23715
rect 9438 23712 9450 23715
rect 9674 23712 9680 23724
rect 9438 23684 9680 23712
rect 9438 23681 9450 23684
rect 9392 23675 9450 23681
rect 9674 23672 9680 23684
rect 9732 23672 9738 23724
rect 10594 23672 10600 23724
rect 10652 23712 10658 23724
rect 10962 23712 10968 23724
rect 10652 23684 10968 23712
rect 10652 23672 10658 23684
rect 10962 23672 10968 23684
rect 11020 23712 11026 23724
rect 12912 23721 12940 23752
rect 14734 23740 14740 23792
rect 14792 23780 14798 23792
rect 14792 23752 15148 23780
rect 14792 23740 14798 23752
rect 11977 23715 12035 23721
rect 11977 23712 11989 23715
rect 11020 23684 11989 23712
rect 11020 23672 11026 23684
rect 11977 23681 11989 23684
rect 12023 23681 12035 23715
rect 11977 23675 12035 23681
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23681 12679 23715
rect 12621 23675 12679 23681
rect 12897 23715 12955 23721
rect 12897 23681 12909 23715
rect 12943 23681 12955 23715
rect 12897 23675 12955 23681
rect 7282 23644 7288 23656
rect 7243 23616 7288 23644
rect 7282 23604 7288 23616
rect 7340 23604 7346 23656
rect 11885 23647 11943 23653
rect 11885 23613 11897 23647
rect 11931 23644 11943 23647
rect 12434 23644 12440 23656
rect 11931 23616 12440 23644
rect 11931 23613 11943 23616
rect 11885 23607 11943 23613
rect 12434 23604 12440 23616
rect 12492 23604 12498 23656
rect 10870 23536 10876 23588
rect 10928 23576 10934 23588
rect 12161 23579 12219 23585
rect 12161 23576 12173 23579
rect 10928 23548 12173 23576
rect 10928 23536 10934 23548
rect 12161 23545 12173 23548
rect 12207 23545 12219 23579
rect 12636 23576 12664 23675
rect 13354 23672 13360 23724
rect 13412 23712 13418 23724
rect 13633 23715 13691 23721
rect 13633 23712 13645 23715
rect 13412 23684 13645 23712
rect 13412 23672 13418 23684
rect 13633 23681 13645 23684
rect 13679 23712 13691 23715
rect 15010 23712 15016 23724
rect 13679 23684 15016 23712
rect 13679 23681 13691 23684
rect 13633 23675 13691 23681
rect 15010 23672 15016 23684
rect 15068 23672 15074 23724
rect 15120 23712 15148 23752
rect 15470 23740 15476 23792
rect 15528 23780 15534 23792
rect 16666 23780 16672 23792
rect 15528 23752 16672 23780
rect 15528 23740 15534 23752
rect 16666 23740 16672 23752
rect 16724 23780 16730 23792
rect 18141 23783 18199 23789
rect 16724 23752 17172 23780
rect 16724 23740 16730 23752
rect 17144 23721 17172 23752
rect 17236 23752 17816 23780
rect 17236 23721 17264 23752
rect 16117 23715 16175 23721
rect 15120 23684 15240 23712
rect 12986 23644 12992 23656
rect 12947 23616 12992 23644
rect 12986 23604 12992 23616
rect 13044 23604 13050 23656
rect 14458 23604 14464 23656
rect 14516 23644 14522 23656
rect 15102 23644 15108 23656
rect 14516 23616 15108 23644
rect 14516 23604 14522 23616
rect 15102 23604 15108 23616
rect 15160 23604 15166 23656
rect 15212 23653 15240 23684
rect 16117 23681 16129 23715
rect 16163 23681 16175 23715
rect 16117 23675 16175 23681
rect 17129 23715 17187 23721
rect 17129 23681 17141 23715
rect 17175 23681 17187 23715
rect 17129 23675 17187 23681
rect 17221 23715 17279 23721
rect 17221 23681 17233 23715
rect 17267 23681 17279 23715
rect 17494 23712 17500 23724
rect 17455 23684 17500 23712
rect 17221 23675 17279 23681
rect 15197 23647 15255 23653
rect 15197 23613 15209 23647
rect 15243 23613 15255 23647
rect 16132 23644 16160 23675
rect 17494 23672 17500 23684
rect 17552 23672 17558 23724
rect 17788 23644 17816 23752
rect 18141 23749 18153 23783
rect 18187 23780 18199 23783
rect 18322 23780 18328 23792
rect 18187 23752 18328 23780
rect 18187 23749 18199 23752
rect 18141 23743 18199 23749
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 17954 23712 17960 23724
rect 17867 23684 17960 23712
rect 17954 23672 17960 23684
rect 18012 23712 18018 23724
rect 18785 23715 18843 23721
rect 18064 23712 18276 23713
rect 18785 23712 18797 23715
rect 18012 23685 18797 23712
rect 18012 23684 18092 23685
rect 18248 23684 18797 23685
rect 18012 23672 18018 23684
rect 18785 23681 18797 23684
rect 18831 23681 18843 23715
rect 18785 23675 18843 23681
rect 18877 23715 18935 23721
rect 18877 23681 18889 23715
rect 18923 23712 18935 23715
rect 19058 23712 19064 23724
rect 18923 23684 19064 23712
rect 18923 23681 18935 23684
rect 18877 23675 18935 23681
rect 19058 23672 19064 23684
rect 19116 23672 19122 23724
rect 19334 23672 19340 23724
rect 19392 23712 19398 23724
rect 20272 23721 20300 23820
rect 24305 23817 24317 23851
rect 24351 23848 24363 23851
rect 24486 23848 24492 23860
rect 24351 23820 24492 23848
rect 24351 23817 24363 23820
rect 24305 23811 24363 23817
rect 24486 23808 24492 23820
rect 24544 23808 24550 23860
rect 26326 23848 26332 23860
rect 24872 23820 26332 23848
rect 22186 23740 22192 23792
rect 22244 23780 22250 23792
rect 22281 23783 22339 23789
rect 22281 23780 22293 23783
rect 22244 23752 22293 23780
rect 22244 23740 22250 23752
rect 22281 23749 22293 23752
rect 22327 23749 22339 23783
rect 22281 23743 22339 23749
rect 23017 23783 23075 23789
rect 23017 23749 23029 23783
rect 23063 23780 23075 23783
rect 24872 23780 24900 23820
rect 26326 23808 26332 23820
rect 26384 23808 26390 23860
rect 27706 23808 27712 23860
rect 27764 23848 27770 23860
rect 29273 23851 29331 23857
rect 29273 23848 29285 23851
rect 27764 23820 29285 23848
rect 27764 23808 27770 23820
rect 29273 23817 29285 23820
rect 29319 23817 29331 23851
rect 29273 23811 29331 23817
rect 28442 23780 28448 23792
rect 23063 23752 24900 23780
rect 24964 23752 28448 23780
rect 23063 23749 23075 23752
rect 23017 23743 23075 23749
rect 19889 23715 19947 23721
rect 19889 23712 19901 23715
rect 19392 23684 19901 23712
rect 19392 23672 19398 23684
rect 19889 23681 19901 23684
rect 19935 23712 19947 23715
rect 20165 23715 20223 23721
rect 20165 23712 20177 23715
rect 19935 23684 20177 23712
rect 19935 23681 19947 23684
rect 19889 23675 19947 23681
rect 20165 23681 20177 23684
rect 20211 23681 20223 23715
rect 20165 23675 20223 23681
rect 20257 23715 20315 23721
rect 20257 23681 20269 23715
rect 20303 23681 20315 23715
rect 22922 23712 22928 23724
rect 22883 23684 22928 23712
rect 20257 23675 20315 23681
rect 19797 23647 19855 23653
rect 16132 23616 17540 23644
rect 17788 23616 19748 23644
rect 15197 23607 15255 23613
rect 14826 23576 14832 23588
rect 12636 23548 14832 23576
rect 12161 23539 12219 23545
rect 14826 23536 14832 23548
rect 14884 23536 14890 23588
rect 17034 23536 17040 23588
rect 17092 23576 17098 23588
rect 17405 23579 17463 23585
rect 17405 23576 17417 23579
rect 17092 23548 17417 23576
rect 17092 23536 17098 23548
rect 17405 23545 17417 23548
rect 17451 23545 17463 23579
rect 17512 23576 17540 23616
rect 17512 23548 18184 23576
rect 17405 23539 17463 23545
rect 10410 23468 10416 23520
rect 10468 23508 10474 23520
rect 10505 23511 10563 23517
rect 10505 23508 10517 23511
rect 10468 23480 10517 23508
rect 10468 23468 10474 23480
rect 10505 23477 10517 23480
rect 10551 23477 10563 23511
rect 11974 23508 11980 23520
rect 11935 23480 11980 23508
rect 10505 23471 10563 23477
rect 11974 23468 11980 23480
rect 12032 23468 12038 23520
rect 12713 23511 12771 23517
rect 12713 23477 12725 23511
rect 12759 23508 12771 23511
rect 13078 23508 13084 23520
rect 12759 23480 13084 23508
rect 12759 23477 12771 23480
rect 12713 23471 12771 23477
rect 13078 23468 13084 23480
rect 13136 23468 13142 23520
rect 13538 23468 13544 23520
rect 13596 23508 13602 23520
rect 13633 23511 13691 23517
rect 13633 23508 13645 23511
rect 13596 23480 13645 23508
rect 13596 23468 13602 23480
rect 13633 23477 13645 23480
rect 13679 23477 13691 23511
rect 14642 23508 14648 23520
rect 14603 23480 14648 23508
rect 13633 23471 13691 23477
rect 14642 23468 14648 23480
rect 14700 23468 14706 23520
rect 15933 23511 15991 23517
rect 15933 23477 15945 23511
rect 15979 23508 15991 23511
rect 16298 23508 16304 23520
rect 15979 23480 16304 23508
rect 15979 23477 15991 23480
rect 15933 23471 15991 23477
rect 16298 23468 16304 23480
rect 16356 23468 16362 23520
rect 16942 23508 16948 23520
rect 16903 23480 16948 23508
rect 16942 23468 16948 23480
rect 17000 23468 17006 23520
rect 17218 23468 17224 23520
rect 17276 23508 17282 23520
rect 17586 23508 17592 23520
rect 17276 23480 17592 23508
rect 17276 23468 17282 23480
rect 17586 23468 17592 23480
rect 17644 23468 17650 23520
rect 18156 23508 18184 23548
rect 18325 23511 18383 23517
rect 18325 23508 18337 23511
rect 18156 23480 18337 23508
rect 18325 23477 18337 23480
rect 18371 23477 18383 23511
rect 18325 23471 18383 23477
rect 18785 23511 18843 23517
rect 18785 23477 18797 23511
rect 18831 23508 18843 23511
rect 19061 23511 19119 23517
rect 19061 23508 19073 23511
rect 18831 23480 19073 23508
rect 18831 23477 18843 23480
rect 18785 23471 18843 23477
rect 19061 23477 19073 23480
rect 19107 23477 19119 23511
rect 19610 23508 19616 23520
rect 19571 23480 19616 23508
rect 19061 23471 19119 23477
rect 19610 23468 19616 23480
rect 19668 23468 19674 23520
rect 19720 23508 19748 23616
rect 19797 23613 19809 23647
rect 19843 23644 19855 23647
rect 20180 23644 20208 23675
rect 22922 23672 22928 23684
rect 22980 23672 22986 23724
rect 23106 23712 23112 23724
rect 23067 23684 23112 23712
rect 23106 23672 23112 23684
rect 23164 23672 23170 23724
rect 24489 23715 24547 23721
rect 24489 23681 24501 23715
rect 24535 23712 24547 23715
rect 24854 23712 24860 23724
rect 24535 23684 24860 23712
rect 24535 23681 24547 23684
rect 24489 23675 24547 23681
rect 24854 23672 24860 23684
rect 24912 23672 24918 23724
rect 24964 23721 24992 23752
rect 24949 23715 25007 23721
rect 24949 23681 24961 23715
rect 24995 23681 25007 23715
rect 24949 23675 25007 23681
rect 25216 23715 25274 23721
rect 25216 23681 25228 23715
rect 25262 23712 25274 23715
rect 25774 23712 25780 23724
rect 25262 23684 25780 23712
rect 25262 23681 25274 23684
rect 25216 23675 25274 23681
rect 25774 23672 25780 23684
rect 25832 23672 25838 23724
rect 27448 23721 27476 23752
rect 28442 23740 28448 23752
rect 28500 23740 28506 23792
rect 27433 23715 27491 23721
rect 27433 23681 27445 23715
rect 27479 23681 27491 23715
rect 27433 23675 27491 23681
rect 27700 23715 27758 23721
rect 27700 23681 27712 23715
rect 27746 23712 27758 23715
rect 27982 23712 27988 23724
rect 27746 23684 27988 23712
rect 27746 23681 27758 23684
rect 27700 23675 27758 23681
rect 27982 23672 27988 23684
rect 28040 23672 28046 23724
rect 28810 23672 28816 23724
rect 28868 23712 28874 23724
rect 29457 23715 29515 23721
rect 29457 23712 29469 23715
rect 28868 23684 29469 23712
rect 28868 23672 28874 23684
rect 29457 23681 29469 23684
rect 29503 23681 29515 23715
rect 30098 23712 30104 23724
rect 30059 23684 30104 23712
rect 29457 23675 29515 23681
rect 30098 23672 30104 23684
rect 30156 23672 30162 23724
rect 20438 23644 20444 23656
rect 19843 23616 19932 23644
rect 20180 23616 20444 23644
rect 19843 23613 19855 23616
rect 19797 23607 19855 23613
rect 19904 23588 19932 23616
rect 20438 23604 20444 23616
rect 20496 23604 20502 23656
rect 22465 23647 22523 23653
rect 22465 23613 22477 23647
rect 22511 23644 22523 23647
rect 22830 23644 22836 23656
rect 22511 23616 22836 23644
rect 22511 23613 22523 23616
rect 22465 23607 22523 23613
rect 22830 23604 22836 23616
rect 22888 23604 22894 23656
rect 19886 23536 19892 23588
rect 19944 23536 19950 23588
rect 22848 23548 23060 23576
rect 22848 23508 22876 23548
rect 19720 23480 22876 23508
rect 23032 23508 23060 23548
rect 25314 23508 25320 23520
rect 23032 23480 25320 23508
rect 25314 23468 25320 23480
rect 25372 23468 25378 23520
rect 25590 23468 25596 23520
rect 25648 23508 25654 23520
rect 26329 23511 26387 23517
rect 26329 23508 26341 23511
rect 25648 23480 26341 23508
rect 25648 23468 25654 23480
rect 26329 23477 26341 23480
rect 26375 23477 26387 23511
rect 26329 23471 26387 23477
rect 27798 23468 27804 23520
rect 27856 23508 27862 23520
rect 28813 23511 28871 23517
rect 28813 23508 28825 23511
rect 27856 23480 28825 23508
rect 27856 23468 27862 23480
rect 28813 23477 28825 23480
rect 28859 23477 28871 23511
rect 28813 23471 28871 23477
rect 29822 23468 29828 23520
rect 29880 23508 29886 23520
rect 29917 23511 29975 23517
rect 29917 23508 29929 23511
rect 29880 23480 29929 23508
rect 29880 23468 29886 23480
rect 29917 23477 29929 23480
rect 29963 23477 29975 23511
rect 29917 23471 29975 23477
rect 1104 23418 30820 23440
rect 1104 23366 5915 23418
rect 5967 23366 5979 23418
rect 6031 23366 6043 23418
rect 6095 23366 6107 23418
rect 6159 23366 6171 23418
rect 6223 23366 15846 23418
rect 15898 23366 15910 23418
rect 15962 23366 15974 23418
rect 16026 23366 16038 23418
rect 16090 23366 16102 23418
rect 16154 23366 25776 23418
rect 25828 23366 25840 23418
rect 25892 23366 25904 23418
rect 25956 23366 25968 23418
rect 26020 23366 26032 23418
rect 26084 23366 30820 23418
rect 1104 23344 30820 23366
rect 8294 23304 8300 23316
rect 8255 23276 8300 23304
rect 8294 23264 8300 23276
rect 8352 23264 8358 23316
rect 9674 23304 9680 23316
rect 9635 23276 9680 23304
rect 9674 23264 9680 23276
rect 9732 23264 9738 23316
rect 11882 23304 11888 23316
rect 11843 23276 11888 23304
rect 11882 23264 11888 23276
rect 11940 23264 11946 23316
rect 12345 23307 12403 23313
rect 12345 23273 12357 23307
rect 12391 23304 12403 23307
rect 12618 23304 12624 23316
rect 12391 23276 12624 23304
rect 12391 23273 12403 23276
rect 12345 23267 12403 23273
rect 12618 23264 12624 23276
rect 12676 23304 12682 23316
rect 12986 23304 12992 23316
rect 12676 23276 12992 23304
rect 12676 23264 12682 23276
rect 12986 23264 12992 23276
rect 13044 23264 13050 23316
rect 16942 23304 16948 23316
rect 13280 23276 16948 23304
rect 13280 23236 13308 23276
rect 16942 23264 16948 23276
rect 17000 23264 17006 23316
rect 17034 23264 17040 23316
rect 17092 23304 17098 23316
rect 18322 23304 18328 23316
rect 17092 23276 18328 23304
rect 17092 23264 17098 23276
rect 18322 23264 18328 23276
rect 18380 23264 18386 23316
rect 18874 23264 18880 23316
rect 18932 23304 18938 23316
rect 18932 23276 19564 23304
rect 18932 23264 18938 23276
rect 2148 23208 13308 23236
rect 2148 23109 2176 23208
rect 14090 23196 14096 23248
rect 14148 23236 14154 23248
rect 14148 23208 14228 23236
rect 14148 23196 14154 23208
rect 8294 23128 8300 23180
rect 8352 23168 8358 23180
rect 9214 23168 9220 23180
rect 8352 23140 9220 23168
rect 8352 23128 8358 23140
rect 9214 23128 9220 23140
rect 9272 23128 9278 23180
rect 9309 23171 9367 23177
rect 9309 23137 9321 23171
rect 9355 23168 9367 23171
rect 9355 23140 10088 23168
rect 9355 23137 9367 23140
rect 9309 23131 9367 23137
rect 1397 23103 1455 23109
rect 1397 23069 1409 23103
rect 1443 23069 1455 23103
rect 1397 23063 1455 23069
rect 2133 23103 2191 23109
rect 2133 23069 2145 23103
rect 2179 23069 2191 23103
rect 2314 23100 2320 23112
rect 2275 23072 2320 23100
rect 2133 23063 2191 23069
rect 1412 23032 1440 23063
rect 2314 23060 2320 23072
rect 2372 23060 2378 23112
rect 8205 23103 8263 23109
rect 8205 23069 8217 23103
rect 8251 23069 8263 23103
rect 8938 23100 8944 23112
rect 8899 23072 8944 23100
rect 8205 23063 8263 23069
rect 2225 23035 2283 23041
rect 2225 23032 2237 23035
rect 1412 23004 2237 23032
rect 2225 23001 2237 23004
rect 2271 23001 2283 23035
rect 8220 23032 8248 23063
rect 8938 23060 8944 23072
rect 8996 23060 9002 23112
rect 9125 23103 9183 23109
rect 9125 23069 9137 23103
rect 9171 23100 9183 23103
rect 9398 23100 9404 23112
rect 9171 23072 9404 23100
rect 9171 23069 9183 23072
rect 9125 23063 9183 23069
rect 9140 23032 9168 23063
rect 9398 23060 9404 23072
rect 9456 23060 9462 23112
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23100 9551 23103
rect 9858 23100 9864 23112
rect 9539 23072 9864 23100
rect 9539 23069 9551 23072
rect 9493 23063 9551 23069
rect 9858 23060 9864 23072
rect 9916 23060 9922 23112
rect 10060 23100 10088 23140
rect 10134 23128 10140 23180
rect 10192 23168 10198 23180
rect 10321 23171 10379 23177
rect 10321 23168 10333 23171
rect 10192 23140 10333 23168
rect 10192 23128 10198 23140
rect 10321 23137 10333 23140
rect 10367 23137 10379 23171
rect 10321 23131 10379 23137
rect 10410 23128 10416 23180
rect 10468 23168 10474 23180
rect 10594 23168 10600 23180
rect 10468 23140 10600 23168
rect 10468 23128 10474 23140
rect 10594 23128 10600 23140
rect 10652 23128 10658 23180
rect 10962 23128 10968 23180
rect 11020 23168 11026 23180
rect 12069 23171 12127 23177
rect 11020 23140 11836 23168
rect 11020 23128 11026 23140
rect 10870 23100 10876 23112
rect 10060 23072 10876 23100
rect 10870 23060 10876 23072
rect 10928 23060 10934 23112
rect 11330 23060 11336 23112
rect 11388 23100 11394 23112
rect 11701 23103 11759 23109
rect 11701 23100 11713 23103
rect 11388 23072 11713 23100
rect 11388 23060 11394 23072
rect 11701 23069 11713 23072
rect 11747 23069 11759 23103
rect 11808 23100 11836 23140
rect 12069 23137 12081 23171
rect 12115 23168 12127 23171
rect 12710 23168 12716 23180
rect 12115 23140 12716 23168
rect 12115 23137 12127 23140
rect 12069 23131 12127 23137
rect 12710 23128 12716 23140
rect 12768 23128 12774 23180
rect 13357 23171 13415 23177
rect 13004 23140 13308 23168
rect 12161 23103 12219 23109
rect 12161 23100 12173 23103
rect 11808 23072 12173 23100
rect 11701 23063 11759 23069
rect 12161 23069 12173 23072
rect 12207 23069 12219 23103
rect 12161 23063 12219 23069
rect 12434 23060 12440 23112
rect 12492 23100 12498 23112
rect 12894 23100 12900 23112
rect 12492 23072 12900 23100
rect 12492 23060 12498 23072
rect 12894 23060 12900 23072
rect 12952 23100 12958 23112
rect 13004 23100 13032 23140
rect 12952 23072 13032 23100
rect 13081 23103 13139 23109
rect 12952 23060 12958 23072
rect 13081 23069 13093 23103
rect 13127 23100 13139 23103
rect 13170 23100 13176 23112
rect 13127 23072 13176 23100
rect 13127 23069 13139 23072
rect 13081 23063 13139 23069
rect 13170 23060 13176 23072
rect 13228 23060 13234 23112
rect 13280 23100 13308 23140
rect 13357 23137 13369 23171
rect 13403 23168 13415 23171
rect 13403 23140 14136 23168
rect 13403 23137 13415 23140
rect 13357 23131 13415 23137
rect 14108 23109 14136 23140
rect 13454 23103 13512 23109
rect 13454 23100 13466 23103
rect 13280 23072 13466 23100
rect 13454 23069 13466 23072
rect 13500 23069 13512 23103
rect 13454 23063 13512 23069
rect 14093 23103 14151 23109
rect 14093 23069 14105 23103
rect 14139 23069 14151 23103
rect 14200 23100 14228 23208
rect 14642 23196 14648 23248
rect 14700 23196 14706 23248
rect 15930 23236 15936 23248
rect 15891 23208 15936 23236
rect 15930 23196 15936 23208
rect 15988 23196 15994 23248
rect 19337 23239 19395 23245
rect 19337 23205 19349 23239
rect 19383 23205 19395 23239
rect 19536 23236 19564 23276
rect 19610 23264 19616 23316
rect 19668 23304 19674 23316
rect 20349 23307 20407 23313
rect 20349 23304 20361 23307
rect 19668 23276 20361 23304
rect 19668 23264 19674 23276
rect 20349 23273 20361 23276
rect 20395 23273 20407 23307
rect 21910 23304 21916 23316
rect 20349 23267 20407 23273
rect 21468 23276 21916 23304
rect 21468 23236 21496 23276
rect 21910 23264 21916 23276
rect 21968 23264 21974 23316
rect 22005 23307 22063 23313
rect 22005 23273 22017 23307
rect 22051 23304 22063 23307
rect 23382 23304 23388 23316
rect 22051 23276 23388 23304
rect 22051 23273 22063 23276
rect 22005 23267 22063 23273
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 23750 23264 23756 23316
rect 23808 23304 23814 23316
rect 24489 23307 24547 23313
rect 24489 23304 24501 23307
rect 23808 23276 24501 23304
rect 23808 23264 23814 23276
rect 24489 23273 24501 23276
rect 24535 23273 24547 23307
rect 24854 23304 24860 23316
rect 24815 23276 24860 23304
rect 24489 23267 24547 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 25317 23307 25375 23313
rect 25317 23273 25329 23307
rect 25363 23304 25375 23307
rect 25406 23304 25412 23316
rect 25363 23276 25412 23304
rect 25363 23273 25375 23276
rect 25317 23267 25375 23273
rect 25406 23264 25412 23276
rect 25464 23264 25470 23316
rect 22830 23236 22836 23248
rect 19536 23208 21496 23236
rect 21560 23208 22836 23236
rect 19337 23199 19395 23205
rect 14360 23168 14366 23180
rect 14273 23140 14366 23168
rect 14360 23128 14366 23140
rect 14418 23168 14424 23180
rect 14418 23140 14587 23168
rect 14418 23128 14424 23140
rect 14277 23103 14335 23109
rect 14277 23100 14289 23103
rect 14200 23072 14289 23100
rect 14093 23063 14151 23069
rect 14277 23069 14289 23072
rect 14323 23069 14335 23103
rect 14277 23063 14335 23069
rect 14461 23103 14519 23109
rect 14461 23069 14473 23103
rect 14507 23069 14519 23103
rect 14461 23063 14519 23069
rect 8220 23004 9168 23032
rect 2225 22995 2283 23001
rect 10318 22992 10324 23044
rect 10376 23032 10382 23044
rect 12066 23032 12072 23044
rect 10376 23004 12072 23032
rect 10376 22992 10382 23004
rect 12066 22992 12072 23004
rect 12124 22992 12130 23044
rect 13262 23032 13268 23044
rect 13223 23004 13268 23032
rect 13262 22992 13268 23004
rect 13320 22992 13326 23044
rect 13357 23035 13415 23041
rect 13357 23001 13369 23035
rect 13403 23032 13415 23035
rect 13538 23032 13544 23044
rect 13403 23004 13544 23032
rect 13403 23001 13415 23004
rect 13357 22995 13415 23001
rect 13538 22992 13544 23004
rect 13596 22992 13602 23044
rect 14366 22992 14372 23044
rect 14424 23032 14430 23044
rect 14476 23032 14504 23063
rect 14424 23004 14504 23032
rect 14559 23032 14587 23140
rect 14660 23109 14688 23196
rect 16206 23168 16212 23180
rect 16040 23140 16212 23168
rect 14645 23103 14703 23109
rect 14645 23069 14657 23103
rect 14691 23069 14703 23103
rect 14645 23063 14703 23069
rect 15194 23060 15200 23112
rect 15252 23100 15258 23112
rect 16040 23100 16068 23140
rect 16206 23128 16212 23140
rect 16264 23168 16270 23180
rect 16485 23171 16543 23177
rect 16485 23168 16497 23171
rect 16264 23140 16497 23168
rect 16264 23128 16270 23140
rect 16485 23137 16497 23140
rect 16531 23137 16543 23171
rect 17310 23168 17316 23180
rect 17271 23140 17316 23168
rect 16485 23131 16543 23137
rect 17310 23128 17316 23140
rect 17368 23128 17374 23180
rect 19352 23168 19380 23199
rect 20714 23168 20720 23180
rect 19352 23140 20116 23168
rect 16298 23100 16304 23112
rect 15252 23072 16068 23100
rect 16259 23072 16304 23100
rect 15252 23060 15258 23072
rect 16298 23060 16304 23072
rect 16356 23060 16362 23112
rect 17328 23100 17356 23128
rect 18322 23100 18328 23112
rect 17328 23072 18328 23100
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 19245 23103 19303 23109
rect 19245 23069 19257 23103
rect 19291 23100 19303 23103
rect 19334 23100 19340 23112
rect 19291 23072 19340 23100
rect 19291 23069 19303 23072
rect 19245 23063 19303 23069
rect 19334 23060 19340 23072
rect 19392 23060 19398 23112
rect 20088 23109 20116 23140
rect 20180 23140 20720 23168
rect 20180 23109 20208 23140
rect 20714 23128 20720 23140
rect 20772 23128 20778 23180
rect 21560 23177 21588 23208
rect 22830 23196 22836 23208
rect 22888 23196 22894 23248
rect 25590 23236 25596 23248
rect 23676 23208 25596 23236
rect 21545 23171 21603 23177
rect 21545 23137 21557 23171
rect 21591 23137 21603 23171
rect 21545 23131 21603 23137
rect 21634 23128 21640 23180
rect 21692 23168 21698 23180
rect 21692 23140 21737 23168
rect 21692 23128 21698 23140
rect 20073 23103 20131 23109
rect 20073 23069 20085 23103
rect 20119 23069 20131 23103
rect 20073 23063 20131 23069
rect 20165 23103 20223 23109
rect 20165 23069 20177 23103
rect 20211 23069 20223 23103
rect 20165 23063 20223 23069
rect 20346 23060 20352 23112
rect 20404 23100 20410 23112
rect 20441 23103 20499 23109
rect 20441 23100 20453 23103
rect 20404 23072 20453 23100
rect 20404 23060 20410 23072
rect 20441 23069 20453 23072
rect 20487 23069 20499 23103
rect 20441 23063 20499 23069
rect 21269 23103 21327 23109
rect 21269 23069 21281 23103
rect 21315 23069 21327 23103
rect 21269 23063 21327 23069
rect 21453 23103 21511 23109
rect 21453 23069 21465 23103
rect 21499 23100 21511 23103
rect 21726 23100 21732 23112
rect 21499 23072 21732 23100
rect 21499 23069 21511 23072
rect 21453 23063 21511 23069
rect 14918 23032 14924 23044
rect 14559 23004 14924 23032
rect 14424 22992 14430 23004
rect 14918 22992 14924 23004
rect 14976 22992 14982 23044
rect 15010 22992 15016 23044
rect 15068 23032 15074 23044
rect 16393 23035 16451 23041
rect 15068 23004 16344 23032
rect 15068 22992 15074 23004
rect 1578 22964 1584 22976
rect 1539 22936 1584 22964
rect 1578 22924 1584 22936
rect 1636 22924 1642 22976
rect 14829 22967 14887 22973
rect 14829 22933 14841 22967
rect 14875 22964 14887 22967
rect 15194 22964 15200 22976
rect 14875 22936 15200 22964
rect 14875 22933 14887 22936
rect 14829 22927 14887 22933
rect 15194 22924 15200 22936
rect 15252 22924 15258 22976
rect 16316 22964 16344 23004
rect 16393 23001 16405 23035
rect 16439 23032 16451 23035
rect 17402 23032 17408 23044
rect 16439 23004 17408 23032
rect 16439 23001 16451 23004
rect 16393 22995 16451 23001
rect 17402 22992 17408 23004
rect 17460 22992 17466 23044
rect 17580 23035 17638 23041
rect 17580 23001 17592 23035
rect 17626 23032 17638 23035
rect 18598 23032 18604 23044
rect 17626 23004 18604 23032
rect 17626 23001 17638 23004
rect 17580 22995 17638 23001
rect 18598 22992 18604 23004
rect 18656 22992 18662 23044
rect 19889 23035 19947 23041
rect 19889 23001 19901 23035
rect 19935 23032 19947 23035
rect 21284 23032 21312 23063
rect 21726 23060 21732 23072
rect 21784 23060 21790 23112
rect 21821 23103 21879 23109
rect 21821 23069 21833 23103
rect 21867 23100 21879 23103
rect 22462 23100 22468 23112
rect 21867 23072 22094 23100
rect 22423 23072 22468 23100
rect 21867 23069 21879 23072
rect 21821 23063 21879 23069
rect 19935 23004 21312 23032
rect 22066 23032 22094 23072
rect 22462 23060 22468 23072
rect 22520 23060 22526 23112
rect 23676 23109 23704 23208
rect 25590 23196 25596 23208
rect 25648 23196 25654 23248
rect 27154 23196 27160 23248
rect 27212 23236 27218 23248
rect 27525 23239 27583 23245
rect 27525 23236 27537 23239
rect 27212 23208 27537 23236
rect 27212 23196 27218 23208
rect 27525 23205 27537 23208
rect 27571 23236 27583 23239
rect 27571 23208 29592 23236
rect 27571 23205 27583 23208
rect 27525 23199 27583 23205
rect 24486 23128 24492 23180
rect 24544 23168 24550 23180
rect 26145 23171 26203 23177
rect 26145 23168 26157 23171
rect 24544 23140 26157 23168
rect 24544 23128 24550 23140
rect 26145 23137 26157 23140
rect 26191 23137 26203 23171
rect 26145 23131 26203 23137
rect 28074 23128 28080 23180
rect 28132 23168 28138 23180
rect 28261 23171 28319 23177
rect 28261 23168 28273 23171
rect 28132 23140 28273 23168
rect 28132 23128 28138 23140
rect 28261 23137 28273 23140
rect 28307 23137 28319 23171
rect 28261 23131 28319 23137
rect 23661 23103 23719 23109
rect 23661 23069 23673 23103
rect 23707 23069 23719 23103
rect 23661 23063 23719 23069
rect 24397 23103 24455 23109
rect 24397 23069 24409 23103
rect 24443 23100 24455 23103
rect 25038 23100 25044 23112
rect 24443 23072 25044 23100
rect 24443 23069 24455 23072
rect 24397 23063 24455 23069
rect 25038 23060 25044 23072
rect 25096 23060 25102 23112
rect 25498 23100 25504 23112
rect 25459 23072 25504 23100
rect 25498 23060 25504 23072
rect 25556 23060 25562 23112
rect 26412 23103 26470 23109
rect 26412 23069 26424 23103
rect 26458 23100 26470 23103
rect 27338 23100 27344 23112
rect 26458 23072 27344 23100
rect 26458 23069 26470 23072
rect 26412 23063 26470 23069
rect 27338 23060 27344 23072
rect 27396 23060 27402 23112
rect 29564 23109 29592 23208
rect 27985 23103 28043 23109
rect 27985 23069 27997 23103
rect 28031 23069 28043 23103
rect 27985 23063 28043 23069
rect 29549 23103 29607 23109
rect 29549 23069 29561 23103
rect 29595 23069 29607 23103
rect 29549 23063 29607 23069
rect 22557 23035 22615 23041
rect 22557 23032 22569 23035
rect 22066 23004 22569 23032
rect 19935 23001 19947 23004
rect 19889 22995 19947 23001
rect 22557 23001 22569 23004
rect 22603 23001 22615 23035
rect 22557 22995 22615 23001
rect 23382 22992 23388 23044
rect 23440 23032 23446 23044
rect 28000 23032 28028 23063
rect 28350 23032 28356 23044
rect 23440 23004 28356 23032
rect 23440 22992 23446 23004
rect 28350 22992 28356 23004
rect 28408 22992 28414 23044
rect 16942 22964 16948 22976
rect 16316 22936 16948 22964
rect 16942 22924 16948 22936
rect 17000 22924 17006 22976
rect 17034 22924 17040 22976
rect 17092 22964 17098 22976
rect 18693 22967 18751 22973
rect 18693 22964 18705 22967
rect 17092 22936 18705 22964
rect 17092 22924 17098 22936
rect 18693 22933 18705 22936
rect 18739 22964 18751 22967
rect 18874 22964 18880 22976
rect 18739 22936 18880 22964
rect 18739 22933 18751 22936
rect 18693 22927 18751 22933
rect 18874 22924 18880 22936
rect 18932 22924 18938 22976
rect 19242 22924 19248 22976
rect 19300 22964 19306 22976
rect 23658 22964 23664 22976
rect 19300 22936 23664 22964
rect 19300 22924 19306 22936
rect 23658 22924 23664 22936
rect 23716 22924 23722 22976
rect 23753 22967 23811 22973
rect 23753 22933 23765 22967
rect 23799 22964 23811 22967
rect 24670 22964 24676 22976
rect 23799 22936 24676 22964
rect 23799 22933 23811 22936
rect 23753 22927 23811 22933
rect 24670 22924 24676 22936
rect 24728 22924 24734 22976
rect 26510 22924 26516 22976
rect 26568 22964 26574 22976
rect 29641 22967 29699 22973
rect 29641 22964 29653 22967
rect 26568 22936 29653 22964
rect 26568 22924 26574 22936
rect 29641 22933 29653 22936
rect 29687 22933 29699 22967
rect 29641 22927 29699 22933
rect 1104 22874 30820 22896
rect 1104 22822 10880 22874
rect 10932 22822 10944 22874
rect 10996 22822 11008 22874
rect 11060 22822 11072 22874
rect 11124 22822 11136 22874
rect 11188 22822 20811 22874
rect 20863 22822 20875 22874
rect 20927 22822 20939 22874
rect 20991 22822 21003 22874
rect 21055 22822 21067 22874
rect 21119 22822 30820 22874
rect 1104 22800 30820 22822
rect 8294 22720 8300 22772
rect 8352 22760 8358 22772
rect 9677 22763 9735 22769
rect 8352 22732 8892 22760
rect 8352 22720 8358 22732
rect 8864 22701 8892 22732
rect 9677 22729 9689 22763
rect 9723 22760 9735 22763
rect 9766 22760 9772 22772
rect 9723 22732 9772 22760
rect 9723 22729 9735 22732
rect 9677 22723 9735 22729
rect 9766 22720 9772 22732
rect 9824 22720 9830 22772
rect 11609 22763 11667 22769
rect 11609 22729 11621 22763
rect 11655 22760 11667 22763
rect 11974 22760 11980 22772
rect 11655 22732 11980 22760
rect 11655 22729 11667 22732
rect 11609 22723 11667 22729
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 13262 22720 13268 22772
rect 13320 22760 13326 22772
rect 14001 22763 14059 22769
rect 14001 22760 14013 22763
rect 13320 22732 14013 22760
rect 13320 22720 13326 22732
rect 14001 22729 14013 22732
rect 14047 22729 14059 22763
rect 14001 22723 14059 22729
rect 14461 22763 14519 22769
rect 14461 22729 14473 22763
rect 14507 22760 14519 22763
rect 17034 22760 17040 22772
rect 14507 22732 17040 22760
rect 14507 22729 14519 22732
rect 14461 22723 14519 22729
rect 17034 22720 17040 22732
rect 17092 22720 17098 22772
rect 17126 22720 17132 22772
rect 17184 22760 17190 22772
rect 19702 22760 19708 22772
rect 17184 22732 19708 22760
rect 17184 22720 17190 22732
rect 19702 22720 19708 22732
rect 19760 22720 19766 22772
rect 22002 22720 22008 22772
rect 22060 22760 22066 22772
rect 23382 22760 23388 22772
rect 22060 22732 23388 22760
rect 22060 22720 22066 22732
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 23658 22720 23664 22772
rect 23716 22760 23722 22772
rect 24673 22763 24731 22769
rect 24673 22760 24685 22763
rect 23716 22732 24685 22760
rect 23716 22720 23722 22732
rect 24673 22729 24685 22732
rect 24719 22760 24731 22763
rect 25130 22760 25136 22772
rect 24719 22732 25136 22760
rect 24719 22729 24731 22732
rect 24673 22723 24731 22729
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 27982 22760 27988 22772
rect 27943 22732 27988 22760
rect 27982 22720 27988 22732
rect 28040 22720 28046 22772
rect 8849 22695 8907 22701
rect 8849 22661 8861 22695
rect 8895 22661 8907 22695
rect 8849 22655 8907 22661
rect 9490 22652 9496 22704
rect 9548 22692 9554 22704
rect 18417 22695 18475 22701
rect 18417 22692 18429 22695
rect 9548 22664 18429 22692
rect 9548 22652 9554 22664
rect 18417 22661 18429 22664
rect 18463 22661 18475 22695
rect 18417 22655 18475 22661
rect 20993 22695 21051 22701
rect 20993 22661 21005 22695
rect 21039 22692 21051 22695
rect 22186 22692 22192 22704
rect 21039 22664 22192 22692
rect 21039 22661 21051 22664
rect 20993 22655 21051 22661
rect 22186 22652 22192 22664
rect 22244 22652 22250 22704
rect 23750 22692 23756 22704
rect 23711 22664 23756 22692
rect 23750 22652 23756 22664
rect 23808 22652 23814 22704
rect 24762 22692 24768 22704
rect 24504 22664 24768 22692
rect 8386 22584 8392 22636
rect 8444 22624 8450 22636
rect 8481 22627 8539 22633
rect 8481 22624 8493 22627
rect 8444 22596 8493 22624
rect 8444 22584 8450 22596
rect 8481 22593 8493 22596
rect 8527 22593 8539 22627
rect 8481 22587 8539 22593
rect 8573 22627 8631 22633
rect 8573 22593 8585 22627
rect 8619 22593 8631 22627
rect 8573 22587 8631 22593
rect 8757 22627 8815 22633
rect 8757 22593 8769 22627
rect 8803 22593 8815 22627
rect 8757 22587 8815 22593
rect 8588 22556 8616 22587
rect 8772 22556 8800 22587
rect 8938 22584 8944 22636
rect 8996 22624 9002 22636
rect 8996 22596 9041 22624
rect 8996 22584 9002 22596
rect 9122 22584 9128 22636
rect 9180 22624 9186 22636
rect 9585 22627 9643 22633
rect 9585 22624 9597 22627
rect 9180 22596 9597 22624
rect 9180 22584 9186 22596
rect 9585 22593 9597 22596
rect 9631 22593 9643 22627
rect 9585 22587 9643 22593
rect 9766 22584 9772 22636
rect 9824 22624 9830 22636
rect 10505 22627 10563 22633
rect 10505 22624 10517 22627
rect 9824 22596 10517 22624
rect 9824 22584 9830 22596
rect 10505 22593 10517 22596
rect 10551 22593 10563 22627
rect 10505 22587 10563 22593
rect 10781 22627 10839 22633
rect 10781 22593 10793 22627
rect 10827 22624 10839 22627
rect 11238 22624 11244 22636
rect 10827 22596 11244 22624
rect 10827 22593 10839 22596
rect 10781 22587 10839 22593
rect 11238 22584 11244 22596
rect 11296 22584 11302 22636
rect 11517 22627 11575 22633
rect 11517 22593 11529 22627
rect 11563 22624 11575 22627
rect 11882 22624 11888 22636
rect 11563 22596 11888 22624
rect 11563 22593 11575 22596
rect 11517 22587 11575 22593
rect 11882 22584 11888 22596
rect 11940 22584 11946 22636
rect 12161 22627 12219 22633
rect 12161 22593 12173 22627
rect 12207 22624 12219 22627
rect 12710 22624 12716 22636
rect 12207 22596 12716 22624
rect 12207 22593 12219 22596
rect 12161 22587 12219 22593
rect 12710 22584 12716 22596
rect 12768 22584 12774 22636
rect 13357 22627 13415 22633
rect 13357 22593 13369 22627
rect 13403 22593 13415 22627
rect 13357 22587 13415 22593
rect 9674 22556 9680 22568
rect 8588 22528 8708 22556
rect 8772 22528 9680 22556
rect 8570 22448 8576 22500
rect 8628 22488 8634 22500
rect 8680 22488 8708 22528
rect 9674 22516 9680 22528
rect 9732 22516 9738 22568
rect 11330 22516 11336 22568
rect 11388 22556 11394 22568
rect 13372 22556 13400 22587
rect 13538 22584 13544 22636
rect 13596 22624 13602 22636
rect 14369 22627 14427 22633
rect 14369 22624 14381 22627
rect 13596 22596 14381 22624
rect 13596 22584 13602 22596
rect 14369 22593 14381 22596
rect 14415 22593 14427 22627
rect 15194 22624 15200 22636
rect 15155 22596 15200 22624
rect 14369 22587 14427 22593
rect 15194 22584 15200 22596
rect 15252 22584 15258 22636
rect 15286 22584 15292 22636
rect 15344 22584 15350 22636
rect 15381 22627 15439 22633
rect 15381 22593 15393 22627
rect 15427 22593 15439 22627
rect 15381 22587 15439 22593
rect 11388 22528 13400 22556
rect 11388 22516 11394 22528
rect 9950 22488 9956 22500
rect 8628 22460 9956 22488
rect 8628 22448 8634 22460
rect 9950 22448 9956 22460
rect 10008 22448 10014 22500
rect 10689 22491 10747 22497
rect 10689 22457 10701 22491
rect 10735 22488 10747 22491
rect 12158 22488 12164 22500
rect 10735 22460 12164 22488
rect 10735 22457 10747 22460
rect 10689 22451 10747 22457
rect 12158 22448 12164 22460
rect 12216 22448 12222 22500
rect 13372 22488 13400 22528
rect 14645 22559 14703 22565
rect 14645 22525 14657 22559
rect 14691 22556 14703 22559
rect 14734 22556 14740 22568
rect 14691 22528 14740 22556
rect 14691 22525 14703 22528
rect 14645 22519 14703 22525
rect 14734 22516 14740 22528
rect 14792 22516 14798 22568
rect 15194 22488 15200 22500
rect 13372 22460 15200 22488
rect 15194 22448 15200 22460
rect 15252 22448 15258 22500
rect 15304 22488 15332 22584
rect 15396 22556 15424 22587
rect 15470 22584 15476 22636
rect 15528 22624 15534 22636
rect 15746 22624 15752 22636
rect 15528 22596 15573 22624
rect 15707 22596 15752 22624
rect 15528 22584 15534 22596
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 16574 22584 16580 22636
rect 16632 22624 16638 22636
rect 16632 22596 16804 22624
rect 16632 22584 16638 22596
rect 16776 22556 16804 22596
rect 16942 22584 16948 22636
rect 17000 22624 17006 22636
rect 17037 22627 17095 22633
rect 17037 22624 17049 22627
rect 17000 22596 17049 22624
rect 17000 22584 17006 22596
rect 17037 22593 17049 22596
rect 17083 22593 17095 22627
rect 17037 22587 17095 22593
rect 17129 22627 17187 22633
rect 17129 22593 17141 22627
rect 17175 22624 17187 22627
rect 17402 22624 17408 22636
rect 17175 22596 17408 22624
rect 17175 22593 17187 22596
rect 17129 22587 17187 22593
rect 17402 22584 17408 22596
rect 17460 22584 17466 22636
rect 20806 22624 20812 22636
rect 20719 22596 20812 22624
rect 20806 22584 20812 22596
rect 20864 22624 20870 22636
rect 21266 22624 21272 22636
rect 20864 22596 21272 22624
rect 20864 22584 20870 22596
rect 21266 22584 21272 22596
rect 21324 22584 21330 22636
rect 21634 22624 21640 22636
rect 21376 22596 21640 22624
rect 17221 22559 17279 22565
rect 17221 22556 17233 22559
rect 15396 22528 16712 22556
rect 16776 22528 17233 22556
rect 15657 22491 15715 22497
rect 15657 22488 15669 22491
rect 15304 22460 15669 22488
rect 15657 22457 15669 22460
rect 15703 22488 15715 22491
rect 15746 22488 15752 22500
rect 15703 22460 15752 22488
rect 15703 22457 15715 22460
rect 15657 22451 15715 22457
rect 15746 22448 15752 22460
rect 15804 22448 15810 22500
rect 16684 22497 16712 22528
rect 17221 22525 17233 22528
rect 17267 22525 17279 22559
rect 17221 22519 17279 22525
rect 17494 22516 17500 22568
rect 17552 22556 17558 22568
rect 19150 22556 19156 22568
rect 17552 22528 19156 22556
rect 17552 22516 17558 22528
rect 19150 22516 19156 22528
rect 19208 22516 19214 22568
rect 20622 22516 20628 22568
rect 20680 22556 20686 22568
rect 21376 22556 21404 22596
rect 21634 22584 21640 22596
rect 21692 22584 21698 22636
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22624 21879 22627
rect 21910 22624 21916 22636
rect 21867 22596 21916 22624
rect 21867 22593 21879 22596
rect 21821 22587 21879 22593
rect 21910 22584 21916 22596
rect 21968 22584 21974 22636
rect 22088 22627 22146 22633
rect 22088 22593 22100 22627
rect 22134 22624 22146 22627
rect 22554 22624 22560 22636
rect 22134 22596 22560 22624
rect 22134 22593 22146 22596
rect 22088 22587 22146 22593
rect 22554 22584 22560 22596
rect 22612 22584 22618 22636
rect 24504 22633 24532 22664
rect 24762 22652 24768 22664
rect 24820 22652 24826 22704
rect 27522 22692 27528 22704
rect 27448 22664 27528 22692
rect 24489 22627 24547 22633
rect 24489 22593 24501 22627
rect 24535 22593 24547 22627
rect 24489 22587 24547 22593
rect 24578 22584 24584 22636
rect 24636 22624 24642 22636
rect 25317 22627 25375 22633
rect 25317 22624 25329 22627
rect 24636 22596 25329 22624
rect 24636 22584 24642 22596
rect 25317 22593 25329 22596
rect 25363 22593 25375 22627
rect 25317 22587 25375 22593
rect 26237 22627 26295 22633
rect 26237 22593 26249 22627
rect 26283 22593 26295 22627
rect 26237 22587 26295 22593
rect 27249 22627 27307 22633
rect 27249 22593 27261 22627
rect 27295 22624 27307 22627
rect 27338 22624 27344 22636
rect 27295 22596 27344 22624
rect 27295 22593 27307 22596
rect 27249 22587 27307 22593
rect 24854 22556 24860 22568
rect 20680 22528 21404 22556
rect 22940 22528 24860 22556
rect 20680 22516 20686 22528
rect 16669 22491 16727 22497
rect 16669 22457 16681 22491
rect 16715 22457 16727 22491
rect 16669 22451 16727 22457
rect 18414 22448 18420 22500
rect 18472 22488 18478 22500
rect 18472 22460 21496 22488
rect 18472 22448 18478 22460
rect 8478 22420 8484 22432
rect 8439 22392 8484 22420
rect 8478 22380 8484 22392
rect 8536 22380 8542 22432
rect 9858 22380 9864 22432
rect 9916 22420 9922 22432
rect 10321 22423 10379 22429
rect 10321 22420 10333 22423
rect 9916 22392 10333 22420
rect 9916 22380 9922 22392
rect 10321 22389 10333 22392
rect 10367 22389 10379 22423
rect 10321 22383 10379 22389
rect 12253 22423 12311 22429
rect 12253 22389 12265 22423
rect 12299 22420 12311 22423
rect 12526 22420 12532 22432
rect 12299 22392 12532 22420
rect 12299 22389 12311 22392
rect 12253 22383 12311 22389
rect 12526 22380 12532 22392
rect 12584 22380 12590 22432
rect 13078 22380 13084 22432
rect 13136 22420 13142 22432
rect 13449 22423 13507 22429
rect 13449 22420 13461 22423
rect 13136 22392 13461 22420
rect 13136 22380 13142 22392
rect 13449 22389 13461 22392
rect 13495 22420 13507 22423
rect 14366 22420 14372 22432
rect 13495 22392 14372 22420
rect 13495 22389 13507 22392
rect 13449 22383 13507 22389
rect 14366 22380 14372 22392
rect 14424 22380 14430 22432
rect 15378 22380 15384 22432
rect 15436 22420 15442 22432
rect 15565 22423 15623 22429
rect 15565 22420 15577 22423
rect 15436 22392 15577 22420
rect 15436 22380 15442 22392
rect 15565 22389 15577 22392
rect 15611 22389 15623 22423
rect 15565 22383 15623 22389
rect 16942 22380 16948 22432
rect 17000 22420 17006 22432
rect 17678 22420 17684 22432
rect 17000 22392 17684 22420
rect 17000 22380 17006 22392
rect 17678 22380 17684 22392
rect 17736 22380 17742 22432
rect 21177 22423 21235 22429
rect 21177 22389 21189 22423
rect 21223 22420 21235 22423
rect 21358 22420 21364 22432
rect 21223 22392 21364 22420
rect 21223 22389 21235 22392
rect 21177 22383 21235 22389
rect 21358 22380 21364 22392
rect 21416 22380 21422 22432
rect 21468 22420 21496 22460
rect 22940 22420 22968 22528
rect 24854 22516 24860 22528
rect 24912 22556 24918 22568
rect 25501 22559 25559 22565
rect 25501 22556 25513 22559
rect 24912 22528 25513 22556
rect 24912 22516 24918 22528
rect 25501 22525 25513 22528
rect 25547 22556 25559 22559
rect 25590 22556 25596 22568
rect 25547 22528 25596 22556
rect 25547 22525 25559 22528
rect 25501 22519 25559 22525
rect 25590 22516 25596 22528
rect 25648 22516 25654 22568
rect 23106 22448 23112 22500
rect 23164 22488 23170 22500
rect 23937 22491 23995 22497
rect 23937 22488 23949 22491
rect 23164 22460 23949 22488
rect 23164 22448 23170 22460
rect 23937 22457 23949 22460
rect 23983 22457 23995 22491
rect 26252 22488 26280 22587
rect 27338 22584 27344 22596
rect 27396 22584 27402 22636
rect 27448 22633 27476 22664
rect 27522 22652 27528 22664
rect 27580 22652 27586 22704
rect 27433 22627 27491 22633
rect 27433 22593 27445 22627
rect 27479 22593 27491 22627
rect 27798 22624 27804 22636
rect 27759 22596 27804 22624
rect 27433 22587 27491 22593
rect 27798 22584 27804 22596
rect 27856 22584 27862 22636
rect 28442 22624 28448 22636
rect 28403 22596 28448 22624
rect 28442 22584 28448 22596
rect 28500 22584 28506 22636
rect 28712 22627 28770 22633
rect 28712 22593 28724 22627
rect 28758 22624 28770 22627
rect 28994 22624 29000 22636
rect 28758 22596 29000 22624
rect 28758 22593 28770 22596
rect 28712 22587 28770 22593
rect 28994 22584 29000 22596
rect 29052 22584 29058 22636
rect 26878 22516 26884 22568
rect 26936 22556 26942 22568
rect 27525 22559 27583 22565
rect 27525 22556 27537 22559
rect 26936 22528 27537 22556
rect 26936 22516 26942 22528
rect 27525 22525 27537 22528
rect 27571 22525 27583 22559
rect 27525 22519 27583 22525
rect 27617 22559 27675 22565
rect 27617 22525 27629 22559
rect 27663 22556 27675 22559
rect 28074 22556 28080 22568
rect 27663 22528 28080 22556
rect 27663 22525 27675 22528
rect 27617 22519 27675 22525
rect 28074 22516 28080 22528
rect 28132 22516 28138 22568
rect 27982 22488 27988 22500
rect 26252 22460 27988 22488
rect 23937 22451 23995 22457
rect 27982 22448 27988 22460
rect 28040 22448 28046 22500
rect 21468 22392 22968 22420
rect 23014 22380 23020 22432
rect 23072 22420 23078 22432
rect 23201 22423 23259 22429
rect 23201 22420 23213 22423
rect 23072 22392 23213 22420
rect 23072 22380 23078 22392
rect 23201 22389 23213 22392
rect 23247 22389 23259 22423
rect 26326 22420 26332 22432
rect 26287 22392 26332 22420
rect 23201 22383 23259 22389
rect 26326 22380 26332 22392
rect 26384 22380 26390 22432
rect 27614 22380 27620 22432
rect 27672 22420 27678 22432
rect 27798 22420 27804 22432
rect 27672 22392 27804 22420
rect 27672 22380 27678 22392
rect 27798 22380 27804 22392
rect 27856 22380 27862 22432
rect 29546 22380 29552 22432
rect 29604 22420 29610 22432
rect 29825 22423 29883 22429
rect 29825 22420 29837 22423
rect 29604 22392 29837 22420
rect 29604 22380 29610 22392
rect 29825 22389 29837 22392
rect 29871 22389 29883 22423
rect 29825 22383 29883 22389
rect 1104 22330 30820 22352
rect 1104 22278 5915 22330
rect 5967 22278 5979 22330
rect 6031 22278 6043 22330
rect 6095 22278 6107 22330
rect 6159 22278 6171 22330
rect 6223 22278 15846 22330
rect 15898 22278 15910 22330
rect 15962 22278 15974 22330
rect 16026 22278 16038 22330
rect 16090 22278 16102 22330
rect 16154 22278 25776 22330
rect 25828 22278 25840 22330
rect 25892 22278 25904 22330
rect 25956 22278 25968 22330
rect 26020 22278 26032 22330
rect 26084 22278 30820 22330
rect 1104 22256 30820 22278
rect 8294 22216 8300 22228
rect 8255 22188 8300 22216
rect 8294 22176 8300 22188
rect 8352 22176 8358 22228
rect 8938 22176 8944 22228
rect 8996 22216 9002 22228
rect 9493 22219 9551 22225
rect 9493 22216 9505 22219
rect 8996 22188 9505 22216
rect 8996 22176 9002 22188
rect 9493 22185 9505 22188
rect 9539 22185 9551 22219
rect 9493 22179 9551 22185
rect 9766 22176 9772 22228
rect 9824 22216 9830 22228
rect 10778 22216 10784 22228
rect 9824 22188 10784 22216
rect 9824 22176 9830 22188
rect 10778 22176 10784 22188
rect 10836 22176 10842 22228
rect 12526 22216 12532 22228
rect 11440 22188 12532 22216
rect 9858 22148 9864 22160
rect 9819 22120 9864 22148
rect 9858 22108 9864 22120
rect 9916 22108 9922 22160
rect 2130 22040 2136 22092
rect 2188 22080 2194 22092
rect 2188 22052 2774 22080
rect 2188 22040 2194 22052
rect 2746 21876 2774 22052
rect 9582 22040 9588 22092
rect 9640 22080 9646 22092
rect 9769 22083 9827 22089
rect 9769 22080 9781 22083
rect 9640 22052 9781 22080
rect 9640 22040 9646 22052
rect 9769 22049 9781 22052
rect 9815 22080 9827 22083
rect 9815 22052 11008 22080
rect 9815 22049 9827 22052
rect 9769 22043 9827 22049
rect 8205 22015 8263 22021
rect 8205 21981 8217 22015
rect 8251 22012 8263 22015
rect 8570 22012 8576 22024
rect 8251 21984 8576 22012
rect 8251 21981 8263 21984
rect 8205 21975 8263 21981
rect 8570 21972 8576 21984
rect 8628 21972 8634 22024
rect 8662 21972 8668 22024
rect 8720 22012 8726 22024
rect 9677 22015 9735 22021
rect 9677 22012 9689 22015
rect 8720 21984 9689 22012
rect 8720 21972 8726 21984
rect 9677 21981 9689 21984
rect 9723 21981 9735 22015
rect 9677 21975 9735 21981
rect 9953 22015 10011 22021
rect 9953 21981 9965 22015
rect 9999 22012 10011 22015
rect 10042 22012 10048 22024
rect 9999 21984 10048 22012
rect 9999 21981 10011 21984
rect 9953 21975 10011 21981
rect 10042 21972 10048 21984
rect 10100 21972 10106 22024
rect 10137 22015 10195 22021
rect 10137 21981 10149 22015
rect 10183 21981 10195 22015
rect 10137 21975 10195 21981
rect 10042 21876 10048 21888
rect 2746 21848 10048 21876
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 10152 21876 10180 21975
rect 10686 21972 10692 22024
rect 10744 22012 10750 22024
rect 10980 22021 11008 22052
rect 10873 22015 10931 22021
rect 10873 22012 10885 22015
rect 10744 21984 10885 22012
rect 10744 21972 10750 21984
rect 10873 21981 10885 21984
rect 10919 21981 10931 22015
rect 10873 21975 10931 21981
rect 10965 22015 11023 22021
rect 10965 21981 10977 22015
rect 11011 21981 11023 22015
rect 10965 21975 11023 21981
rect 11057 22015 11115 22021
rect 11057 21981 11069 22015
rect 11103 22012 11115 22015
rect 11146 22012 11152 22024
rect 11103 21984 11152 22012
rect 11103 21981 11115 21984
rect 11057 21975 11115 21981
rect 11146 21972 11152 21984
rect 11204 21972 11210 22024
rect 11241 22015 11299 22021
rect 11241 21981 11253 22015
rect 11287 22012 11299 22015
rect 11440 22012 11468 22188
rect 12526 22176 12532 22188
rect 12584 22176 12590 22228
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 17218 22216 17224 22228
rect 16632 22188 17224 22216
rect 16632 22176 16638 22188
rect 17218 22176 17224 22188
rect 17276 22176 17282 22228
rect 20714 22176 20720 22228
rect 20772 22216 20778 22228
rect 23017 22219 23075 22225
rect 23017 22216 23029 22219
rect 20772 22188 23029 22216
rect 20772 22176 20778 22188
rect 23017 22185 23029 22188
rect 23063 22185 23075 22219
rect 23017 22179 23075 22185
rect 12986 22148 12992 22160
rect 12176 22120 12992 22148
rect 12176 22080 12204 22120
rect 12986 22108 12992 22120
rect 13044 22108 13050 22160
rect 17034 22148 17040 22160
rect 16684 22120 17040 22148
rect 15562 22080 15568 22092
rect 11900 22052 12204 22080
rect 15212 22052 15568 22080
rect 11900 22021 11928 22052
rect 11287 21984 11468 22012
rect 11885 22015 11943 22021
rect 11287 21981 11299 21984
rect 11241 21975 11299 21981
rect 11885 21981 11897 22015
rect 11931 21981 11943 22015
rect 12069 22015 12127 22021
rect 12069 22012 12081 22015
rect 11885 21975 11943 21981
rect 11992 21984 12081 22012
rect 10597 21947 10655 21953
rect 10597 21913 10609 21947
rect 10643 21944 10655 21947
rect 11992 21944 12020 21984
rect 12069 21981 12081 21984
rect 12115 21981 12127 22015
rect 12069 21975 12127 21981
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 22012 12219 22015
rect 12434 22012 12440 22024
rect 12207 21984 12440 22012
rect 12207 21981 12219 21984
rect 12161 21975 12219 21981
rect 12434 21972 12440 21984
rect 12492 21972 12498 22024
rect 12618 22012 12624 22024
rect 12579 21984 12624 22012
rect 12618 21972 12624 21984
rect 12676 21972 12682 22024
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 22012 12771 22015
rect 15212 22012 15240 22052
rect 15562 22040 15568 22052
rect 15620 22040 15626 22092
rect 15838 22080 15844 22092
rect 15672 22052 15844 22080
rect 15378 22012 15384 22024
rect 12759 21984 15240 22012
rect 15339 21984 15384 22012
rect 12759 21981 12771 21984
rect 12713 21975 12771 21981
rect 15378 21972 15384 21984
rect 15436 21972 15442 22024
rect 15470 21972 15476 22024
rect 15528 22012 15534 22024
rect 15672 22012 15700 22052
rect 15838 22040 15844 22052
rect 15896 22040 15902 22092
rect 16684 22089 16712 22120
rect 17034 22108 17040 22120
rect 17092 22108 17098 22160
rect 17972 22120 18828 22148
rect 16669 22083 16727 22089
rect 16669 22049 16681 22083
rect 16715 22080 16727 22083
rect 16850 22080 16856 22092
rect 16715 22052 16749 22080
rect 16811 22052 16856 22080
rect 16715 22049 16727 22052
rect 16669 22043 16727 22049
rect 16850 22040 16856 22052
rect 16908 22040 16914 22092
rect 17218 22040 17224 22092
rect 17276 22080 17282 22092
rect 17494 22080 17500 22092
rect 17276 22052 17500 22080
rect 17276 22040 17282 22052
rect 17494 22040 17500 22052
rect 17552 22040 17558 22092
rect 15528 21984 15700 22012
rect 15528 21972 15534 21984
rect 15746 21972 15752 22024
rect 15804 22012 15810 22024
rect 17310 22012 17316 22024
rect 15804 21984 17316 22012
rect 15804 21972 15810 21984
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 17972 22021 18000 22120
rect 18800 22080 18828 22120
rect 21450 22108 21456 22160
rect 21508 22148 21514 22160
rect 21821 22151 21879 22157
rect 21821 22148 21833 22151
rect 21508 22120 21833 22148
rect 21508 22108 21514 22120
rect 21821 22117 21833 22120
rect 21867 22148 21879 22151
rect 22462 22148 22468 22160
rect 21867 22120 22468 22148
rect 21867 22117 21879 22120
rect 21821 22111 21879 22117
rect 22462 22108 22468 22120
rect 22520 22108 22526 22160
rect 23032 22148 23060 22179
rect 23106 22176 23112 22228
rect 23164 22216 23170 22228
rect 24489 22219 24547 22225
rect 24489 22216 24501 22219
rect 23164 22188 24501 22216
rect 23164 22176 23170 22188
rect 24489 22185 24501 22188
rect 24535 22185 24547 22219
rect 24489 22179 24547 22185
rect 24857 22219 24915 22225
rect 24857 22185 24869 22219
rect 24903 22216 24915 22219
rect 25498 22216 25504 22228
rect 24903 22188 25504 22216
rect 24903 22185 24915 22188
rect 24857 22179 24915 22185
rect 25498 22176 25504 22188
rect 25556 22176 25562 22228
rect 27614 22176 27620 22228
rect 27672 22216 27678 22228
rect 28350 22216 28356 22228
rect 27672 22188 28356 22216
rect 27672 22176 27678 22188
rect 28350 22176 28356 22188
rect 28408 22176 28414 22228
rect 28626 22176 28632 22228
rect 28684 22216 28690 22228
rect 28902 22216 28908 22228
rect 28684 22188 28908 22216
rect 28684 22176 28690 22188
rect 28902 22176 28908 22188
rect 28960 22176 28966 22228
rect 23750 22148 23756 22160
rect 23032 22120 23756 22148
rect 23750 22108 23756 22120
rect 23808 22108 23814 22160
rect 25590 22108 25596 22160
rect 25648 22148 25654 22160
rect 25648 22120 25820 22148
rect 25648 22108 25654 22120
rect 18800 22052 19196 22080
rect 17957 22015 18015 22021
rect 17957 21981 17969 22015
rect 18003 21981 18015 22015
rect 18138 22012 18144 22024
rect 18099 21984 18144 22012
rect 17957 21975 18015 21981
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 18325 22015 18383 22021
rect 18325 21981 18337 22015
rect 18371 22012 18383 22015
rect 18414 22012 18420 22024
rect 18371 21984 18420 22012
rect 18371 21981 18383 21984
rect 18325 21975 18383 21981
rect 10643 21916 12020 21944
rect 10643 21913 10655 21916
rect 10597 21907 10655 21913
rect 13814 21904 13820 21956
rect 13872 21944 13878 21956
rect 14093 21947 14151 21953
rect 14093 21944 14105 21947
rect 13872 21916 14105 21944
rect 13872 21904 13878 21916
rect 14093 21913 14105 21916
rect 14139 21913 14151 21947
rect 14093 21907 14151 21913
rect 14182 21904 14188 21956
rect 14240 21944 14246 21956
rect 14277 21947 14335 21953
rect 14277 21944 14289 21947
rect 14240 21916 14289 21944
rect 14240 21904 14246 21916
rect 14277 21913 14289 21916
rect 14323 21913 14335 21947
rect 14277 21907 14335 21913
rect 11514 21876 11520 21888
rect 10152 21848 11520 21876
rect 11514 21836 11520 21848
rect 11572 21836 11578 21888
rect 11698 21876 11704 21888
rect 11659 21848 11704 21876
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 14461 21879 14519 21885
rect 14461 21845 14473 21879
rect 14507 21876 14519 21879
rect 14826 21876 14832 21888
rect 14507 21848 14832 21876
rect 14507 21845 14519 21848
rect 14461 21839 14519 21845
rect 14826 21836 14832 21848
rect 14884 21836 14890 21888
rect 15010 21876 15016 21888
rect 14971 21848 15016 21876
rect 15010 21836 15016 21848
rect 15068 21836 15074 21888
rect 15473 21879 15531 21885
rect 15473 21845 15485 21879
rect 15519 21876 15531 21879
rect 16209 21879 16267 21885
rect 16209 21876 16221 21879
rect 15519 21848 16221 21876
rect 15519 21845 15531 21848
rect 15473 21839 15531 21845
rect 16209 21845 16221 21848
rect 16255 21845 16267 21879
rect 16574 21876 16580 21888
rect 16535 21848 16580 21876
rect 16209 21839 16267 21845
rect 16574 21836 16580 21848
rect 16632 21836 16638 21888
rect 18248 21876 18276 21975
rect 18414 21972 18420 21984
rect 18472 21972 18478 22024
rect 18509 22015 18567 22021
rect 18509 21981 18521 22015
rect 18555 22012 18567 22015
rect 18782 22012 18788 22024
rect 18555 21984 18788 22012
rect 18555 21981 18567 21984
rect 18509 21975 18567 21981
rect 18782 21972 18788 21984
rect 18840 21972 18846 22024
rect 18598 21904 18604 21956
rect 18656 21944 18662 21956
rect 18693 21947 18751 21953
rect 18693 21944 18705 21947
rect 18656 21916 18705 21944
rect 18656 21904 18662 21916
rect 18693 21913 18705 21916
rect 18739 21913 18751 21947
rect 19168 21944 19196 22052
rect 21910 22040 21916 22092
rect 21968 22080 21974 22092
rect 25682 22080 25688 22092
rect 21968 22052 25688 22080
rect 21968 22040 21974 22052
rect 25682 22040 25688 22052
rect 25740 22040 25746 22092
rect 25792 22089 25820 22120
rect 26804 22120 29132 22148
rect 25777 22083 25835 22089
rect 25777 22049 25789 22083
rect 25823 22049 25835 22083
rect 26804 22080 26832 22120
rect 27430 22080 27436 22092
rect 25777 22043 25835 22049
rect 25976 22052 26832 22080
rect 26896 22052 27436 22080
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 22012 19671 22015
rect 20441 22015 20499 22021
rect 19659 21984 19932 22012
rect 19659 21981 19671 21984
rect 19613 21975 19671 21981
rect 19168 21916 19840 21944
rect 18693 21907 18751 21913
rect 19812 21888 19840 21916
rect 19058 21876 19064 21888
rect 18248 21848 19064 21876
rect 19058 21836 19064 21848
rect 19116 21836 19122 21888
rect 19794 21876 19800 21888
rect 19755 21848 19800 21876
rect 19794 21836 19800 21848
rect 19852 21836 19858 21888
rect 19904 21876 19932 21984
rect 20441 21981 20453 22015
rect 20487 22012 20499 22015
rect 22002 22012 22008 22024
rect 20487 21984 22008 22012
rect 20487 21981 20499 21984
rect 20441 21975 20499 21981
rect 22002 21972 22008 21984
rect 22060 21972 22066 22024
rect 22925 22015 22983 22021
rect 22925 21981 22937 22015
rect 22971 22012 22983 22015
rect 23382 22012 23388 22024
rect 22971 21984 23388 22012
rect 22971 21981 22983 21984
rect 22925 21975 22983 21981
rect 23382 21972 23388 21984
rect 23440 21972 23446 22024
rect 24210 21972 24216 22024
rect 24268 22012 24274 22024
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 24268 21984 24409 22012
rect 24268 21972 24274 21984
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 25406 22012 25412 22024
rect 25367 21984 25412 22012
rect 24397 21975 24455 21981
rect 25406 21972 25412 21984
rect 25464 21972 25470 22024
rect 25590 22012 25596 22024
rect 25551 21984 25596 22012
rect 25590 21972 25596 21984
rect 25648 21972 25654 22024
rect 25976 22021 26004 22052
rect 26896 22021 26924 22052
rect 27430 22040 27436 22052
rect 27488 22040 27494 22092
rect 28718 22080 28724 22092
rect 28460 22052 28724 22080
rect 27154 22021 27160 22024
rect 25961 22015 26019 22021
rect 25961 21981 25973 22015
rect 26007 21981 26019 22015
rect 25961 21975 26019 21981
rect 26697 22015 26755 22021
rect 26697 21981 26709 22015
rect 26743 21981 26755 22015
rect 26697 21975 26755 21981
rect 26881 22015 26939 22021
rect 26881 21981 26893 22015
rect 26927 21981 26939 22015
rect 26881 21975 26939 21981
rect 26967 22015 27025 22021
rect 26967 21981 26979 22015
rect 27013 21981 27025 22015
rect 26967 21975 27025 21981
rect 27111 22015 27160 22021
rect 27111 21981 27123 22015
rect 27157 21981 27160 22015
rect 27111 21975 27160 21981
rect 20708 21947 20766 21953
rect 20708 21913 20720 21947
rect 20754 21944 20766 21947
rect 21266 21944 21272 21956
rect 20754 21916 21272 21944
rect 20754 21913 20766 21916
rect 20708 21907 20766 21913
rect 21266 21904 21272 21916
rect 21324 21904 21330 21956
rect 23934 21944 23940 21956
rect 21376 21916 23940 21944
rect 19978 21876 19984 21888
rect 19904 21848 19984 21876
rect 19978 21836 19984 21848
rect 20036 21876 20042 21888
rect 21376 21876 21404 21916
rect 23934 21904 23940 21916
rect 23992 21904 23998 21956
rect 25314 21904 25320 21956
rect 25372 21944 25378 21956
rect 26145 21947 26203 21953
rect 26145 21944 26157 21947
rect 25372 21916 26157 21944
rect 25372 21904 25378 21916
rect 26145 21913 26157 21916
rect 26191 21913 26203 21947
rect 26145 21907 26203 21913
rect 20036 21848 21404 21876
rect 20036 21836 20042 21848
rect 22094 21836 22100 21888
rect 22152 21876 22158 21888
rect 22738 21876 22744 21888
rect 22152 21848 22744 21876
rect 22152 21836 22158 21848
rect 22738 21836 22744 21848
rect 22796 21836 22802 21888
rect 22922 21836 22928 21888
rect 22980 21876 22986 21888
rect 23385 21879 23443 21885
rect 23385 21876 23397 21879
rect 22980 21848 23397 21876
rect 22980 21836 22986 21848
rect 23385 21845 23397 21848
rect 23431 21845 23443 21879
rect 26712 21876 26740 21975
rect 26786 21904 26792 21956
rect 26844 21944 26850 21956
rect 26988 21944 27016 21975
rect 27154 21972 27160 21975
rect 27212 21972 27218 22024
rect 27249 22015 27307 22021
rect 27249 21981 27261 22015
rect 27295 22012 27307 22015
rect 28074 22012 28080 22024
rect 27295 21984 28080 22012
rect 27295 21981 27307 21984
rect 27249 21975 27307 21981
rect 28074 21972 28080 21984
rect 28132 21972 28138 22024
rect 28460 22021 28488 22052
rect 28718 22040 28724 22052
rect 28776 22040 28782 22092
rect 28994 22080 29000 22092
rect 28955 22052 29000 22080
rect 28994 22040 29000 22052
rect 29052 22040 29058 22092
rect 29104 22080 29132 22120
rect 29641 22083 29699 22089
rect 29641 22080 29653 22083
rect 29104 22052 29653 22080
rect 29641 22049 29653 22052
rect 29687 22049 29699 22083
rect 29641 22043 29699 22049
rect 28261 22015 28319 22021
rect 28261 21981 28273 22015
rect 28307 21981 28319 22015
rect 28261 21975 28319 21981
rect 28445 22015 28503 22021
rect 28445 21981 28457 22015
rect 28491 21981 28503 22015
rect 28445 21975 28503 21981
rect 28537 22015 28595 22021
rect 28537 21981 28549 22015
rect 28583 21981 28595 22015
rect 28537 21975 28595 21981
rect 26844 21916 27016 21944
rect 26844 21904 26850 21916
rect 27338 21904 27344 21956
rect 27396 21944 27402 21956
rect 28276 21944 28304 21975
rect 27396 21916 28304 21944
rect 27396 21904 27402 21916
rect 28350 21904 28356 21956
rect 28408 21944 28414 21956
rect 28552 21944 28580 21975
rect 28626 21972 28632 22024
rect 28684 22012 28690 22024
rect 28813 22015 28871 22021
rect 28684 21984 28729 22012
rect 28684 21972 28690 21984
rect 28813 21981 28825 22015
rect 28859 22012 28871 22015
rect 29546 22012 29552 22024
rect 28859 21984 29552 22012
rect 28859 21981 28871 21984
rect 28813 21975 28871 21981
rect 29546 21972 29552 21984
rect 29604 21972 29610 22024
rect 28408 21916 28580 21944
rect 28408 21904 28414 21916
rect 27062 21876 27068 21888
rect 26712 21848 27068 21876
rect 23385 21839 23443 21845
rect 27062 21836 27068 21848
rect 27120 21836 27126 21888
rect 27246 21836 27252 21888
rect 27304 21876 27310 21888
rect 27433 21879 27491 21885
rect 27433 21876 27445 21879
rect 27304 21848 27445 21876
rect 27304 21836 27310 21848
rect 27433 21845 27445 21848
rect 27479 21845 27491 21879
rect 27433 21839 27491 21845
rect 1104 21786 30820 21808
rect 1104 21734 10880 21786
rect 10932 21734 10944 21786
rect 10996 21734 11008 21786
rect 11060 21734 11072 21786
rect 11124 21734 11136 21786
rect 11188 21734 20811 21786
rect 20863 21734 20875 21786
rect 20927 21734 20939 21786
rect 20991 21734 21003 21786
rect 21055 21734 21067 21786
rect 21119 21734 30820 21786
rect 1104 21712 30820 21734
rect 8662 21632 8668 21684
rect 8720 21672 8726 21684
rect 9125 21675 9183 21681
rect 9125 21672 9137 21675
rect 8720 21644 9137 21672
rect 8720 21632 8726 21644
rect 9125 21641 9137 21644
rect 9171 21672 9183 21675
rect 10686 21672 10692 21684
rect 9171 21644 10692 21672
rect 9171 21641 9183 21644
rect 9125 21635 9183 21641
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 11238 21632 11244 21684
rect 11296 21672 11302 21684
rect 12158 21672 12164 21684
rect 11296 21644 12164 21672
rect 11296 21632 11302 21644
rect 12158 21632 12164 21644
rect 12216 21632 12222 21684
rect 13357 21675 13415 21681
rect 13357 21641 13369 21675
rect 13403 21672 13415 21675
rect 13446 21672 13452 21684
rect 13403 21644 13452 21672
rect 13403 21641 13415 21644
rect 13357 21635 13415 21641
rect 13446 21632 13452 21644
rect 13504 21632 13510 21684
rect 16574 21632 16580 21684
rect 16632 21672 16638 21684
rect 16853 21675 16911 21681
rect 16853 21672 16865 21675
rect 16632 21644 16865 21672
rect 16632 21632 16638 21644
rect 16853 21641 16865 21644
rect 16899 21641 16911 21675
rect 20530 21672 20536 21684
rect 16853 21635 16911 21641
rect 19628 21644 20536 21672
rect 2225 21607 2283 21613
rect 2225 21604 2237 21607
rect 1412 21576 2237 21604
rect 1412 21545 1440 21576
rect 2225 21573 2237 21576
rect 2271 21573 2283 21607
rect 2225 21567 2283 21573
rect 8012 21607 8070 21613
rect 8012 21573 8024 21607
rect 8058 21604 8070 21607
rect 8478 21604 8484 21616
rect 8058 21576 8484 21604
rect 8058 21573 8070 21576
rect 8012 21567 8070 21573
rect 8478 21564 8484 21576
rect 8536 21564 8542 21616
rect 9968 21576 11928 21604
rect 1397 21539 1455 21545
rect 1397 21505 1409 21539
rect 1443 21505 1455 21539
rect 2130 21536 2136 21548
rect 2091 21508 2136 21536
rect 1397 21499 1455 21505
rect 2130 21496 2136 21508
rect 2188 21496 2194 21548
rect 2314 21536 2320 21548
rect 2275 21508 2320 21536
rect 2314 21496 2320 21508
rect 2372 21496 2378 21548
rect 7282 21496 7288 21548
rect 7340 21536 7346 21548
rect 9968 21545 9996 21576
rect 7745 21539 7803 21545
rect 7745 21536 7757 21539
rect 7340 21508 7757 21536
rect 7340 21496 7346 21508
rect 7745 21505 7757 21508
rect 7791 21505 7803 21539
rect 7745 21499 7803 21505
rect 9953 21539 10011 21545
rect 9953 21505 9965 21539
rect 9999 21505 10011 21539
rect 9953 21499 10011 21505
rect 10321 21539 10379 21545
rect 10321 21505 10333 21539
rect 10367 21536 10379 21539
rect 10410 21536 10416 21548
rect 10367 21508 10416 21536
rect 10367 21505 10379 21508
rect 10321 21499 10379 21505
rect 10410 21496 10416 21508
rect 10468 21496 10474 21548
rect 11422 21496 11428 21548
rect 11480 21536 11486 21548
rect 11782 21539 11840 21545
rect 11782 21536 11794 21539
rect 11480 21508 11794 21536
rect 11480 21496 11486 21508
rect 11782 21505 11794 21508
rect 11828 21505 11840 21539
rect 11782 21499 11840 21505
rect 10045 21471 10103 21477
rect 10045 21437 10057 21471
rect 10091 21437 10103 21471
rect 11900 21468 11928 21576
rect 12986 21564 12992 21616
rect 13044 21604 13050 21616
rect 14645 21607 14703 21613
rect 14645 21604 14657 21607
rect 13044 21576 14657 21604
rect 13044 21564 13050 21576
rect 14645 21573 14657 21576
rect 14691 21573 14703 21607
rect 14826 21604 14832 21616
rect 14787 21576 14832 21604
rect 14645 21567 14703 21573
rect 14826 21564 14832 21576
rect 14884 21604 14890 21616
rect 14884 21576 15516 21604
rect 14884 21564 14890 21576
rect 13814 21496 13820 21548
rect 13872 21536 13878 21548
rect 15488 21545 15516 21576
rect 19426 21564 19432 21616
rect 19484 21604 19490 21616
rect 19628 21613 19656 21644
rect 20530 21632 20536 21644
rect 20588 21672 20594 21684
rect 21177 21675 21235 21681
rect 21177 21672 21189 21675
rect 20588 21644 21189 21672
rect 20588 21632 20594 21644
rect 21177 21641 21189 21644
rect 21223 21641 21235 21675
rect 21177 21635 21235 21641
rect 22002 21632 22008 21684
rect 22060 21632 22066 21684
rect 22462 21632 22468 21684
rect 22520 21672 22526 21684
rect 23382 21672 23388 21684
rect 22520 21644 23388 21672
rect 22520 21632 22526 21644
rect 23382 21632 23388 21644
rect 23440 21632 23446 21684
rect 24946 21632 24952 21684
rect 25004 21672 25010 21684
rect 25682 21672 25688 21684
rect 25004 21644 25688 21672
rect 25004 21632 25010 21644
rect 25682 21632 25688 21644
rect 25740 21672 25746 21684
rect 26237 21675 26295 21681
rect 26237 21672 26249 21675
rect 25740 21644 26249 21672
rect 25740 21632 25746 21644
rect 26237 21641 26249 21644
rect 26283 21641 26295 21675
rect 26237 21635 26295 21641
rect 19613 21607 19671 21613
rect 19613 21604 19625 21607
rect 19484 21576 19625 21604
rect 19484 21564 19490 21576
rect 19613 21573 19625 21576
rect 19659 21573 19671 21607
rect 19613 21567 19671 21573
rect 19797 21607 19855 21613
rect 19797 21573 19809 21607
rect 19843 21604 19855 21607
rect 19978 21604 19984 21616
rect 19843 21576 19984 21604
rect 19843 21573 19855 21576
rect 19797 21567 19855 21573
rect 19978 21564 19984 21576
rect 20036 21564 20042 21616
rect 20254 21604 20260 21616
rect 20215 21576 20260 21604
rect 20254 21564 20260 21576
rect 20312 21564 20318 21616
rect 20346 21564 20352 21616
rect 20404 21604 20410 21616
rect 20441 21607 20499 21613
rect 20441 21604 20453 21607
rect 20404 21576 20453 21604
rect 20404 21564 20410 21576
rect 20441 21573 20453 21576
rect 20487 21573 20499 21607
rect 20441 21567 20499 21573
rect 20625 21607 20683 21613
rect 20625 21573 20637 21607
rect 20671 21604 20683 21607
rect 21821 21607 21879 21613
rect 21821 21604 21833 21607
rect 20671 21576 21833 21604
rect 20671 21573 20683 21576
rect 20625 21567 20683 21573
rect 21821 21573 21833 21576
rect 21867 21604 21879 21607
rect 21910 21604 21916 21616
rect 21867 21576 21916 21604
rect 21867 21573 21879 21576
rect 21821 21567 21879 21573
rect 21910 21564 21916 21576
rect 21968 21564 21974 21616
rect 22020 21604 22048 21632
rect 26142 21604 26148 21616
rect 22020 21576 22692 21604
rect 14001 21539 14059 21545
rect 14001 21536 14013 21539
rect 13872 21508 14013 21536
rect 13872 21496 13878 21508
rect 14001 21505 14013 21508
rect 14047 21505 14059 21539
rect 14001 21499 14059 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21505 15531 21539
rect 15473 21499 15531 21505
rect 16298 21496 16304 21548
rect 16356 21536 16362 21548
rect 16669 21539 16727 21545
rect 16669 21536 16681 21539
rect 16356 21508 16681 21536
rect 16356 21496 16362 21508
rect 16669 21505 16681 21508
rect 16715 21505 16727 21539
rect 16669 21499 16727 21505
rect 17586 21496 17592 21548
rect 17644 21536 17650 21548
rect 17681 21539 17739 21545
rect 17681 21536 17693 21539
rect 17644 21508 17693 21536
rect 17644 21496 17650 21508
rect 17681 21505 17693 21508
rect 17727 21505 17739 21539
rect 17681 21499 17739 21505
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 17862 21536 17868 21548
rect 17819 21508 17868 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 17862 21496 17868 21508
rect 17920 21496 17926 21548
rect 17954 21496 17960 21548
rect 18012 21536 18018 21548
rect 18049 21539 18107 21545
rect 18049 21536 18061 21539
rect 18012 21508 18061 21536
rect 18012 21496 18018 21508
rect 18049 21505 18061 21508
rect 18095 21505 18107 21539
rect 18049 21499 18107 21505
rect 18598 21496 18604 21548
rect 18656 21536 18662 21548
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 18656 21508 18705 21536
rect 18656 21496 18662 21508
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 18782 21496 18788 21548
rect 18840 21536 18846 21548
rect 19061 21539 19119 21545
rect 18840 21508 18885 21536
rect 18840 21496 18846 21508
rect 19061 21505 19073 21539
rect 19107 21536 19119 21539
rect 19150 21536 19156 21548
rect 19107 21508 19156 21536
rect 19107 21505 19119 21508
rect 19061 21499 19119 21505
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 20162 21496 20168 21548
rect 20220 21536 20226 21548
rect 22664 21545 22692 21576
rect 25056 21576 26148 21604
rect 25056 21545 25084 21576
rect 26142 21564 26148 21576
rect 26200 21604 26206 21616
rect 27154 21604 27160 21616
rect 26200 21576 27160 21604
rect 26200 21564 26206 21576
rect 27154 21564 27160 21576
rect 27212 21564 27218 21616
rect 28166 21604 28172 21616
rect 27724 21576 28172 21604
rect 21085 21539 21143 21545
rect 21085 21536 21097 21539
rect 20220 21508 21097 21536
rect 20220 21496 20226 21508
rect 21085 21505 21097 21508
rect 21131 21505 21143 21539
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 21085 21499 21143 21505
rect 21928 21508 22017 21536
rect 12066 21468 12072 21480
rect 10045 21431 10103 21437
rect 11808 21440 11928 21468
rect 12027 21440 12072 21468
rect 9950 21400 9956 21412
rect 9911 21372 9956 21400
rect 9950 21360 9956 21372
rect 10008 21360 10014 21412
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 10060 21332 10088 21431
rect 10962 21360 10968 21412
rect 11020 21400 11026 21412
rect 11020 21372 11560 21400
rect 11020 21360 11026 21372
rect 11422 21332 11428 21344
rect 10060 21304 11428 21332
rect 11422 21292 11428 21304
rect 11480 21292 11486 21344
rect 11532 21332 11560 21372
rect 11698 21360 11704 21412
rect 11756 21400 11762 21412
rect 11808 21400 11836 21440
rect 12066 21428 12072 21440
rect 12124 21428 12130 21480
rect 12250 21428 12256 21480
rect 12308 21468 12314 21480
rect 18509 21471 18567 21477
rect 18509 21468 18521 21471
rect 12308 21440 18521 21468
rect 12308 21428 12314 21440
rect 18509 21437 18521 21440
rect 18555 21437 18567 21471
rect 18966 21468 18972 21480
rect 18927 21440 18972 21468
rect 18509 21431 18567 21437
rect 18966 21428 18972 21440
rect 19024 21428 19030 21480
rect 20714 21428 20720 21480
rect 20772 21468 20778 21480
rect 21928 21468 21956 21508
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21505 22707 21539
rect 22905 21539 22963 21545
rect 22905 21536 22917 21539
rect 22649 21499 22707 21505
rect 22756 21508 22917 21536
rect 22186 21468 22192 21480
rect 20772 21440 21956 21468
rect 22147 21440 22192 21468
rect 20772 21428 20778 21440
rect 22186 21428 22192 21440
rect 22244 21428 22250 21480
rect 22756 21468 22784 21508
rect 22905 21505 22917 21508
rect 22951 21505 22963 21539
rect 22905 21499 22963 21505
rect 25041 21539 25099 21545
rect 25041 21505 25053 21539
rect 25087 21505 25099 21539
rect 25041 21499 25099 21505
rect 27246 21496 27252 21548
rect 27304 21536 27310 21548
rect 27724 21545 27752 21576
rect 28166 21564 28172 21576
rect 28224 21564 28230 21616
rect 28261 21607 28319 21613
rect 28261 21573 28273 21607
rect 28307 21604 28319 21607
rect 28966 21607 29024 21613
rect 28966 21604 28978 21607
rect 28307 21576 28978 21604
rect 28307 21573 28319 21576
rect 28261 21567 28319 21573
rect 28966 21573 28978 21576
rect 29012 21573 29024 21607
rect 28966 21567 29024 21573
rect 27525 21539 27583 21545
rect 27525 21536 27537 21539
rect 27304 21508 27537 21536
rect 27304 21496 27310 21508
rect 27525 21505 27537 21508
rect 27571 21505 27583 21539
rect 27525 21499 27583 21505
rect 27709 21539 27767 21545
rect 27709 21505 27721 21539
rect 27755 21505 27767 21539
rect 27890 21536 27896 21548
rect 27851 21508 27896 21536
rect 27709 21499 27767 21505
rect 27890 21496 27896 21508
rect 27948 21496 27954 21548
rect 27982 21496 27988 21548
rect 28040 21536 28046 21548
rect 28077 21539 28135 21545
rect 28077 21536 28089 21539
rect 28040 21508 28089 21536
rect 28040 21496 28046 21508
rect 28077 21505 28089 21508
rect 28123 21536 28135 21539
rect 28123 21508 28396 21536
rect 28123 21505 28135 21508
rect 28077 21499 28135 21505
rect 24762 21468 24768 21480
rect 22664 21440 22784 21468
rect 24723 21440 24768 21468
rect 22664 21412 22692 21440
rect 24762 21428 24768 21440
rect 24820 21428 24826 21480
rect 27801 21471 27859 21477
rect 27801 21437 27813 21471
rect 27847 21468 27859 21471
rect 28166 21468 28172 21480
rect 27847 21440 28172 21468
rect 27847 21437 27859 21440
rect 27801 21431 27859 21437
rect 28166 21428 28172 21440
rect 28224 21428 28230 21480
rect 11756 21372 11836 21400
rect 11756 21360 11762 21372
rect 12986 21360 12992 21412
rect 13044 21400 13050 21412
rect 15565 21403 15623 21409
rect 15565 21400 15577 21403
rect 13044 21372 15577 21400
rect 13044 21360 13050 21372
rect 15565 21369 15577 21372
rect 15611 21400 15623 21403
rect 16850 21400 16856 21412
rect 15611 21372 16856 21400
rect 15611 21369 15623 21372
rect 15565 21363 15623 21369
rect 16850 21360 16856 21372
rect 16908 21360 16914 21412
rect 18138 21360 18144 21412
rect 18196 21400 18202 21412
rect 18196 21372 19748 21400
rect 18196 21360 18202 21372
rect 12710 21332 12716 21344
rect 11532 21304 12716 21332
rect 12710 21292 12716 21304
rect 12768 21292 12774 21344
rect 14093 21335 14151 21341
rect 14093 21301 14105 21335
rect 14139 21332 14151 21335
rect 14642 21332 14648 21344
rect 14139 21304 14648 21332
rect 14139 21301 14151 21304
rect 14093 21295 14151 21301
rect 14642 21292 14648 21304
rect 14700 21292 14706 21344
rect 14826 21292 14832 21344
rect 14884 21332 14890 21344
rect 14921 21335 14979 21341
rect 14921 21332 14933 21335
rect 14884 21304 14933 21332
rect 14884 21292 14890 21304
rect 14921 21301 14933 21304
rect 14967 21301 14979 21335
rect 14921 21295 14979 21301
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 17497 21335 17555 21341
rect 17497 21332 17509 21335
rect 16632 21304 17509 21332
rect 16632 21292 16638 21304
rect 17497 21301 17509 21304
rect 17543 21301 17555 21335
rect 17497 21295 17555 21301
rect 17957 21335 18015 21341
rect 17957 21301 17969 21335
rect 18003 21332 18015 21335
rect 19610 21332 19616 21344
rect 18003 21304 19616 21332
rect 18003 21301 18015 21304
rect 17957 21295 18015 21301
rect 19610 21292 19616 21304
rect 19668 21292 19674 21344
rect 19720 21332 19748 21372
rect 19794 21360 19800 21412
rect 19852 21400 19858 21412
rect 22094 21400 22100 21412
rect 19852 21372 22100 21400
rect 19852 21360 19858 21372
rect 22094 21360 22100 21372
rect 22152 21360 22158 21412
rect 22646 21360 22652 21412
rect 22704 21360 22710 21412
rect 21450 21332 21456 21344
rect 19720 21304 21456 21332
rect 21450 21292 21456 21304
rect 21508 21292 21514 21344
rect 21726 21292 21732 21344
rect 21784 21332 21790 21344
rect 24029 21335 24087 21341
rect 24029 21332 24041 21335
rect 21784 21304 24041 21332
rect 21784 21292 21790 21304
rect 24029 21301 24041 21304
rect 24075 21332 24087 21335
rect 24210 21332 24216 21344
rect 24075 21304 24216 21332
rect 24075 21301 24087 21304
rect 24029 21295 24087 21301
rect 24210 21292 24216 21304
rect 24268 21292 24274 21344
rect 28368 21332 28396 21508
rect 28442 21496 28448 21548
rect 28500 21536 28506 21548
rect 28721 21539 28779 21545
rect 28721 21536 28733 21539
rect 28500 21508 28733 21536
rect 28500 21496 28506 21508
rect 28721 21505 28733 21508
rect 28767 21505 28779 21539
rect 28721 21499 28779 21505
rect 30101 21335 30159 21341
rect 30101 21332 30113 21335
rect 28368 21304 30113 21332
rect 30101 21301 30113 21304
rect 30147 21301 30159 21335
rect 30101 21295 30159 21301
rect 1104 21242 30820 21264
rect 1104 21190 5915 21242
rect 5967 21190 5979 21242
rect 6031 21190 6043 21242
rect 6095 21190 6107 21242
rect 6159 21190 6171 21242
rect 6223 21190 15846 21242
rect 15898 21190 15910 21242
rect 15962 21190 15974 21242
rect 16026 21190 16038 21242
rect 16090 21190 16102 21242
rect 16154 21190 25776 21242
rect 25828 21190 25840 21242
rect 25892 21190 25904 21242
rect 25956 21190 25968 21242
rect 26020 21190 26032 21242
rect 26084 21190 30820 21242
rect 1104 21168 30820 21190
rect 10502 21088 10508 21140
rect 10560 21128 10566 21140
rect 12158 21128 12164 21140
rect 10560 21100 11836 21128
rect 12119 21100 12164 21128
rect 10560 21088 10566 21100
rect 2406 21020 2412 21072
rect 2464 21060 2470 21072
rect 11054 21060 11060 21072
rect 2464 21032 11060 21060
rect 2464 21020 2470 21032
rect 11054 21020 11060 21032
rect 11112 21020 11118 21072
rect 10318 20992 10324 21004
rect 8956 20964 10324 20992
rect 8956 20933 8984 20964
rect 10318 20952 10324 20964
rect 10376 20952 10382 21004
rect 11808 21001 11836 21100
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 13446 21128 13452 21140
rect 12268 21100 13452 21128
rect 11701 20995 11759 21001
rect 11701 20992 11713 20995
rect 11256 20964 11713 20992
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20893 8999 20927
rect 9950 20924 9956 20936
rect 9863 20896 9956 20924
rect 8941 20887 8999 20893
rect 9950 20884 9956 20896
rect 10008 20924 10014 20936
rect 10410 20924 10416 20936
rect 10008 20896 10416 20924
rect 10008 20884 10014 20896
rect 10410 20884 10416 20896
rect 10468 20884 10474 20936
rect 10594 20924 10600 20936
rect 10555 20896 10600 20924
rect 10594 20884 10600 20896
rect 10652 20884 10658 20936
rect 10686 20884 10692 20936
rect 10744 20924 10750 20936
rect 10781 20927 10839 20933
rect 10781 20924 10793 20927
rect 10744 20896 10793 20924
rect 10744 20884 10750 20896
rect 10781 20893 10793 20896
rect 10827 20893 10839 20927
rect 11256 20924 11284 20964
rect 11701 20961 11713 20964
rect 11747 20961 11759 20995
rect 11701 20955 11759 20961
rect 11793 20995 11851 21001
rect 11793 20961 11805 20995
rect 11839 20961 11851 20995
rect 12268 20992 12296 21100
rect 13446 21088 13452 21100
rect 13504 21088 13510 21140
rect 14182 21088 14188 21140
rect 14240 21128 14246 21140
rect 14369 21131 14427 21137
rect 14369 21128 14381 21131
rect 14240 21100 14381 21128
rect 14240 21088 14246 21100
rect 14369 21097 14381 21100
rect 14415 21097 14427 21131
rect 14369 21091 14427 21097
rect 14737 21131 14795 21137
rect 14737 21097 14749 21131
rect 14783 21128 14795 21131
rect 15286 21128 15292 21140
rect 14783 21100 15292 21128
rect 14783 21097 14795 21100
rect 14737 21091 14795 21097
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 16301 21131 16359 21137
rect 16301 21128 16313 21131
rect 15580 21100 16313 21128
rect 12526 21020 12532 21072
rect 12584 21060 12590 21072
rect 13722 21060 13728 21072
rect 12584 21032 13728 21060
rect 12584 21020 12590 21032
rect 13722 21020 13728 21032
rect 13780 21060 13786 21072
rect 15580 21060 15608 21100
rect 16301 21097 16313 21100
rect 16347 21097 16359 21131
rect 16301 21091 16359 21097
rect 17034 21088 17040 21140
rect 17092 21128 17098 21140
rect 22462 21128 22468 21140
rect 17092 21100 22468 21128
rect 17092 21088 17098 21100
rect 22462 21088 22468 21100
rect 22520 21088 22526 21140
rect 22646 21128 22652 21140
rect 22607 21100 22652 21128
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 23845 21131 23903 21137
rect 23845 21097 23857 21131
rect 23891 21128 23903 21131
rect 24394 21128 24400 21140
rect 23891 21100 24400 21128
rect 23891 21097 23903 21100
rect 23845 21091 23903 21097
rect 24394 21088 24400 21100
rect 24452 21088 24458 21140
rect 24578 21088 24584 21140
rect 24636 21128 24642 21140
rect 24762 21128 24768 21140
rect 24636 21100 24768 21128
rect 24636 21088 24642 21100
rect 24762 21088 24768 21100
rect 24820 21128 24826 21140
rect 24820 21100 25544 21128
rect 24820 21088 24826 21100
rect 13780 21032 15608 21060
rect 15657 21063 15715 21069
rect 13780 21020 13786 21032
rect 15657 21029 15669 21063
rect 15703 21060 15715 21063
rect 18230 21060 18236 21072
rect 15703 21032 18236 21060
rect 15703 21029 15715 21032
rect 15657 21023 15715 21029
rect 18230 21020 18236 21032
rect 18288 21020 18294 21072
rect 18782 21020 18788 21072
rect 18840 21060 18846 21072
rect 25225 21063 25283 21069
rect 25225 21060 25237 21063
rect 18840 21032 25237 21060
rect 18840 21020 18846 21032
rect 25225 21029 25237 21032
rect 25271 21029 25283 21063
rect 25225 21023 25283 21029
rect 15010 20992 15016 21004
rect 11793 20955 11851 20961
rect 11900 20964 12296 20992
rect 12406 20964 15016 20992
rect 10781 20887 10839 20893
rect 10888 20896 11284 20924
rect 11425 20905 11483 20911
rect 10318 20816 10324 20868
rect 10376 20856 10382 20868
rect 10888 20856 10916 20896
rect 11425 20871 11437 20905
rect 11471 20871 11483 20905
rect 11606 20884 11612 20936
rect 11664 20924 11670 20936
rect 11900 20924 11928 20964
rect 11664 20896 11928 20924
rect 11977 20927 12035 20933
rect 11664 20884 11670 20896
rect 11977 20893 11989 20927
rect 12023 20924 12035 20927
rect 12406 20924 12434 20964
rect 15010 20952 15016 20964
rect 15068 20952 15074 21004
rect 18046 20992 18052 21004
rect 15580 20964 18052 20992
rect 12710 20924 12716 20936
rect 12023 20896 12434 20924
rect 12671 20896 12716 20924
rect 12023 20893 12035 20896
rect 11977 20887 12035 20893
rect 12710 20884 12716 20896
rect 12768 20884 12774 20936
rect 14366 20924 14372 20936
rect 14327 20896 14372 20924
rect 14366 20884 14372 20896
rect 14424 20884 14430 20936
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20893 14519 20927
rect 14461 20887 14519 20893
rect 10376 20828 10916 20856
rect 10376 20816 10382 20828
rect 10962 20816 10968 20868
rect 11020 20856 11026 20868
rect 11425 20865 11483 20871
rect 11020 20828 11065 20856
rect 11020 20816 11026 20828
rect 9122 20788 9128 20800
rect 9083 20760 9128 20788
rect 9122 20748 9128 20760
rect 9180 20748 9186 20800
rect 10042 20788 10048 20800
rect 10003 20760 10048 20788
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 10134 20748 10140 20800
rect 10192 20788 10198 20800
rect 10410 20788 10416 20800
rect 10192 20760 10416 20788
rect 10192 20748 10198 20760
rect 10410 20748 10416 20760
rect 10468 20748 10474 20800
rect 10686 20748 10692 20800
rect 10744 20788 10750 20800
rect 10980 20788 11008 20816
rect 10744 20760 11008 20788
rect 11440 20788 11468 20865
rect 12894 20816 12900 20868
rect 12952 20856 12958 20868
rect 12989 20859 13047 20865
rect 12989 20856 13001 20859
rect 12952 20828 13001 20856
rect 12952 20816 12958 20828
rect 12989 20825 13001 20828
rect 13035 20856 13047 20859
rect 13446 20856 13452 20868
rect 13035 20828 13452 20856
rect 13035 20825 13047 20828
rect 12989 20819 13047 20825
rect 13446 20816 13452 20828
rect 13504 20816 13510 20868
rect 13906 20816 13912 20868
rect 13964 20856 13970 20868
rect 14476 20856 14504 20887
rect 15102 20884 15108 20936
rect 15160 20924 15166 20936
rect 15473 20927 15531 20933
rect 15473 20924 15485 20927
rect 15160 20896 15485 20924
rect 15160 20884 15166 20896
rect 15473 20893 15485 20896
rect 15519 20893 15531 20927
rect 15473 20887 15531 20893
rect 13964 20828 14504 20856
rect 15289 20859 15347 20865
rect 13964 20816 13970 20828
rect 15289 20825 15301 20859
rect 15335 20856 15347 20859
rect 15378 20856 15384 20868
rect 15335 20828 15384 20856
rect 15335 20825 15347 20828
rect 15289 20819 15347 20825
rect 15378 20816 15384 20828
rect 15436 20816 15442 20868
rect 15580 20788 15608 20964
rect 18046 20952 18052 20964
rect 18104 20952 18110 21004
rect 19978 20992 19984 21004
rect 18524 20964 19984 20992
rect 16301 20927 16359 20933
rect 16301 20893 16313 20927
rect 16347 20924 16359 20927
rect 16485 20927 16543 20933
rect 16485 20924 16497 20927
rect 16347 20896 16497 20924
rect 16347 20893 16359 20896
rect 16301 20887 16359 20893
rect 16485 20893 16497 20896
rect 16531 20924 16543 20927
rect 17129 20927 17187 20933
rect 17129 20924 17141 20927
rect 16531 20896 17141 20924
rect 16531 20893 16543 20896
rect 16485 20887 16543 20893
rect 17129 20893 17141 20896
rect 17175 20893 17187 20927
rect 17129 20887 17187 20893
rect 17405 20927 17463 20933
rect 17405 20893 17417 20927
rect 17451 20924 17463 20927
rect 17954 20924 17960 20936
rect 17451 20896 17960 20924
rect 17451 20893 17463 20896
rect 17405 20887 17463 20893
rect 17954 20884 17960 20896
rect 18012 20884 18018 20936
rect 18524 20933 18552 20964
rect 19978 20952 19984 20964
rect 20036 20952 20042 21004
rect 21542 20952 21548 21004
rect 21600 20992 21606 21004
rect 21600 20964 22048 20992
rect 21600 20952 21606 20964
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20893 18567 20927
rect 19426 20924 19432 20936
rect 19387 20896 19432 20924
rect 18509 20887 18567 20893
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 20714 20924 20720 20936
rect 20675 20896 20720 20924
rect 20714 20884 20720 20896
rect 20772 20884 20778 20936
rect 22020 20933 22048 20964
rect 22278 20952 22284 21004
rect 22336 20992 22342 21004
rect 23198 20992 23204 21004
rect 22336 20964 23204 20992
rect 22336 20952 22342 20964
rect 23198 20952 23204 20964
rect 23256 20952 23262 21004
rect 23477 20995 23535 21001
rect 23477 20961 23489 20995
rect 23523 20992 23535 20995
rect 23750 20992 23756 21004
rect 23523 20964 23756 20992
rect 23523 20961 23535 20964
rect 23477 20955 23535 20961
rect 23750 20952 23756 20964
rect 23808 20952 23814 21004
rect 24854 20992 24860 21004
rect 24815 20964 24860 20992
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 25516 20992 25544 21100
rect 27338 21020 27344 21072
rect 27396 21060 27402 21072
rect 29917 21063 29975 21069
rect 29917 21060 29929 21063
rect 27396 21032 29929 21060
rect 27396 21020 27402 21032
rect 29917 21029 29929 21032
rect 29963 21029 29975 21063
rect 29917 21023 29975 21029
rect 25685 20995 25743 21001
rect 25685 20992 25697 20995
rect 25056 20964 25452 20992
rect 25516 20964 25697 20992
rect 21361 20927 21419 20933
rect 21361 20893 21373 20927
rect 21407 20893 21419 20927
rect 21361 20887 21419 20893
rect 22005 20927 22063 20933
rect 22005 20893 22017 20927
rect 22051 20893 22063 20927
rect 22005 20887 22063 20893
rect 16666 20856 16672 20868
rect 16579 20828 16672 20856
rect 16666 20816 16672 20828
rect 16724 20856 16730 20868
rect 17218 20856 17224 20868
rect 16724 20828 17224 20856
rect 16724 20816 16730 20828
rect 17218 20816 17224 20828
rect 17276 20856 17282 20868
rect 18598 20856 18604 20868
rect 17276 20828 18604 20856
rect 17276 20816 17282 20828
rect 18598 20816 18604 20828
rect 18656 20816 18662 20868
rect 18693 20859 18751 20865
rect 18693 20825 18705 20859
rect 18739 20856 18751 20859
rect 18782 20856 18788 20868
rect 18739 20828 18788 20856
rect 18739 20825 18751 20828
rect 18693 20819 18751 20825
rect 18782 20816 18788 20828
rect 18840 20816 18846 20868
rect 20162 20856 20168 20868
rect 19306 20828 20168 20856
rect 11440 20760 15608 20788
rect 10744 20748 10750 20760
rect 18230 20748 18236 20800
rect 18288 20788 18294 20800
rect 19306 20788 19334 20828
rect 20162 20816 20168 20828
rect 20220 20816 20226 20868
rect 20533 20859 20591 20865
rect 20533 20825 20545 20859
rect 20579 20856 20591 20859
rect 20622 20856 20628 20868
rect 20579 20828 20628 20856
rect 20579 20825 20591 20828
rect 20533 20819 20591 20825
rect 20622 20816 20628 20828
rect 20680 20816 20686 20868
rect 20901 20859 20959 20865
rect 20901 20825 20913 20859
rect 20947 20856 20959 20859
rect 21376 20856 21404 20887
rect 22094 20884 22100 20936
rect 22152 20933 22158 20936
rect 22152 20927 22211 20933
rect 22152 20893 22165 20927
rect 22199 20924 22211 20927
rect 22296 20924 22324 20952
rect 22199 20896 22324 20924
rect 22199 20893 22211 20896
rect 22152 20887 22211 20893
rect 22152 20884 22158 20887
rect 22462 20884 22468 20936
rect 22520 20933 22526 20936
rect 22520 20924 22528 20933
rect 22520 20896 22565 20924
rect 22520 20887 22528 20896
rect 22520 20884 22526 20887
rect 22922 20884 22928 20936
rect 22980 20924 22986 20936
rect 23109 20927 23167 20933
rect 23109 20924 23121 20927
rect 22980 20896 23121 20924
rect 22980 20884 22986 20896
rect 23109 20893 23121 20896
rect 23155 20893 23167 20927
rect 23290 20924 23296 20936
rect 23251 20896 23296 20924
rect 23109 20887 23167 20893
rect 23290 20884 23296 20896
rect 23348 20884 23354 20936
rect 23385 20927 23443 20933
rect 23385 20893 23397 20927
rect 23431 20893 23443 20927
rect 23385 20887 23443 20893
rect 23661 20927 23719 20933
rect 23661 20893 23673 20927
rect 23707 20924 23719 20927
rect 24026 20924 24032 20936
rect 23707 20896 24032 20924
rect 23707 20893 23719 20896
rect 23661 20887 23719 20893
rect 20947 20828 21404 20856
rect 20947 20825 20959 20828
rect 20901 20819 20959 20825
rect 18288 20760 19334 20788
rect 19613 20791 19671 20797
rect 18288 20748 18294 20760
rect 19613 20757 19625 20791
rect 19659 20788 19671 20791
rect 20070 20788 20076 20800
rect 19659 20760 20076 20788
rect 19659 20757 19671 20760
rect 19613 20751 19671 20757
rect 20070 20748 20076 20760
rect 20128 20788 20134 20800
rect 20254 20788 20260 20800
rect 20128 20760 20260 20788
rect 20128 20748 20134 20760
rect 20254 20748 20260 20760
rect 20312 20748 20318 20800
rect 20438 20748 20444 20800
rect 20496 20788 20502 20800
rect 20916 20788 20944 20819
rect 21726 20816 21732 20868
rect 21784 20856 21790 20868
rect 22281 20859 22339 20865
rect 22281 20856 22293 20859
rect 21784 20828 22293 20856
rect 21784 20816 21790 20828
rect 22281 20825 22293 20828
rect 22327 20825 22339 20859
rect 22281 20819 22339 20825
rect 22373 20859 22431 20865
rect 22373 20825 22385 20859
rect 22419 20856 22431 20859
rect 22646 20856 22652 20868
rect 22419 20828 22652 20856
rect 22419 20825 22431 20828
rect 22373 20819 22431 20825
rect 22646 20816 22652 20828
rect 22704 20816 22710 20868
rect 22738 20816 22744 20868
rect 22796 20856 22802 20868
rect 23400 20856 23428 20887
rect 24026 20884 24032 20896
rect 24084 20884 24090 20936
rect 24394 20884 24400 20936
rect 24452 20924 24458 20936
rect 24489 20927 24547 20933
rect 24489 20924 24501 20927
rect 24452 20896 24501 20924
rect 24452 20884 24458 20896
rect 24489 20893 24501 20896
rect 24535 20893 24547 20927
rect 24489 20887 24547 20893
rect 24673 20927 24731 20933
rect 24673 20893 24685 20927
rect 24719 20893 24731 20927
rect 24673 20887 24731 20893
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20924 24823 20927
rect 24946 20924 24952 20936
rect 24811 20896 24952 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 22796 20828 23428 20856
rect 22796 20816 22802 20828
rect 20496 20760 20944 20788
rect 20496 20748 20502 20760
rect 21174 20748 21180 20800
rect 21232 20788 21238 20800
rect 21453 20791 21511 20797
rect 21453 20788 21465 20791
rect 21232 20760 21465 20788
rect 21232 20748 21238 20760
rect 21453 20757 21465 20760
rect 21499 20757 21511 20791
rect 21453 20751 21511 20757
rect 22186 20748 22192 20800
rect 22244 20788 22250 20800
rect 22922 20788 22928 20800
rect 22244 20760 22928 20788
rect 22244 20748 22250 20760
rect 22922 20748 22928 20760
rect 22980 20748 22986 20800
rect 24688 20788 24716 20887
rect 24946 20884 24952 20896
rect 25004 20884 25010 20936
rect 25056 20933 25084 20964
rect 25041 20927 25099 20933
rect 25041 20893 25053 20927
rect 25087 20893 25099 20927
rect 25041 20887 25099 20893
rect 25130 20884 25136 20936
rect 25188 20924 25194 20936
rect 25314 20924 25320 20936
rect 25188 20896 25320 20924
rect 25188 20884 25194 20896
rect 25314 20884 25320 20896
rect 25372 20884 25378 20936
rect 25130 20788 25136 20800
rect 24688 20760 25136 20788
rect 25130 20748 25136 20760
rect 25188 20748 25194 20800
rect 25424 20788 25452 20964
rect 25685 20961 25697 20964
rect 25731 20961 25743 20995
rect 25958 20992 25964 21004
rect 25871 20964 25964 20992
rect 25685 20955 25743 20961
rect 25958 20952 25964 20964
rect 26016 20992 26022 21004
rect 26786 20992 26792 21004
rect 26016 20964 26792 20992
rect 26016 20952 26022 20964
rect 26786 20952 26792 20964
rect 26844 20952 26850 21004
rect 27798 20952 27804 21004
rect 27856 20992 27862 21004
rect 27985 20995 28043 21001
rect 27985 20992 27997 20995
rect 27856 20964 27997 20992
rect 27856 20952 27862 20964
rect 27985 20961 27997 20964
rect 28031 20961 28043 20995
rect 27985 20955 28043 20961
rect 27341 20927 27399 20933
rect 27341 20893 27353 20927
rect 27387 20924 27399 20927
rect 27614 20924 27620 20936
rect 27387 20896 27620 20924
rect 27387 20893 27399 20896
rect 27341 20887 27399 20893
rect 27614 20884 27620 20896
rect 27672 20884 27678 20936
rect 28166 20884 28172 20936
rect 28224 20924 28230 20936
rect 28261 20927 28319 20933
rect 28261 20924 28273 20927
rect 28224 20896 28273 20924
rect 28224 20884 28230 20896
rect 28261 20893 28273 20896
rect 28307 20924 28319 20927
rect 28350 20924 28356 20936
rect 28307 20896 28356 20924
rect 28307 20893 28319 20896
rect 28261 20887 28319 20893
rect 28350 20884 28356 20896
rect 28408 20884 28414 20936
rect 29086 20884 29092 20936
rect 29144 20924 29150 20936
rect 30101 20927 30159 20933
rect 30101 20924 30113 20927
rect 29144 20896 30113 20924
rect 29144 20884 29150 20896
rect 30101 20893 30113 20896
rect 30147 20893 30159 20927
rect 30101 20887 30159 20893
rect 26326 20788 26332 20800
rect 25424 20760 26332 20788
rect 26326 20748 26332 20760
rect 26384 20748 26390 20800
rect 27430 20788 27436 20800
rect 27391 20760 27436 20788
rect 27430 20748 27436 20760
rect 27488 20748 27494 20800
rect 1104 20698 30820 20720
rect 1104 20646 10880 20698
rect 10932 20646 10944 20698
rect 10996 20646 11008 20698
rect 11060 20646 11072 20698
rect 11124 20646 11136 20698
rect 11188 20646 20811 20698
rect 20863 20646 20875 20698
rect 20927 20646 20939 20698
rect 20991 20646 21003 20698
rect 21055 20646 21067 20698
rect 21119 20646 30820 20698
rect 1104 20624 30820 20646
rect 8849 20587 8907 20593
rect 8849 20553 8861 20587
rect 8895 20584 8907 20587
rect 9674 20584 9680 20596
rect 8895 20556 9680 20584
rect 8895 20553 8907 20556
rect 8849 20547 8907 20553
rect 9674 20544 9680 20556
rect 9732 20584 9738 20596
rect 12710 20584 12716 20596
rect 9732 20556 12716 20584
rect 9732 20544 9738 20556
rect 12710 20544 12716 20556
rect 12768 20544 12774 20596
rect 12989 20587 13047 20593
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 13814 20584 13820 20596
rect 13035 20556 13820 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 13814 20544 13820 20556
rect 13872 20544 13878 20596
rect 14090 20544 14096 20596
rect 14148 20584 14154 20596
rect 14148 20556 15700 20584
rect 14148 20544 14154 20556
rect 9493 20519 9551 20525
rect 9493 20485 9505 20519
rect 9539 20516 9551 20519
rect 9950 20516 9956 20528
rect 9539 20488 9956 20516
rect 9539 20485 9551 20488
rect 9493 20479 9551 20485
rect 9950 20476 9956 20488
rect 10008 20476 10014 20528
rect 10042 20476 10048 20528
rect 10100 20516 10106 20528
rect 10229 20519 10287 20525
rect 10229 20516 10241 20519
rect 10100 20488 10241 20516
rect 10100 20476 10106 20488
rect 10229 20485 10241 20488
rect 10275 20485 10287 20519
rect 10229 20479 10287 20485
rect 10413 20519 10471 20525
rect 10413 20485 10425 20519
rect 10459 20516 10471 20519
rect 10502 20516 10508 20528
rect 10459 20488 10508 20516
rect 10459 20485 10471 20488
rect 10413 20479 10471 20485
rect 10502 20476 10508 20488
rect 10560 20476 10566 20528
rect 11606 20476 11612 20528
rect 11664 20516 11670 20528
rect 11701 20519 11759 20525
rect 11701 20516 11713 20519
rect 11664 20488 11713 20516
rect 11664 20476 11670 20488
rect 11701 20485 11713 20488
rect 11747 20485 11759 20519
rect 11701 20479 11759 20485
rect 11790 20476 11796 20528
rect 11848 20516 11854 20528
rect 11885 20519 11943 20525
rect 11885 20516 11897 20519
rect 11848 20488 11897 20516
rect 11848 20476 11854 20488
rect 11885 20485 11897 20488
rect 11931 20485 11943 20519
rect 11885 20479 11943 20485
rect 12069 20519 12127 20525
rect 12069 20485 12081 20519
rect 12115 20516 12127 20519
rect 12434 20516 12440 20528
rect 12115 20488 12440 20516
rect 12115 20485 12127 20488
rect 12069 20479 12127 20485
rect 12434 20476 12440 20488
rect 12492 20476 12498 20528
rect 12529 20519 12587 20525
rect 12529 20485 12541 20519
rect 12575 20516 12587 20519
rect 12805 20519 12863 20525
rect 12805 20516 12817 20519
rect 12575 20488 12817 20516
rect 12575 20485 12587 20488
rect 12529 20479 12587 20485
rect 12805 20485 12817 20488
rect 12851 20516 12863 20519
rect 15010 20516 15016 20528
rect 12851 20488 14412 20516
rect 14971 20488 15016 20516
rect 12851 20485 12863 20488
rect 12805 20479 12863 20485
rect 8386 20408 8392 20460
rect 8444 20448 8450 20460
rect 8665 20451 8723 20457
rect 8665 20448 8677 20451
rect 8444 20420 8677 20448
rect 8444 20408 8450 20420
rect 8665 20417 8677 20420
rect 8711 20448 8723 20451
rect 9122 20448 9128 20460
rect 8711 20420 9128 20448
rect 8711 20417 8723 20420
rect 8665 20411 8723 20417
rect 9122 20408 9128 20420
rect 9180 20408 9186 20460
rect 12158 20408 12164 20460
rect 12216 20448 12222 20460
rect 12621 20451 12679 20457
rect 12621 20448 12633 20451
rect 12216 20420 12633 20448
rect 12216 20408 12222 20420
rect 12621 20417 12633 20420
rect 12667 20417 12679 20451
rect 13814 20448 13820 20460
rect 13775 20420 13820 20448
rect 12621 20411 12679 20417
rect 13814 20408 13820 20420
rect 13872 20408 13878 20460
rect 14182 20448 14188 20460
rect 14143 20420 14188 20448
rect 14182 20408 14188 20420
rect 14240 20408 14246 20460
rect 14384 20457 14412 20488
rect 15010 20476 15016 20488
rect 15068 20476 15074 20528
rect 15672 20525 15700 20556
rect 19518 20544 19524 20596
rect 19576 20584 19582 20596
rect 19705 20587 19763 20593
rect 19705 20584 19717 20587
rect 19576 20556 19717 20584
rect 19576 20544 19582 20556
rect 19705 20553 19717 20556
rect 19751 20584 19763 20587
rect 19794 20584 19800 20596
rect 19751 20556 19800 20584
rect 19751 20553 19763 20556
rect 19705 20547 19763 20553
rect 19794 20544 19800 20556
rect 19852 20544 19858 20596
rect 20162 20544 20168 20596
rect 20220 20584 20226 20596
rect 24762 20584 24768 20596
rect 20220 20556 24768 20584
rect 20220 20544 20226 20556
rect 24762 20544 24768 20556
rect 24820 20544 24826 20596
rect 25222 20584 25228 20596
rect 25183 20556 25228 20584
rect 25222 20544 25228 20556
rect 25280 20544 25286 20596
rect 26142 20584 26148 20596
rect 25608 20556 26148 20584
rect 15657 20519 15715 20525
rect 15657 20485 15669 20519
rect 15703 20485 15715 20519
rect 15657 20479 15715 20485
rect 17129 20519 17187 20525
rect 17129 20485 17141 20519
rect 17175 20516 17187 20519
rect 20070 20516 20076 20528
rect 17175 20488 20076 20516
rect 17175 20485 17187 20488
rect 17129 20479 17187 20485
rect 20070 20476 20076 20488
rect 20128 20476 20134 20528
rect 20438 20476 20444 20528
rect 20496 20516 20502 20528
rect 21174 20516 21180 20528
rect 20496 20488 20852 20516
rect 20496 20476 20502 20488
rect 14369 20451 14427 20457
rect 14369 20417 14381 20451
rect 14415 20417 14427 20451
rect 14369 20411 14427 20417
rect 14550 20408 14556 20460
rect 14608 20448 14614 20460
rect 14737 20451 14795 20457
rect 14737 20448 14749 20451
rect 14608 20420 14749 20448
rect 14608 20408 14614 20420
rect 14737 20417 14749 20420
rect 14783 20417 14795 20451
rect 15470 20448 15476 20460
rect 15431 20420 15476 20448
rect 14737 20411 14795 20417
rect 15470 20408 15476 20420
rect 15528 20408 15534 20460
rect 17034 20448 17040 20460
rect 16995 20420 17040 20448
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 18322 20448 18328 20460
rect 18283 20420 18328 20448
rect 18322 20408 18328 20420
rect 18380 20408 18386 20460
rect 18592 20451 18650 20457
rect 18592 20417 18604 20451
rect 18638 20448 18650 20451
rect 19978 20448 19984 20460
rect 18638 20420 19984 20448
rect 18638 20417 18650 20420
rect 18592 20411 18650 20417
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20448 20591 20451
rect 20622 20448 20628 20460
rect 20579 20420 20628 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 20622 20408 20628 20420
rect 20680 20408 20686 20460
rect 20824 20457 20852 20488
rect 20916 20488 21180 20516
rect 20916 20457 20944 20488
rect 21174 20476 21180 20488
rect 21232 20476 21238 20528
rect 21266 20476 21272 20528
rect 21324 20516 21330 20528
rect 21324 20488 21369 20516
rect 21324 20476 21330 20488
rect 21910 20476 21916 20528
rect 21968 20516 21974 20528
rect 23109 20519 23167 20525
rect 23109 20516 23121 20519
rect 21968 20488 23121 20516
rect 21968 20476 21974 20488
rect 23109 20485 23121 20488
rect 23155 20485 23167 20519
rect 23109 20479 23167 20485
rect 20717 20451 20775 20457
rect 20717 20417 20729 20451
rect 20763 20417 20775 20451
rect 20717 20411 20775 20417
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 20901 20451 20959 20457
rect 20901 20417 20913 20451
rect 20947 20417 20959 20451
rect 20901 20411 20959 20417
rect 21068 20451 21126 20457
rect 21068 20417 21080 20451
rect 21114 20448 21126 20451
rect 21821 20451 21879 20457
rect 21114 20417 21128 20448
rect 21068 20411 21128 20417
rect 21821 20417 21833 20451
rect 21867 20417 21879 20451
rect 21821 20411 21879 20417
rect 22005 20451 22063 20457
rect 22005 20417 22017 20451
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 1578 20340 1584 20392
rect 1636 20380 1642 20392
rect 16574 20380 16580 20392
rect 1636 20352 16580 20380
rect 1636 20340 1642 20352
rect 16574 20340 16580 20352
rect 16632 20340 16638 20392
rect 16850 20340 16856 20392
rect 16908 20380 16914 20392
rect 17221 20383 17279 20389
rect 17221 20380 17233 20383
rect 16908 20352 17233 20380
rect 16908 20340 16914 20352
rect 17221 20349 17233 20352
rect 17267 20349 17279 20383
rect 17221 20343 17279 20349
rect 20070 20340 20076 20392
rect 20128 20380 20134 20392
rect 20438 20380 20444 20392
rect 20128 20352 20444 20380
rect 20128 20340 20134 20352
rect 20438 20340 20444 20352
rect 20496 20340 20502 20392
rect 9122 20272 9128 20324
rect 9180 20312 9186 20324
rect 9180 20284 10456 20312
rect 9180 20272 9186 20284
rect 9585 20247 9643 20253
rect 9585 20213 9597 20247
rect 9631 20244 9643 20247
rect 9950 20244 9956 20256
rect 9631 20216 9956 20244
rect 9631 20213 9643 20216
rect 9585 20207 9643 20213
rect 9950 20204 9956 20216
rect 10008 20244 10014 20256
rect 10318 20244 10324 20256
rect 10008 20216 10324 20244
rect 10008 20204 10014 20216
rect 10318 20204 10324 20216
rect 10376 20204 10382 20256
rect 10428 20244 10456 20284
rect 11238 20272 11244 20324
rect 11296 20312 11302 20324
rect 11698 20312 11704 20324
rect 11296 20284 11704 20312
rect 11296 20272 11302 20284
rect 11698 20272 11704 20284
rect 11756 20272 11762 20324
rect 12342 20272 12348 20324
rect 12400 20312 12406 20324
rect 12529 20315 12587 20321
rect 12529 20312 12541 20315
rect 12400 20284 12541 20312
rect 12400 20272 12406 20284
rect 12529 20281 12541 20284
rect 12575 20281 12587 20315
rect 12529 20275 12587 20281
rect 15841 20315 15899 20321
rect 15841 20281 15853 20315
rect 15887 20312 15899 20315
rect 17402 20312 17408 20324
rect 15887 20284 17408 20312
rect 15887 20281 15899 20284
rect 15841 20275 15899 20281
rect 17402 20272 17408 20284
rect 17460 20272 17466 20324
rect 19426 20272 19432 20324
rect 19484 20312 19490 20324
rect 20162 20312 20168 20324
rect 19484 20284 20168 20312
rect 19484 20272 19490 20284
rect 20162 20272 20168 20284
rect 20220 20272 20226 20324
rect 16482 20244 16488 20256
rect 10428 20216 16488 20244
rect 16482 20204 16488 20216
rect 16540 20204 16546 20256
rect 16666 20244 16672 20256
rect 16627 20216 16672 20244
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 17126 20204 17132 20256
rect 17184 20244 17190 20256
rect 19518 20244 19524 20256
rect 17184 20216 19524 20244
rect 17184 20204 17190 20216
rect 19518 20204 19524 20216
rect 19576 20204 19582 20256
rect 20732 20244 20760 20411
rect 21100 20380 21128 20411
rect 21450 20380 21456 20392
rect 21100 20352 21456 20380
rect 21450 20340 21456 20352
rect 21508 20340 21514 20392
rect 21836 20380 21864 20411
rect 21910 20380 21916 20392
rect 21836 20352 21916 20380
rect 21910 20340 21916 20352
rect 21968 20340 21974 20392
rect 21634 20244 21640 20256
rect 20732 20216 21640 20244
rect 21634 20204 21640 20216
rect 21692 20244 21698 20256
rect 22020 20244 22048 20411
rect 22094 20408 22100 20460
rect 22152 20448 22158 20460
rect 22152 20420 22197 20448
rect 22152 20408 22158 20420
rect 22278 20408 22284 20460
rect 22336 20448 22342 20460
rect 22373 20451 22431 20457
rect 22373 20448 22385 20451
rect 22336 20420 22385 20448
rect 22336 20408 22342 20420
rect 22373 20417 22385 20420
rect 22419 20448 22431 20451
rect 23014 20448 23020 20460
rect 22419 20420 23020 20448
rect 22419 20417 22431 20420
rect 22373 20411 22431 20417
rect 23014 20408 23020 20420
rect 23072 20408 23078 20460
rect 23198 20408 23204 20460
rect 23256 20448 23262 20460
rect 23753 20451 23811 20457
rect 23753 20448 23765 20451
rect 23256 20420 23765 20448
rect 23256 20408 23262 20420
rect 23753 20417 23765 20420
rect 23799 20417 23811 20451
rect 23753 20411 23811 20417
rect 24489 20451 24547 20457
rect 24489 20417 24501 20451
rect 24535 20417 24547 20451
rect 24670 20448 24676 20460
rect 24631 20420 24676 20448
rect 24489 20411 24547 20417
rect 22189 20383 22247 20389
rect 22189 20349 22201 20383
rect 22235 20380 22247 20383
rect 22462 20380 22468 20392
rect 22235 20352 22468 20380
rect 22235 20349 22247 20352
rect 22189 20343 22247 20349
rect 22462 20340 22468 20352
rect 22520 20380 22526 20392
rect 23845 20383 23903 20389
rect 23845 20380 23857 20383
rect 22520 20352 23857 20380
rect 22520 20340 22526 20352
rect 23845 20349 23857 20352
rect 23891 20349 23903 20383
rect 24504 20380 24532 20411
rect 24670 20408 24676 20420
rect 24728 20408 24734 20460
rect 24762 20408 24768 20460
rect 24820 20448 24826 20460
rect 25038 20448 25044 20460
rect 24820 20420 24865 20448
rect 24999 20420 25044 20448
rect 24820 20408 24826 20420
rect 25038 20408 25044 20420
rect 25096 20408 25102 20460
rect 25608 20448 25636 20556
rect 26142 20544 26148 20556
rect 26200 20544 26206 20596
rect 26234 20544 26240 20596
rect 26292 20584 26298 20596
rect 26421 20587 26479 20593
rect 26421 20584 26433 20587
rect 26292 20556 26433 20584
rect 26292 20544 26298 20556
rect 26421 20553 26433 20556
rect 26467 20553 26479 20587
rect 26421 20547 26479 20553
rect 27614 20544 27620 20596
rect 27672 20584 27678 20596
rect 30101 20587 30159 20593
rect 30101 20584 30113 20587
rect 27672 20556 30113 20584
rect 27672 20544 27678 20556
rect 27430 20516 27436 20528
rect 25884 20488 27436 20516
rect 25884 20457 25912 20488
rect 27430 20476 27436 20488
rect 27488 20476 27494 20528
rect 25516 20420 25636 20448
rect 25685 20451 25743 20457
rect 24578 20380 24584 20392
rect 24504 20352 24584 20380
rect 23845 20343 23903 20349
rect 24578 20340 24584 20352
rect 24636 20340 24642 20392
rect 24857 20383 24915 20389
rect 24857 20349 24869 20383
rect 24903 20380 24915 20383
rect 25516 20380 25544 20420
rect 25685 20417 25697 20451
rect 25731 20417 25743 20451
rect 25685 20411 25743 20417
rect 25869 20451 25927 20457
rect 25869 20417 25881 20451
rect 25915 20417 25927 20451
rect 26234 20448 26240 20460
rect 26195 20420 26240 20448
rect 25869 20411 25927 20417
rect 24903 20352 25544 20380
rect 25700 20380 25728 20411
rect 26234 20408 26240 20420
rect 26292 20408 26298 20460
rect 27246 20408 27252 20460
rect 27304 20448 27310 20460
rect 27525 20451 27583 20457
rect 27525 20448 27537 20451
rect 27304 20420 27537 20448
rect 27304 20408 27310 20420
rect 27525 20417 27537 20420
rect 27571 20417 27583 20451
rect 27525 20411 27583 20417
rect 27713 20449 27771 20455
rect 27713 20415 27725 20449
rect 27759 20415 27771 20449
rect 27890 20448 27896 20460
rect 27851 20420 27896 20448
rect 25958 20380 25964 20392
rect 25700 20352 25820 20380
rect 25919 20352 25964 20380
rect 24903 20349 24915 20352
rect 24857 20343 24915 20349
rect 22554 20312 22560 20324
rect 22515 20284 22560 20312
rect 22554 20272 22560 20284
rect 22612 20272 22618 20324
rect 22738 20272 22744 20324
rect 22796 20312 22802 20324
rect 23293 20315 23351 20321
rect 23293 20312 23305 20315
rect 22796 20284 23305 20312
rect 22796 20272 22802 20284
rect 23293 20281 23305 20284
rect 23339 20281 23351 20315
rect 23293 20275 23351 20281
rect 21692 20216 22048 20244
rect 21692 20204 21698 20216
rect 22830 20204 22836 20256
rect 22888 20244 22894 20256
rect 23750 20244 23756 20256
rect 22888 20216 23756 20244
rect 22888 20204 22894 20216
rect 23750 20204 23756 20216
rect 23808 20204 23814 20256
rect 25792 20244 25820 20352
rect 25958 20340 25964 20352
rect 26016 20340 26022 20392
rect 26053 20383 26111 20389
rect 26053 20349 26065 20383
rect 26099 20380 26111 20383
rect 26142 20380 26148 20392
rect 26099 20352 26148 20380
rect 26099 20349 26111 20352
rect 26053 20343 26111 20349
rect 26142 20340 26148 20352
rect 26200 20340 26206 20392
rect 27540 20256 27568 20411
rect 27713 20409 27771 20415
rect 27715 20324 27743 20409
rect 27890 20408 27896 20420
rect 27948 20408 27954 20460
rect 28092 20457 28120 20556
rect 30101 20553 30113 20556
rect 30147 20553 30159 20587
rect 30101 20547 30159 20553
rect 28261 20519 28319 20525
rect 28261 20485 28273 20519
rect 28307 20516 28319 20519
rect 28966 20519 29024 20525
rect 28966 20516 28978 20519
rect 28307 20488 28978 20516
rect 28307 20485 28319 20488
rect 28261 20479 28319 20485
rect 28966 20485 28978 20488
rect 29012 20485 29024 20519
rect 28966 20479 29024 20485
rect 28077 20451 28135 20457
rect 28077 20417 28089 20451
rect 28123 20417 28135 20451
rect 28077 20411 28135 20417
rect 28442 20408 28448 20460
rect 28500 20448 28506 20460
rect 28721 20451 28779 20457
rect 28721 20448 28733 20451
rect 28500 20420 28733 20448
rect 28500 20408 28506 20420
rect 28721 20417 28733 20420
rect 28767 20417 28779 20451
rect 28721 20411 28779 20417
rect 27801 20383 27859 20389
rect 27801 20349 27813 20383
rect 27847 20380 27859 20383
rect 28166 20380 28172 20392
rect 27847 20352 28172 20380
rect 27847 20349 27859 20352
rect 27801 20343 27859 20349
rect 28166 20340 28172 20352
rect 28224 20340 28230 20392
rect 27706 20272 27712 20324
rect 27764 20272 27770 20324
rect 26602 20244 26608 20256
rect 25792 20216 26608 20244
rect 26602 20204 26608 20216
rect 26660 20204 26666 20256
rect 27522 20204 27528 20256
rect 27580 20204 27586 20256
rect 1104 20154 30820 20176
rect 1104 20102 5915 20154
rect 5967 20102 5979 20154
rect 6031 20102 6043 20154
rect 6095 20102 6107 20154
rect 6159 20102 6171 20154
rect 6223 20102 15846 20154
rect 15898 20102 15910 20154
rect 15962 20102 15974 20154
rect 16026 20102 16038 20154
rect 16090 20102 16102 20154
rect 16154 20102 25776 20154
rect 25828 20102 25840 20154
rect 25892 20102 25904 20154
rect 25956 20102 25968 20154
rect 26020 20102 26032 20154
rect 26084 20102 30820 20154
rect 1104 20080 30820 20102
rect 11701 20043 11759 20049
rect 11701 20009 11713 20043
rect 11747 20040 11759 20043
rect 11793 20043 11851 20049
rect 11793 20040 11805 20043
rect 11747 20012 11805 20040
rect 11747 20009 11759 20012
rect 11701 20003 11759 20009
rect 11793 20009 11805 20012
rect 11839 20009 11851 20043
rect 12158 20040 12164 20052
rect 12119 20012 12164 20040
rect 11793 20003 11851 20009
rect 11808 19972 11836 20003
rect 12158 20000 12164 20012
rect 12216 20000 12222 20052
rect 13357 20043 13415 20049
rect 13357 20009 13369 20043
rect 13403 20040 13415 20043
rect 13538 20040 13544 20052
rect 13403 20012 13544 20040
rect 13403 20009 13415 20012
rect 13357 20003 13415 20009
rect 13538 20000 13544 20012
rect 13596 20040 13602 20052
rect 14090 20040 14096 20052
rect 13596 20012 14096 20040
rect 13596 20000 13602 20012
rect 14090 20000 14096 20012
rect 14148 20000 14154 20052
rect 14185 20043 14243 20049
rect 14185 20009 14197 20043
rect 14231 20009 14243 20043
rect 14185 20003 14243 20009
rect 14553 20043 14611 20049
rect 14553 20009 14565 20043
rect 14599 20040 14611 20043
rect 15470 20040 15476 20052
rect 14599 20012 15476 20040
rect 14599 20009 14611 20012
rect 14553 20003 14611 20009
rect 14200 19972 14228 20003
rect 15470 20000 15476 20012
rect 15528 20000 15534 20052
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 17310 20040 17316 20052
rect 16632 20012 17316 20040
rect 16632 20000 16638 20012
rect 17310 20000 17316 20012
rect 17368 20000 17374 20052
rect 17402 20000 17408 20052
rect 17460 20040 17466 20052
rect 19426 20040 19432 20052
rect 17460 20012 19432 20040
rect 17460 20000 17466 20012
rect 19426 20000 19432 20012
rect 19484 20000 19490 20052
rect 19978 20040 19984 20052
rect 19939 20012 19984 20040
rect 19978 20000 19984 20012
rect 20036 20000 20042 20052
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 23106 20040 23112 20052
rect 20680 20012 23112 20040
rect 20680 20000 20686 20012
rect 23106 20000 23112 20012
rect 23164 20000 23170 20052
rect 23382 20000 23388 20052
rect 23440 20040 23446 20052
rect 25777 20043 25835 20049
rect 25777 20040 25789 20043
rect 23440 20012 25789 20040
rect 23440 20000 23446 20012
rect 14918 19972 14924 19984
rect 11808 19944 14924 19972
rect 14918 19932 14924 19944
rect 14976 19932 14982 19984
rect 16666 19972 16672 19984
rect 15488 19944 16672 19972
rect 10778 19864 10784 19916
rect 10836 19904 10842 19916
rect 11885 19907 11943 19913
rect 11885 19904 11897 19907
rect 10836 19876 11897 19904
rect 10836 19864 10842 19876
rect 11885 19873 11897 19876
rect 11931 19904 11943 19907
rect 13814 19904 13820 19916
rect 11931 19876 13820 19904
rect 11931 19873 11943 19876
rect 11885 19867 11943 19873
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 14090 19864 14096 19916
rect 14148 19904 14154 19916
rect 15488 19913 15516 19944
rect 16666 19932 16672 19944
rect 16724 19932 16730 19984
rect 22278 19972 22284 19984
rect 19444 19944 22284 19972
rect 14185 19907 14243 19913
rect 14185 19904 14197 19907
rect 14148 19876 14197 19904
rect 14148 19864 14154 19876
rect 14185 19873 14197 19876
rect 14231 19873 14243 19907
rect 14185 19867 14243 19873
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 15562 19864 15568 19916
rect 15620 19904 15626 19916
rect 16298 19904 16304 19916
rect 15620 19876 16304 19904
rect 15620 19864 15626 19876
rect 16298 19864 16304 19876
rect 16356 19864 16362 19916
rect 16853 19907 16911 19913
rect 16853 19873 16865 19907
rect 16899 19904 16911 19907
rect 17494 19904 17500 19916
rect 16899 19876 17500 19904
rect 16899 19873 16911 19876
rect 16853 19867 16911 19873
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 17865 19907 17923 19913
rect 17865 19873 17877 19907
rect 17911 19904 17923 19907
rect 19150 19904 19156 19916
rect 17911 19876 19156 19904
rect 17911 19873 17923 19876
rect 17865 19867 17923 19873
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 1578 19836 1584 19848
rect 1539 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 2314 19836 2320 19848
rect 1820 19808 2320 19836
rect 1820 19796 1826 19808
rect 2314 19796 2320 19808
rect 2372 19796 2378 19848
rect 8941 19839 8999 19845
rect 8941 19805 8953 19839
rect 8987 19836 8999 19839
rect 11793 19839 11851 19845
rect 8987 19808 9352 19836
rect 8987 19805 8999 19808
rect 8941 19799 8999 19805
rect 9324 19780 9352 19808
rect 11793 19805 11805 19839
rect 11839 19805 11851 19839
rect 11793 19799 11851 19805
rect 9214 19777 9220 19780
rect 9208 19768 9220 19777
rect 9175 19740 9220 19768
rect 9208 19731 9220 19740
rect 9214 19728 9220 19731
rect 9272 19728 9278 19780
rect 9306 19728 9312 19780
rect 9364 19728 9370 19780
rect 11808 19768 11836 19799
rect 12342 19796 12348 19848
rect 12400 19836 12406 19848
rect 13173 19839 13231 19845
rect 13173 19836 13185 19839
rect 12400 19808 13185 19836
rect 12400 19796 12406 19808
rect 13173 19805 13185 19808
rect 13219 19805 13231 19839
rect 13354 19836 13360 19848
rect 13315 19808 13360 19836
rect 13173 19799 13231 19805
rect 12434 19768 12440 19780
rect 11808 19740 12440 19768
rect 12434 19728 12440 19740
rect 12492 19768 12498 19780
rect 13078 19768 13084 19780
rect 12492 19740 13084 19768
rect 12492 19728 12498 19740
rect 13078 19728 13084 19740
rect 13136 19728 13142 19780
rect 13188 19768 13216 19799
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 13832 19836 13860 19864
rect 14369 19839 14427 19845
rect 14369 19836 14381 19839
rect 13832 19808 14381 19836
rect 14369 19805 14381 19808
rect 14415 19805 14427 19839
rect 14369 19799 14427 19805
rect 16206 19796 16212 19848
rect 16264 19836 16270 19848
rect 16482 19836 16488 19848
rect 16264 19808 16488 19836
rect 16264 19796 16270 19808
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 16577 19839 16635 19845
rect 16577 19805 16589 19839
rect 16623 19836 16635 19839
rect 17126 19836 17132 19848
rect 16623 19808 17132 19836
rect 16623 19805 16635 19808
rect 16577 19799 16635 19805
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 17586 19836 17592 19848
rect 17547 19808 17592 19836
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19805 17739 19839
rect 17954 19836 17960 19848
rect 17915 19808 17960 19836
rect 17681 19799 17739 19805
rect 14093 19771 14151 19777
rect 14093 19768 14105 19771
rect 13188 19740 14105 19768
rect 14093 19737 14105 19740
rect 14139 19737 14151 19771
rect 14093 19731 14151 19737
rect 14182 19728 14188 19780
rect 14240 19768 14246 19780
rect 15562 19768 15568 19780
rect 14240 19740 15568 19768
rect 14240 19728 14246 19740
rect 15562 19728 15568 19740
rect 15620 19768 15626 19780
rect 16669 19771 16727 19777
rect 16669 19768 16681 19771
rect 15620 19740 16681 19768
rect 15620 19728 15626 19740
rect 16669 19737 16681 19740
rect 16715 19737 16727 19771
rect 16669 19731 16727 19737
rect 16758 19728 16764 19780
rect 16816 19768 16822 19780
rect 17696 19768 17724 19799
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 18782 19796 18788 19848
rect 18840 19836 18846 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 18840 19808 19257 19836
rect 18840 19796 18846 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 19444 19845 19472 19944
rect 22278 19932 22284 19944
rect 22336 19932 22342 19984
rect 20162 19864 20168 19916
rect 20220 19904 20226 19916
rect 21174 19904 21180 19916
rect 20220 19876 21180 19904
rect 20220 19864 20226 19876
rect 21174 19864 21180 19876
rect 21232 19864 21238 19916
rect 22094 19904 22100 19916
rect 21652 19876 22100 19904
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 19392 19808 19441 19836
rect 19392 19796 19398 19808
rect 19429 19805 19441 19808
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 19521 19839 19579 19845
rect 19521 19805 19533 19839
rect 19567 19805 19579 19839
rect 19521 19799 19579 19805
rect 16816 19740 17724 19768
rect 16816 19728 16822 19740
rect 18874 19728 18880 19780
rect 18932 19768 18938 19780
rect 19536 19768 19564 19799
rect 19610 19796 19616 19848
rect 19668 19836 19674 19848
rect 19794 19836 19800 19848
rect 19668 19808 19713 19836
rect 19755 19808 19800 19836
rect 19668 19796 19674 19808
rect 19794 19796 19800 19808
rect 19852 19796 19858 19848
rect 19978 19796 19984 19848
rect 20036 19836 20042 19848
rect 20346 19836 20352 19848
rect 20036 19808 20352 19836
rect 20036 19796 20042 19808
rect 20346 19796 20352 19808
rect 20404 19796 20410 19848
rect 20530 19836 20536 19848
rect 20491 19808 20536 19836
rect 20530 19796 20536 19808
rect 20588 19796 20594 19848
rect 20990 19796 20996 19848
rect 21048 19836 21054 19848
rect 21266 19836 21272 19848
rect 21048 19808 21272 19836
rect 21048 19796 21054 19808
rect 21266 19796 21272 19808
rect 21324 19836 21330 19848
rect 21652 19845 21680 19876
rect 22094 19864 22100 19876
rect 22152 19864 22158 19916
rect 22554 19864 22560 19916
rect 22612 19904 22618 19916
rect 23477 19907 23535 19913
rect 22612 19876 23336 19904
rect 22612 19864 22618 19876
rect 21453 19839 21511 19845
rect 21453 19836 21465 19839
rect 21324 19808 21465 19836
rect 21324 19796 21330 19808
rect 21453 19805 21465 19808
rect 21499 19805 21511 19839
rect 21453 19799 21511 19805
rect 21601 19839 21680 19845
rect 21601 19805 21613 19839
rect 21647 19808 21680 19839
rect 21647 19805 21659 19808
rect 21601 19799 21659 19805
rect 21726 19796 21732 19848
rect 21784 19836 21790 19848
rect 21959 19839 22017 19845
rect 21784 19808 21829 19836
rect 21784 19796 21790 19808
rect 21959 19805 21971 19839
rect 22005 19836 22017 19839
rect 22462 19836 22468 19848
rect 22005 19808 22468 19836
rect 22005 19805 22017 19808
rect 21959 19799 22017 19805
rect 22462 19796 22468 19808
rect 22520 19796 22526 19848
rect 23106 19836 23112 19848
rect 23067 19808 23112 19836
rect 23106 19796 23112 19808
rect 23164 19796 23170 19848
rect 23308 19845 23336 19876
rect 23477 19873 23489 19907
rect 23523 19904 23535 19907
rect 23750 19904 23756 19916
rect 23523 19876 23756 19904
rect 23523 19873 23535 19876
rect 23477 19867 23535 19873
rect 23750 19864 23756 19876
rect 23808 19864 23814 19916
rect 23293 19839 23351 19845
rect 23293 19805 23305 19839
rect 23339 19805 23351 19839
rect 23293 19799 23351 19805
rect 23382 19796 23388 19848
rect 23440 19836 23446 19848
rect 23661 19839 23719 19845
rect 23440 19808 23485 19836
rect 23440 19796 23446 19808
rect 23661 19805 23673 19839
rect 23707 19836 23719 19839
rect 23860 19836 23888 20012
rect 25777 20009 25789 20012
rect 25823 20009 25835 20043
rect 25777 20003 25835 20009
rect 26142 20000 26148 20052
rect 26200 20040 26206 20052
rect 26200 20012 26832 20040
rect 26200 20000 26206 20012
rect 25590 19932 25596 19984
rect 25648 19972 25654 19984
rect 26050 19972 26056 19984
rect 25648 19944 26056 19972
rect 25648 19932 25654 19944
rect 26050 19932 26056 19944
rect 26108 19932 26114 19984
rect 26694 19972 26700 19984
rect 26436 19944 26700 19972
rect 23707 19808 23888 19836
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 23934 19796 23940 19848
rect 23992 19836 23998 19848
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 23992 19808 24409 19836
rect 23992 19796 23998 19808
rect 24397 19805 24409 19808
rect 24443 19836 24455 19839
rect 24486 19836 24492 19848
rect 24443 19808 24492 19836
rect 24443 19805 24455 19808
rect 24397 19799 24455 19805
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 26436 19845 26464 19944
rect 26694 19932 26700 19944
rect 26752 19932 26758 19984
rect 26804 19913 26832 20012
rect 27172 20012 28028 20040
rect 26970 19932 26976 19984
rect 27028 19932 27034 19984
rect 26789 19907 26847 19913
rect 26789 19873 26801 19907
rect 26835 19873 26847 19907
rect 26988 19904 27016 19932
rect 26789 19867 26847 19873
rect 26896 19876 27016 19904
rect 26421 19839 26479 19845
rect 26421 19805 26433 19839
rect 26467 19805 26479 19839
rect 26421 19799 26479 19805
rect 26510 19796 26516 19848
rect 26568 19836 26574 19848
rect 26605 19839 26663 19845
rect 26605 19836 26617 19839
rect 26568 19808 26617 19836
rect 26568 19796 26574 19808
rect 26605 19805 26617 19808
rect 26651 19805 26663 19839
rect 26605 19799 26663 19805
rect 26697 19839 26755 19845
rect 26697 19805 26709 19839
rect 26743 19836 26755 19839
rect 26896 19836 26924 19876
rect 26743 19808 26924 19836
rect 26973 19839 27031 19845
rect 26743 19805 26755 19808
rect 26697 19799 26755 19805
rect 26973 19805 26985 19839
rect 27019 19836 27031 19839
rect 27172 19836 27200 20012
rect 27430 19932 27436 19984
rect 27488 19972 27494 19984
rect 28000 19972 28028 20012
rect 28074 20000 28080 20052
rect 28132 20040 28138 20052
rect 28905 20043 28963 20049
rect 28905 20040 28917 20043
rect 28132 20012 28917 20040
rect 28132 20000 28138 20012
rect 28905 20009 28917 20012
rect 28951 20009 28963 20043
rect 28905 20003 28963 20009
rect 29641 19975 29699 19981
rect 29641 19972 29653 19975
rect 27488 19944 27936 19972
rect 28000 19944 29653 19972
rect 27488 19932 27494 19944
rect 27019 19808 27200 19836
rect 27019 19805 27031 19808
rect 26973 19799 27031 19805
rect 27246 19796 27252 19848
rect 27304 19836 27310 19848
rect 27617 19839 27675 19845
rect 27617 19836 27629 19839
rect 27304 19808 27629 19836
rect 27304 19796 27310 19808
rect 27617 19805 27629 19808
rect 27663 19805 27675 19839
rect 27617 19799 27675 19805
rect 27706 19796 27712 19848
rect 27764 19836 27770 19848
rect 27908 19845 27936 19944
rect 29641 19941 29653 19944
rect 29687 19941 29699 19975
rect 29641 19935 29699 19941
rect 27801 19839 27859 19845
rect 27801 19836 27813 19839
rect 27764 19808 27813 19836
rect 27764 19796 27770 19808
rect 27801 19805 27813 19808
rect 27847 19805 27859 19839
rect 27801 19799 27859 19805
rect 27893 19839 27951 19845
rect 27893 19805 27905 19839
rect 27939 19805 27951 19839
rect 27893 19799 27951 19805
rect 27982 19796 27988 19848
rect 28040 19836 28046 19848
rect 28169 19839 28227 19845
rect 28040 19808 28085 19836
rect 28040 19796 28046 19808
rect 28169 19805 28181 19839
rect 28215 19805 28227 19839
rect 28169 19799 28227 19805
rect 28813 19839 28871 19845
rect 28813 19805 28825 19839
rect 28859 19836 28871 19839
rect 29454 19836 29460 19848
rect 28859 19808 29460 19836
rect 28859 19805 28871 19808
rect 28813 19799 28871 19805
rect 18932 19740 19564 19768
rect 20717 19771 20775 19777
rect 18932 19728 18938 19740
rect 20717 19737 20729 19771
rect 20763 19768 20775 19771
rect 20806 19768 20812 19780
rect 20763 19740 20812 19768
rect 20763 19737 20775 19740
rect 20717 19731 20775 19737
rect 20806 19728 20812 19740
rect 20864 19728 20870 19780
rect 21821 19771 21879 19777
rect 21821 19768 21833 19771
rect 20916 19740 21833 19768
rect 1394 19660 1400 19712
rect 1452 19700 1458 19712
rect 1673 19703 1731 19709
rect 1673 19700 1685 19703
rect 1452 19672 1685 19700
rect 1452 19660 1458 19672
rect 1673 19669 1685 19672
rect 1719 19669 1731 19703
rect 1673 19663 1731 19669
rect 10042 19660 10048 19712
rect 10100 19700 10106 19712
rect 10321 19703 10379 19709
rect 10321 19700 10333 19703
rect 10100 19672 10333 19700
rect 10100 19660 10106 19672
rect 10321 19669 10333 19672
rect 10367 19700 10379 19703
rect 11701 19703 11759 19709
rect 11701 19700 11713 19703
rect 10367 19672 11713 19700
rect 10367 19669 10379 19672
rect 10321 19663 10379 19669
rect 11701 19669 11713 19672
rect 11747 19669 11759 19703
rect 11701 19663 11759 19669
rect 12066 19660 12072 19712
rect 12124 19700 12130 19712
rect 12618 19700 12624 19712
rect 12124 19672 12624 19700
rect 12124 19660 12130 19672
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 13541 19703 13599 19709
rect 13541 19669 13553 19703
rect 13587 19700 13599 19703
rect 14366 19700 14372 19712
rect 13587 19672 14372 19700
rect 13587 19669 13599 19672
rect 13541 19663 13599 19669
rect 14366 19660 14372 19672
rect 14424 19700 14430 19712
rect 14734 19700 14740 19712
rect 14424 19672 14740 19700
rect 14424 19660 14430 19672
rect 14734 19660 14740 19672
rect 14792 19660 14798 19712
rect 15010 19700 15016 19712
rect 14971 19672 15016 19700
rect 15010 19660 15016 19672
rect 15068 19660 15074 19712
rect 15378 19700 15384 19712
rect 15339 19672 15384 19700
rect 15378 19660 15384 19672
rect 15436 19660 15442 19712
rect 16206 19700 16212 19712
rect 16167 19672 16212 19700
rect 16206 19660 16212 19672
rect 16264 19660 16270 19712
rect 16850 19660 16856 19712
rect 16908 19700 16914 19712
rect 17405 19703 17463 19709
rect 17405 19700 17417 19703
rect 16908 19672 17417 19700
rect 16908 19660 16914 19672
rect 17405 19669 17417 19672
rect 17451 19669 17463 19703
rect 17405 19663 17463 19669
rect 17770 19660 17776 19712
rect 17828 19700 17834 19712
rect 19426 19700 19432 19712
rect 17828 19672 19432 19700
rect 17828 19660 17834 19672
rect 19426 19660 19432 19672
rect 19484 19660 19490 19712
rect 20346 19660 20352 19712
rect 20404 19700 20410 19712
rect 20916 19700 20944 19740
rect 21821 19737 21833 19740
rect 21867 19737 21879 19771
rect 21821 19731 21879 19737
rect 23845 19771 23903 19777
rect 23845 19737 23857 19771
rect 23891 19768 23903 19771
rect 24642 19771 24700 19777
rect 24642 19768 24654 19771
rect 23891 19740 24654 19768
rect 23891 19737 23903 19740
rect 23845 19731 23903 19737
rect 24642 19737 24654 19740
rect 24688 19737 24700 19771
rect 24642 19731 24700 19737
rect 24762 19728 24768 19780
rect 24820 19768 24826 19780
rect 27157 19771 27215 19777
rect 27157 19768 27169 19771
rect 24820 19740 27169 19768
rect 24820 19728 24826 19740
rect 27157 19737 27169 19740
rect 27203 19737 27215 19771
rect 28184 19768 28212 19799
rect 29454 19796 29460 19808
rect 29512 19796 29518 19848
rect 29549 19839 29607 19845
rect 29549 19805 29561 19839
rect 29595 19805 29607 19839
rect 29549 19799 29607 19805
rect 28534 19768 28540 19780
rect 28184 19740 28540 19768
rect 27157 19731 27215 19737
rect 28534 19728 28540 19740
rect 28592 19768 28598 19780
rect 29564 19768 29592 19799
rect 28592 19740 29592 19768
rect 28592 19728 28598 19740
rect 22094 19700 22100 19712
rect 20404 19672 20944 19700
rect 22055 19672 22100 19700
rect 20404 19660 20410 19672
rect 22094 19660 22100 19672
rect 22152 19660 22158 19712
rect 25590 19660 25596 19712
rect 25648 19700 25654 19712
rect 26970 19700 26976 19712
rect 25648 19672 26976 19700
rect 25648 19660 25654 19672
rect 26970 19660 26976 19672
rect 27028 19660 27034 19712
rect 28350 19700 28356 19712
rect 28311 19672 28356 19700
rect 28350 19660 28356 19672
rect 28408 19660 28414 19712
rect 1104 19610 30820 19632
rect 1104 19558 10880 19610
rect 10932 19558 10944 19610
rect 10996 19558 11008 19610
rect 11060 19558 11072 19610
rect 11124 19558 11136 19610
rect 11188 19558 20811 19610
rect 20863 19558 20875 19610
rect 20927 19558 20939 19610
rect 20991 19558 21003 19610
rect 21055 19558 21067 19610
rect 21119 19558 30820 19610
rect 1104 19536 30820 19558
rect 9214 19456 9220 19508
rect 9272 19496 9278 19508
rect 10321 19499 10379 19505
rect 10321 19496 10333 19499
rect 9272 19468 10333 19496
rect 9272 19456 9278 19468
rect 10321 19465 10333 19468
rect 10367 19465 10379 19499
rect 10321 19459 10379 19465
rect 12526 19456 12532 19508
rect 12584 19496 12590 19508
rect 13449 19499 13507 19505
rect 13449 19496 13461 19499
rect 12584 19468 13461 19496
rect 12584 19456 12590 19468
rect 13449 19465 13461 19468
rect 13495 19465 13507 19499
rect 13449 19459 13507 19465
rect 13538 19456 13544 19508
rect 13596 19496 13602 19508
rect 14182 19496 14188 19508
rect 13596 19468 14188 19496
rect 13596 19456 13602 19468
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 14829 19499 14887 19505
rect 14829 19465 14841 19499
rect 14875 19496 14887 19499
rect 22002 19496 22008 19508
rect 14875 19468 22008 19496
rect 14875 19465 14887 19468
rect 14829 19459 14887 19465
rect 22002 19456 22008 19468
rect 22060 19456 22066 19508
rect 22278 19456 22284 19508
rect 22336 19496 22342 19508
rect 22738 19496 22744 19508
rect 22336 19468 22744 19496
rect 22336 19456 22342 19468
rect 22738 19456 22744 19468
rect 22796 19456 22802 19508
rect 24946 19456 24952 19508
rect 25004 19496 25010 19508
rect 25317 19499 25375 19505
rect 25317 19496 25329 19499
rect 25004 19468 25329 19496
rect 25004 19456 25010 19468
rect 25317 19465 25329 19468
rect 25363 19465 25375 19499
rect 25317 19459 25375 19465
rect 26234 19456 26240 19508
rect 26292 19496 26298 19508
rect 28166 19496 28172 19508
rect 26292 19468 28172 19496
rect 26292 19456 26298 19468
rect 28166 19456 28172 19468
rect 28224 19456 28230 19508
rect 29178 19456 29184 19508
rect 29236 19496 29242 19508
rect 30101 19499 30159 19505
rect 30101 19496 30113 19499
rect 29236 19468 30113 19496
rect 29236 19456 29242 19468
rect 30101 19465 30113 19468
rect 30147 19465 30159 19499
rect 30101 19459 30159 19465
rect 9953 19431 10011 19437
rect 9953 19397 9965 19431
rect 9999 19428 10011 19431
rect 15010 19428 15016 19440
rect 9999 19400 15016 19428
rect 9999 19397 10011 19400
rect 9953 19391 10011 19397
rect 15010 19388 15016 19400
rect 15068 19388 15074 19440
rect 15562 19428 15568 19440
rect 15523 19400 15568 19428
rect 15562 19388 15568 19400
rect 15620 19388 15626 19440
rect 16945 19431 17003 19437
rect 16945 19397 16957 19431
rect 16991 19428 17003 19431
rect 17034 19428 17040 19440
rect 16991 19400 17040 19428
rect 16991 19397 17003 19400
rect 16945 19391 17003 19397
rect 17034 19388 17040 19400
rect 17092 19388 17098 19440
rect 17957 19431 18015 19437
rect 17957 19397 17969 19431
rect 18003 19428 18015 19431
rect 21174 19428 21180 19440
rect 18003 19400 21180 19428
rect 18003 19397 18015 19400
rect 17957 19391 18015 19397
rect 21174 19388 21180 19400
rect 21232 19388 21238 19440
rect 23658 19428 23664 19440
rect 21836 19400 23664 19428
rect 1394 19360 1400 19372
rect 1355 19332 1400 19360
rect 1394 19320 1400 19332
rect 1452 19320 1458 19372
rect 9674 19360 9680 19372
rect 9635 19332 9680 19360
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 9858 19369 9864 19372
rect 9825 19363 9864 19369
rect 9825 19329 9837 19363
rect 9825 19323 9864 19329
rect 9858 19320 9864 19323
rect 9916 19320 9922 19372
rect 10042 19360 10048 19372
rect 10003 19332 10048 19360
rect 10042 19320 10048 19332
rect 10100 19320 10106 19372
rect 10134 19320 10140 19372
rect 10192 19369 10198 19372
rect 10192 19360 10200 19369
rect 11977 19363 12035 19369
rect 10192 19332 10237 19360
rect 10192 19323 10200 19332
rect 11977 19329 11989 19363
rect 12023 19360 12035 19363
rect 12437 19363 12495 19369
rect 12023 19332 12296 19360
rect 12023 19329 12035 19332
rect 11977 19323 12035 19329
rect 10192 19320 10198 19323
rect 11882 19252 11888 19304
rect 11940 19252 11946 19304
rect 10042 19184 10048 19236
rect 10100 19224 10106 19236
rect 11900 19224 11928 19252
rect 10100 19196 11928 19224
rect 10100 19184 10106 19196
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 11606 19116 11612 19168
rect 11664 19156 11670 19168
rect 11882 19156 11888 19168
rect 11664 19128 11888 19156
rect 11664 19116 11670 19128
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 12268 19156 12296 19332
rect 12437 19329 12449 19363
rect 12483 19360 12495 19363
rect 13078 19360 13084 19372
rect 12483 19332 13084 19360
rect 12483 19329 12495 19332
rect 12437 19323 12495 19329
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 13265 19363 13323 19369
rect 13265 19360 13277 19363
rect 13188 19332 13277 19360
rect 12345 19295 12403 19301
rect 12345 19261 12357 19295
rect 12391 19292 12403 19295
rect 13188 19292 13216 19332
rect 13265 19329 13277 19332
rect 13311 19360 13323 19363
rect 13311 19332 13860 19360
rect 13311 19329 13323 19332
rect 13265 19323 13323 19329
rect 12391 19264 13216 19292
rect 12391 19261 12403 19264
rect 12345 19255 12403 19261
rect 13832 19168 13860 19332
rect 13906 19320 13912 19372
rect 13964 19360 13970 19372
rect 13964 19332 14009 19360
rect 13964 19320 13970 19332
rect 14182 19320 14188 19372
rect 14240 19360 14246 19372
rect 14734 19360 14740 19372
rect 14240 19346 14596 19360
rect 14240 19332 14372 19346
rect 14240 19320 14246 19332
rect 14366 19294 14372 19332
rect 14424 19306 14596 19346
rect 14695 19332 14740 19360
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 14918 19360 14924 19372
rect 14879 19332 14924 19360
rect 14918 19320 14924 19332
rect 14976 19360 14982 19372
rect 15473 19363 15531 19369
rect 15473 19360 15485 19363
rect 14976 19332 15485 19360
rect 14976 19320 14982 19332
rect 15473 19329 15485 19332
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 16206 19320 16212 19372
rect 16264 19360 16270 19372
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 16264 19332 16681 19360
rect 16264 19320 16270 19332
rect 16669 19329 16681 19332
rect 16715 19329 16727 19363
rect 16669 19323 16727 19329
rect 17310 19320 17316 19372
rect 17368 19360 17374 19372
rect 17770 19369 17776 19372
rect 17589 19363 17647 19369
rect 17589 19360 17601 19363
rect 17368 19332 17601 19360
rect 17368 19320 17374 19332
rect 17589 19329 17601 19332
rect 17635 19329 17647 19363
rect 17589 19323 17647 19329
rect 17737 19363 17776 19369
rect 17737 19329 17749 19363
rect 17737 19323 17776 19329
rect 17770 19320 17776 19323
rect 17828 19320 17834 19372
rect 17865 19363 17923 19369
rect 17865 19329 17877 19363
rect 17911 19329 17923 19363
rect 17865 19323 17923 19329
rect 14424 19294 14430 19306
rect 14936 19292 14964 19320
rect 15010 19292 15016 19304
rect 14936 19264 15016 19292
rect 15010 19252 15016 19264
rect 15068 19252 15074 19304
rect 17880 19292 17908 19323
rect 18046 19320 18052 19372
rect 18104 19369 18110 19372
rect 18104 19360 18112 19369
rect 19521 19363 19579 19369
rect 18104 19332 18149 19360
rect 18104 19323 18112 19332
rect 19521 19329 19533 19363
rect 19567 19360 19579 19363
rect 20530 19360 20536 19372
rect 19567 19332 20536 19360
rect 19567 19329 19579 19332
rect 19521 19323 19579 19329
rect 18104 19320 18110 19323
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 20714 19320 20720 19372
rect 20772 19360 20778 19372
rect 21836 19369 21864 19400
rect 23658 19388 23664 19400
rect 23716 19388 23722 19440
rect 20809 19363 20867 19369
rect 20809 19360 20821 19363
rect 20772 19332 20821 19360
rect 20772 19320 20778 19332
rect 20809 19329 20821 19332
rect 20855 19329 20867 19363
rect 20809 19323 20867 19329
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 21910 19320 21916 19372
rect 21968 19320 21974 19372
rect 22094 19369 22100 19372
rect 22088 19360 22100 19369
rect 22055 19332 22100 19360
rect 22088 19323 22100 19332
rect 22094 19320 22100 19323
rect 22152 19320 22158 19372
rect 24210 19369 24216 19372
rect 24204 19323 24216 19369
rect 24268 19360 24274 19372
rect 26234 19360 26240 19372
rect 24268 19332 24304 19360
rect 26195 19332 26240 19360
rect 24210 19320 24216 19323
rect 24268 19320 24274 19332
rect 26234 19320 26240 19332
rect 26292 19320 26298 19372
rect 27433 19363 27491 19369
rect 27433 19329 27445 19363
rect 27479 19360 27491 19363
rect 27479 19332 27513 19360
rect 27479 19329 27491 19332
rect 27433 19323 27491 19329
rect 17696 19264 17908 19292
rect 20993 19295 21051 19301
rect 17696 19236 17724 19264
rect 20993 19261 21005 19295
rect 21039 19292 21051 19295
rect 21928 19292 21956 19320
rect 21039 19264 21956 19292
rect 21039 19261 21051 19264
rect 20993 19255 21051 19261
rect 23658 19252 23664 19304
rect 23716 19292 23722 19304
rect 23934 19292 23940 19304
rect 23716 19264 23940 19292
rect 23716 19252 23722 19264
rect 23934 19252 23940 19264
rect 23992 19252 23998 19304
rect 25682 19252 25688 19304
rect 25740 19292 25746 19304
rect 27157 19295 27215 19301
rect 27157 19292 27169 19295
rect 25740 19264 27169 19292
rect 25740 19252 25746 19264
rect 27157 19261 27169 19264
rect 27203 19261 27215 19295
rect 27448 19292 27476 19323
rect 28442 19320 28448 19372
rect 28500 19360 28506 19372
rect 28994 19369 29000 19372
rect 28721 19363 28779 19369
rect 28721 19360 28733 19363
rect 28500 19332 28733 19360
rect 28500 19320 28506 19332
rect 28721 19329 28733 19332
rect 28767 19329 28779 19363
rect 28721 19323 28779 19329
rect 28988 19323 29000 19369
rect 29052 19360 29058 19372
rect 29052 19332 29088 19360
rect 28994 19320 29000 19323
rect 29052 19320 29058 19332
rect 27522 19292 27528 19304
rect 27435 19264 27528 19292
rect 27157 19255 27215 19261
rect 27522 19252 27528 19264
rect 27580 19292 27586 19304
rect 27580 19264 28764 19292
rect 27580 19252 27586 19264
rect 28736 19236 28764 19264
rect 17678 19184 17684 19236
rect 17736 19184 17742 19236
rect 19150 19184 19156 19236
rect 19208 19224 19214 19236
rect 20898 19224 20904 19236
rect 19208 19196 20904 19224
rect 19208 19184 19214 19196
rect 20898 19184 20904 19196
rect 20956 19184 20962 19236
rect 26326 19224 26332 19236
rect 25240 19196 26332 19224
rect 12526 19156 12532 19168
rect 12268 19128 12532 19156
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 12621 19159 12679 19165
rect 12621 19125 12633 19159
rect 12667 19156 12679 19159
rect 13170 19156 13176 19168
rect 12667 19128 13176 19156
rect 12667 19125 12679 19128
rect 12621 19119 12679 19125
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 13814 19116 13820 19168
rect 13872 19116 13878 19168
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 18233 19159 18291 19165
rect 18233 19156 18245 19159
rect 18012 19128 18245 19156
rect 18012 19116 18018 19128
rect 18233 19125 18245 19128
rect 18279 19125 18291 19159
rect 18233 19119 18291 19125
rect 19518 19116 19524 19168
rect 19576 19156 19582 19168
rect 19705 19159 19763 19165
rect 19705 19156 19717 19159
rect 19576 19128 19717 19156
rect 19576 19116 19582 19128
rect 19705 19125 19717 19128
rect 19751 19125 19763 19159
rect 19705 19119 19763 19125
rect 21726 19116 21732 19168
rect 21784 19156 21790 19168
rect 22002 19156 22008 19168
rect 21784 19128 22008 19156
rect 21784 19116 21790 19128
rect 22002 19116 22008 19128
rect 22060 19156 22066 19168
rect 23201 19159 23259 19165
rect 23201 19156 23213 19159
rect 22060 19128 23213 19156
rect 22060 19116 22066 19128
rect 23201 19125 23213 19128
rect 23247 19125 23259 19159
rect 23201 19119 23259 19125
rect 23658 19116 23664 19168
rect 23716 19156 23722 19168
rect 25240 19156 25268 19196
rect 26326 19184 26332 19196
rect 26384 19184 26390 19236
rect 26421 19227 26479 19233
rect 26421 19193 26433 19227
rect 26467 19224 26479 19227
rect 28442 19224 28448 19236
rect 26467 19196 28448 19224
rect 26467 19193 26479 19196
rect 26421 19187 26479 19193
rect 28442 19184 28448 19196
rect 28500 19184 28506 19236
rect 28718 19184 28724 19236
rect 28776 19184 28782 19236
rect 23716 19128 25268 19156
rect 23716 19116 23722 19128
rect 1104 19066 30820 19088
rect 1104 19014 5915 19066
rect 5967 19014 5979 19066
rect 6031 19014 6043 19066
rect 6095 19014 6107 19066
rect 6159 19014 6171 19066
rect 6223 19014 15846 19066
rect 15898 19014 15910 19066
rect 15962 19014 15974 19066
rect 16026 19014 16038 19066
rect 16090 19014 16102 19066
rect 16154 19014 25776 19066
rect 25828 19014 25840 19066
rect 25892 19014 25904 19066
rect 25956 19014 25968 19066
rect 26020 19014 26032 19066
rect 26084 19014 30820 19066
rect 1104 18992 30820 19014
rect 10134 18912 10140 18964
rect 10192 18952 10198 18964
rect 10502 18952 10508 18964
rect 10192 18924 10508 18952
rect 10192 18912 10198 18924
rect 10502 18912 10508 18924
rect 10560 18952 10566 18964
rect 11241 18955 11299 18961
rect 10560 18924 11100 18952
rect 10560 18912 10566 18924
rect 11072 18816 11100 18924
rect 11241 18921 11253 18955
rect 11287 18952 11299 18955
rect 11790 18952 11796 18964
rect 11287 18924 11796 18952
rect 11287 18921 11299 18924
rect 11241 18915 11299 18921
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 11882 18912 11888 18964
rect 11940 18952 11946 18964
rect 15378 18952 15384 18964
rect 11940 18924 14596 18952
rect 15339 18924 15384 18952
rect 11940 18912 11946 18924
rect 11808 18884 11836 18912
rect 13354 18884 13360 18896
rect 11808 18856 13360 18884
rect 13354 18844 13360 18856
rect 13412 18844 13418 18896
rect 14182 18844 14188 18896
rect 14240 18884 14246 18896
rect 14458 18884 14464 18896
rect 14240 18856 14464 18884
rect 14240 18844 14246 18856
rect 14458 18844 14464 18856
rect 14516 18844 14522 18896
rect 14568 18884 14596 18924
rect 15378 18912 15384 18924
rect 15436 18912 15442 18964
rect 19981 18955 20039 18961
rect 19981 18921 19993 18955
rect 20027 18952 20039 18955
rect 21726 18952 21732 18964
rect 20027 18924 21732 18952
rect 20027 18921 20039 18924
rect 19981 18915 20039 18921
rect 21726 18912 21732 18924
rect 21784 18912 21790 18964
rect 23753 18955 23811 18961
rect 23753 18921 23765 18955
rect 23799 18952 23811 18955
rect 25038 18952 25044 18964
rect 23799 18924 25044 18952
rect 23799 18921 23811 18924
rect 23753 18915 23811 18921
rect 25038 18912 25044 18924
rect 25096 18912 25102 18964
rect 25314 18912 25320 18964
rect 25372 18952 25378 18964
rect 25498 18952 25504 18964
rect 25372 18924 25504 18952
rect 25372 18912 25378 18924
rect 25498 18912 25504 18924
rect 25556 18912 25562 18964
rect 26510 18912 26516 18964
rect 26568 18952 26574 18964
rect 29917 18955 29975 18961
rect 29917 18952 29929 18955
rect 26568 18924 29929 18952
rect 26568 18912 26574 18924
rect 29917 18921 29929 18924
rect 29963 18921 29975 18955
rect 29917 18915 29975 18921
rect 16390 18884 16396 18896
rect 14568 18856 16396 18884
rect 16390 18844 16396 18856
rect 16448 18844 16454 18896
rect 20714 18844 20720 18896
rect 20772 18884 20778 18896
rect 21453 18887 21511 18893
rect 21453 18884 21465 18887
rect 20772 18856 21465 18884
rect 20772 18844 20778 18856
rect 21453 18853 21465 18856
rect 21499 18853 21511 18887
rect 25869 18887 25927 18893
rect 25869 18884 25881 18887
rect 21453 18847 21511 18853
rect 22066 18856 25881 18884
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 11072 18788 12173 18816
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12161 18779 12219 18785
rect 13078 18776 13084 18828
rect 13136 18816 13142 18828
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 13136 18788 14381 18816
rect 13136 18776 13142 18788
rect 14369 18785 14381 18788
rect 14415 18816 14427 18819
rect 14550 18816 14556 18828
rect 14415 18788 14556 18816
rect 14415 18785 14427 18788
rect 14369 18779 14427 18785
rect 14550 18776 14556 18788
rect 14608 18776 14614 18828
rect 15378 18776 15384 18828
rect 15436 18816 15442 18828
rect 16022 18816 16028 18828
rect 15436 18788 16028 18816
rect 15436 18776 15442 18788
rect 16022 18776 16028 18788
rect 16080 18776 16086 18828
rect 16853 18819 16911 18825
rect 16853 18785 16865 18819
rect 16899 18816 16911 18819
rect 17494 18816 17500 18828
rect 16899 18788 17500 18816
rect 16899 18785 16911 18788
rect 16853 18779 16911 18785
rect 17494 18776 17500 18788
rect 17552 18776 17558 18828
rect 19536 18788 20668 18816
rect 9306 18708 9312 18760
rect 9364 18748 9370 18760
rect 9861 18751 9919 18757
rect 9861 18748 9873 18751
rect 9364 18720 9873 18748
rect 9364 18708 9370 18720
rect 9861 18717 9873 18720
rect 9907 18717 9919 18751
rect 9861 18711 9919 18717
rect 11606 18708 11612 18760
rect 11664 18748 11670 18760
rect 11793 18751 11851 18757
rect 11793 18748 11805 18751
rect 11664 18720 11805 18748
rect 11664 18708 11670 18720
rect 11793 18717 11805 18720
rect 11839 18717 11851 18751
rect 11793 18711 11851 18717
rect 11882 18708 11888 18760
rect 11940 18748 11946 18760
rect 11977 18751 12035 18757
rect 11977 18748 11989 18751
rect 11940 18720 11989 18748
rect 11940 18708 11946 18720
rect 11977 18717 11989 18720
rect 12023 18717 12035 18751
rect 11977 18711 12035 18717
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18748 12127 18751
rect 12250 18748 12256 18760
rect 12115 18720 12256 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 12345 18751 12403 18757
rect 12345 18717 12357 18751
rect 12391 18748 12403 18751
rect 12710 18748 12716 18760
rect 12391 18720 12716 18748
rect 12391 18717 12403 18720
rect 12345 18711 12403 18717
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 13354 18748 13360 18760
rect 13315 18720 13360 18748
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 13449 18751 13507 18757
rect 13449 18717 13461 18751
rect 13495 18748 13507 18751
rect 14090 18748 14096 18760
rect 13495 18720 14096 18748
rect 13495 18717 13507 18720
rect 13449 18711 13507 18717
rect 14090 18708 14096 18720
rect 14148 18708 14154 18760
rect 14185 18751 14243 18757
rect 14185 18717 14197 18751
rect 14231 18748 14243 18751
rect 14734 18748 14740 18760
rect 14231 18720 14740 18748
rect 14231 18717 14243 18720
rect 14185 18711 14243 18717
rect 14734 18708 14740 18720
rect 14792 18708 14798 18760
rect 15197 18751 15255 18757
rect 15197 18717 15209 18751
rect 15243 18717 15255 18751
rect 15197 18711 15255 18717
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18717 15347 18751
rect 15470 18748 15476 18760
rect 15431 18720 15476 18748
rect 15289 18711 15347 18717
rect 10128 18683 10186 18689
rect 10128 18649 10140 18683
rect 10174 18680 10186 18683
rect 12529 18683 12587 18689
rect 12529 18680 12541 18683
rect 10174 18652 12541 18680
rect 10174 18649 10186 18652
rect 10128 18643 10186 18649
rect 12529 18649 12541 18652
rect 12575 18649 12587 18683
rect 15212 18680 15240 18711
rect 12529 18643 12587 18649
rect 13372 18652 15240 18680
rect 15304 18680 15332 18711
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 15562 18708 15568 18760
rect 15620 18748 15626 18760
rect 15620 18720 15665 18748
rect 15620 18708 15626 18720
rect 16114 18708 16120 18760
rect 16172 18748 16178 18760
rect 16577 18751 16635 18757
rect 16577 18748 16589 18751
rect 16172 18720 16589 18748
rect 16172 18708 16178 18720
rect 16577 18717 16589 18720
rect 16623 18717 16635 18751
rect 16577 18711 16635 18717
rect 17310 18708 17316 18760
rect 17368 18748 17374 18760
rect 17770 18757 17776 18760
rect 17589 18751 17647 18757
rect 17589 18748 17601 18751
rect 17368 18720 17601 18748
rect 17368 18708 17374 18720
rect 17589 18717 17601 18720
rect 17635 18717 17647 18751
rect 17589 18711 17647 18717
rect 17737 18751 17776 18757
rect 17737 18717 17749 18751
rect 17737 18711 17776 18717
rect 17770 18708 17776 18711
rect 17828 18708 17834 18760
rect 18046 18748 18052 18760
rect 18005 18720 18052 18748
rect 18046 18708 18052 18720
rect 18104 18757 18110 18760
rect 18104 18751 18153 18757
rect 18104 18717 18107 18751
rect 18141 18748 18153 18751
rect 18690 18748 18696 18760
rect 18141 18720 18696 18748
rect 18141 18717 18153 18720
rect 18104 18711 18153 18717
rect 18104 18708 18110 18711
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 19536 18757 19564 18788
rect 19521 18751 19579 18757
rect 19521 18717 19533 18751
rect 19567 18717 19579 18751
rect 19521 18711 19579 18717
rect 19794 18708 19800 18760
rect 19852 18748 19858 18760
rect 20165 18751 20223 18757
rect 20165 18748 20177 18751
rect 19852 18720 20177 18748
rect 19852 18708 19858 18720
rect 20165 18717 20177 18720
rect 20211 18717 20223 18751
rect 20165 18711 20223 18717
rect 17126 18680 17132 18692
rect 15304 18652 17132 18680
rect 12250 18572 12256 18624
rect 12308 18612 12314 18624
rect 13372 18612 13400 18652
rect 17126 18640 17132 18652
rect 17184 18640 17190 18692
rect 17862 18680 17868 18692
rect 17823 18652 17868 18680
rect 17862 18640 17868 18652
rect 17920 18640 17926 18692
rect 17957 18683 18015 18689
rect 17957 18649 17969 18683
rect 18003 18680 18015 18683
rect 20438 18680 20444 18692
rect 18003 18652 20444 18680
rect 18003 18649 18015 18652
rect 17957 18643 18015 18649
rect 20438 18640 20444 18652
rect 20496 18640 20502 18692
rect 20640 18680 20668 18788
rect 20732 18757 20760 18844
rect 20898 18776 20904 18828
rect 20956 18816 20962 18828
rect 22066 18816 22094 18856
rect 25869 18853 25881 18856
rect 25915 18853 25927 18887
rect 25869 18847 25927 18853
rect 20956 18788 22094 18816
rect 20956 18776 20962 18788
rect 22186 18776 22192 18828
rect 22244 18816 22250 18828
rect 22373 18819 22431 18825
rect 22373 18816 22385 18819
rect 22244 18788 22385 18816
rect 22244 18776 22250 18788
rect 22373 18785 22385 18788
rect 22419 18785 22431 18819
rect 22373 18779 22431 18785
rect 22649 18819 22707 18825
rect 22649 18785 22661 18819
rect 22695 18816 22707 18819
rect 23198 18816 23204 18828
rect 22695 18788 23204 18816
rect 22695 18785 22707 18788
rect 22649 18779 22707 18785
rect 23198 18776 23204 18788
rect 23256 18816 23262 18828
rect 23382 18816 23388 18828
rect 23256 18788 23388 18816
rect 23256 18776 23262 18788
rect 23382 18776 23388 18788
rect 23440 18776 23446 18828
rect 25498 18816 25504 18828
rect 25459 18788 25504 18816
rect 25498 18776 25504 18788
rect 25556 18776 25562 18828
rect 26418 18816 26424 18828
rect 25700 18788 26424 18816
rect 20717 18751 20775 18757
rect 20717 18717 20729 18751
rect 20763 18717 20775 18751
rect 20717 18711 20775 18717
rect 21266 18708 21272 18760
rect 21324 18748 21330 18760
rect 21361 18751 21419 18757
rect 21361 18748 21373 18751
rect 21324 18720 21373 18748
rect 21324 18708 21330 18720
rect 21361 18717 21373 18720
rect 21407 18717 21419 18751
rect 23658 18748 23664 18760
rect 23619 18720 23664 18748
rect 21361 18711 21419 18717
rect 23658 18708 23664 18720
rect 23716 18708 23722 18760
rect 24854 18748 24860 18760
rect 24412 18720 24860 18748
rect 24412 18680 24440 18720
rect 24854 18708 24860 18720
rect 24912 18708 24918 18760
rect 25130 18748 25136 18760
rect 25091 18720 25136 18748
rect 25130 18708 25136 18720
rect 25188 18708 25194 18760
rect 25314 18748 25320 18760
rect 25275 18720 25320 18748
rect 25314 18708 25320 18720
rect 25372 18708 25378 18760
rect 25409 18751 25467 18757
rect 25409 18717 25421 18751
rect 25455 18748 25467 18751
rect 25590 18748 25596 18760
rect 25455 18720 25596 18748
rect 25455 18717 25467 18720
rect 25409 18711 25467 18717
rect 25590 18708 25596 18720
rect 25648 18708 25654 18760
rect 25700 18757 25728 18788
rect 26418 18776 26424 18788
rect 26476 18776 26482 18828
rect 28994 18776 29000 18828
rect 29052 18816 29058 18828
rect 29362 18816 29368 18828
rect 29052 18788 29368 18816
rect 29052 18776 29058 18788
rect 29362 18776 29368 18788
rect 29420 18776 29426 18828
rect 25685 18751 25743 18757
rect 25685 18717 25697 18751
rect 25731 18717 25743 18751
rect 25685 18711 25743 18717
rect 25866 18708 25872 18760
rect 25924 18748 25930 18760
rect 26329 18751 26387 18757
rect 26329 18748 26341 18751
rect 25924 18720 26341 18748
rect 25924 18708 25930 18720
rect 26329 18717 26341 18720
rect 26375 18717 26387 18751
rect 26329 18711 26387 18717
rect 26605 18751 26663 18757
rect 26605 18717 26617 18751
rect 26651 18748 26663 18751
rect 27154 18748 27160 18760
rect 26651 18720 27160 18748
rect 26651 18717 26663 18720
rect 26605 18711 26663 18717
rect 27154 18708 27160 18720
rect 27212 18708 27218 18760
rect 27614 18748 27620 18760
rect 27527 18720 27620 18748
rect 27614 18708 27620 18720
rect 27672 18748 27678 18760
rect 28442 18748 28448 18760
rect 27672 18720 28448 18748
rect 27672 18708 27678 18720
rect 28442 18708 28448 18720
rect 28500 18708 28506 18760
rect 28626 18708 28632 18760
rect 28684 18748 28690 18760
rect 30101 18751 30159 18757
rect 30101 18748 30113 18751
rect 28684 18720 30113 18748
rect 28684 18708 28690 18720
rect 30101 18717 30113 18720
rect 30147 18717 30159 18751
rect 30101 18711 30159 18717
rect 20640 18652 24440 18680
rect 24489 18683 24547 18689
rect 24489 18649 24501 18683
rect 24535 18680 24547 18683
rect 26234 18680 26240 18692
rect 24535 18652 26240 18680
rect 24535 18649 24547 18652
rect 24489 18643 24547 18649
rect 26234 18640 26240 18652
rect 26292 18640 26298 18692
rect 27884 18683 27942 18689
rect 27884 18649 27896 18683
rect 27930 18680 27942 18683
rect 29730 18680 29736 18692
rect 27930 18652 29736 18680
rect 27930 18649 27942 18652
rect 27884 18643 27942 18649
rect 29730 18640 29736 18652
rect 29788 18640 29794 18692
rect 12308 18584 13400 18612
rect 12308 18572 12314 18584
rect 14274 18572 14280 18624
rect 14332 18612 14338 18624
rect 14369 18615 14427 18621
rect 14369 18612 14381 18615
rect 14332 18584 14381 18612
rect 14332 18572 14338 18584
rect 14369 18581 14381 18584
rect 14415 18581 14427 18615
rect 14369 18575 14427 18581
rect 15194 18572 15200 18624
rect 15252 18612 15258 18624
rect 16209 18615 16267 18621
rect 16209 18612 16221 18615
rect 15252 18584 16221 18612
rect 15252 18572 15258 18584
rect 16209 18581 16221 18584
rect 16255 18581 16267 18615
rect 16209 18575 16267 18581
rect 16669 18615 16727 18621
rect 16669 18581 16681 18615
rect 16715 18612 16727 18615
rect 17678 18612 17684 18624
rect 16715 18584 17684 18612
rect 16715 18581 16727 18584
rect 16669 18575 16727 18581
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 18230 18612 18236 18624
rect 18191 18584 18236 18612
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 19334 18572 19340 18624
rect 19392 18612 19398 18624
rect 19392 18584 19437 18612
rect 19392 18572 19398 18584
rect 20622 18572 20628 18624
rect 20680 18612 20686 18624
rect 20809 18615 20867 18621
rect 20809 18612 20821 18615
rect 20680 18584 20821 18612
rect 20680 18572 20686 18584
rect 20809 18581 20821 18584
rect 20855 18581 20867 18615
rect 20809 18575 20867 18581
rect 22738 18572 22744 18624
rect 22796 18612 22802 18624
rect 23014 18612 23020 18624
rect 22796 18584 23020 18612
rect 22796 18572 22802 18584
rect 23014 18572 23020 18584
rect 23072 18572 23078 18624
rect 23934 18572 23940 18624
rect 23992 18612 23998 18624
rect 24581 18615 24639 18621
rect 24581 18612 24593 18615
rect 23992 18584 24593 18612
rect 23992 18572 23998 18584
rect 24581 18581 24593 18584
rect 24627 18612 24639 18615
rect 24854 18612 24860 18624
rect 24627 18584 24860 18612
rect 24627 18581 24639 18584
rect 24581 18575 24639 18581
rect 24854 18572 24860 18584
rect 24912 18572 24918 18624
rect 28997 18615 29055 18621
rect 28997 18581 29009 18615
rect 29043 18612 29055 18615
rect 29454 18612 29460 18624
rect 29043 18584 29460 18612
rect 29043 18581 29055 18584
rect 28997 18575 29055 18581
rect 29454 18572 29460 18584
rect 29512 18572 29518 18624
rect 1104 18522 30820 18544
rect 1104 18470 10880 18522
rect 10932 18470 10944 18522
rect 10996 18470 11008 18522
rect 11060 18470 11072 18522
rect 11124 18470 11136 18522
rect 11188 18470 20811 18522
rect 20863 18470 20875 18522
rect 20927 18470 20939 18522
rect 20991 18470 21003 18522
rect 21055 18470 21067 18522
rect 21119 18470 30820 18522
rect 1104 18448 30820 18470
rect 10686 18368 10692 18420
rect 10744 18408 10750 18420
rect 12250 18408 12256 18420
rect 10744 18380 12256 18408
rect 10744 18368 10750 18380
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 12989 18411 13047 18417
rect 12989 18377 13001 18411
rect 13035 18408 13047 18411
rect 15473 18411 15531 18417
rect 13035 18380 15424 18408
rect 13035 18377 13047 18380
rect 12989 18371 13047 18377
rect 2682 18300 2688 18352
rect 2740 18340 2746 18352
rect 13078 18340 13084 18352
rect 2740 18312 13084 18340
rect 2740 18300 2746 18312
rect 13078 18300 13084 18312
rect 13136 18300 13142 18352
rect 15102 18300 15108 18352
rect 15160 18300 15166 18352
rect 7742 18272 7748 18284
rect 7703 18244 7748 18272
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 8018 18281 8024 18284
rect 8012 18235 8024 18281
rect 8076 18272 8082 18284
rect 11698 18272 11704 18284
rect 8076 18244 8112 18272
rect 11659 18244 11704 18272
rect 8018 18232 8024 18235
rect 8076 18232 8082 18244
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 12253 18275 12311 18281
rect 12253 18241 12265 18275
rect 12299 18241 12311 18275
rect 13170 18272 13176 18284
rect 13131 18244 13176 18272
rect 12253 18235 12311 18241
rect 10778 18164 10784 18216
rect 10836 18204 10842 18216
rect 12268 18204 12296 18235
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 14734 18272 14740 18284
rect 14695 18244 14740 18272
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 14925 18273 14983 18279
rect 14925 18239 14937 18273
rect 14971 18239 14983 18273
rect 14925 18233 14983 18239
rect 15013 18275 15071 18281
rect 15013 18241 15025 18275
rect 15059 18272 15071 18275
rect 15120 18272 15148 18300
rect 15286 18272 15292 18284
rect 15059 18244 15148 18272
rect 15247 18244 15292 18272
rect 15059 18241 15071 18244
rect 15013 18235 15071 18241
rect 10836 18176 12296 18204
rect 10836 18164 10842 18176
rect 9766 18096 9772 18148
rect 9824 18136 9830 18148
rect 13538 18136 13544 18148
rect 9824 18108 13544 18136
rect 9824 18096 9830 18108
rect 13538 18096 13544 18108
rect 13596 18136 13602 18148
rect 14936 18136 14964 18233
rect 15286 18232 15292 18244
rect 15344 18232 15350 18284
rect 15396 18272 15424 18380
rect 15473 18377 15485 18411
rect 15519 18408 15531 18411
rect 15562 18408 15568 18420
rect 15519 18380 15568 18408
rect 15519 18377 15531 18380
rect 15473 18371 15531 18377
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 16025 18411 16083 18417
rect 16025 18377 16037 18411
rect 16071 18408 16083 18411
rect 17126 18408 17132 18420
rect 16071 18380 17132 18408
rect 16071 18377 16083 18380
rect 16025 18371 16083 18377
rect 17126 18368 17132 18380
rect 17184 18368 17190 18420
rect 17678 18368 17684 18420
rect 17736 18408 17742 18420
rect 19061 18411 19119 18417
rect 19061 18408 19073 18411
rect 17736 18380 19073 18408
rect 17736 18368 17742 18380
rect 19061 18377 19073 18380
rect 19107 18377 19119 18411
rect 19061 18371 19119 18377
rect 20438 18368 20444 18420
rect 20496 18408 20502 18420
rect 21913 18411 21971 18417
rect 21913 18408 21925 18411
rect 20496 18380 21925 18408
rect 20496 18368 20502 18380
rect 21913 18377 21925 18380
rect 21959 18408 21971 18411
rect 22002 18408 22008 18420
rect 21959 18380 22008 18408
rect 21959 18377 21971 18380
rect 21913 18371 21971 18377
rect 22002 18368 22008 18380
rect 22060 18368 22066 18420
rect 24121 18411 24179 18417
rect 24121 18377 24133 18411
rect 24167 18408 24179 18411
rect 24210 18408 24216 18420
rect 24167 18380 24216 18408
rect 24167 18377 24179 18380
rect 24121 18371 24179 18377
rect 24210 18368 24216 18380
rect 24268 18368 24274 18420
rect 29730 18408 29736 18420
rect 24320 18380 29408 18408
rect 29691 18380 29736 18408
rect 16666 18340 16672 18352
rect 16627 18312 16672 18340
rect 16666 18300 16672 18312
rect 16724 18300 16730 18352
rect 18322 18340 18328 18352
rect 17696 18312 18328 18340
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 15396 18244 15945 18272
rect 15933 18241 15945 18244
rect 15979 18272 15991 18275
rect 16114 18272 16120 18284
rect 15979 18244 16120 18272
rect 15979 18241 15991 18244
rect 15933 18235 15991 18241
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16592 18244 16865 18272
rect 15102 18204 15108 18216
rect 15063 18176 15108 18204
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 16022 18164 16028 18216
rect 16080 18204 16086 18216
rect 16482 18204 16488 18216
rect 16080 18176 16488 18204
rect 16080 18164 16086 18176
rect 16482 18164 16488 18176
rect 16540 18204 16546 18216
rect 16592 18204 16620 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 16942 18232 16948 18284
rect 17000 18272 17006 18284
rect 17000 18244 17045 18272
rect 17000 18232 17006 18244
rect 17218 18232 17224 18284
rect 17276 18272 17282 18284
rect 17696 18281 17724 18312
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 19334 18300 19340 18352
rect 19392 18340 19398 18352
rect 24320 18340 24348 18380
rect 27614 18340 27620 18352
rect 19392 18312 24348 18340
rect 25056 18312 27620 18340
rect 19392 18300 19398 18312
rect 17954 18281 17960 18284
rect 17681 18275 17739 18281
rect 17276 18244 17369 18272
rect 17276 18232 17282 18244
rect 17681 18241 17693 18275
rect 17727 18241 17739 18275
rect 17948 18272 17960 18281
rect 17915 18244 17960 18272
rect 17681 18235 17739 18241
rect 17948 18235 17960 18244
rect 17954 18232 17960 18235
rect 18012 18232 18018 18284
rect 19788 18275 19846 18281
rect 19788 18241 19800 18275
rect 19834 18272 19846 18275
rect 20806 18272 20812 18284
rect 19834 18244 20812 18272
rect 19834 18241 19846 18244
rect 19788 18235 19846 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 21913 18275 21971 18281
rect 21913 18241 21925 18275
rect 21959 18272 21971 18275
rect 22005 18275 22063 18281
rect 22005 18272 22017 18275
rect 21959 18244 22017 18272
rect 21959 18241 21971 18244
rect 21913 18235 21971 18241
rect 22005 18241 22017 18244
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 22462 18232 22468 18284
rect 22520 18272 22526 18284
rect 22741 18275 22799 18281
rect 22741 18272 22753 18275
rect 22520 18244 22753 18272
rect 22520 18232 22526 18244
rect 22741 18241 22753 18244
rect 22787 18241 22799 18275
rect 22741 18235 22799 18241
rect 23106 18232 23112 18284
rect 23164 18272 23170 18284
rect 23382 18272 23388 18284
rect 23164 18244 23388 18272
rect 23164 18232 23170 18244
rect 23382 18232 23388 18244
rect 23440 18232 23446 18284
rect 23569 18275 23627 18281
rect 23569 18241 23581 18275
rect 23615 18272 23627 18275
rect 23842 18272 23848 18284
rect 23615 18244 23848 18272
rect 23615 18241 23627 18244
rect 23569 18235 23627 18241
rect 23842 18232 23848 18244
rect 23900 18232 23906 18284
rect 23934 18232 23940 18284
rect 23992 18272 23998 18284
rect 24946 18272 24952 18284
rect 23992 18244 24952 18272
rect 23992 18232 23998 18244
rect 24946 18232 24952 18244
rect 25004 18232 25010 18284
rect 25056 18281 25084 18312
rect 27614 18300 27620 18312
rect 27672 18300 27678 18352
rect 27982 18300 27988 18352
rect 28040 18340 28046 18352
rect 29086 18340 29092 18352
rect 28040 18312 29092 18340
rect 28040 18300 28046 18312
rect 29086 18300 29092 18312
rect 29144 18300 29150 18352
rect 29380 18294 29408 18380
rect 29730 18368 29736 18380
rect 29788 18368 29794 18420
rect 25041 18275 25099 18281
rect 25041 18241 25053 18275
rect 25087 18241 25099 18275
rect 25041 18235 25099 18241
rect 25308 18275 25366 18281
rect 25308 18241 25320 18275
rect 25354 18272 25366 18275
rect 27246 18272 27252 18284
rect 25354 18244 27252 18272
rect 25354 18241 25366 18244
rect 25308 18235 25366 18241
rect 27246 18232 27252 18244
rect 27304 18232 27310 18284
rect 27424 18275 27482 18281
rect 27424 18241 27436 18275
rect 27470 18272 27482 18275
rect 28350 18272 28356 18284
rect 27470 18244 28356 18272
rect 27470 18241 27482 18244
rect 27424 18235 27482 18241
rect 28350 18232 28356 18244
rect 28408 18232 28414 18284
rect 28718 18232 28724 18284
rect 28776 18272 28782 18284
rect 29196 18281 29408 18294
rect 28985 18275 29043 18281
rect 28985 18272 28997 18275
rect 28776 18244 28997 18272
rect 28776 18232 28782 18244
rect 28985 18241 28997 18244
rect 29031 18241 29043 18275
rect 28985 18235 29043 18241
rect 29181 18275 29408 18281
rect 29181 18241 29193 18275
rect 29227 18266 29408 18275
rect 29227 18241 29239 18266
rect 29181 18235 29239 18241
rect 29454 18232 29460 18284
rect 29512 18272 29518 18284
rect 29549 18275 29607 18281
rect 29549 18272 29561 18275
rect 29512 18244 29561 18272
rect 29512 18232 29518 18244
rect 29549 18241 29561 18244
rect 29595 18241 29607 18275
rect 29549 18235 29607 18241
rect 16540 18176 16620 18204
rect 16540 18164 16546 18176
rect 16758 18164 16764 18216
rect 16816 18204 16822 18216
rect 17236 18204 17264 18232
rect 16816 18176 17264 18204
rect 16816 18164 16822 18176
rect 19334 18164 19340 18216
rect 19392 18204 19398 18216
rect 19521 18207 19579 18213
rect 19521 18204 19533 18207
rect 19392 18176 19533 18204
rect 19392 18164 19398 18176
rect 19521 18173 19533 18176
rect 19567 18173 19579 18207
rect 19521 18167 19579 18173
rect 23198 18164 23204 18216
rect 23256 18204 23262 18216
rect 23661 18207 23719 18213
rect 23661 18204 23673 18207
rect 23256 18176 23673 18204
rect 23256 18164 23262 18176
rect 23661 18173 23673 18176
rect 23707 18173 23719 18207
rect 23661 18167 23719 18173
rect 23750 18164 23756 18216
rect 23808 18204 23814 18216
rect 27157 18207 27215 18213
rect 27157 18204 27169 18207
rect 23808 18176 23853 18204
rect 26068 18176 27169 18204
rect 23808 18164 23814 18176
rect 15746 18136 15752 18148
rect 13596 18108 14872 18136
rect 14936 18108 15752 18136
rect 13596 18096 13602 18108
rect 8386 18028 8392 18080
rect 8444 18068 8450 18080
rect 9125 18071 9183 18077
rect 9125 18068 9137 18071
rect 8444 18040 9137 18068
rect 8444 18028 8450 18040
rect 9125 18037 9137 18040
rect 9171 18037 9183 18071
rect 11514 18068 11520 18080
rect 11475 18040 11520 18068
rect 9125 18031 9183 18037
rect 11514 18028 11520 18040
rect 11572 18028 11578 18080
rect 11790 18028 11796 18080
rect 11848 18068 11854 18080
rect 12250 18068 12256 18080
rect 11848 18040 12256 18068
rect 11848 18028 11854 18040
rect 12250 18028 12256 18040
rect 12308 18028 12314 18080
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 14844 18068 14872 18108
rect 15746 18096 15752 18108
rect 15804 18096 15810 18148
rect 15838 18096 15844 18148
rect 15896 18096 15902 18148
rect 19426 18136 19432 18148
rect 18984 18108 19432 18136
rect 15102 18068 15108 18080
rect 12492 18040 12537 18068
rect 14844 18040 15108 18068
rect 12492 18028 12498 18040
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 15654 18028 15660 18080
rect 15712 18068 15718 18080
rect 15856 18068 15884 18096
rect 15712 18040 15884 18068
rect 17129 18071 17187 18077
rect 15712 18028 15718 18040
rect 17129 18037 17141 18071
rect 17175 18068 17187 18071
rect 18984 18068 19012 18108
rect 19426 18096 19432 18108
rect 19484 18096 19490 18148
rect 22925 18139 22983 18145
rect 22925 18105 22937 18139
rect 22971 18136 22983 18139
rect 23014 18136 23020 18148
rect 22971 18108 23020 18136
rect 22971 18105 22983 18108
rect 22925 18099 22983 18105
rect 23014 18096 23020 18108
rect 23072 18136 23078 18148
rect 23768 18136 23796 18164
rect 23072 18108 23796 18136
rect 23072 18096 23078 18108
rect 17175 18040 19012 18068
rect 20901 18071 20959 18077
rect 17175 18037 17187 18040
rect 17129 18031 17187 18037
rect 20901 18037 20913 18071
rect 20947 18068 20959 18071
rect 21174 18068 21180 18080
rect 20947 18040 21180 18068
rect 20947 18037 20959 18040
rect 20901 18031 20959 18037
rect 21174 18028 21180 18040
rect 21232 18068 21238 18080
rect 21450 18068 21456 18080
rect 21232 18040 21456 18068
rect 21232 18028 21238 18040
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 22097 18071 22155 18077
rect 22097 18037 22109 18071
rect 22143 18068 22155 18071
rect 22186 18068 22192 18080
rect 22143 18040 22192 18068
rect 22143 18037 22155 18040
rect 22097 18031 22155 18037
rect 22186 18028 22192 18040
rect 22244 18028 22250 18080
rect 24854 18028 24860 18080
rect 24912 18068 24918 18080
rect 26068 18068 26096 18176
rect 27157 18173 27169 18176
rect 27203 18173 27215 18207
rect 27157 18167 27215 18173
rect 28258 18164 28264 18216
rect 28316 18204 28322 18216
rect 29273 18207 29331 18213
rect 29273 18204 29285 18207
rect 28316 18176 29285 18204
rect 28316 18164 28322 18176
rect 29273 18173 29285 18176
rect 29319 18173 29331 18207
rect 29273 18167 29331 18173
rect 29365 18207 29423 18213
rect 29365 18173 29377 18207
rect 29411 18173 29423 18207
rect 29365 18167 29423 18173
rect 26326 18096 26332 18148
rect 26384 18136 26390 18148
rect 26421 18139 26479 18145
rect 26421 18136 26433 18139
rect 26384 18108 26433 18136
rect 26384 18096 26390 18108
rect 26421 18105 26433 18108
rect 26467 18105 26479 18139
rect 28534 18136 28540 18148
rect 28495 18108 28540 18136
rect 26421 18099 26479 18105
rect 24912 18040 26096 18068
rect 26436 18068 26464 18099
rect 28534 18096 28540 18108
rect 28592 18096 28598 18148
rect 29086 18096 29092 18148
rect 29144 18136 29150 18148
rect 29380 18136 29408 18167
rect 29144 18108 29408 18136
rect 29144 18096 29150 18108
rect 28074 18068 28080 18080
rect 26436 18040 28080 18068
rect 24912 18028 24918 18040
rect 28074 18028 28080 18040
rect 28132 18028 28138 18080
rect 1104 17978 30820 18000
rect 1104 17926 5915 17978
rect 5967 17926 5979 17978
rect 6031 17926 6043 17978
rect 6095 17926 6107 17978
rect 6159 17926 6171 17978
rect 6223 17926 15846 17978
rect 15898 17926 15910 17978
rect 15962 17926 15974 17978
rect 16026 17926 16038 17978
rect 16090 17926 16102 17978
rect 16154 17926 25776 17978
rect 25828 17926 25840 17978
rect 25892 17926 25904 17978
rect 25956 17926 25968 17978
rect 26020 17926 26032 17978
rect 26084 17926 30820 17978
rect 1104 17904 30820 17926
rect 8018 17824 8024 17876
rect 8076 17864 8082 17876
rect 8205 17867 8263 17873
rect 8205 17864 8217 17867
rect 8076 17836 8217 17864
rect 8076 17824 8082 17836
rect 8205 17833 8217 17836
rect 8251 17833 8263 17867
rect 12710 17864 12716 17876
rect 12671 17836 12716 17864
rect 8205 17827 8263 17833
rect 12710 17824 12716 17836
rect 12768 17824 12774 17876
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15746 17824 15752 17876
rect 15804 17864 15810 17876
rect 15841 17867 15899 17873
rect 15841 17864 15853 17867
rect 15804 17836 15853 17864
rect 15804 17824 15810 17836
rect 15841 17833 15853 17836
rect 15887 17833 15899 17867
rect 15841 17827 15899 17833
rect 15948 17836 20116 17864
rect 10045 17799 10103 17805
rect 10045 17765 10057 17799
rect 10091 17765 10103 17799
rect 10045 17759 10103 17765
rect 12621 17799 12679 17805
rect 12621 17765 12633 17799
rect 12667 17796 12679 17799
rect 15948 17796 15976 17836
rect 19518 17796 19524 17808
rect 12667 17768 15976 17796
rect 19479 17768 19524 17796
rect 12667 17765 12679 17768
rect 12621 17759 12679 17765
rect 10060 17728 10088 17759
rect 19518 17756 19524 17768
rect 19576 17756 19582 17808
rect 20088 17796 20116 17836
rect 20162 17824 20168 17876
rect 20220 17864 20226 17876
rect 20622 17864 20628 17876
rect 20220 17836 20628 17864
rect 20220 17824 20226 17836
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 20806 17864 20812 17876
rect 20767 17836 20812 17864
rect 20806 17824 20812 17836
rect 20864 17824 20870 17876
rect 21726 17824 21732 17876
rect 21784 17824 21790 17876
rect 22370 17864 22376 17876
rect 22331 17836 22376 17864
rect 22370 17824 22376 17836
rect 22428 17824 22434 17876
rect 22738 17864 22744 17876
rect 22480 17836 22744 17864
rect 21082 17796 21088 17808
rect 20088 17768 21088 17796
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 21174 17756 21180 17808
rect 21232 17796 21238 17808
rect 21542 17796 21548 17808
rect 21232 17768 21548 17796
rect 21232 17756 21238 17768
rect 21542 17756 21548 17768
rect 21600 17756 21606 17808
rect 8404 17700 10088 17728
rect 1578 17660 1584 17672
rect 1539 17632 1584 17660
rect 1578 17620 1584 17632
rect 1636 17620 1642 17672
rect 1762 17660 1768 17672
rect 1723 17632 1768 17660
rect 1762 17620 1768 17632
rect 1820 17620 1826 17672
rect 8404 17669 8432 17700
rect 11422 17688 11428 17740
rect 11480 17728 11486 17740
rect 11790 17728 11796 17740
rect 11480 17700 11796 17728
rect 11480 17688 11486 17700
rect 11790 17688 11796 17700
rect 11848 17688 11854 17740
rect 11882 17688 11888 17740
rect 11940 17728 11946 17740
rect 13354 17728 13360 17740
rect 11940 17700 13360 17728
rect 11940 17688 11946 17700
rect 13354 17688 13360 17700
rect 13412 17688 13418 17740
rect 14369 17731 14427 17737
rect 14369 17728 14381 17731
rect 14200 17700 14381 17728
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17629 8447 17663
rect 8389 17623 8447 17629
rect 9401 17663 9459 17669
rect 9401 17629 9413 17663
rect 9447 17660 9459 17663
rect 10226 17660 10232 17672
rect 9447 17632 10232 17660
rect 9447 17629 9459 17632
rect 9401 17623 9459 17629
rect 10226 17620 10232 17632
rect 10284 17620 10290 17672
rect 10689 17663 10747 17669
rect 10689 17629 10701 17663
rect 10735 17629 10747 17663
rect 10689 17623 10747 17629
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17660 10839 17663
rect 11238 17660 11244 17672
rect 10827 17632 11244 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 9674 17552 9680 17604
rect 9732 17592 9738 17604
rect 9886 17595 9944 17601
rect 9732 17564 9777 17592
rect 9732 17552 9738 17564
rect 9886 17561 9898 17595
rect 9932 17592 9944 17595
rect 10594 17592 10600 17604
rect 9932 17564 10600 17592
rect 9932 17561 9944 17564
rect 9886 17555 9944 17561
rect 10594 17552 10600 17564
rect 10652 17552 10658 17604
rect 10704 17592 10732 17623
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 11514 17620 11520 17672
rect 11572 17660 11578 17672
rect 11609 17663 11667 17669
rect 11609 17660 11621 17663
rect 11572 17632 11621 17660
rect 11572 17620 11578 17632
rect 11609 17629 11621 17632
rect 11655 17629 11667 17663
rect 11609 17623 11667 17629
rect 11701 17663 11759 17669
rect 11701 17629 11713 17663
rect 11747 17660 11759 17663
rect 12621 17663 12679 17669
rect 12621 17660 12633 17663
rect 11747 17632 12633 17660
rect 11747 17629 11759 17632
rect 11701 17623 11759 17629
rect 12621 17629 12633 17632
rect 12667 17629 12679 17663
rect 12621 17623 12679 17629
rect 13446 17620 13452 17672
rect 13504 17660 13510 17672
rect 14200 17660 14228 17700
rect 14369 17697 14381 17700
rect 14415 17697 14427 17731
rect 14369 17691 14427 17697
rect 14461 17731 14519 17737
rect 14461 17697 14473 17731
rect 14507 17728 14519 17731
rect 14642 17728 14648 17740
rect 14507 17700 14648 17728
rect 14507 17697 14519 17700
rect 14461 17691 14519 17697
rect 14642 17688 14648 17700
rect 14700 17688 14706 17740
rect 16390 17728 16396 17740
rect 16351 17700 16396 17728
rect 16390 17688 16396 17700
rect 16448 17688 16454 17740
rect 19242 17688 19248 17740
rect 19300 17728 19306 17740
rect 20346 17728 20352 17740
rect 19300 17700 20352 17728
rect 19300 17688 19306 17700
rect 13504 17632 14228 17660
rect 13504 17620 13510 17632
rect 14274 17620 14280 17672
rect 14332 17660 14338 17672
rect 14332 17632 14377 17660
rect 14332 17620 14338 17632
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 15194 17660 15200 17672
rect 14608 17632 14653 17660
rect 15155 17632 15200 17660
rect 14608 17620 14614 17632
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 16206 17660 16212 17672
rect 16167 17632 16212 17660
rect 16206 17620 16212 17632
rect 16264 17620 16270 17672
rect 17313 17663 17371 17669
rect 17313 17629 17325 17663
rect 17359 17660 17371 17663
rect 18322 17660 18328 17672
rect 17359 17632 18328 17660
rect 17359 17629 17371 17632
rect 17313 17623 17371 17629
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 20180 17669 20208 17700
rect 20346 17688 20352 17700
rect 20404 17688 20410 17740
rect 21450 17728 21456 17740
rect 20548 17700 21456 17728
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17629 19763 17663
rect 19705 17623 19763 17629
rect 20165 17663 20223 17669
rect 20165 17629 20177 17663
rect 20211 17629 20223 17663
rect 20165 17623 20223 17629
rect 20258 17663 20316 17669
rect 20258 17629 20270 17663
rect 20304 17629 20316 17663
rect 20258 17623 20316 17629
rect 20441 17663 20499 17669
rect 20441 17629 20453 17663
rect 20487 17662 20499 17663
rect 20548 17662 20576 17700
rect 21450 17688 21456 17700
rect 21508 17688 21514 17740
rect 21744 17672 21772 17824
rect 22002 17756 22008 17808
rect 22060 17796 22066 17808
rect 22480 17796 22508 17836
rect 22738 17824 22744 17836
rect 22796 17864 22802 17876
rect 23566 17864 23572 17876
rect 22796 17836 23244 17864
rect 23527 17836 23572 17864
rect 22796 17824 22802 17836
rect 22060 17768 22508 17796
rect 22060 17756 22066 17768
rect 22830 17756 22836 17808
rect 22888 17756 22894 17808
rect 21913 17731 21971 17737
rect 21913 17697 21925 17731
rect 21959 17728 21971 17731
rect 22848 17728 22876 17756
rect 23216 17737 23244 17836
rect 23566 17824 23572 17836
rect 23624 17824 23630 17876
rect 25314 17824 25320 17876
rect 25372 17864 25378 17876
rect 25593 17867 25651 17873
rect 25593 17864 25605 17867
rect 25372 17836 25605 17864
rect 25372 17824 25378 17836
rect 25593 17833 25605 17836
rect 25639 17833 25651 17867
rect 25593 17827 25651 17833
rect 25682 17824 25688 17876
rect 25740 17864 25746 17876
rect 26881 17867 26939 17873
rect 26881 17864 26893 17867
rect 25740 17836 26893 17864
rect 25740 17824 25746 17836
rect 26881 17833 26893 17836
rect 26927 17833 26939 17867
rect 26881 17827 26939 17833
rect 26436 17768 26556 17796
rect 23109 17731 23167 17737
rect 23109 17728 23121 17731
rect 21959 17700 23121 17728
rect 21959 17697 21971 17700
rect 21913 17691 21971 17697
rect 23109 17697 23121 17700
rect 23155 17697 23167 17731
rect 23109 17691 23167 17697
rect 23201 17731 23259 17737
rect 23201 17697 23213 17731
rect 23247 17728 23259 17731
rect 23566 17728 23572 17740
rect 23247 17700 23572 17728
rect 23247 17697 23259 17700
rect 23201 17691 23259 17697
rect 23566 17688 23572 17700
rect 23624 17688 23630 17740
rect 25590 17688 25596 17740
rect 25648 17728 25654 17740
rect 26436 17728 26464 17768
rect 26528 17737 26556 17768
rect 27614 17756 27620 17808
rect 27672 17796 27678 17808
rect 29454 17796 29460 17808
rect 27672 17768 29460 17796
rect 27672 17756 27678 17768
rect 29454 17756 29460 17768
rect 29512 17756 29518 17808
rect 25648 17700 26464 17728
rect 26513 17731 26571 17737
rect 25648 17688 25654 17700
rect 26513 17697 26525 17731
rect 26559 17697 26571 17731
rect 26970 17728 26976 17740
rect 26513 17691 26571 17697
rect 26620 17700 26976 17728
rect 20487 17634 20576 17662
rect 20487 17629 20499 17634
rect 20441 17623 20499 17629
rect 13081 17595 13139 17601
rect 10704 17564 11560 17592
rect 11532 17536 11560 17564
rect 13081 17561 13093 17595
rect 13127 17592 13139 17595
rect 17580 17595 17638 17601
rect 13127 17564 14136 17592
rect 13127 17561 13139 17564
rect 13081 17555 13139 17561
rect 1394 17484 1400 17536
rect 1452 17524 1458 17536
rect 1673 17527 1731 17533
rect 1673 17524 1685 17527
rect 1452 17496 1685 17524
rect 1452 17484 1458 17496
rect 1673 17493 1685 17496
rect 1719 17493 1731 17527
rect 1673 17487 1731 17493
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 11241 17527 11299 17533
rect 9824 17496 9869 17524
rect 9824 17484 9830 17496
rect 11241 17493 11253 17527
rect 11287 17524 11299 17527
rect 11330 17524 11336 17536
rect 11287 17496 11336 17524
rect 11287 17493 11299 17496
rect 11241 17487 11299 17493
rect 11330 17484 11336 17496
rect 11388 17484 11394 17536
rect 11514 17484 11520 17536
rect 11572 17484 11578 17536
rect 13173 17527 13231 17533
rect 13173 17493 13185 17527
rect 13219 17524 13231 17527
rect 13722 17524 13728 17536
rect 13219 17496 13728 17524
rect 13219 17493 13231 17496
rect 13173 17487 13231 17493
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 14108 17533 14136 17564
rect 17580 17561 17592 17595
rect 17626 17592 17638 17595
rect 18230 17592 18236 17604
rect 17626 17564 18236 17592
rect 17626 17561 17638 17564
rect 17580 17555 17638 17561
rect 18230 17552 18236 17564
rect 18288 17552 18294 17604
rect 14093 17527 14151 17533
rect 14093 17493 14105 17527
rect 14139 17493 14151 17527
rect 14093 17487 14151 17493
rect 16301 17527 16359 17533
rect 16301 17493 16313 17527
rect 16347 17524 16359 17527
rect 17126 17524 17132 17536
rect 16347 17496 17132 17524
rect 16347 17493 16359 17496
rect 16301 17487 16359 17493
rect 17126 17484 17132 17496
rect 17184 17484 17190 17536
rect 17862 17484 17868 17536
rect 17920 17524 17926 17536
rect 18693 17527 18751 17533
rect 18693 17524 18705 17527
rect 17920 17496 18705 17524
rect 17920 17484 17926 17496
rect 18693 17493 18705 17496
rect 18739 17493 18751 17527
rect 19720 17524 19748 17623
rect 20070 17552 20076 17604
rect 20128 17592 20134 17604
rect 20273 17592 20301 17623
rect 20622 17620 20628 17672
rect 20680 17669 20686 17672
rect 20680 17663 20707 17669
rect 20695 17629 20707 17663
rect 21634 17660 21640 17672
rect 21595 17632 21640 17660
rect 20680 17623 20707 17629
rect 20680 17620 20686 17623
rect 21634 17620 21640 17632
rect 21692 17620 21698 17672
rect 21726 17620 21732 17672
rect 21784 17620 21790 17672
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17629 21879 17663
rect 22002 17660 22008 17672
rect 21963 17632 22008 17660
rect 21821 17623 21879 17629
rect 20128 17564 20301 17592
rect 20541 17595 20599 17601
rect 20128 17552 20134 17564
rect 20541 17561 20553 17595
rect 20587 17592 20599 17595
rect 20806 17592 20812 17604
rect 20587 17564 20812 17592
rect 20587 17561 20599 17564
rect 20541 17555 20599 17561
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 21542 17552 21548 17604
rect 21600 17592 21606 17604
rect 21836 17592 21864 17623
rect 22002 17620 22008 17632
rect 22060 17620 22066 17672
rect 22186 17620 22192 17672
rect 22244 17660 22250 17672
rect 22830 17660 22836 17672
rect 22244 17632 22289 17660
rect 22791 17632 22836 17660
rect 22244 17620 22250 17632
rect 22830 17620 22836 17632
rect 22888 17620 22894 17672
rect 23385 17663 23443 17669
rect 23021 17657 23079 17663
rect 23021 17623 23033 17657
rect 23067 17654 23079 17657
rect 23067 17626 23152 17654
rect 23067 17623 23079 17626
rect 23021 17617 23079 17623
rect 21600 17564 21864 17592
rect 23124 17592 23152 17626
rect 23385 17629 23397 17663
rect 23431 17660 23443 17663
rect 24210 17660 24216 17672
rect 23431 17632 24216 17660
rect 23431 17629 23443 17632
rect 23385 17623 23443 17629
rect 24210 17620 24216 17632
rect 24268 17620 24274 17672
rect 24397 17663 24455 17669
rect 24397 17629 24409 17663
rect 24443 17629 24455 17663
rect 24397 17623 24455 17629
rect 25501 17663 25559 17669
rect 25501 17629 25513 17663
rect 25547 17660 25559 17663
rect 26050 17660 26056 17672
rect 25547 17632 26056 17660
rect 25547 17629 25559 17632
rect 25501 17623 25559 17629
rect 23658 17592 23664 17604
rect 23124 17564 23664 17592
rect 21600 17552 21606 17564
rect 23658 17552 23664 17564
rect 23716 17552 23722 17604
rect 24412 17592 24440 17623
rect 26050 17620 26056 17632
rect 26108 17620 26114 17672
rect 26145 17663 26203 17669
rect 26145 17629 26157 17663
rect 26191 17629 26203 17663
rect 26333 17663 26391 17669
rect 26333 17660 26345 17663
rect 26145 17623 26203 17629
rect 26252 17632 26345 17660
rect 25038 17592 25044 17604
rect 24412 17564 25044 17592
rect 21266 17524 21272 17536
rect 19720 17496 21272 17524
rect 18693 17487 18751 17493
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 23106 17484 23112 17536
rect 23164 17524 23170 17536
rect 24412 17524 24440 17564
rect 25038 17552 25044 17564
rect 25096 17552 25102 17604
rect 23164 17496 24440 17524
rect 24489 17527 24547 17533
rect 23164 17484 23170 17496
rect 24489 17493 24501 17527
rect 24535 17524 24547 17527
rect 24946 17524 24952 17536
rect 24535 17496 24952 17524
rect 24535 17493 24547 17496
rect 24489 17487 24547 17493
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 26160 17524 26188 17623
rect 26252 17592 26280 17632
rect 26333 17629 26345 17632
rect 26379 17629 26391 17663
rect 26333 17623 26391 17629
rect 26421 17663 26479 17669
rect 26421 17629 26433 17663
rect 26467 17658 26479 17663
rect 26620 17660 26648 17700
rect 26970 17688 26976 17700
rect 27028 17688 27034 17740
rect 27522 17728 27528 17740
rect 27483 17700 27528 17728
rect 27522 17688 27528 17700
rect 27580 17688 27586 17740
rect 27801 17731 27859 17737
rect 27801 17697 27813 17731
rect 27847 17728 27859 17731
rect 27982 17728 27988 17740
rect 27847 17700 27988 17728
rect 27847 17697 27859 17700
rect 27801 17691 27859 17697
rect 27982 17688 27988 17700
rect 28040 17688 28046 17740
rect 28810 17688 28816 17740
rect 28868 17728 28874 17740
rect 28868 17700 30144 17728
rect 28868 17688 28874 17700
rect 26528 17658 26648 17660
rect 26467 17632 26648 17658
rect 26697 17663 26755 17669
rect 26467 17630 26556 17632
rect 26467 17629 26479 17630
rect 26421 17623 26479 17629
rect 26697 17629 26709 17663
rect 26743 17660 26755 17663
rect 27614 17660 27620 17672
rect 26743 17632 27620 17660
rect 26743 17629 26755 17632
rect 26697 17623 26755 17629
rect 27614 17620 27620 17632
rect 27672 17620 27678 17672
rect 28534 17620 28540 17672
rect 28592 17660 28598 17672
rect 30116 17669 30144 17700
rect 28997 17663 29055 17669
rect 28997 17660 29009 17663
rect 28592 17632 29009 17660
rect 28592 17620 28598 17632
rect 28997 17629 29009 17632
rect 29043 17629 29055 17663
rect 28997 17623 29055 17629
rect 30101 17663 30159 17669
rect 30101 17629 30113 17663
rect 30147 17629 30159 17663
rect 30101 17623 30159 17629
rect 26252 17564 26464 17592
rect 26436 17536 26464 17564
rect 28350 17552 28356 17604
rect 28408 17592 28414 17604
rect 28408 17564 29960 17592
rect 28408 17552 28414 17564
rect 26326 17524 26332 17536
rect 26160 17496 26332 17524
rect 26326 17484 26332 17496
rect 26384 17484 26390 17536
rect 26418 17484 26424 17536
rect 26476 17484 26482 17536
rect 27890 17484 27896 17536
rect 27948 17524 27954 17536
rect 29932 17533 29960 17564
rect 28813 17527 28871 17533
rect 28813 17524 28825 17527
rect 27948 17496 28825 17524
rect 27948 17484 27954 17496
rect 28813 17493 28825 17496
rect 28859 17493 28871 17527
rect 28813 17487 28871 17493
rect 29917 17527 29975 17533
rect 29917 17493 29929 17527
rect 29963 17493 29975 17527
rect 29917 17487 29975 17493
rect 1104 17434 30820 17456
rect 1104 17382 10880 17434
rect 10932 17382 10944 17434
rect 10996 17382 11008 17434
rect 11060 17382 11072 17434
rect 11124 17382 11136 17434
rect 11188 17382 20811 17434
rect 20863 17382 20875 17434
rect 20927 17382 20939 17434
rect 20991 17382 21003 17434
rect 21055 17382 21067 17434
rect 21119 17382 30820 17434
rect 1104 17360 30820 17382
rect 1578 17280 1584 17332
rect 1636 17320 1642 17332
rect 1636 17292 10548 17320
rect 1636 17280 1642 17292
rect 1394 17184 1400 17196
rect 1355 17156 1400 17184
rect 1394 17144 1400 17156
rect 1452 17144 1458 17196
rect 1486 17144 1492 17196
rect 1544 17184 1550 17196
rect 2133 17187 2191 17193
rect 2133 17184 2145 17187
rect 1544 17156 2145 17184
rect 1544 17144 1550 17156
rect 2133 17153 2145 17156
rect 2179 17184 2191 17187
rect 8386 17184 8392 17196
rect 2179 17156 8392 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17184 8815 17187
rect 9306 17184 9312 17196
rect 8803 17156 9312 17184
rect 8803 17153 8815 17156
rect 8757 17147 8815 17153
rect 9306 17144 9312 17156
rect 9364 17144 9370 17196
rect 9033 17119 9091 17125
rect 9033 17085 9045 17119
rect 9079 17116 9091 17119
rect 10410 17116 10416 17128
rect 9079 17088 10416 17116
rect 9079 17085 9091 17088
rect 9033 17079 9091 17085
rect 10410 17076 10416 17088
rect 10468 17076 10474 17128
rect 10520 17116 10548 17292
rect 11698 17280 11704 17332
rect 11756 17320 11762 17332
rect 11977 17323 12035 17329
rect 11977 17320 11989 17323
rect 11756 17292 11989 17320
rect 11756 17280 11762 17292
rect 11977 17289 11989 17292
rect 12023 17289 12035 17323
rect 11977 17283 12035 17289
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 13722 17320 13728 17332
rect 12492 17292 12537 17320
rect 13683 17292 13728 17320
rect 12492 17280 12498 17292
rect 13722 17280 13728 17292
rect 13780 17280 13786 17332
rect 14185 17323 14243 17329
rect 14185 17289 14197 17323
rect 14231 17320 14243 17323
rect 15378 17320 15384 17332
rect 14231 17292 15384 17320
rect 14231 17289 14243 17292
rect 14185 17283 14243 17289
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 15470 17280 15476 17332
rect 15528 17320 15534 17332
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 15528 17292 15577 17320
rect 15528 17280 15534 17292
rect 15565 17289 15577 17292
rect 15611 17289 15623 17323
rect 17126 17320 17132 17332
rect 17087 17292 17132 17320
rect 15565 17283 15623 17289
rect 17126 17280 17132 17292
rect 17184 17320 17190 17332
rect 17957 17323 18015 17329
rect 17957 17320 17969 17323
rect 17184 17292 17969 17320
rect 17184 17280 17190 17292
rect 17957 17289 17969 17292
rect 18003 17289 18015 17323
rect 17957 17283 18015 17289
rect 20717 17323 20775 17329
rect 20717 17289 20729 17323
rect 20763 17320 20775 17323
rect 21634 17320 21640 17332
rect 20763 17292 21640 17320
rect 20763 17289 20775 17292
rect 20717 17283 20775 17289
rect 21634 17280 21640 17292
rect 21692 17280 21698 17332
rect 21726 17280 21732 17332
rect 21784 17320 21790 17332
rect 21784 17292 24808 17320
rect 21784 17280 21790 17292
rect 11790 17212 11796 17264
rect 11848 17252 11854 17264
rect 16758 17252 16764 17264
rect 11848 17224 14320 17252
rect 11848 17212 11854 17224
rect 12345 17187 12403 17193
rect 12345 17153 12357 17187
rect 12391 17184 12403 17187
rect 12391 17156 12664 17184
rect 12391 17153 12403 17156
rect 12345 17147 12403 17153
rect 12636 17128 12664 17156
rect 13446 17144 13452 17196
rect 13504 17184 13510 17196
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 13504 17156 14105 17184
rect 13504 17144 13510 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 12529 17119 12587 17125
rect 10520 17088 12434 17116
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 1854 16940 1860 16992
rect 1912 16980 1918 16992
rect 2225 16983 2283 16989
rect 2225 16980 2237 16983
rect 1912 16952 2237 16980
rect 1912 16940 1918 16952
rect 2225 16949 2237 16952
rect 2271 16980 2283 16983
rect 9766 16980 9772 16992
rect 2271 16952 9772 16980
rect 2271 16949 2283 16952
rect 2225 16943 2283 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 10137 16983 10195 16989
rect 10137 16980 10149 16983
rect 9916 16952 10149 16980
rect 9916 16940 9922 16952
rect 10137 16949 10149 16952
rect 10183 16949 10195 16983
rect 10137 16943 10195 16949
rect 10502 16940 10508 16992
rect 10560 16980 10566 16992
rect 11606 16980 11612 16992
rect 10560 16952 11612 16980
rect 10560 16940 10566 16952
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 12406 16980 12434 17088
rect 12529 17085 12541 17119
rect 12575 17085 12587 17119
rect 12529 17079 12587 17085
rect 12544 17048 12572 17079
rect 12618 17076 12624 17128
rect 12676 17076 12682 17128
rect 14292 17125 14320 17224
rect 16040 17224 16764 17252
rect 14366 17144 14372 17196
rect 14424 17184 14430 17196
rect 14921 17187 14979 17193
rect 14921 17184 14933 17187
rect 14424 17156 14933 17184
rect 14424 17144 14430 17156
rect 14921 17153 14933 17156
rect 14967 17153 14979 17187
rect 15746 17184 15752 17196
rect 15707 17156 15752 17184
rect 14921 17147 14979 17153
rect 15746 17144 15752 17156
rect 15804 17144 15810 17196
rect 15841 17187 15899 17193
rect 15841 17153 15853 17187
rect 15887 17184 15899 17187
rect 16040 17184 16068 17224
rect 16758 17212 16764 17224
rect 16816 17212 16822 17264
rect 17034 17252 17040 17264
rect 16995 17224 17040 17252
rect 17034 17212 17040 17224
rect 17092 17212 17098 17264
rect 21913 17255 21971 17261
rect 21913 17252 21925 17255
rect 21376 17224 21925 17252
rect 15887 17156 16068 17184
rect 16117 17187 16175 17193
rect 15887 17153 15899 17156
rect 15841 17147 15899 17153
rect 16117 17153 16129 17187
rect 16163 17184 16175 17187
rect 16666 17184 16672 17196
rect 16163 17156 16672 17184
rect 16163 17153 16175 17156
rect 16117 17147 16175 17153
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 17862 17184 17868 17196
rect 17823 17156 17868 17184
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 19426 17184 19432 17196
rect 19387 17156 19432 17184
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 20073 17187 20131 17193
rect 20073 17184 20085 17187
rect 19996 17156 20085 17184
rect 19996 17128 20024 17156
rect 20073 17153 20085 17156
rect 20119 17153 20131 17187
rect 20898 17184 20904 17196
rect 20859 17156 20904 17184
rect 20073 17147 20131 17153
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 20990 17144 20996 17196
rect 21048 17184 21054 17196
rect 21269 17187 21327 17193
rect 21048 17156 21093 17184
rect 21048 17144 21054 17156
rect 21269 17153 21281 17187
rect 21315 17182 21327 17187
rect 21376 17182 21404 17224
rect 21913 17221 21925 17224
rect 21959 17221 21971 17255
rect 23198 17252 23204 17264
rect 21913 17215 21971 17221
rect 22848 17224 23204 17252
rect 21315 17154 21404 17182
rect 21315 17153 21327 17154
rect 21269 17147 21327 17153
rect 21450 17144 21456 17196
rect 21508 17184 21514 17196
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 21508 17156 21833 17184
rect 21508 17144 21514 17156
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 22370 17144 22376 17196
rect 22428 17184 22434 17196
rect 22848 17193 22876 17224
rect 23198 17212 23204 17224
rect 23256 17212 23262 17264
rect 23293 17255 23351 17261
rect 23293 17221 23305 17255
rect 23339 17252 23351 17255
rect 23998 17255 24056 17261
rect 23998 17252 24010 17255
rect 23339 17224 24010 17252
rect 23339 17221 23351 17224
rect 23293 17215 23351 17221
rect 23998 17221 24010 17224
rect 24044 17221 24056 17255
rect 24780 17252 24808 17292
rect 25038 17280 25044 17332
rect 25096 17320 25102 17332
rect 25133 17323 25191 17329
rect 25133 17320 25145 17323
rect 25096 17292 25145 17320
rect 25096 17280 25102 17292
rect 25133 17289 25145 17292
rect 25179 17289 25191 17323
rect 25133 17283 25191 17289
rect 26234 17280 26240 17332
rect 26292 17320 26298 17332
rect 26329 17323 26387 17329
rect 26329 17320 26341 17323
rect 26292 17292 26341 17320
rect 26292 17280 26298 17292
rect 26329 17289 26341 17292
rect 26375 17289 26387 17323
rect 26329 17283 26387 17289
rect 27246 17280 27252 17332
rect 27304 17320 27310 17332
rect 28077 17323 28135 17329
rect 28077 17320 28089 17323
rect 27304 17292 28089 17320
rect 27304 17280 27310 17292
rect 28077 17289 28089 17292
rect 28123 17289 28135 17323
rect 28077 17283 28135 17289
rect 24780 17224 27568 17252
rect 23998 17215 24056 17221
rect 22557 17187 22615 17193
rect 22557 17184 22569 17187
rect 22428 17156 22569 17184
rect 22428 17144 22434 17156
rect 22557 17153 22569 17156
rect 22603 17153 22615 17187
rect 22557 17147 22615 17153
rect 22741 17187 22799 17193
rect 22741 17153 22753 17187
rect 22787 17153 22799 17187
rect 22741 17147 22799 17153
rect 22833 17187 22891 17193
rect 22833 17153 22845 17187
rect 22879 17153 22891 17187
rect 23106 17184 23112 17196
rect 23067 17156 23112 17184
rect 22833 17147 22891 17153
rect 14277 17119 14335 17125
rect 14277 17085 14289 17119
rect 14323 17085 14335 17119
rect 16850 17116 16856 17128
rect 14277 17079 14335 17085
rect 14384 17088 16856 17116
rect 12710 17048 12716 17060
rect 12544 17020 12716 17048
rect 12710 17008 12716 17020
rect 12768 17008 12774 17060
rect 14384 16980 14412 17088
rect 16850 17076 16856 17088
rect 16908 17076 16914 17128
rect 17313 17119 17371 17125
rect 17313 17085 17325 17119
rect 17359 17116 17371 17119
rect 17494 17116 17500 17128
rect 17359 17088 17500 17116
rect 17359 17085 17371 17088
rect 17313 17079 17371 17085
rect 17494 17076 17500 17088
rect 17552 17076 17558 17128
rect 19978 17076 19984 17128
rect 20036 17076 20042 17128
rect 21174 17116 21180 17128
rect 21135 17088 21180 17116
rect 21174 17076 21180 17088
rect 21232 17076 21238 17128
rect 22462 17076 22468 17128
rect 22520 17116 22526 17128
rect 22756 17116 22784 17147
rect 23106 17144 23112 17156
rect 23164 17144 23170 17196
rect 25498 17144 25504 17196
rect 25556 17184 25562 17196
rect 26237 17187 26295 17193
rect 26237 17184 26249 17187
rect 25556 17156 26249 17184
rect 25556 17144 25562 17156
rect 26237 17153 26249 17156
rect 26283 17153 26295 17187
rect 26237 17147 26295 17153
rect 27154 17144 27160 17196
rect 27212 17184 27218 17196
rect 27540 17193 27568 17224
rect 27341 17187 27399 17193
rect 27341 17184 27353 17187
rect 27212 17156 27353 17184
rect 27212 17144 27218 17156
rect 27341 17153 27353 17156
rect 27387 17153 27399 17187
rect 27341 17147 27399 17153
rect 27525 17187 27583 17193
rect 27525 17153 27537 17187
rect 27571 17153 27583 17187
rect 27525 17147 27583 17153
rect 27893 17187 27951 17193
rect 27893 17153 27905 17187
rect 27939 17184 27951 17187
rect 28074 17184 28080 17196
rect 27939 17156 28080 17184
rect 27939 17153 27951 17156
rect 27893 17147 27951 17153
rect 28074 17144 28080 17156
rect 28132 17144 28138 17196
rect 28442 17144 28448 17196
rect 28500 17184 28506 17196
rect 28629 17187 28687 17193
rect 28629 17184 28641 17187
rect 28500 17156 28641 17184
rect 28500 17144 28506 17156
rect 28629 17153 28641 17156
rect 28675 17153 28687 17187
rect 28629 17147 28687 17153
rect 28718 17144 28724 17196
rect 28776 17184 28782 17196
rect 28885 17187 28943 17193
rect 28885 17184 28897 17187
rect 28776 17156 28897 17184
rect 28776 17144 28782 17156
rect 28885 17153 28897 17156
rect 28931 17153 28943 17187
rect 28885 17147 28943 17153
rect 22520 17088 22784 17116
rect 22925 17119 22983 17125
rect 22520 17076 22526 17088
rect 22925 17085 22937 17119
rect 22971 17116 22983 17119
rect 23014 17116 23020 17128
rect 22971 17088 23020 17116
rect 22971 17085 22983 17088
rect 22925 17079 22983 17085
rect 23014 17076 23020 17088
rect 23072 17076 23078 17128
rect 23750 17116 23756 17128
rect 23711 17088 23756 17116
rect 23750 17076 23756 17088
rect 23808 17076 23814 17128
rect 27430 17076 27436 17128
rect 27488 17116 27494 17128
rect 27617 17119 27675 17125
rect 27617 17116 27629 17119
rect 27488 17088 27629 17116
rect 27488 17076 27494 17088
rect 27617 17085 27629 17088
rect 27663 17085 27675 17119
rect 27617 17079 27675 17085
rect 27709 17119 27767 17125
rect 27709 17085 27721 17119
rect 27755 17116 27767 17119
rect 27982 17116 27988 17128
rect 27755 17088 27988 17116
rect 27755 17085 27767 17088
rect 27709 17079 27767 17085
rect 27982 17076 27988 17088
rect 28040 17076 28046 17128
rect 15930 17008 15936 17060
rect 15988 17048 15994 17060
rect 16669 17051 16727 17057
rect 16669 17048 16681 17051
rect 15988 17020 16681 17048
rect 15988 17008 15994 17020
rect 16669 17017 16681 17020
rect 16715 17017 16727 17051
rect 16669 17011 16727 17017
rect 20165 17051 20223 17057
rect 20165 17017 20177 17051
rect 20211 17048 20223 17051
rect 21634 17048 21640 17060
rect 20211 17020 21640 17048
rect 20211 17017 20223 17020
rect 20165 17011 20223 17017
rect 21634 17008 21640 17020
rect 21692 17008 21698 17060
rect 22370 17008 22376 17060
rect 22428 17048 22434 17060
rect 23382 17048 23388 17060
rect 22428 17020 23388 17048
rect 22428 17008 22434 17020
rect 23382 17008 23388 17020
rect 23440 17008 23446 17060
rect 15010 16980 15016 16992
rect 12406 16952 14412 16980
rect 14971 16952 15016 16980
rect 15010 16940 15016 16952
rect 15068 16940 15074 16992
rect 15654 16940 15660 16992
rect 15712 16980 15718 16992
rect 16025 16983 16083 16989
rect 16025 16980 16037 16983
rect 15712 16952 16037 16980
rect 15712 16940 15718 16952
rect 16025 16949 16037 16952
rect 16071 16949 16083 16983
rect 16025 16943 16083 16949
rect 19521 16983 19579 16989
rect 19521 16949 19533 16983
rect 19567 16980 19579 16983
rect 20346 16980 20352 16992
rect 19567 16952 20352 16980
rect 19567 16949 19579 16952
rect 19521 16943 19579 16949
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 20898 16940 20904 16992
rect 20956 16980 20962 16992
rect 21726 16980 21732 16992
rect 20956 16952 21732 16980
rect 20956 16940 20962 16952
rect 21726 16940 21732 16952
rect 21784 16940 21790 16992
rect 25682 16940 25688 16992
rect 25740 16980 25746 16992
rect 29270 16980 29276 16992
rect 25740 16952 29276 16980
rect 25740 16940 25746 16952
rect 29270 16940 29276 16952
rect 29328 16940 29334 16992
rect 29546 16940 29552 16992
rect 29604 16980 29610 16992
rect 30009 16983 30067 16989
rect 30009 16980 30021 16983
rect 29604 16952 30021 16980
rect 29604 16940 29610 16952
rect 30009 16949 30021 16952
rect 30055 16949 30067 16983
rect 30009 16943 30067 16949
rect 1104 16890 30820 16912
rect 1104 16838 5915 16890
rect 5967 16838 5979 16890
rect 6031 16838 6043 16890
rect 6095 16838 6107 16890
rect 6159 16838 6171 16890
rect 6223 16838 15846 16890
rect 15898 16838 15910 16890
rect 15962 16838 15974 16890
rect 16026 16838 16038 16890
rect 16090 16838 16102 16890
rect 16154 16838 25776 16890
rect 25828 16838 25840 16890
rect 25892 16838 25904 16890
rect 25956 16838 25968 16890
rect 26020 16838 26032 16890
rect 26084 16838 30820 16890
rect 1104 16816 30820 16838
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10410 16776 10416 16788
rect 9916 16748 10272 16776
rect 10371 16748 10416 16776
rect 9916 16736 9922 16748
rect 9950 16640 9956 16652
rect 9911 16612 9956 16640
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10244 16640 10272 16748
rect 10410 16736 10416 16748
rect 10468 16736 10474 16788
rect 10686 16736 10692 16788
rect 10744 16776 10750 16788
rect 11790 16776 11796 16788
rect 10744 16748 11796 16776
rect 10744 16736 10750 16748
rect 11790 16736 11796 16748
rect 11848 16736 11854 16788
rect 13446 16776 13452 16788
rect 13407 16748 13452 16776
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 14734 16736 14740 16788
rect 14792 16776 14798 16788
rect 15657 16779 15715 16785
rect 15657 16776 15669 16779
rect 14792 16748 15669 16776
rect 14792 16736 14798 16748
rect 15657 16745 15669 16748
rect 15703 16745 15715 16779
rect 23106 16776 23112 16788
rect 15657 16739 15715 16745
rect 18156 16748 23112 16776
rect 11606 16668 11612 16720
rect 11664 16708 11670 16720
rect 12710 16708 12716 16720
rect 11664 16680 12716 16708
rect 11664 16668 11670 16680
rect 12710 16668 12716 16680
rect 12768 16708 12774 16720
rect 12768 16680 14780 16708
rect 12768 16668 12774 16680
rect 10778 16640 10784 16652
rect 10244 16612 10784 16640
rect 10778 16600 10784 16612
rect 10836 16640 10842 16652
rect 11330 16640 11336 16652
rect 10836 16612 11008 16640
rect 11291 16612 11336 16640
rect 10836 16600 10842 16612
rect 9674 16572 9680 16584
rect 9635 16544 9680 16572
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 9858 16572 9864 16584
rect 9819 16544 9864 16572
rect 9858 16532 9864 16544
rect 9916 16532 9922 16584
rect 10045 16575 10103 16581
rect 10045 16541 10057 16575
rect 10091 16572 10103 16575
rect 10134 16572 10140 16584
rect 10091 16544 10140 16572
rect 10091 16541 10103 16544
rect 10045 16535 10103 16541
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 10229 16575 10287 16581
rect 10229 16541 10241 16575
rect 10275 16572 10287 16575
rect 10275 16544 10916 16572
rect 10275 16541 10287 16544
rect 10229 16535 10287 16541
rect 9692 16504 9720 16532
rect 10502 16504 10508 16516
rect 9692 16476 10508 16504
rect 10502 16464 10508 16476
rect 10560 16464 10566 16516
rect 10888 16445 10916 16544
rect 10980 16504 11008 16612
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16640 11575 16643
rect 11882 16640 11888 16652
rect 11563 16612 11888 16640
rect 11563 16609 11575 16612
rect 11517 16603 11575 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16640 12127 16643
rect 12434 16640 12440 16652
rect 12115 16612 12440 16640
rect 12115 16609 12127 16612
rect 12069 16603 12127 16609
rect 12434 16600 12440 16612
rect 12492 16600 12498 16652
rect 12618 16640 12624 16652
rect 12579 16612 12624 16640
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 14090 16600 14096 16652
rect 14148 16640 14154 16652
rect 14752 16649 14780 16680
rect 15378 16668 15384 16720
rect 15436 16708 15442 16720
rect 18156 16708 18184 16748
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 23293 16779 23351 16785
rect 23293 16745 23305 16779
rect 23339 16776 23351 16779
rect 23474 16776 23480 16788
rect 23339 16748 23480 16776
rect 23339 16745 23351 16748
rect 23293 16739 23351 16745
rect 23474 16736 23480 16748
rect 23532 16736 23538 16788
rect 24302 16736 24308 16788
rect 24360 16776 24366 16788
rect 24397 16779 24455 16785
rect 24397 16776 24409 16779
rect 24360 16748 24409 16776
rect 24360 16736 24366 16748
rect 24397 16745 24409 16748
rect 24443 16745 24455 16779
rect 24397 16739 24455 16745
rect 26513 16779 26571 16785
rect 26513 16745 26525 16779
rect 26559 16776 26571 16779
rect 27522 16776 27528 16788
rect 26559 16748 27528 16776
rect 26559 16745 26571 16748
rect 26513 16739 26571 16745
rect 27522 16736 27528 16748
rect 27580 16736 27586 16788
rect 27801 16779 27859 16785
rect 27801 16745 27813 16779
rect 27847 16776 27859 16779
rect 28718 16776 28724 16788
rect 27847 16748 28724 16776
rect 27847 16745 27859 16748
rect 27801 16739 27859 16745
rect 28718 16736 28724 16748
rect 28776 16736 28782 16788
rect 28997 16779 29055 16785
rect 28997 16745 29009 16779
rect 29043 16776 29055 16779
rect 29362 16776 29368 16788
rect 29043 16748 29368 16776
rect 29043 16745 29055 16748
rect 28997 16739 29055 16745
rect 29362 16736 29368 16748
rect 29420 16736 29426 16788
rect 15436 16680 18184 16708
rect 21085 16711 21143 16717
rect 15436 16668 15442 16680
rect 21085 16677 21097 16711
rect 21131 16708 21143 16711
rect 21131 16680 22600 16708
rect 21131 16677 21143 16680
rect 21085 16671 21143 16677
rect 14553 16643 14611 16649
rect 14553 16640 14565 16643
rect 14148 16612 14565 16640
rect 14148 16600 14154 16612
rect 14553 16609 14565 16612
rect 14599 16609 14611 16643
rect 14553 16603 14611 16609
rect 14737 16643 14795 16649
rect 14737 16609 14749 16643
rect 14783 16640 14795 16643
rect 16574 16640 16580 16652
rect 14783 16612 16580 16640
rect 14783 16609 14795 16612
rect 14737 16603 14795 16609
rect 16574 16600 16580 16612
rect 16632 16600 16638 16652
rect 19245 16643 19303 16649
rect 19245 16609 19257 16643
rect 19291 16640 19303 16643
rect 19291 16612 19380 16640
rect 19291 16609 19303 16612
rect 19245 16603 19303 16609
rect 19352 16584 19380 16612
rect 20346 16600 20352 16652
rect 20404 16640 20410 16652
rect 20404 16612 20944 16640
rect 20404 16600 20410 16612
rect 11238 16572 11244 16584
rect 11199 16544 11244 16572
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 12253 16575 12311 16581
rect 12253 16541 12265 16575
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 13449 16575 13507 16581
rect 13449 16541 13461 16575
rect 13495 16541 13507 16575
rect 15286 16572 15292 16584
rect 15247 16544 15292 16572
rect 13449 16535 13507 16541
rect 12268 16504 12296 16535
rect 10980 16476 12296 16504
rect 10873 16439 10931 16445
rect 10873 16405 10885 16439
rect 10919 16405 10931 16439
rect 10873 16399 10931 16405
rect 12253 16439 12311 16445
rect 12253 16405 12265 16439
rect 12299 16436 12311 16439
rect 12434 16436 12440 16448
rect 12299 16408 12440 16436
rect 12299 16405 12311 16408
rect 12253 16399 12311 16405
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 13464 16436 13492 16535
rect 15286 16532 15292 16544
rect 15344 16532 15350 16584
rect 15930 16532 15936 16584
rect 15988 16572 15994 16584
rect 16482 16572 16488 16584
rect 15988 16544 16488 16572
rect 15988 16532 15994 16544
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 19334 16572 19340 16584
rect 19247 16544 19340 16572
rect 19334 16532 19340 16544
rect 19392 16572 19398 16584
rect 19886 16572 19892 16584
rect 19392 16544 19892 16572
rect 19392 16532 19398 16544
rect 19886 16532 19892 16544
rect 19944 16532 19950 16584
rect 15378 16464 15384 16516
rect 15436 16504 15442 16516
rect 19518 16513 19524 16516
rect 15473 16507 15531 16513
rect 15473 16504 15485 16507
rect 15436 16476 15485 16504
rect 15436 16464 15442 16476
rect 15473 16473 15485 16476
rect 15519 16473 15531 16507
rect 19512 16504 19524 16513
rect 19479 16476 19524 16504
rect 15473 16467 15531 16473
rect 19512 16467 19524 16476
rect 19518 16464 19524 16467
rect 19576 16464 19582 16516
rect 20916 16504 20944 16612
rect 20990 16600 20996 16652
rect 21048 16640 21054 16652
rect 21048 16612 21404 16640
rect 21048 16600 21054 16612
rect 21266 16572 21272 16584
rect 21227 16544 21272 16572
rect 21266 16532 21272 16544
rect 21324 16532 21330 16584
rect 21376 16581 21404 16612
rect 21450 16600 21456 16652
rect 21508 16640 21514 16652
rect 21545 16643 21603 16649
rect 21545 16640 21557 16643
rect 21508 16612 21557 16640
rect 21508 16600 21514 16612
rect 21545 16609 21557 16612
rect 21591 16609 21603 16643
rect 21545 16603 21603 16609
rect 21361 16575 21419 16581
rect 21361 16541 21373 16575
rect 21407 16541 21419 16575
rect 21634 16572 21640 16584
rect 21595 16544 21640 16572
rect 21361 16535 21419 16541
rect 21174 16504 21180 16516
rect 19628 16476 20760 16504
rect 20916 16476 21180 16504
rect 14090 16436 14096 16448
rect 13464 16408 14096 16436
rect 14090 16396 14096 16408
rect 14148 16396 14154 16448
rect 14461 16439 14519 16445
rect 14461 16405 14473 16439
rect 14507 16436 14519 16439
rect 15010 16436 15016 16448
rect 14507 16408 15016 16436
rect 14507 16405 14519 16408
rect 14461 16399 14519 16405
rect 15010 16396 15016 16408
rect 15068 16396 15074 16448
rect 18506 16396 18512 16448
rect 18564 16436 18570 16448
rect 19628 16436 19656 16476
rect 18564 16408 19656 16436
rect 18564 16396 18570 16408
rect 20346 16396 20352 16448
rect 20404 16436 20410 16448
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20404 16408 20637 16436
rect 20404 16396 20410 16408
rect 20625 16405 20637 16408
rect 20671 16405 20683 16439
rect 20732 16436 20760 16476
rect 21174 16464 21180 16476
rect 21232 16464 21238 16516
rect 21376 16504 21404 16535
rect 21634 16532 21640 16544
rect 21692 16532 21698 16584
rect 22572 16581 22600 16680
rect 22738 16668 22744 16720
rect 22796 16668 22802 16720
rect 23382 16668 23388 16720
rect 23440 16708 23446 16720
rect 27430 16708 27436 16720
rect 23440 16680 24716 16708
rect 23440 16668 23446 16680
rect 22756 16640 22784 16668
rect 22833 16643 22891 16649
rect 22833 16640 22845 16643
rect 22756 16612 22845 16640
rect 22833 16609 22845 16612
rect 22879 16609 22891 16643
rect 22833 16603 22891 16609
rect 22925 16643 22983 16649
rect 22925 16609 22937 16643
rect 22971 16640 22983 16643
rect 23566 16640 23572 16652
rect 22971 16612 23572 16640
rect 22971 16609 22983 16612
rect 22925 16603 22983 16609
rect 22557 16575 22615 16581
rect 22557 16541 22569 16575
rect 22603 16541 22615 16575
rect 22738 16572 22744 16584
rect 22699 16544 22744 16572
rect 22557 16535 22615 16541
rect 22738 16532 22744 16544
rect 22796 16532 22802 16584
rect 23106 16572 23112 16584
rect 23067 16544 23112 16572
rect 23106 16532 23112 16544
rect 23164 16532 23170 16584
rect 22278 16504 22284 16516
rect 21376 16476 22284 16504
rect 22278 16464 22284 16476
rect 22336 16504 22342 16516
rect 23382 16504 23388 16516
rect 22336 16476 23388 16504
rect 22336 16464 22342 16476
rect 23382 16464 23388 16476
rect 23440 16464 23446 16516
rect 23492 16504 23520 16612
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 24302 16600 24308 16652
rect 24360 16640 24366 16652
rect 24360 16612 24624 16640
rect 24360 16600 24366 16612
rect 24596 16581 24624 16612
rect 24688 16581 24716 16680
rect 27356 16680 27436 16708
rect 27356 16649 27384 16680
rect 27430 16668 27436 16680
rect 27488 16668 27494 16720
rect 27614 16668 27620 16720
rect 27672 16708 27678 16720
rect 28074 16708 28080 16720
rect 27672 16680 28080 16708
rect 27672 16668 27678 16680
rect 28074 16668 28080 16680
rect 28132 16668 28138 16720
rect 28258 16668 28264 16720
rect 28316 16708 28322 16720
rect 28316 16680 28764 16708
rect 28316 16668 28322 16680
rect 24857 16643 24915 16649
rect 24857 16640 24869 16643
rect 24771 16612 24869 16640
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 24673 16575 24731 16581
rect 24673 16541 24685 16575
rect 24719 16541 24731 16575
rect 24673 16535 24731 16541
rect 24771 16504 24799 16612
rect 24857 16609 24869 16612
rect 24903 16609 24915 16643
rect 24857 16603 24915 16609
rect 27341 16643 27399 16649
rect 27341 16609 27353 16643
rect 27387 16609 27399 16643
rect 27982 16640 27988 16652
rect 27341 16603 27399 16609
rect 27448 16612 27988 16640
rect 24946 16572 24952 16584
rect 24907 16544 24952 16572
rect 24946 16532 24952 16544
rect 25004 16532 25010 16584
rect 25682 16572 25688 16584
rect 25643 16544 25688 16572
rect 25682 16532 25688 16544
rect 25740 16532 25746 16584
rect 26329 16575 26387 16581
rect 26329 16541 26341 16575
rect 26375 16572 26387 16575
rect 27065 16575 27123 16581
rect 26375 16544 26556 16572
rect 26375 16541 26387 16544
rect 26329 16535 26387 16541
rect 23492 16476 24799 16504
rect 25777 16507 25835 16513
rect 25777 16473 25789 16507
rect 25823 16504 25835 16507
rect 26418 16504 26424 16516
rect 25823 16476 26424 16504
rect 25823 16473 25835 16476
rect 25777 16467 25835 16473
rect 26418 16464 26424 16476
rect 26476 16464 26482 16516
rect 24118 16436 24124 16448
rect 20732 16408 24124 16436
rect 20625 16399 20683 16405
rect 24118 16396 24124 16408
rect 24176 16396 24182 16448
rect 26528 16436 26556 16544
rect 27065 16541 27077 16575
rect 27111 16572 27123 16575
rect 27154 16572 27160 16584
rect 27111 16544 27160 16572
rect 27111 16541 27123 16544
rect 27065 16535 27123 16541
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 27246 16532 27252 16584
rect 27304 16572 27310 16584
rect 27448 16581 27476 16612
rect 27982 16600 27988 16612
rect 28040 16640 28046 16652
rect 28629 16643 28687 16649
rect 28629 16640 28641 16643
rect 28040 16612 28641 16640
rect 28040 16600 28046 16612
rect 28629 16609 28641 16612
rect 28675 16609 28687 16643
rect 28629 16603 28687 16609
rect 27433 16575 27491 16581
rect 27304 16544 27349 16572
rect 27304 16532 27310 16544
rect 27433 16541 27445 16575
rect 27479 16541 27491 16575
rect 27433 16535 27491 16541
rect 27617 16575 27675 16581
rect 27617 16541 27629 16575
rect 27663 16541 27675 16575
rect 28258 16572 28264 16584
rect 28219 16544 28264 16572
rect 27617 16535 27675 16541
rect 27338 16436 27344 16448
rect 26528 16408 27344 16436
rect 27338 16396 27344 16408
rect 27396 16396 27402 16448
rect 27632 16436 27660 16535
rect 28258 16532 28264 16544
rect 28316 16532 28322 16584
rect 28445 16575 28503 16581
rect 28445 16541 28457 16575
rect 28491 16541 28503 16575
rect 28445 16535 28503 16541
rect 28537 16575 28595 16581
rect 28537 16541 28549 16575
rect 28583 16572 28595 16575
rect 28736 16572 28764 16680
rect 28994 16600 29000 16652
rect 29052 16640 29058 16652
rect 29052 16612 29592 16640
rect 29052 16600 29058 16612
rect 28583 16544 28764 16572
rect 28813 16575 28871 16581
rect 28583 16541 28595 16544
rect 28537 16535 28595 16541
rect 28813 16541 28825 16575
rect 28859 16572 28871 16575
rect 29178 16572 29184 16584
rect 28859 16544 29184 16572
rect 28859 16541 28871 16544
rect 28813 16535 28871 16541
rect 28460 16504 28488 16535
rect 29178 16532 29184 16544
rect 29236 16532 29242 16584
rect 29564 16581 29592 16612
rect 29549 16575 29607 16581
rect 29549 16541 29561 16575
rect 29595 16541 29607 16575
rect 29549 16535 29607 16541
rect 29822 16504 29828 16516
rect 28460 16476 29828 16504
rect 29822 16464 29828 16476
rect 29880 16464 29886 16516
rect 29546 16436 29552 16448
rect 27632 16408 29552 16436
rect 29546 16396 29552 16408
rect 29604 16396 29610 16448
rect 29638 16396 29644 16448
rect 29696 16436 29702 16448
rect 29696 16408 29741 16436
rect 29696 16396 29702 16408
rect 1104 16346 30820 16368
rect 1104 16294 10880 16346
rect 10932 16294 10944 16346
rect 10996 16294 11008 16346
rect 11060 16294 11072 16346
rect 11124 16294 11136 16346
rect 11188 16294 20811 16346
rect 20863 16294 20875 16346
rect 20927 16294 20939 16346
rect 20991 16294 21003 16346
rect 21055 16294 21067 16346
rect 21119 16294 30820 16346
rect 1104 16272 30820 16294
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 11974 16232 11980 16244
rect 11388 16204 11980 16232
rect 11388 16192 11394 16204
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 12069 16235 12127 16241
rect 12069 16201 12081 16235
rect 12115 16201 12127 16235
rect 15102 16232 15108 16244
rect 12069 16195 12127 16201
rect 13648 16204 15108 16232
rect 12084 16164 12112 16195
rect 10612 16136 12112 16164
rect 10612 16105 10640 16136
rect 10597 16099 10655 16105
rect 10597 16065 10609 16099
rect 10643 16065 10655 16099
rect 10597 16059 10655 16065
rect 10689 16099 10747 16105
rect 10689 16065 10701 16099
rect 10735 16065 10747 16099
rect 10689 16059 10747 16065
rect 10965 16099 11023 16105
rect 10965 16065 10977 16099
rect 11011 16065 11023 16099
rect 10965 16059 11023 16065
rect 10318 15988 10324 16040
rect 10376 16028 10382 16040
rect 10704 16028 10732 16059
rect 10376 16000 10732 16028
rect 10980 16028 11008 16059
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 13648 16105 13676 16204
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 15378 16232 15384 16244
rect 15339 16204 15384 16232
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 15749 16235 15807 16241
rect 15749 16201 15761 16235
rect 15795 16232 15807 16235
rect 17034 16232 17040 16244
rect 15795 16204 17040 16232
rect 15795 16201 15807 16204
rect 15749 16195 15807 16201
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 19518 16232 19524 16244
rect 19479 16204 19524 16232
rect 19518 16192 19524 16204
rect 19576 16192 19582 16244
rect 20346 16232 20352 16244
rect 19628 16204 20352 16232
rect 13722 16124 13728 16176
rect 13780 16164 13786 16176
rect 17957 16167 18015 16173
rect 17957 16164 17969 16167
rect 13780 16136 17969 16164
rect 13780 16124 13786 16136
rect 17957 16133 17969 16136
rect 18003 16133 18015 16167
rect 17957 16127 18015 16133
rect 18046 16124 18052 16176
rect 18104 16164 18110 16176
rect 19628 16164 19656 16204
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 21821 16235 21879 16241
rect 21821 16201 21833 16235
rect 21867 16232 21879 16235
rect 22830 16232 22836 16244
rect 21867 16204 22836 16232
rect 21867 16201 21879 16204
rect 21821 16195 21879 16201
rect 22830 16192 22836 16204
rect 22888 16192 22894 16244
rect 23106 16232 23112 16244
rect 23067 16204 23112 16232
rect 23106 16192 23112 16204
rect 23164 16192 23170 16244
rect 24118 16192 24124 16244
rect 24176 16232 24182 16244
rect 24305 16235 24363 16241
rect 24305 16232 24317 16235
rect 24176 16204 24317 16232
rect 24176 16192 24182 16204
rect 24305 16201 24317 16204
rect 24351 16201 24363 16235
rect 24305 16195 24363 16201
rect 27154 16192 27160 16244
rect 27212 16232 27218 16244
rect 28258 16232 28264 16244
rect 27212 16204 28264 16232
rect 27212 16192 27218 16204
rect 28258 16192 28264 16204
rect 28316 16192 28322 16244
rect 18104 16136 19656 16164
rect 18104 16124 18110 16136
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 11756 16068 12449 16096
rect 11756 16056 11762 16068
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16096 12587 16099
rect 13633 16099 13691 16105
rect 12575 16068 13584 16096
rect 12575 16065 12587 16068
rect 12529 16059 12587 16065
rect 11882 16028 11888 16040
rect 10980 16000 11888 16028
rect 10376 15988 10382 16000
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 12713 16031 12771 16037
rect 12713 15997 12725 16031
rect 12759 16028 12771 16031
rect 13354 16028 13360 16040
rect 12759 16000 13360 16028
rect 12759 15997 12771 16000
rect 12713 15991 12771 15997
rect 13354 15988 13360 16000
rect 13412 15988 13418 16040
rect 13556 16028 13584 16068
rect 13633 16065 13645 16099
rect 13679 16065 13691 16099
rect 13814 16096 13820 16108
rect 13775 16068 13820 16096
rect 13633 16059 13691 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16065 13967 16099
rect 14182 16096 14188 16108
rect 14143 16068 14188 16096
rect 13909 16059 13967 16065
rect 13722 16028 13728 16040
rect 13556 16000 13728 16028
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 13924 16028 13952 16059
rect 14182 16056 14188 16068
rect 14240 16056 14246 16108
rect 15841 16099 15899 16105
rect 15841 16065 15853 16099
rect 15887 16096 15899 16099
rect 16942 16096 16948 16108
rect 15887 16068 16948 16096
rect 15887 16065 15899 16068
rect 15841 16059 15899 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16096 17923 16099
rect 18506 16096 18512 16108
rect 17911 16068 18512 16096
rect 17911 16065 17923 16068
rect 17865 16059 17923 16065
rect 18506 16056 18512 16068
rect 18564 16056 18570 16108
rect 18782 16096 18788 16108
rect 18743 16068 18788 16096
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 18969 16099 19027 16105
rect 18969 16065 18981 16099
rect 19015 16065 19027 16099
rect 18969 16059 19027 16065
rect 15930 16028 15936 16040
rect 13832 16000 15936 16028
rect 10413 15963 10471 15969
rect 10413 15929 10425 15963
rect 10459 15960 10471 15963
rect 11698 15960 11704 15972
rect 10459 15932 11704 15960
rect 10459 15929 10471 15932
rect 10413 15923 10471 15929
rect 11698 15920 11704 15932
rect 11756 15920 11762 15972
rect 12526 15920 12532 15972
rect 12584 15960 12590 15972
rect 13832 15960 13860 16000
rect 15930 15988 15936 16000
rect 15988 15988 15994 16040
rect 16025 16031 16083 16037
rect 16025 15997 16037 16031
rect 16071 15997 16083 16031
rect 16025 15991 16083 15997
rect 12584 15932 13860 15960
rect 14001 15963 14059 15969
rect 12584 15920 12590 15932
rect 14001 15929 14013 15963
rect 14047 15960 14059 15963
rect 14550 15960 14556 15972
rect 14047 15932 14556 15960
rect 14047 15929 14059 15932
rect 14001 15923 14059 15929
rect 14550 15920 14556 15932
rect 14608 15920 14614 15972
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 10873 15895 10931 15901
rect 10873 15892 10885 15895
rect 10560 15864 10885 15892
rect 10560 15852 10566 15864
rect 10873 15861 10885 15864
rect 10919 15892 10931 15895
rect 12986 15892 12992 15904
rect 10919 15864 12992 15892
rect 10919 15861 10931 15864
rect 10873 15855 10931 15861
rect 12986 15852 12992 15864
rect 13044 15852 13050 15904
rect 14093 15895 14151 15901
rect 14093 15861 14105 15895
rect 14139 15892 14151 15895
rect 14918 15892 14924 15904
rect 14139 15864 14924 15892
rect 14139 15861 14151 15864
rect 14093 15855 14151 15861
rect 14918 15852 14924 15864
rect 14976 15852 14982 15904
rect 16040 15892 16068 15991
rect 16390 15988 16396 16040
rect 16448 16028 16454 16040
rect 17129 16031 17187 16037
rect 17129 16028 17141 16031
rect 16448 16000 17141 16028
rect 16448 15988 16454 16000
rect 17129 15997 17141 16000
rect 17175 15997 17187 16031
rect 17129 15991 17187 15997
rect 17313 16031 17371 16037
rect 17313 15997 17325 16031
rect 17359 16028 17371 16031
rect 17494 16028 17500 16040
rect 17359 16000 17500 16028
rect 17359 15997 17371 16000
rect 17313 15991 17371 15997
rect 16666 15960 16672 15972
rect 16627 15932 16672 15960
rect 16666 15920 16672 15932
rect 16724 15920 16730 15972
rect 16574 15892 16580 15904
rect 16040 15864 16580 15892
rect 16574 15852 16580 15864
rect 16632 15892 16638 15904
rect 17328 15892 17356 15991
rect 17494 15988 17500 16000
rect 17552 15988 17558 16040
rect 18984 16028 19012 16059
rect 19058 16056 19064 16108
rect 19116 16096 19122 16108
rect 19352 16105 19380 16136
rect 19702 16124 19708 16176
rect 19760 16164 19766 16176
rect 21085 16167 21143 16173
rect 21085 16164 21097 16167
rect 19760 16136 21097 16164
rect 19760 16124 19766 16136
rect 21085 16133 21097 16136
rect 21131 16133 21143 16167
rect 21085 16127 21143 16133
rect 21174 16124 21180 16176
rect 21232 16164 21238 16176
rect 27338 16164 27344 16176
rect 21232 16136 22416 16164
rect 21232 16124 21238 16136
rect 19337 16099 19395 16105
rect 19116 16068 19161 16096
rect 19116 16056 19122 16068
rect 19337 16065 19349 16099
rect 19383 16065 19395 16099
rect 20346 16096 20352 16108
rect 20307 16068 20352 16096
rect 19337 16059 19395 16065
rect 20346 16056 20352 16068
rect 20404 16056 20410 16108
rect 21634 16056 21640 16108
rect 21692 16096 21698 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21692 16068 22017 16096
rect 21692 16056 21698 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 22097 16099 22155 16105
rect 22097 16065 22109 16099
rect 22143 16096 22155 16099
rect 22186 16096 22192 16108
rect 22143 16068 22192 16096
rect 22143 16065 22155 16068
rect 22097 16059 22155 16065
rect 22186 16056 22192 16068
rect 22244 16056 22250 16108
rect 22388 16105 22416 16136
rect 24136 16136 27344 16164
rect 22373 16099 22431 16105
rect 22373 16065 22385 16099
rect 22419 16065 22431 16099
rect 22373 16059 22431 16065
rect 23017 16099 23075 16105
rect 23017 16065 23029 16099
rect 23063 16096 23075 16099
rect 23382 16096 23388 16108
rect 23063 16068 23388 16096
rect 23063 16065 23075 16068
rect 23017 16059 23075 16065
rect 23382 16056 23388 16068
rect 23440 16056 23446 16108
rect 24136 16105 24164 16136
rect 27338 16124 27344 16136
rect 27396 16124 27402 16176
rect 27614 16124 27620 16176
rect 27672 16164 27678 16176
rect 28966 16167 29024 16173
rect 28966 16164 28978 16167
rect 27672 16136 28978 16164
rect 27672 16124 27678 16136
rect 28966 16133 28978 16136
rect 29012 16133 29024 16167
rect 28966 16127 29024 16133
rect 29638 16124 29644 16176
rect 29696 16124 29702 16176
rect 25130 16105 25136 16108
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16065 24179 16099
rect 24121 16059 24179 16065
rect 25124 16059 25136 16105
rect 25188 16096 25194 16108
rect 27433 16099 27491 16105
rect 25188 16068 25224 16096
rect 25130 16056 25136 16059
rect 25188 16056 25194 16068
rect 27433 16065 27445 16099
rect 27479 16096 27491 16099
rect 27522 16096 27528 16108
rect 27479 16068 27528 16096
rect 27479 16065 27491 16068
rect 27433 16059 27491 16065
rect 27522 16056 27528 16068
rect 27580 16056 27586 16108
rect 27632 16068 28396 16096
rect 19153 16031 19211 16037
rect 18984 16000 19104 16028
rect 19076 15960 19104 16000
rect 19153 15997 19165 16031
rect 19199 16028 19211 16031
rect 19610 16028 19616 16040
rect 19199 16000 19616 16028
rect 19199 15997 19211 16000
rect 19153 15991 19211 15997
rect 19610 15988 19616 16000
rect 19668 15988 19674 16040
rect 20438 15988 20444 16040
rect 20496 16028 20502 16040
rect 21358 16028 21364 16040
rect 20496 16000 21364 16028
rect 20496 15988 20502 16000
rect 21358 15988 21364 16000
rect 21416 15988 21422 16040
rect 21450 15988 21456 16040
rect 21508 16028 21514 16040
rect 22281 16031 22339 16037
rect 22281 16028 22293 16031
rect 21508 16000 22293 16028
rect 21508 15988 21514 16000
rect 22281 15997 22293 16000
rect 22327 15997 22339 16031
rect 22281 15991 22339 15997
rect 23750 15988 23756 16040
rect 23808 16028 23814 16040
rect 24854 16028 24860 16040
rect 23808 16000 24860 16028
rect 23808 15988 23814 16000
rect 24854 15988 24860 16000
rect 24912 15988 24918 16040
rect 26142 15988 26148 16040
rect 26200 16028 26206 16040
rect 27632 16028 27660 16068
rect 26200 16000 27660 16028
rect 27709 16031 27767 16037
rect 26200 15988 26206 16000
rect 27709 15997 27721 16031
rect 27755 16028 27767 16031
rect 27982 16028 27988 16040
rect 27755 16000 27988 16028
rect 27755 15997 27767 16000
rect 27709 15991 27767 15997
rect 27982 15988 27988 16000
rect 28040 15988 28046 16040
rect 28368 16028 28396 16068
rect 28442 16056 28448 16108
rect 28500 16096 28506 16108
rect 28721 16099 28779 16105
rect 28721 16096 28733 16099
rect 28500 16068 28733 16096
rect 28500 16056 28506 16068
rect 28721 16065 28733 16068
rect 28767 16065 28779 16099
rect 29656 16096 29684 16124
rect 28721 16059 28779 16065
rect 28828 16068 29684 16096
rect 28828 16028 28856 16068
rect 28368 16000 28856 16028
rect 19518 15960 19524 15972
rect 19076 15932 19524 15960
rect 19518 15920 19524 15932
rect 19576 15960 19582 15972
rect 19978 15960 19984 15972
rect 19576 15932 19984 15960
rect 19576 15920 19582 15932
rect 19978 15920 19984 15932
rect 20036 15920 20042 15972
rect 28074 15920 28080 15972
rect 28132 15960 28138 15972
rect 28258 15960 28264 15972
rect 28132 15932 28264 15960
rect 28132 15920 28138 15932
rect 28258 15920 28264 15932
rect 28316 15920 28322 15972
rect 16632 15864 17356 15892
rect 16632 15852 16638 15864
rect 19886 15852 19892 15904
rect 19944 15892 19950 15904
rect 20441 15895 20499 15901
rect 20441 15892 20453 15895
rect 19944 15864 20453 15892
rect 19944 15852 19950 15864
rect 20441 15861 20453 15864
rect 20487 15861 20499 15895
rect 21174 15892 21180 15904
rect 21135 15864 21180 15892
rect 20441 15855 20499 15861
rect 21174 15852 21180 15864
rect 21232 15852 21238 15904
rect 22370 15852 22376 15904
rect 22428 15892 22434 15904
rect 22830 15892 22836 15904
rect 22428 15864 22836 15892
rect 22428 15852 22434 15864
rect 22830 15852 22836 15864
rect 22888 15852 22894 15904
rect 26142 15852 26148 15904
rect 26200 15892 26206 15904
rect 26237 15895 26295 15901
rect 26237 15892 26249 15895
rect 26200 15864 26249 15892
rect 26200 15852 26206 15864
rect 26237 15861 26249 15864
rect 26283 15861 26295 15895
rect 26237 15855 26295 15861
rect 27246 15852 27252 15904
rect 27304 15892 27310 15904
rect 30101 15895 30159 15901
rect 30101 15892 30113 15895
rect 27304 15864 30113 15892
rect 27304 15852 27310 15864
rect 30101 15861 30113 15864
rect 30147 15861 30159 15895
rect 30101 15855 30159 15861
rect 1104 15802 30820 15824
rect 1104 15750 5915 15802
rect 5967 15750 5979 15802
rect 6031 15750 6043 15802
rect 6095 15750 6107 15802
rect 6159 15750 6171 15802
rect 6223 15750 15846 15802
rect 15898 15750 15910 15802
rect 15962 15750 15974 15802
rect 16026 15750 16038 15802
rect 16090 15750 16102 15802
rect 16154 15750 25776 15802
rect 25828 15750 25840 15802
rect 25892 15750 25904 15802
rect 25956 15750 25968 15802
rect 26020 15750 26032 15802
rect 26084 15750 30820 15802
rect 1104 15728 30820 15750
rect 11241 15691 11299 15697
rect 11241 15657 11253 15691
rect 11287 15688 11299 15691
rect 11514 15688 11520 15700
rect 11287 15660 11520 15688
rect 11287 15657 11299 15660
rect 11241 15651 11299 15657
rect 11514 15648 11520 15660
rect 11572 15648 11578 15700
rect 11974 15648 11980 15700
rect 12032 15688 12038 15700
rect 13541 15691 13599 15697
rect 13541 15688 13553 15691
rect 12032 15660 13553 15688
rect 12032 15648 12038 15660
rect 13541 15657 13553 15660
rect 13587 15657 13599 15691
rect 14182 15688 14188 15700
rect 14143 15660 14188 15688
rect 13541 15651 13599 15657
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 18506 15688 18512 15700
rect 18467 15660 18512 15688
rect 18506 15648 18512 15660
rect 18564 15688 18570 15700
rect 19058 15688 19064 15700
rect 18564 15660 19064 15688
rect 18564 15648 18570 15660
rect 19058 15648 19064 15660
rect 19116 15648 19122 15700
rect 23750 15688 23756 15700
rect 20916 15660 23756 15688
rect 10594 15580 10600 15632
rect 10652 15620 10658 15632
rect 11609 15623 11667 15629
rect 10652 15592 11560 15620
rect 10652 15580 10658 15592
rect 2682 15552 2688 15564
rect 1596 15524 2688 15552
rect 1596 15493 1624 15524
rect 2682 15512 2688 15524
rect 2740 15512 2746 15564
rect 11532 15561 11560 15592
rect 11609 15589 11621 15623
rect 11655 15620 11667 15623
rect 12434 15620 12440 15632
rect 11655 15592 12440 15620
rect 11655 15589 11667 15592
rect 11609 15583 11667 15589
rect 12434 15580 12440 15592
rect 12492 15620 12498 15632
rect 13262 15620 13268 15632
rect 12492 15592 13268 15620
rect 12492 15580 12498 15592
rect 13262 15580 13268 15592
rect 13320 15580 13326 15632
rect 13354 15580 13360 15632
rect 13412 15620 13418 15632
rect 16298 15620 16304 15632
rect 13412 15592 16304 15620
rect 13412 15580 13418 15592
rect 11517 15555 11575 15561
rect 11517 15521 11529 15555
rect 11563 15521 11575 15555
rect 11517 15515 11575 15521
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 13081 15555 13139 15561
rect 13081 15552 13093 15555
rect 12759 15524 13093 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 13081 15521 13093 15524
rect 13127 15552 13139 15555
rect 13906 15552 13912 15564
rect 13127 15524 13912 15552
rect 13127 15521 13139 15524
rect 13081 15515 13139 15521
rect 13906 15512 13912 15524
rect 13964 15512 13970 15564
rect 14844 15561 14872 15592
rect 16298 15580 16304 15592
rect 16356 15580 16362 15632
rect 14829 15555 14887 15561
rect 14829 15521 14841 15555
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 16025 15555 16083 15561
rect 16025 15521 16037 15555
rect 16071 15552 16083 15555
rect 16574 15552 16580 15564
rect 16071 15524 16580 15552
rect 16071 15521 16083 15524
rect 16025 15515 16083 15521
rect 16574 15512 16580 15524
rect 16632 15512 16638 15564
rect 18230 15512 18236 15564
rect 18288 15552 18294 15564
rect 19150 15552 19156 15564
rect 18288 15524 19156 15552
rect 18288 15512 18294 15524
rect 19150 15512 19156 15524
rect 19208 15552 19214 15564
rect 20916 15561 20944 15660
rect 23750 15648 23756 15660
rect 23808 15648 23814 15700
rect 25130 15648 25136 15700
rect 25188 15688 25194 15700
rect 25317 15691 25375 15697
rect 25317 15688 25329 15691
rect 25188 15660 25329 15688
rect 25188 15648 25194 15660
rect 25317 15657 25329 15660
rect 25363 15657 25375 15691
rect 25317 15651 25375 15657
rect 28166 15648 28172 15700
rect 28224 15688 28230 15700
rect 28629 15691 28687 15697
rect 28629 15688 28641 15691
rect 28224 15660 28641 15688
rect 28224 15648 28230 15660
rect 28629 15657 28641 15660
rect 28675 15657 28687 15691
rect 28629 15651 28687 15657
rect 23014 15580 23020 15632
rect 23072 15620 23078 15632
rect 28074 15620 28080 15632
rect 23072 15592 23152 15620
rect 27987 15592 28080 15620
rect 23072 15580 23078 15592
rect 19521 15555 19579 15561
rect 19521 15552 19533 15555
rect 19208 15524 19533 15552
rect 19208 15512 19214 15524
rect 19521 15521 19533 15524
rect 19567 15521 19579 15555
rect 19521 15515 19579 15521
rect 20901 15555 20959 15561
rect 20901 15521 20913 15555
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 22278 15512 22284 15564
rect 22336 15552 22342 15564
rect 23124 15561 23152 15592
rect 28074 15580 28080 15592
rect 28132 15620 28138 15632
rect 28902 15620 28908 15632
rect 28132 15592 28908 15620
rect 28132 15580 28138 15592
rect 28902 15580 28908 15592
rect 28960 15580 28966 15632
rect 23109 15555 23167 15561
rect 22336 15524 22968 15552
rect 22336 15512 22342 15524
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15453 1639 15487
rect 1762 15484 1768 15496
rect 1723 15456 1768 15484
rect 1581 15447 1639 15453
rect 1762 15444 1768 15456
rect 1820 15444 1826 15496
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 10042 15484 10048 15496
rect 9916 15456 10048 15484
rect 9916 15444 9922 15456
rect 10042 15444 10048 15456
rect 10100 15484 10106 15496
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 10100 15456 10609 15484
rect 10100 15444 10106 15456
rect 10597 15453 10609 15456
rect 10643 15453 10655 15487
rect 11422 15484 11428 15496
rect 11383 15456 11428 15484
rect 10597 15447 10655 15453
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 11698 15484 11704 15496
rect 11659 15456 11704 15484
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15484 11943 15487
rect 11974 15484 11980 15496
rect 11931 15456 11980 15484
rect 11931 15453 11943 15456
rect 11885 15447 11943 15453
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 12802 15484 12808 15496
rect 12763 15456 12808 15484
rect 12802 15444 12808 15456
rect 12860 15444 12866 15496
rect 12986 15484 12992 15496
rect 12947 15456 12992 15484
rect 12986 15444 12992 15456
rect 13044 15444 13050 15496
rect 13173 15487 13231 15493
rect 13173 15484 13185 15487
rect 13096 15456 13185 15484
rect 10781 15419 10839 15425
rect 10781 15385 10793 15419
rect 10827 15416 10839 15419
rect 13096 15416 13124 15456
rect 13173 15453 13185 15456
rect 13219 15453 13231 15487
rect 13354 15484 13360 15496
rect 13315 15456 13360 15484
rect 13173 15447 13231 15453
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 14090 15444 14096 15496
rect 14148 15484 14154 15496
rect 14553 15487 14611 15493
rect 14553 15484 14565 15487
rect 14148 15456 14565 15484
rect 14148 15444 14154 15456
rect 14553 15453 14565 15456
rect 14599 15453 14611 15487
rect 15654 15484 15660 15496
rect 14553 15447 14611 15453
rect 14936 15456 15660 15484
rect 14936 15416 14964 15456
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 17126 15484 17132 15496
rect 17087 15456 17132 15484
rect 17126 15444 17132 15456
rect 17184 15444 17190 15496
rect 18782 15444 18788 15496
rect 18840 15484 18846 15496
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 18840 15456 19257 15484
rect 18840 15444 18846 15456
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 19426 15484 19432 15496
rect 19387 15456 19432 15484
rect 19245 15447 19303 15453
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 19610 15484 19616 15496
rect 19571 15456 19616 15484
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 19702 15444 19708 15496
rect 19760 15484 19766 15496
rect 19797 15487 19855 15493
rect 19797 15484 19809 15487
rect 19760 15456 19809 15484
rect 19760 15444 19766 15456
rect 19797 15453 19809 15456
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 22940 15493 22968 15524
rect 23109 15521 23121 15555
rect 23155 15552 23167 15555
rect 23155 15524 23520 15552
rect 23155 15521 23167 15524
rect 23109 15515 23167 15521
rect 23492 15496 23520 15524
rect 24118 15512 24124 15564
rect 24176 15552 24182 15564
rect 24949 15555 25007 15561
rect 24949 15552 24961 15555
rect 24176 15524 24961 15552
rect 24176 15512 24182 15524
rect 24949 15521 24961 15524
rect 24995 15521 25007 15555
rect 26142 15552 26148 15564
rect 24949 15515 25007 15521
rect 25148 15524 26148 15552
rect 22741 15487 22799 15493
rect 22741 15484 22753 15487
rect 22152 15456 22753 15484
rect 22152 15444 22158 15456
rect 22741 15453 22753 15456
rect 22787 15453 22799 15487
rect 22741 15447 22799 15453
rect 22925 15487 22983 15493
rect 22925 15453 22937 15487
rect 22971 15453 22983 15487
rect 22925 15447 22983 15453
rect 23017 15487 23075 15493
rect 23017 15453 23029 15487
rect 23063 15484 23075 15487
rect 23198 15484 23204 15496
rect 23063 15456 23204 15484
rect 23063 15453 23075 15456
rect 23017 15447 23075 15453
rect 23198 15444 23204 15456
rect 23256 15444 23262 15496
rect 23293 15487 23351 15493
rect 23293 15453 23305 15487
rect 23339 15484 23351 15487
rect 23382 15484 23388 15496
rect 23339 15456 23388 15484
rect 23339 15453 23351 15456
rect 23293 15447 23351 15453
rect 23382 15444 23388 15456
rect 23440 15444 23446 15496
rect 23474 15444 23480 15496
rect 23532 15444 23538 15496
rect 24394 15444 24400 15496
rect 24452 15484 24458 15496
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 24452 15456 24593 15484
rect 24452 15444 24458 15456
rect 24581 15453 24593 15456
rect 24627 15453 24639 15487
rect 24581 15447 24639 15453
rect 24765 15487 24823 15493
rect 24765 15453 24777 15487
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 10827 15388 11560 15416
rect 13096 15388 14964 15416
rect 10827 15385 10839 15388
rect 10781 15379 10839 15385
rect 1394 15308 1400 15360
rect 1452 15348 1458 15360
rect 1673 15351 1731 15357
rect 1673 15348 1685 15351
rect 1452 15320 1685 15348
rect 1452 15308 1458 15320
rect 1673 15317 1685 15320
rect 1719 15317 1731 15351
rect 1673 15311 1731 15317
rect 9950 15308 9956 15360
rect 10008 15348 10014 15360
rect 11422 15348 11428 15360
rect 10008 15320 11428 15348
rect 10008 15308 10014 15320
rect 11422 15308 11428 15320
rect 11480 15308 11486 15360
rect 11532 15348 11560 15388
rect 15010 15376 15016 15428
rect 15068 15416 15074 15428
rect 15749 15419 15807 15425
rect 15749 15416 15761 15419
rect 15068 15388 15761 15416
rect 15068 15376 15074 15388
rect 15749 15385 15761 15388
rect 15795 15385 15807 15419
rect 15749 15379 15807 15385
rect 17396 15419 17454 15425
rect 17396 15385 17408 15419
rect 17442 15416 17454 15419
rect 19150 15416 19156 15428
rect 17442 15388 19156 15416
rect 17442 15385 17454 15388
rect 17396 15379 17454 15385
rect 19150 15376 19156 15388
rect 19208 15376 19214 15428
rect 19444 15416 19472 15444
rect 21168 15419 21226 15425
rect 19444 15388 20760 15416
rect 12713 15351 12771 15357
rect 12713 15348 12725 15351
rect 11532 15320 12725 15348
rect 12713 15317 12725 15320
rect 12759 15317 12771 15351
rect 12713 15311 12771 15317
rect 14645 15351 14703 15357
rect 14645 15317 14657 15351
rect 14691 15348 14703 15351
rect 15194 15348 15200 15360
rect 14691 15320 15200 15348
rect 14691 15317 14703 15320
rect 14645 15311 14703 15317
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 15378 15348 15384 15360
rect 15339 15320 15384 15348
rect 15378 15308 15384 15320
rect 15436 15308 15442 15360
rect 15841 15351 15899 15357
rect 15841 15317 15853 15351
rect 15887 15348 15899 15351
rect 16574 15348 16580 15360
rect 15887 15320 16580 15348
rect 15887 15317 15899 15320
rect 15841 15311 15899 15317
rect 16574 15308 16580 15320
rect 16632 15308 16638 15360
rect 19978 15348 19984 15360
rect 19939 15320 19984 15348
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 20732 15348 20760 15388
rect 21168 15385 21180 15419
rect 21214 15416 21226 15419
rect 21818 15416 21824 15428
rect 21214 15388 21824 15416
rect 21214 15385 21226 15388
rect 21168 15379 21226 15385
rect 21818 15376 21824 15388
rect 21876 15376 21882 15428
rect 23934 15416 23940 15428
rect 23032 15388 23940 15416
rect 23032 15360 23060 15388
rect 23934 15376 23940 15388
rect 23992 15416 23998 15428
rect 24780 15416 24808 15447
rect 24854 15444 24860 15496
rect 24912 15484 24918 15496
rect 25148 15493 25176 15524
rect 26142 15512 26148 15524
rect 26200 15512 26206 15564
rect 25133 15487 25191 15493
rect 24912 15456 24957 15484
rect 24912 15444 24918 15456
rect 25133 15453 25145 15487
rect 25179 15453 25191 15487
rect 25133 15447 25191 15453
rect 26053 15487 26111 15493
rect 26053 15453 26065 15487
rect 26099 15484 26111 15487
rect 26697 15487 26755 15493
rect 26099 15456 26648 15484
rect 26099 15453 26111 15456
rect 26053 15447 26111 15453
rect 23992 15388 24808 15416
rect 23992 15376 23998 15388
rect 25314 15376 25320 15428
rect 25372 15416 25378 15428
rect 26145 15419 26203 15425
rect 26145 15416 26157 15419
rect 25372 15388 26157 15416
rect 25372 15376 25378 15388
rect 26145 15385 26157 15388
rect 26191 15385 26203 15419
rect 26145 15379 26203 15385
rect 22002 15348 22008 15360
rect 20732 15320 22008 15348
rect 22002 15308 22008 15320
rect 22060 15348 22066 15360
rect 22281 15351 22339 15357
rect 22281 15348 22293 15351
rect 22060 15320 22293 15348
rect 22060 15308 22066 15320
rect 22281 15317 22293 15320
rect 22327 15317 22339 15351
rect 22281 15311 22339 15317
rect 23014 15308 23020 15360
rect 23072 15308 23078 15360
rect 23477 15351 23535 15357
rect 23477 15317 23489 15351
rect 23523 15348 23535 15351
rect 23566 15348 23572 15360
rect 23523 15320 23572 15348
rect 23523 15317 23535 15320
rect 23477 15311 23535 15317
rect 23566 15308 23572 15320
rect 23624 15308 23630 15360
rect 26620 15348 26648 15456
rect 26697 15453 26709 15487
rect 26743 15484 26755 15487
rect 28442 15484 28448 15496
rect 26743 15456 28448 15484
rect 26743 15453 26755 15456
rect 26697 15447 26755 15453
rect 28442 15444 28448 15456
rect 28500 15444 28506 15496
rect 28537 15487 28595 15493
rect 28537 15453 28549 15487
rect 28583 15453 28595 15487
rect 28537 15447 28595 15453
rect 26964 15419 27022 15425
rect 26964 15385 26976 15419
rect 27010 15416 27022 15419
rect 28166 15416 28172 15428
rect 27010 15388 28172 15416
rect 27010 15385 27022 15388
rect 26964 15379 27022 15385
rect 28166 15376 28172 15388
rect 28224 15376 28230 15428
rect 28552 15416 28580 15447
rect 28902 15444 28908 15496
rect 28960 15484 28966 15496
rect 30101 15487 30159 15493
rect 30101 15484 30113 15487
rect 28960 15456 30113 15484
rect 28960 15444 28966 15456
rect 30101 15453 30113 15456
rect 30147 15453 30159 15487
rect 30101 15447 30159 15453
rect 29086 15416 29092 15428
rect 28552 15388 29092 15416
rect 29086 15376 29092 15388
rect 29144 15376 29150 15428
rect 27246 15348 27252 15360
rect 26620 15320 27252 15348
rect 27246 15308 27252 15320
rect 27304 15308 27310 15360
rect 29178 15308 29184 15360
rect 29236 15348 29242 15360
rect 29917 15351 29975 15357
rect 29917 15348 29929 15351
rect 29236 15320 29929 15348
rect 29236 15308 29242 15320
rect 29917 15317 29929 15320
rect 29963 15317 29975 15351
rect 29917 15311 29975 15317
rect 1104 15258 30820 15280
rect 1104 15206 10880 15258
rect 10932 15206 10944 15258
rect 10996 15206 11008 15258
rect 11060 15206 11072 15258
rect 11124 15206 11136 15258
rect 11188 15206 20811 15258
rect 20863 15206 20875 15258
rect 20927 15206 20939 15258
rect 20991 15206 21003 15258
rect 21055 15206 21067 15258
rect 21119 15206 30820 15258
rect 1104 15184 30820 15206
rect 12253 15147 12311 15153
rect 12253 15144 12265 15147
rect 10980 15116 12265 15144
rect 9668 15079 9726 15085
rect 9668 15045 9680 15079
rect 9714 15076 9726 15079
rect 10980 15076 11008 15116
rect 12253 15113 12265 15116
rect 12299 15113 12311 15147
rect 12253 15107 12311 15113
rect 12897 15147 12955 15153
rect 12897 15113 12909 15147
rect 12943 15144 12955 15147
rect 12986 15144 12992 15156
rect 12943 15116 12992 15144
rect 12943 15113 12955 15116
rect 12897 15107 12955 15113
rect 12986 15104 12992 15116
rect 13044 15104 13050 15156
rect 13357 15147 13415 15153
rect 13357 15113 13369 15147
rect 13403 15144 13415 15147
rect 13722 15144 13728 15156
rect 13403 15116 13728 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 18138 15104 18144 15156
rect 18196 15144 18202 15156
rect 18874 15144 18880 15156
rect 18196 15116 18880 15144
rect 18196 15104 18202 15116
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 19150 15104 19156 15156
rect 19208 15144 19214 15156
rect 19337 15147 19395 15153
rect 19337 15144 19349 15147
rect 19208 15116 19349 15144
rect 19208 15104 19214 15116
rect 19337 15113 19349 15116
rect 19383 15113 19395 15147
rect 19337 15107 19395 15113
rect 19518 15104 19524 15156
rect 19576 15144 19582 15156
rect 22557 15147 22615 15153
rect 22557 15144 22569 15147
rect 19576 15116 20944 15144
rect 19576 15104 19582 15116
rect 20916 15088 20944 15116
rect 21100 15116 22569 15144
rect 13170 15076 13176 15088
rect 9714 15048 11008 15076
rect 11532 15048 13176 15076
rect 9714 15045 9726 15048
rect 9668 15039 9726 15045
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 14968 1458 15020
rect 11532 15017 11560 15048
rect 13170 15036 13176 15048
rect 13228 15036 13234 15088
rect 15378 15076 15384 15088
rect 14844 15048 15384 15076
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 14977 11575 15011
rect 11705 15011 11763 15017
rect 11705 15008 11717 15011
rect 11517 14971 11575 14977
rect 11624 14980 11717 15008
rect 11624 14952 11652 14980
rect 11705 14977 11717 14980
rect 11751 14977 11763 15011
rect 12066 15008 12072 15020
rect 12027 14980 12072 15008
rect 11705 14971 11763 14977
rect 12066 14968 12072 14980
rect 12124 14968 12130 15020
rect 13262 15008 13268 15020
rect 13175 14980 13268 15008
rect 13262 14968 13268 14980
rect 13320 15008 13326 15020
rect 13722 15008 13728 15020
rect 13320 14980 13728 15008
rect 13320 14968 13326 14980
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 14645 15011 14703 15017
rect 14645 14977 14657 15011
rect 14691 15008 14703 15011
rect 14734 15008 14740 15020
rect 14691 14980 14740 15008
rect 14691 14977 14703 14980
rect 14645 14971 14703 14977
rect 14734 14968 14740 14980
rect 14792 14968 14798 15020
rect 14844 15017 14872 15048
rect 15378 15036 15384 15048
rect 15436 15036 15442 15088
rect 15933 15079 15991 15085
rect 15933 15045 15945 15079
rect 15979 15076 15991 15079
rect 20346 15076 20352 15088
rect 15979 15048 20352 15076
rect 15979 15045 15991 15048
rect 15933 15039 15991 15045
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 20898 15036 20904 15088
rect 20956 15036 20962 15088
rect 14829 15011 14887 15017
rect 14829 14977 14841 15011
rect 14875 14977 14887 15011
rect 14829 14971 14887 14977
rect 15197 15011 15255 15017
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 15286 15008 15292 15020
rect 15243 14980 15292 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 17028 15011 17086 15017
rect 17028 14977 17040 15011
rect 17074 15008 17086 15011
rect 18506 15008 18512 15020
rect 17074 14980 18512 15008
rect 17074 14977 17086 14980
rect 17028 14971 17086 14977
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 18601 15011 18659 15017
rect 18601 14977 18613 15011
rect 18647 14977 18659 15011
rect 18601 14971 18659 14977
rect 18785 15011 18843 15017
rect 18785 14977 18797 15011
rect 18831 14977 18843 15011
rect 18785 14971 18843 14977
rect 9306 14900 9312 14952
rect 9364 14940 9370 14952
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 9364 14912 9413 14940
rect 9364 14900 9370 14912
rect 9401 14909 9413 14912
rect 9447 14909 9459 14943
rect 11606 14940 11612 14952
rect 9401 14903 9459 14909
rect 10796 14912 11612 14940
rect 1578 14872 1584 14884
rect 1539 14844 1584 14872
rect 1578 14832 1584 14844
rect 1636 14832 1642 14884
rect 10796 14881 10824 14912
rect 11606 14900 11612 14912
rect 11664 14900 11670 14952
rect 11793 14943 11851 14949
rect 11793 14909 11805 14943
rect 11839 14909 11851 14943
rect 11793 14903 11851 14909
rect 11885 14943 11943 14949
rect 11885 14909 11897 14943
rect 11931 14909 11943 14943
rect 11885 14903 11943 14909
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 10781 14875 10839 14881
rect 10781 14841 10793 14875
rect 10827 14841 10839 14875
rect 10781 14835 10839 14841
rect 11422 14832 11428 14884
rect 11480 14872 11486 14884
rect 11808 14872 11836 14903
rect 11480 14844 11836 14872
rect 11480 14832 11486 14844
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 11900 14804 11928 14903
rect 10192 14776 11928 14804
rect 13464 14804 13492 14903
rect 13538 14900 13544 14952
rect 13596 14940 13602 14952
rect 14921 14943 14979 14949
rect 14921 14940 14933 14943
rect 13596 14912 14933 14940
rect 13596 14900 13602 14912
rect 14921 14909 14933 14912
rect 14967 14909 14979 14943
rect 14921 14903 14979 14909
rect 15013 14943 15071 14949
rect 15013 14909 15025 14943
rect 15059 14909 15071 14943
rect 15013 14903 15071 14909
rect 13906 14832 13912 14884
rect 13964 14872 13970 14884
rect 15028 14872 15056 14903
rect 15102 14900 15108 14952
rect 15160 14940 15166 14952
rect 15381 14943 15439 14949
rect 15381 14940 15393 14943
rect 15160 14912 15393 14940
rect 15160 14900 15166 14912
rect 15381 14909 15393 14912
rect 15427 14909 15439 14943
rect 16758 14940 16764 14952
rect 16719 14912 16764 14940
rect 15381 14903 15439 14909
rect 16758 14900 16764 14912
rect 16816 14900 16822 14952
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18616 14940 18644 14971
rect 18012 14912 18644 14940
rect 18012 14900 18018 14912
rect 13964 14844 15056 14872
rect 13964 14832 13970 14844
rect 14090 14804 14096 14816
rect 13464 14776 14096 14804
rect 10192 14764 10198 14776
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 16025 14807 16083 14813
rect 16025 14804 16037 14807
rect 15804 14776 16037 14804
rect 15804 14764 15810 14776
rect 16025 14773 16037 14776
rect 16071 14804 16083 14807
rect 16666 14804 16672 14816
rect 16071 14776 16672 14804
rect 16071 14773 16083 14776
rect 16025 14767 16083 14773
rect 16666 14764 16672 14776
rect 16724 14804 16730 14816
rect 17126 14804 17132 14816
rect 16724 14776 17132 14804
rect 16724 14764 16730 14776
rect 17126 14764 17132 14776
rect 17184 14764 17190 14816
rect 18141 14807 18199 14813
rect 18141 14773 18153 14807
rect 18187 14804 18199 14807
rect 18598 14804 18604 14816
rect 18187 14776 18604 14804
rect 18187 14773 18199 14776
rect 18141 14767 18199 14773
rect 18598 14764 18604 14776
rect 18656 14764 18662 14816
rect 18800 14804 18828 14971
rect 18874 14968 18880 15020
rect 18932 15008 18938 15020
rect 18932 14980 18977 15008
rect 18932 14968 18938 14980
rect 19058 14968 19064 15020
rect 19116 15008 19122 15020
rect 19153 15011 19211 15017
rect 19153 15008 19165 15011
rect 19116 14980 19165 15008
rect 19116 14968 19122 14980
rect 19153 14977 19165 14980
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 20156 15011 20214 15017
rect 20156 14977 20168 15011
rect 20202 15008 20214 15011
rect 21100 15008 21128 15116
rect 22557 15113 22569 15116
rect 22603 15113 22615 15147
rect 22557 15107 22615 15113
rect 24210 15104 24216 15156
rect 24268 15144 24274 15156
rect 24305 15147 24363 15153
rect 24305 15144 24317 15147
rect 24268 15116 24317 15144
rect 24268 15104 24274 15116
rect 24305 15113 24317 15116
rect 24351 15113 24363 15147
rect 24305 15107 24363 15113
rect 26510 15104 26516 15156
rect 26568 15144 26574 15156
rect 26786 15144 26792 15156
rect 26568 15116 26792 15144
rect 26568 15104 26574 15116
rect 26786 15104 26792 15116
rect 26844 15104 26850 15156
rect 21174 15036 21180 15088
rect 21232 15076 21238 15088
rect 25317 15079 25375 15085
rect 25317 15076 25329 15079
rect 21232 15048 25329 15076
rect 21232 15036 21238 15048
rect 25317 15045 25329 15048
rect 25363 15045 25375 15079
rect 25498 15076 25504 15088
rect 25459 15048 25504 15076
rect 25317 15039 25375 15045
rect 25498 15036 25504 15048
rect 25556 15036 25562 15088
rect 26142 15076 26148 15088
rect 26103 15048 26148 15076
rect 26142 15036 26148 15048
rect 26200 15036 26206 15088
rect 27430 15036 27436 15088
rect 27488 15036 27494 15088
rect 21358 15008 21364 15020
rect 20202 14980 21128 15008
rect 21183 14980 21364 15008
rect 20202 14977 20214 14980
rect 20156 14971 20214 14977
rect 18966 14900 18972 14952
rect 19024 14940 19030 14952
rect 19024 14912 19069 14940
rect 19024 14900 19030 14912
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 19886 14940 19892 14952
rect 19392 14912 19892 14940
rect 19392 14900 19398 14912
rect 19886 14900 19892 14912
rect 19944 14900 19950 14952
rect 21082 14900 21088 14952
rect 21140 14940 21146 14952
rect 21183 14940 21211 14980
rect 21358 14968 21364 14980
rect 21416 15008 21422 15020
rect 21821 15011 21879 15017
rect 21821 15008 21833 15011
rect 21416 14980 21833 15008
rect 21416 14968 21422 14980
rect 21821 14977 21833 14980
rect 21867 14977 21879 15011
rect 21821 14971 21879 14977
rect 22005 15014 22063 15017
rect 22005 15011 22232 15014
rect 22005 14977 22017 15011
rect 22051 15008 22232 15011
rect 22278 15008 22284 15020
rect 22051 14986 22284 15008
rect 22051 14977 22063 14986
rect 22204 14980 22284 14986
rect 22005 14971 22063 14977
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 22370 14968 22376 15020
rect 22428 15008 22434 15020
rect 22428 14980 22473 15008
rect 22428 14968 22434 14980
rect 22830 14968 22836 15020
rect 22888 15008 22894 15020
rect 23017 15011 23075 15017
rect 23017 15008 23029 15011
rect 22888 14980 23029 15008
rect 22888 14968 22894 14980
rect 23017 14977 23029 14980
rect 23063 14977 23075 15011
rect 23198 15008 23204 15020
rect 23159 14980 23204 15008
rect 23017 14971 23075 14977
rect 23198 14968 23204 14980
rect 23256 14968 23262 15020
rect 23385 15011 23443 15017
rect 23385 14977 23397 15011
rect 23431 15008 23443 15011
rect 23474 15008 23480 15020
rect 23431 14980 23480 15008
rect 23431 14977 23443 14980
rect 23385 14971 23443 14977
rect 23474 14968 23480 14980
rect 23532 14968 23538 15020
rect 23569 15011 23627 15017
rect 23569 14977 23581 15011
rect 23615 15008 23627 15011
rect 24210 15008 24216 15020
rect 23615 14980 24216 15008
rect 23615 14977 23627 14980
rect 23569 14971 23627 14977
rect 21140 14912 21211 14940
rect 21140 14900 21146 14912
rect 21266 14900 21272 14952
rect 21324 14940 21330 14952
rect 22097 14943 22155 14949
rect 22097 14940 22109 14943
rect 21324 14912 22109 14940
rect 21324 14900 21330 14912
rect 22097 14909 22109 14912
rect 22143 14909 22155 14943
rect 22097 14903 22155 14909
rect 22186 14900 22192 14952
rect 22244 14940 22250 14952
rect 22244 14912 22289 14940
rect 22244 14900 22250 14912
rect 23106 14900 23112 14952
rect 23164 14940 23170 14952
rect 23293 14943 23351 14949
rect 23293 14940 23305 14943
rect 23164 14912 23305 14940
rect 23164 14900 23170 14912
rect 23293 14909 23305 14912
rect 23339 14909 23351 14943
rect 23293 14903 23351 14909
rect 23584 14872 23612 14971
rect 24210 14968 24216 14980
rect 24268 14968 24274 15020
rect 25590 14968 25596 15020
rect 25648 15008 25654 15020
rect 25961 15011 26019 15017
rect 25961 15008 25973 15011
rect 25648 14980 25973 15008
rect 25648 14968 25654 14980
rect 25961 14977 25973 14980
rect 26007 14977 26019 15011
rect 25961 14971 26019 14977
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 26365 15011 26423 15017
rect 26365 14977 26377 15011
rect 26411 15008 26423 15011
rect 26510 15008 26516 15020
rect 26411 14980 26516 15008
rect 26411 14977 26423 14980
rect 26365 14971 26423 14977
rect 26145 14943 26203 14949
rect 26145 14909 26157 14943
rect 26191 14909 26203 14943
rect 26252 14940 26280 14971
rect 26510 14968 26516 14980
rect 26568 14968 26574 15020
rect 27448 15008 27476 15036
rect 27709 15011 27767 15017
rect 27709 15008 27721 15011
rect 27448 14980 27721 15008
rect 27709 14977 27721 14980
rect 27755 14977 27767 15011
rect 27709 14971 27767 14977
rect 28442 14968 28448 15020
rect 28500 15008 28506 15020
rect 28994 15017 29000 15020
rect 28721 15011 28779 15017
rect 28721 15008 28733 15011
rect 28500 14980 28733 15008
rect 28500 14968 28506 14980
rect 28721 14977 28733 14980
rect 28767 14977 28779 15011
rect 28721 14971 28779 14977
rect 28988 14971 29000 15017
rect 29052 15008 29058 15020
rect 29052 14980 29088 15008
rect 28994 14968 29000 14971
rect 29052 14968 29058 14980
rect 27433 14943 27491 14949
rect 26252 14912 26464 14940
rect 26145 14903 26203 14909
rect 20824 14844 23612 14872
rect 26160 14872 26188 14903
rect 26436 14884 26464 14912
rect 27433 14909 27445 14943
rect 27479 14940 27491 14943
rect 27479 14912 27752 14940
rect 27479 14909 27491 14912
rect 27433 14903 27491 14909
rect 27724 14884 27752 14912
rect 26326 14872 26332 14884
rect 26160 14844 26332 14872
rect 20824 14804 20852 14844
rect 26326 14832 26332 14844
rect 26384 14832 26390 14884
rect 26418 14832 26424 14884
rect 26476 14832 26482 14884
rect 27706 14832 27712 14884
rect 27764 14832 27770 14884
rect 18800 14776 20852 14804
rect 20898 14764 20904 14816
rect 20956 14804 20962 14816
rect 21269 14807 21327 14813
rect 21269 14804 21281 14807
rect 20956 14776 21281 14804
rect 20956 14764 20962 14776
rect 21269 14773 21281 14776
rect 21315 14804 21327 14807
rect 22370 14804 22376 14816
rect 21315 14776 22376 14804
rect 21315 14773 21327 14776
rect 21269 14767 21327 14773
rect 22370 14764 22376 14776
rect 22428 14764 22434 14816
rect 23750 14804 23756 14816
rect 23711 14776 23756 14804
rect 23750 14764 23756 14776
rect 23808 14764 23814 14816
rect 29086 14764 29092 14816
rect 29144 14804 29150 14816
rect 30101 14807 30159 14813
rect 30101 14804 30113 14807
rect 29144 14776 30113 14804
rect 29144 14764 29150 14776
rect 30101 14773 30113 14776
rect 30147 14773 30159 14807
rect 30101 14767 30159 14773
rect 1104 14714 30820 14736
rect 1104 14662 5915 14714
rect 5967 14662 5979 14714
rect 6031 14662 6043 14714
rect 6095 14662 6107 14714
rect 6159 14662 6171 14714
rect 6223 14662 15846 14714
rect 15898 14662 15910 14714
rect 15962 14662 15974 14714
rect 16026 14662 16038 14714
rect 16090 14662 16102 14714
rect 16154 14662 25776 14714
rect 25828 14662 25840 14714
rect 25892 14662 25904 14714
rect 25956 14662 25968 14714
rect 26020 14662 26032 14714
rect 26084 14662 30820 14714
rect 1104 14640 30820 14662
rect 9306 14600 9312 14612
rect 8956 14572 9312 14600
rect 8956 14473 8984 14572
rect 9306 14560 9312 14572
rect 9364 14600 9370 14612
rect 9364 14572 9904 14600
rect 9364 14560 9370 14572
rect 9876 14532 9904 14572
rect 11422 14560 11428 14612
rect 11480 14600 11486 14612
rect 12158 14600 12164 14612
rect 11480 14572 12164 14600
rect 11480 14560 11486 14572
rect 12158 14560 12164 14572
rect 12216 14560 12222 14612
rect 12342 14600 12348 14612
rect 12303 14572 12348 14600
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 13265 14603 13323 14609
rect 13265 14600 13277 14603
rect 12860 14572 13277 14600
rect 12860 14560 12866 14572
rect 13265 14569 13277 14572
rect 13311 14569 13323 14603
rect 15286 14600 15292 14612
rect 15247 14572 15292 14600
rect 13265 14563 13323 14569
rect 15286 14560 15292 14572
rect 15344 14560 15350 14612
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 16669 14603 16727 14609
rect 16669 14600 16681 14603
rect 16632 14572 16681 14600
rect 16632 14560 16638 14572
rect 16669 14569 16681 14572
rect 16715 14569 16727 14603
rect 16669 14563 16727 14569
rect 16758 14560 16764 14612
rect 16816 14600 16822 14612
rect 17310 14600 17316 14612
rect 16816 14572 17316 14600
rect 16816 14560 16822 14572
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 18196 14572 18276 14600
rect 18196 14560 18202 14572
rect 15746 14532 15752 14544
rect 9876 14504 15752 14532
rect 15746 14492 15752 14504
rect 15804 14492 15810 14544
rect 18046 14532 18052 14544
rect 16592 14504 18052 14532
rect 8941 14467 8999 14473
rect 8941 14433 8953 14467
rect 8987 14433 8999 14467
rect 8941 14427 8999 14433
rect 11517 14467 11575 14473
rect 11517 14433 11529 14467
rect 11563 14464 11575 14467
rect 12618 14464 12624 14476
rect 11563 14436 12624 14464
rect 11563 14433 11575 14436
rect 11517 14427 11575 14433
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 14090 14424 14096 14476
rect 14148 14464 14154 14476
rect 14737 14467 14795 14473
rect 14737 14464 14749 14467
rect 14148 14436 14749 14464
rect 14148 14424 14154 14436
rect 14737 14433 14749 14436
rect 14783 14464 14795 14467
rect 15010 14464 15016 14476
rect 14783 14436 15016 14464
rect 14783 14433 14795 14436
rect 14737 14427 14795 14433
rect 15010 14424 15016 14436
rect 15068 14464 15074 14476
rect 15933 14467 15991 14473
rect 15933 14464 15945 14467
rect 15068 14436 15945 14464
rect 15068 14424 15074 14436
rect 15933 14433 15945 14436
rect 15979 14464 15991 14467
rect 16482 14464 16488 14476
rect 15979 14436 16488 14464
rect 15979 14433 15991 14436
rect 15933 14427 15991 14433
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 11422 14396 11428 14408
rect 11383 14368 11428 14396
rect 11422 14356 11428 14368
rect 11480 14356 11486 14408
rect 11606 14356 11612 14408
rect 11664 14396 11670 14408
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 11664 14368 12265 14396
rect 11664 14356 11670 14368
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 12897 14399 12955 14405
rect 12897 14365 12909 14399
rect 12943 14396 12955 14399
rect 13538 14396 13544 14408
rect 12943 14368 13544 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 13722 14356 13728 14408
rect 13780 14396 13786 14408
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 13780 14368 14473 14396
rect 13780 14356 13786 14368
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 15194 14356 15200 14408
rect 15252 14396 15258 14408
rect 15654 14396 15660 14408
rect 15252 14368 15660 14396
rect 15252 14356 15258 14368
rect 15654 14356 15660 14368
rect 15712 14396 15718 14408
rect 16592 14405 16620 14504
rect 18046 14492 18052 14504
rect 18104 14492 18110 14544
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15712 14368 15761 14396
rect 15712 14356 15718 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14365 16635 14399
rect 16577 14359 16635 14365
rect 17221 14399 17279 14405
rect 17221 14365 17233 14399
rect 17267 14396 17279 14399
rect 17954 14396 17960 14408
rect 17267 14368 17816 14396
rect 17915 14368 17960 14396
rect 17267 14365 17279 14368
rect 17221 14359 17279 14365
rect 9208 14331 9266 14337
rect 9208 14297 9220 14331
rect 9254 14328 9266 14331
rect 10226 14328 10232 14340
rect 9254 14300 10232 14328
rect 9254 14297 9266 14300
rect 9208 14291 9266 14297
rect 10226 14288 10232 14300
rect 10284 14288 10290 14340
rect 11790 14328 11796 14340
rect 10336 14300 11796 14328
rect 10336 14269 10364 14300
rect 11790 14288 11796 14300
rect 11848 14328 11854 14340
rect 12069 14331 12127 14337
rect 12069 14328 12081 14331
rect 11848 14300 12081 14328
rect 11848 14288 11854 14300
rect 12069 14297 12081 14300
rect 12115 14297 12127 14331
rect 12069 14291 12127 14297
rect 13081 14331 13139 14337
rect 13081 14297 13093 14331
rect 13127 14328 13139 14331
rect 14553 14331 14611 14337
rect 13127 14300 14136 14328
rect 13127 14297 13139 14300
rect 13081 14291 13139 14297
rect 14108 14269 14136 14300
rect 14553 14297 14565 14331
rect 14599 14328 14611 14331
rect 17313 14331 17371 14337
rect 17313 14328 17325 14331
rect 14599 14300 17325 14328
rect 14599 14297 14611 14300
rect 14553 14291 14611 14297
rect 17313 14297 17325 14300
rect 17359 14297 17371 14331
rect 17313 14291 17371 14297
rect 10321 14263 10379 14269
rect 10321 14229 10333 14263
rect 10367 14229 10379 14263
rect 10321 14223 10379 14229
rect 14093 14263 14151 14269
rect 14093 14229 14105 14263
rect 14139 14229 14151 14263
rect 14093 14223 14151 14229
rect 15102 14220 15108 14272
rect 15160 14260 15166 14272
rect 15657 14263 15715 14269
rect 15657 14260 15669 14263
rect 15160 14232 15669 14260
rect 15160 14220 15166 14232
rect 15657 14229 15669 14232
rect 15703 14229 15715 14263
rect 17788 14260 17816 14368
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 18248 14405 18276 14572
rect 18506 14560 18512 14612
rect 18564 14600 18570 14612
rect 18693 14603 18751 14609
rect 18693 14600 18705 14603
rect 18564 14572 18705 14600
rect 18564 14560 18570 14572
rect 18693 14569 18705 14572
rect 18739 14569 18751 14603
rect 18693 14563 18751 14569
rect 20622 14560 20628 14612
rect 20680 14600 20686 14612
rect 22002 14600 22008 14612
rect 20680 14572 21404 14600
rect 20680 14560 20686 14572
rect 18322 14492 18328 14544
rect 18380 14532 18386 14544
rect 18966 14532 18972 14544
rect 18380 14504 18972 14532
rect 18380 14492 18386 14504
rect 18966 14492 18972 14504
rect 19024 14492 19030 14544
rect 21266 14492 21272 14544
rect 21324 14492 21330 14544
rect 21376 14532 21404 14572
rect 21744 14572 22008 14600
rect 21376 14504 21496 14532
rect 21284 14464 21312 14492
rect 21468 14473 21496 14504
rect 21361 14467 21419 14473
rect 21361 14464 21373 14467
rect 20916 14436 21373 14464
rect 18141 14399 18199 14405
rect 18141 14365 18153 14399
rect 18187 14365 18199 14399
rect 18141 14359 18199 14365
rect 18236 14399 18294 14405
rect 18236 14365 18248 14399
rect 18282 14365 18294 14399
rect 18236 14359 18294 14365
rect 18156 14328 18184 14359
rect 18322 14356 18328 14408
rect 18380 14396 18386 14408
rect 18380 14368 18425 14396
rect 18380 14356 18386 14368
rect 18506 14356 18512 14408
rect 18564 14396 18570 14408
rect 19245 14399 19303 14405
rect 18564 14368 18609 14396
rect 18564 14356 18570 14368
rect 19245 14365 19257 14399
rect 19291 14396 19303 14399
rect 19334 14396 19340 14408
rect 19291 14368 19340 14396
rect 19291 14365 19303 14368
rect 19245 14359 19303 14365
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 19512 14399 19570 14405
rect 19512 14365 19524 14399
rect 19558 14396 19570 14399
rect 19978 14396 19984 14408
rect 19558 14368 19984 14396
rect 19558 14365 19570 14368
rect 19512 14359 19570 14365
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 20070 14356 20076 14408
rect 20128 14396 20134 14408
rect 20916 14396 20944 14436
rect 21361 14433 21373 14436
rect 21407 14433 21419 14467
rect 21361 14427 21419 14433
rect 21453 14467 21511 14473
rect 21453 14433 21465 14467
rect 21499 14433 21511 14467
rect 21453 14427 21511 14433
rect 21082 14396 21088 14408
rect 20128 14368 20944 14396
rect 21043 14368 21088 14396
rect 20128 14356 20134 14368
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 21266 14396 21272 14408
rect 21227 14368 21272 14396
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 21637 14399 21695 14405
rect 21637 14365 21649 14399
rect 21683 14396 21695 14399
rect 21744 14396 21772 14572
rect 22002 14560 22008 14572
rect 22060 14560 22066 14612
rect 26970 14560 26976 14612
rect 27028 14560 27034 14612
rect 27433 14603 27491 14609
rect 27433 14569 27445 14603
rect 27479 14600 27491 14603
rect 27614 14600 27620 14612
rect 27479 14572 27620 14600
rect 27479 14569 27491 14572
rect 27433 14563 27491 14569
rect 27614 14560 27620 14572
rect 27672 14560 27678 14612
rect 26988 14532 27016 14560
rect 29641 14535 29699 14541
rect 29641 14532 29653 14535
rect 26988 14504 29653 14532
rect 29641 14501 29653 14504
rect 29687 14501 29699 14535
rect 29641 14495 29699 14501
rect 26973 14467 27031 14473
rect 26973 14433 26985 14467
rect 27019 14464 27031 14467
rect 27430 14464 27436 14476
rect 27019 14436 27436 14464
rect 27019 14433 27031 14436
rect 26973 14427 27031 14433
rect 27430 14424 27436 14436
rect 27488 14424 27494 14476
rect 27706 14424 27712 14476
rect 27764 14464 27770 14476
rect 27893 14467 27951 14473
rect 27893 14464 27905 14467
rect 27764 14436 27905 14464
rect 27764 14424 27770 14436
rect 27893 14433 27905 14436
rect 27939 14433 27951 14467
rect 27893 14427 27951 14433
rect 21683 14368 21772 14396
rect 22465 14399 22523 14405
rect 21683 14365 21695 14368
rect 21637 14359 21695 14365
rect 22465 14365 22477 14399
rect 22511 14396 22523 14399
rect 23474 14396 23480 14408
rect 22511 14368 23480 14396
rect 22511 14365 22523 14368
rect 22465 14359 22523 14365
rect 23474 14356 23480 14368
rect 23532 14396 23538 14408
rect 24489 14399 24547 14405
rect 24489 14396 24501 14399
rect 23532 14368 24501 14396
rect 23532 14356 23538 14368
rect 24489 14365 24501 14368
rect 24535 14365 24547 14399
rect 24489 14359 24547 14365
rect 26697 14399 26755 14405
rect 26697 14365 26709 14399
rect 26743 14365 26755 14399
rect 26697 14359 26755 14365
rect 22732 14331 22790 14337
rect 18156 14300 22407 14328
rect 19702 14260 19708 14272
rect 17788 14232 19708 14260
rect 15657 14223 15715 14229
rect 19702 14220 19708 14232
rect 19760 14260 19766 14272
rect 20625 14263 20683 14269
rect 20625 14260 20637 14263
rect 19760 14232 20637 14260
rect 19760 14220 19766 14232
rect 20625 14229 20637 14232
rect 20671 14229 20683 14263
rect 21818 14260 21824 14272
rect 21779 14232 21824 14260
rect 20625 14223 20683 14229
rect 21818 14220 21824 14232
rect 21876 14220 21882 14272
rect 22379 14260 22407 14300
rect 22732 14297 22744 14331
rect 22778 14328 22790 14331
rect 23566 14328 23572 14340
rect 22778 14300 23572 14328
rect 22778 14297 22790 14300
rect 22732 14291 22790 14297
rect 23566 14288 23572 14300
rect 23624 14288 23630 14340
rect 24756 14331 24814 14337
rect 24756 14297 24768 14331
rect 24802 14328 24814 14331
rect 25130 14328 25136 14340
rect 24802 14300 25136 14328
rect 24802 14297 24814 14300
rect 24756 14291 24814 14297
rect 25130 14288 25136 14300
rect 25188 14288 25194 14340
rect 26712 14328 26740 14359
rect 26786 14356 26792 14408
rect 26844 14396 26850 14408
rect 26881 14399 26939 14405
rect 26881 14396 26893 14399
rect 26844 14368 26893 14396
rect 26844 14356 26850 14368
rect 26881 14365 26893 14368
rect 26927 14365 26939 14399
rect 26881 14359 26939 14365
rect 27065 14399 27123 14405
rect 27065 14365 27077 14399
rect 27111 14365 27123 14399
rect 27246 14396 27252 14408
rect 27207 14368 27252 14396
rect 27065 14359 27123 14365
rect 26970 14328 26976 14340
rect 26712 14300 26976 14328
rect 26970 14288 26976 14300
rect 27028 14288 27034 14340
rect 27080 14328 27108 14359
rect 27246 14356 27252 14368
rect 27304 14356 27310 14408
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14396 28227 14399
rect 28534 14396 28540 14408
rect 28215 14368 28540 14396
rect 28215 14365 28227 14368
rect 28169 14359 28227 14365
rect 28534 14356 28540 14368
rect 28592 14356 28598 14408
rect 29549 14399 29607 14405
rect 29549 14365 29561 14399
rect 29595 14396 29607 14399
rect 30098 14396 30104 14408
rect 29595 14368 30104 14396
rect 29595 14365 29607 14368
rect 29549 14359 29607 14365
rect 30098 14356 30104 14368
rect 30156 14356 30162 14408
rect 27982 14328 27988 14340
rect 27080 14300 27988 14328
rect 27982 14288 27988 14300
rect 28040 14288 28046 14340
rect 23382 14260 23388 14272
rect 22379 14232 23388 14260
rect 23382 14220 23388 14232
rect 23440 14260 23446 14272
rect 23845 14263 23903 14269
rect 23845 14260 23857 14263
rect 23440 14232 23857 14260
rect 23440 14220 23446 14232
rect 23845 14229 23857 14232
rect 23891 14229 23903 14263
rect 23845 14223 23903 14229
rect 25682 14220 25688 14272
rect 25740 14260 25746 14272
rect 25869 14263 25927 14269
rect 25869 14260 25881 14263
rect 25740 14232 25881 14260
rect 25740 14220 25746 14232
rect 25869 14229 25881 14232
rect 25915 14229 25927 14263
rect 25869 14223 25927 14229
rect 1104 14170 30820 14192
rect 1104 14118 10880 14170
rect 10932 14118 10944 14170
rect 10996 14118 11008 14170
rect 11060 14118 11072 14170
rect 11124 14118 11136 14170
rect 11188 14118 20811 14170
rect 20863 14118 20875 14170
rect 20927 14118 20939 14170
rect 20991 14118 21003 14170
rect 21055 14118 21067 14170
rect 21119 14118 30820 14170
rect 1104 14096 30820 14118
rect 10226 14056 10232 14068
rect 10187 14028 10232 14056
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 14734 14056 14740 14068
rect 14695 14028 14740 14056
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 15654 14056 15660 14068
rect 15615 14028 15660 14056
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 16942 14016 16948 14068
rect 17000 14056 17006 14068
rect 17313 14059 17371 14065
rect 17313 14056 17325 14059
rect 17000 14028 17325 14056
rect 17000 14016 17006 14028
rect 17313 14025 17325 14028
rect 17359 14025 17371 14059
rect 18506 14056 18512 14068
rect 17313 14019 17371 14025
rect 18340 14028 18512 14056
rect 14369 13991 14427 13997
rect 9692 13960 10732 13988
rect 9490 13920 9496 13932
rect 9451 13892 9496 13920
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 9692 13929 9720 13960
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13889 9735 13923
rect 10042 13920 10048 13932
rect 10003 13892 10048 13920
rect 9677 13883 9735 13889
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10704 13929 10732 13960
rect 14369 13957 14381 13991
rect 14415 13988 14427 13991
rect 15470 13988 15476 14000
rect 14415 13960 15476 13988
rect 14415 13957 14427 13960
rect 14369 13951 14427 13957
rect 15470 13948 15476 13960
rect 15528 13948 15534 14000
rect 18340 13988 18368 14028
rect 18506 14016 18512 14028
rect 18564 14016 18570 14068
rect 21910 14056 21916 14068
rect 21871 14028 21916 14056
rect 21910 14016 21916 14028
rect 21968 14016 21974 14068
rect 24210 14016 24216 14068
rect 24268 14056 24274 14068
rect 24305 14059 24363 14065
rect 24305 14056 24317 14059
rect 24268 14028 24317 14056
rect 24268 14016 24274 14028
rect 24305 14025 24317 14028
rect 24351 14025 24363 14059
rect 28166 14056 28172 14068
rect 28127 14028 28172 14056
rect 24305 14019 24363 14025
rect 28166 14016 28172 14028
rect 28224 14016 28230 14068
rect 15580 13960 18368 13988
rect 18417 13991 18475 13997
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13920 10747 13923
rect 11790 13920 11796 13932
rect 10735 13892 11796 13920
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12158 13920 12164 13932
rect 11931 13892 12164 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 14550 13920 14556 13932
rect 14511 13892 14556 13920
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 15580 13929 15608 13960
rect 18417 13957 18429 13991
rect 18463 13988 18475 13991
rect 20346 13988 20352 14000
rect 18463 13960 20352 13988
rect 18463 13957 18475 13960
rect 18417 13951 18475 13957
rect 20346 13948 20352 13960
rect 20404 13948 20410 14000
rect 23474 13988 23480 14000
rect 22940 13960 23480 13988
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 16574 13880 16580 13932
rect 16632 13920 16638 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16632 13892 16681 13920
rect 16632 13880 16638 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 16853 13923 16911 13929
rect 16853 13889 16865 13923
rect 16899 13889 16911 13923
rect 17494 13920 17500 13932
rect 17455 13892 17500 13920
rect 16853 13883 16911 13889
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 9861 13855 9919 13861
rect 9861 13821 9873 13855
rect 9907 13852 9919 13855
rect 10134 13852 10140 13864
rect 9907 13824 10140 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 9784 13784 9812 13815
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 10778 13852 10784 13864
rect 10739 13824 10784 13852
rect 10778 13812 10784 13824
rect 10836 13812 10842 13864
rect 11606 13812 11612 13864
rect 11664 13852 11670 13864
rect 12069 13855 12127 13861
rect 12069 13852 12081 13855
rect 11664 13824 12081 13852
rect 11664 13812 11670 13824
rect 12069 13821 12081 13824
rect 12115 13821 12127 13855
rect 12069 13815 12127 13821
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 16761 13855 16819 13861
rect 16761 13852 16773 13855
rect 15252 13824 16773 13852
rect 15252 13812 15258 13824
rect 16761 13821 16773 13824
rect 16807 13821 16819 13855
rect 16761 13815 16819 13821
rect 9950 13784 9956 13796
rect 9784 13756 9956 13784
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 15654 13744 15660 13796
rect 15712 13784 15718 13796
rect 16868 13784 16896 13883
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 18233 13923 18291 13929
rect 18233 13889 18245 13923
rect 18279 13920 18291 13923
rect 19886 13920 19892 13932
rect 18279 13892 19892 13920
rect 18279 13889 18291 13892
rect 18233 13883 18291 13889
rect 19886 13880 19892 13892
rect 19944 13880 19950 13932
rect 20070 13880 20076 13932
rect 20128 13920 20134 13932
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 20128 13892 21833 13920
rect 20128 13880 20134 13892
rect 21821 13889 21833 13892
rect 21867 13920 21879 13923
rect 22370 13920 22376 13932
rect 21867 13892 22376 13920
rect 21867 13889 21879 13892
rect 21821 13883 21879 13889
rect 22370 13880 22376 13892
rect 22428 13880 22434 13932
rect 22940 13929 22968 13960
rect 23474 13948 23480 13960
rect 23532 13988 23538 14000
rect 23934 13988 23940 14000
rect 23532 13960 23940 13988
rect 23532 13948 23538 13960
rect 23934 13948 23940 13960
rect 23992 13948 23998 14000
rect 24486 13948 24492 14000
rect 24544 13988 24550 14000
rect 25961 13991 26019 13997
rect 25961 13988 25973 13991
rect 24544 13960 25973 13988
rect 24544 13948 24550 13960
rect 25961 13957 25973 13960
rect 26007 13957 26019 13991
rect 29914 13988 29920 14000
rect 25961 13951 26019 13957
rect 26160 13960 29920 13988
rect 22925 13923 22983 13929
rect 22925 13889 22937 13923
rect 22971 13889 22983 13923
rect 22925 13883 22983 13889
rect 23192 13923 23250 13929
rect 23192 13889 23204 13923
rect 23238 13920 23250 13923
rect 23750 13920 23756 13932
rect 23238 13892 23756 13920
rect 23238 13889 23250 13892
rect 23192 13883 23250 13889
rect 23750 13880 23756 13892
rect 23808 13880 23814 13932
rect 24670 13880 24676 13932
rect 24728 13920 24734 13932
rect 24949 13923 25007 13929
rect 24949 13920 24961 13923
rect 24728 13892 24961 13920
rect 24728 13880 24734 13892
rect 24949 13889 24961 13892
rect 24995 13889 25007 13923
rect 25590 13920 25596 13932
rect 25551 13892 25596 13920
rect 24949 13883 25007 13889
rect 17310 13812 17316 13864
rect 17368 13852 17374 13864
rect 19334 13852 19340 13864
rect 17368 13824 19340 13852
rect 17368 13812 17374 13824
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 24964 13852 24992 13883
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 25682 13880 25688 13932
rect 25740 13920 25746 13932
rect 26160 13929 26188 13960
rect 29914 13948 29920 13960
rect 29972 13948 29978 14000
rect 25777 13923 25835 13929
rect 25777 13920 25789 13923
rect 25740 13892 25789 13920
rect 25740 13880 25746 13892
rect 25777 13889 25789 13892
rect 25823 13889 25835 13923
rect 25777 13883 25835 13889
rect 26145 13923 26203 13929
rect 26145 13889 26157 13923
rect 26191 13889 26203 13923
rect 26326 13920 26332 13932
rect 26287 13892 26332 13920
rect 26145 13883 26203 13889
rect 26326 13880 26332 13892
rect 26384 13920 26390 13932
rect 26510 13920 26516 13932
rect 26384 13892 26516 13920
rect 26384 13880 26390 13892
rect 26510 13880 26516 13892
rect 26568 13880 26574 13932
rect 27154 13880 27160 13932
rect 27212 13920 27218 13932
rect 27433 13923 27491 13929
rect 27433 13920 27445 13923
rect 27212 13892 27445 13920
rect 27212 13880 27218 13892
rect 27433 13889 27445 13892
rect 27479 13889 27491 13923
rect 27433 13883 27491 13889
rect 27617 13923 27675 13929
rect 27617 13889 27629 13923
rect 27663 13920 27675 13923
rect 27890 13920 27896 13932
rect 27663 13892 27896 13920
rect 27663 13889 27675 13892
rect 27617 13883 27675 13889
rect 27890 13880 27896 13892
rect 27948 13880 27954 13932
rect 27985 13923 28043 13929
rect 27985 13889 27997 13923
rect 28031 13920 28043 13923
rect 28074 13920 28080 13932
rect 28031 13892 28080 13920
rect 28031 13889 28043 13892
rect 27985 13883 28043 13889
rect 28074 13880 28080 13892
rect 28132 13880 28138 13932
rect 28988 13923 29046 13929
rect 28988 13889 29000 13923
rect 29034 13920 29046 13923
rect 29730 13920 29736 13932
rect 29034 13892 29736 13920
rect 29034 13889 29046 13892
rect 28988 13883 29046 13889
rect 29730 13880 29736 13892
rect 29788 13880 29794 13932
rect 25133 13855 25191 13861
rect 24964 13824 25084 13852
rect 15712 13756 16896 13784
rect 15712 13744 15718 13756
rect 21726 13744 21732 13796
rect 21784 13784 21790 13796
rect 22094 13784 22100 13796
rect 21784 13756 22100 13784
rect 21784 13744 21790 13756
rect 22094 13744 22100 13756
rect 22152 13744 22158 13796
rect 11977 13719 12035 13725
rect 11977 13685 11989 13719
rect 12023 13716 12035 13719
rect 12250 13716 12256 13728
rect 12023 13688 12256 13716
rect 12023 13685 12035 13688
rect 11977 13679 12035 13685
rect 12250 13676 12256 13688
rect 12308 13676 12314 13728
rect 25056 13716 25084 13824
rect 25133 13821 25145 13855
rect 25179 13852 25191 13855
rect 26344 13852 26372 13880
rect 25179 13824 26372 13852
rect 25179 13821 25191 13824
rect 25133 13815 25191 13821
rect 27522 13812 27528 13864
rect 27580 13852 27586 13864
rect 27709 13855 27767 13861
rect 27709 13852 27721 13855
rect 27580 13824 27721 13852
rect 27580 13812 27586 13824
rect 27709 13821 27721 13824
rect 27755 13821 27767 13855
rect 27709 13815 27767 13821
rect 27801 13855 27859 13861
rect 27801 13821 27813 13855
rect 27847 13821 27859 13855
rect 28718 13852 28724 13864
rect 28679 13824 28724 13852
rect 27801 13815 27859 13821
rect 27614 13744 27620 13796
rect 27672 13784 27678 13796
rect 27816 13784 27844 13815
rect 28718 13812 28724 13824
rect 28776 13812 28782 13864
rect 27982 13784 27988 13796
rect 27672 13756 27988 13784
rect 27672 13744 27678 13756
rect 27982 13744 27988 13756
rect 28040 13744 28046 13796
rect 28166 13744 28172 13796
rect 28224 13784 28230 13796
rect 28626 13784 28632 13796
rect 28224 13756 28632 13784
rect 28224 13744 28230 13756
rect 28626 13744 28632 13756
rect 28684 13744 28690 13796
rect 26602 13716 26608 13728
rect 25056 13688 26608 13716
rect 26602 13676 26608 13688
rect 26660 13676 26666 13728
rect 26970 13676 26976 13728
rect 27028 13716 27034 13728
rect 27706 13716 27712 13728
rect 27028 13688 27712 13716
rect 27028 13676 27034 13688
rect 27706 13676 27712 13688
rect 27764 13716 27770 13728
rect 28258 13716 28264 13728
rect 27764 13688 28264 13716
rect 27764 13676 27770 13688
rect 28258 13676 28264 13688
rect 28316 13676 28322 13728
rect 30098 13716 30104 13728
rect 30059 13688 30104 13716
rect 30098 13676 30104 13688
rect 30156 13676 30162 13728
rect 1104 13626 30820 13648
rect 1104 13574 5915 13626
rect 5967 13574 5979 13626
rect 6031 13574 6043 13626
rect 6095 13574 6107 13626
rect 6159 13574 6171 13626
rect 6223 13574 15846 13626
rect 15898 13574 15910 13626
rect 15962 13574 15974 13626
rect 16026 13574 16038 13626
rect 16090 13574 16102 13626
rect 16154 13574 25776 13626
rect 25828 13574 25840 13626
rect 25892 13574 25904 13626
rect 25956 13574 25968 13626
rect 26020 13574 26032 13626
rect 26084 13574 30820 13626
rect 1104 13552 30820 13574
rect 11422 13512 11428 13524
rect 11383 13484 11428 13512
rect 11422 13472 11428 13484
rect 11480 13472 11486 13524
rect 11606 13472 11612 13524
rect 11664 13512 11670 13524
rect 12342 13512 12348 13524
rect 11664 13484 12348 13512
rect 11664 13472 11670 13484
rect 12342 13472 12348 13484
rect 12400 13512 12406 13524
rect 12437 13515 12495 13521
rect 12437 13512 12449 13515
rect 12400 13484 12449 13512
rect 12400 13472 12406 13484
rect 12437 13481 12449 13484
rect 12483 13481 12495 13515
rect 12437 13475 12495 13481
rect 14550 13472 14556 13524
rect 14608 13512 14614 13524
rect 14737 13515 14795 13521
rect 14737 13512 14749 13515
rect 14608 13484 14749 13512
rect 14608 13472 14614 13484
rect 14737 13481 14749 13484
rect 14783 13481 14795 13515
rect 14737 13475 14795 13481
rect 16301 13515 16359 13521
rect 16301 13481 16313 13515
rect 16347 13512 16359 13515
rect 17494 13512 17500 13524
rect 16347 13484 17500 13512
rect 16347 13481 16359 13484
rect 16301 13475 16359 13481
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 19886 13512 19892 13524
rect 19847 13484 19892 13512
rect 19886 13472 19892 13484
rect 19944 13472 19950 13524
rect 22738 13472 22744 13524
rect 22796 13512 22802 13524
rect 22833 13515 22891 13521
rect 22833 13512 22845 13515
rect 22796 13484 22845 13512
rect 22796 13472 22802 13484
rect 22833 13481 22845 13484
rect 22879 13481 22891 13515
rect 22833 13475 22891 13481
rect 23477 13515 23535 13521
rect 23477 13481 23489 13515
rect 23523 13512 23535 13515
rect 23658 13512 23664 13524
rect 23523 13484 23664 13512
rect 23523 13481 23535 13484
rect 23477 13475 23535 13481
rect 23658 13472 23664 13484
rect 23716 13472 23722 13524
rect 24854 13472 24860 13524
rect 24912 13472 24918 13524
rect 25130 13512 25136 13524
rect 25091 13484 25136 13512
rect 25130 13472 25136 13484
rect 25188 13472 25194 13524
rect 25222 13472 25228 13524
rect 25280 13512 25286 13524
rect 25869 13515 25927 13521
rect 25869 13512 25881 13515
rect 25280 13484 25881 13512
rect 25280 13472 25286 13484
rect 25869 13481 25881 13484
rect 25915 13481 25927 13515
rect 28166 13512 28172 13524
rect 25869 13475 25927 13481
rect 27264 13484 28172 13512
rect 11974 13444 11980 13456
rect 10336 13416 11980 13444
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 1762 13308 1768 13320
rect 1443 13280 1768 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 1762 13268 1768 13280
rect 1820 13268 1826 13320
rect 10134 13308 10140 13320
rect 10095 13280 10140 13308
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10336 13308 10364 13416
rect 11974 13404 11980 13416
rect 12032 13404 12038 13456
rect 15010 13404 15016 13456
rect 15068 13444 15074 13456
rect 18230 13444 18236 13456
rect 15068 13416 15332 13444
rect 18191 13416 18236 13444
rect 15068 13404 15074 13416
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13376 10471 13379
rect 10686 13376 10692 13388
rect 10459 13348 10692 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 10686 13336 10692 13348
rect 10744 13376 10750 13388
rect 10965 13379 11023 13385
rect 10965 13376 10977 13379
rect 10744 13348 10977 13376
rect 10744 13336 10750 13348
rect 10965 13345 10977 13348
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 12342 13336 12348 13388
rect 12400 13376 12406 13388
rect 15194 13376 15200 13388
rect 12400 13336 12434 13376
rect 15155 13348 15200 13376
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 15304 13385 15332 13416
rect 18230 13404 18236 13416
rect 18288 13404 18294 13456
rect 20162 13404 20168 13456
rect 20220 13444 20226 13456
rect 21450 13444 21456 13456
rect 20220 13416 21456 13444
rect 20220 13404 20226 13416
rect 21450 13404 21456 13416
rect 21508 13404 21514 13456
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13345 15347 13379
rect 15289 13339 15347 13345
rect 19886 13336 19892 13388
rect 19944 13376 19950 13388
rect 20530 13376 20536 13388
rect 19944 13348 20536 13376
rect 19944 13336 19950 13348
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 21085 13379 21143 13385
rect 21085 13345 21097 13379
rect 21131 13376 21143 13379
rect 21726 13376 21732 13388
rect 21131 13348 21732 13376
rect 21131 13345 21143 13348
rect 21085 13339 21143 13345
rect 21726 13336 21732 13348
rect 21784 13336 21790 13388
rect 23198 13336 23204 13388
rect 23256 13376 23262 13388
rect 23256 13348 24624 13376
rect 23256 13336 23262 13348
rect 10505 13311 10563 13317
rect 10505 13308 10517 13311
rect 10336 13280 10517 13308
rect 10229 13271 10287 13277
rect 10505 13277 10517 13280
rect 10551 13277 10563 13311
rect 10505 13271 10563 13277
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 9950 13172 9956 13184
rect 9911 13144 9956 13172
rect 9950 13132 9956 13144
rect 10008 13132 10014 13184
rect 10244 13172 10272 13271
rect 10778 13268 10784 13320
rect 10836 13308 10842 13320
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 10836 13280 11161 13308
rect 10836 13268 10842 13280
rect 11149 13277 11161 13280
rect 11195 13277 11207 13311
rect 11149 13271 11207 13277
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13277 11299 13311
rect 11241 13271 11299 13277
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 11790 13308 11796 13320
rect 11563 13280 11796 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 11256 13240 11284 13271
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 11974 13268 11980 13320
rect 12032 13308 12038 13320
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 12032 13280 12173 13308
rect 12032 13268 12038 13280
rect 12161 13277 12173 13280
rect 12207 13277 12219 13311
rect 12161 13271 12219 13277
rect 12250 13268 12256 13320
rect 12308 13308 12314 13320
rect 12406 13308 12434 13336
rect 12529 13311 12587 13317
rect 12529 13308 12541 13311
rect 12308 13280 12353 13308
rect 12406 13280 12541 13308
rect 12308 13268 12314 13280
rect 12529 13277 12541 13280
rect 12575 13277 12587 13311
rect 12529 13271 12587 13277
rect 13906 13268 13912 13320
rect 13964 13308 13970 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 13964 13280 14105 13308
rect 13964 13268 13970 13280
rect 14093 13277 14105 13280
rect 14139 13308 14151 13311
rect 14642 13308 14648 13320
rect 14139 13280 14648 13308
rect 14139 13277 14151 13280
rect 14093 13271 14151 13277
rect 14642 13268 14648 13280
rect 14700 13268 14706 13320
rect 15654 13268 15660 13320
rect 15712 13308 15718 13320
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 15712 13280 16129 13308
rect 15712 13268 15718 13280
rect 16117 13277 16129 13280
rect 16163 13277 16175 13311
rect 16117 13271 16175 13277
rect 19242 13268 19248 13320
rect 19300 13308 19306 13320
rect 20346 13308 20352 13320
rect 19300 13280 20352 13308
rect 19300 13268 19306 13280
rect 20346 13268 20352 13280
rect 20404 13268 20410 13320
rect 20438 13268 20444 13320
rect 20496 13308 20502 13320
rect 21358 13308 21364 13320
rect 20496 13280 20541 13308
rect 21319 13280 21364 13308
rect 20496 13268 20502 13280
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 21450 13268 21456 13320
rect 21508 13308 21514 13320
rect 22741 13311 22799 13317
rect 22741 13308 22753 13311
rect 21508 13280 22753 13308
rect 21508 13268 21514 13280
rect 22741 13277 22753 13280
rect 22787 13277 22799 13311
rect 22741 13271 22799 13277
rect 23385 13311 23443 13317
rect 23385 13277 23397 13311
rect 23431 13277 23443 13311
rect 24394 13308 24400 13320
rect 24355 13280 24400 13308
rect 23385 13271 23443 13277
rect 12618 13240 12624 13252
rect 11256 13212 12624 13240
rect 12618 13200 12624 13212
rect 12676 13200 12682 13252
rect 14185 13243 14243 13249
rect 14185 13209 14197 13243
rect 14231 13240 14243 13243
rect 14231 13212 15424 13240
rect 14231 13209 14243 13212
rect 14185 13203 14243 13209
rect 15396 13184 15424 13212
rect 15562 13200 15568 13252
rect 15620 13240 15626 13252
rect 15933 13243 15991 13249
rect 15933 13240 15945 13243
rect 15620 13212 15945 13240
rect 15620 13200 15626 13212
rect 15933 13209 15945 13212
rect 15979 13209 15991 13243
rect 15933 13203 15991 13209
rect 17954 13200 17960 13252
rect 18012 13240 18018 13252
rect 18049 13243 18107 13249
rect 18049 13240 18061 13243
rect 18012 13212 18061 13240
rect 18012 13200 18018 13212
rect 18049 13209 18061 13212
rect 18095 13209 18107 13243
rect 18049 13203 18107 13209
rect 19797 13243 19855 13249
rect 19797 13209 19809 13243
rect 19843 13240 19855 13243
rect 21174 13240 21180 13252
rect 19843 13212 21180 13240
rect 19843 13209 19855 13212
rect 19797 13203 19855 13209
rect 21174 13200 21180 13212
rect 21232 13200 21238 13252
rect 21818 13200 21824 13252
rect 21876 13240 21882 13252
rect 23400 13240 23428 13271
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 24596 13317 24624 13348
rect 24670 13336 24676 13388
rect 24728 13376 24734 13388
rect 24872 13376 24900 13472
rect 24728 13348 24900 13376
rect 24728 13336 24734 13348
rect 24581 13311 24639 13317
rect 24581 13277 24593 13311
rect 24627 13277 24639 13311
rect 24762 13308 24768 13320
rect 24723 13280 24768 13308
rect 24581 13271 24639 13277
rect 24762 13268 24768 13280
rect 24820 13268 24826 13320
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13308 25007 13311
rect 25682 13308 25688 13320
rect 24995 13280 25688 13308
rect 24995 13277 25007 13280
rect 24949 13271 25007 13277
rect 25682 13268 25688 13280
rect 25740 13268 25746 13320
rect 26326 13317 26332 13320
rect 26273 13311 26332 13317
rect 26273 13277 26285 13311
rect 26319 13277 26332 13311
rect 26273 13271 26332 13277
rect 26326 13268 26332 13271
rect 26384 13308 26390 13320
rect 26786 13308 26792 13320
rect 26384 13280 26792 13308
rect 26384 13268 26390 13280
rect 26786 13268 26792 13280
rect 26844 13268 26850 13320
rect 26970 13268 26976 13320
rect 27028 13308 27034 13320
rect 27264 13317 27292 13484
rect 28166 13472 28172 13484
rect 28224 13472 28230 13524
rect 28534 13472 28540 13524
rect 28592 13472 28598 13524
rect 28994 13512 29000 13524
rect 28955 13484 29000 13512
rect 28994 13472 29000 13484
rect 29052 13472 29058 13524
rect 28552 13444 28580 13472
rect 27356 13416 28580 13444
rect 27356 13385 27384 13416
rect 27341 13379 27399 13385
rect 27341 13345 27353 13379
rect 27387 13345 27399 13379
rect 28552 13376 28580 13416
rect 28626 13404 28632 13456
rect 28684 13444 28690 13456
rect 29641 13447 29699 13453
rect 29641 13444 29653 13447
rect 28684 13416 29653 13444
rect 28684 13404 28690 13416
rect 29641 13413 29653 13416
rect 29687 13413 29699 13447
rect 29641 13407 29699 13413
rect 28552 13348 28589 13376
rect 27341 13339 27399 13345
rect 27065 13311 27123 13317
rect 27065 13308 27077 13311
rect 27028 13280 27077 13308
rect 27028 13268 27034 13280
rect 27065 13277 27077 13280
rect 27111 13277 27123 13311
rect 27065 13271 27123 13277
rect 27249 13311 27307 13317
rect 27249 13277 27261 13311
rect 27295 13277 27307 13311
rect 27430 13308 27436 13320
rect 27391 13280 27436 13308
rect 27249 13271 27307 13277
rect 27430 13268 27436 13280
rect 27488 13268 27494 13320
rect 27614 13308 27620 13320
rect 27575 13280 27620 13308
rect 27614 13268 27620 13280
rect 27672 13268 27678 13320
rect 28258 13308 28264 13320
rect 28219 13280 28264 13308
rect 28258 13268 28264 13280
rect 28316 13268 28322 13320
rect 28442 13308 28448 13320
rect 28500 13317 28506 13320
rect 28561 13317 28589 13348
rect 28407 13280 28448 13308
rect 28442 13268 28448 13280
rect 28500 13271 28507 13317
rect 28540 13311 28598 13317
rect 28540 13277 28552 13311
rect 28586 13277 28598 13311
rect 28540 13271 28598 13277
rect 28629 13311 28687 13317
rect 28629 13277 28641 13311
rect 28675 13277 28687 13311
rect 28629 13271 28687 13277
rect 28813 13311 28871 13317
rect 28813 13277 28825 13311
rect 28859 13308 28871 13311
rect 29086 13308 29092 13320
rect 28859 13280 29092 13308
rect 28859 13277 28871 13280
rect 28813 13271 28871 13277
rect 28500 13268 28506 13271
rect 21876 13212 23428 13240
rect 21876 13200 21882 13212
rect 25590 13200 25596 13252
rect 25648 13240 25654 13252
rect 25869 13243 25927 13249
rect 25869 13240 25881 13243
rect 25648 13212 25881 13240
rect 25648 13200 25654 13212
rect 25869 13209 25881 13212
rect 25915 13209 25927 13243
rect 25869 13203 25927 13209
rect 26053 13243 26111 13249
rect 26053 13209 26065 13243
rect 26099 13209 26111 13243
rect 26053 13203 26111 13209
rect 26145 13243 26203 13249
rect 26145 13209 26157 13243
rect 26191 13240 26203 13243
rect 27890 13240 27896 13252
rect 26191 13212 27896 13240
rect 26191 13209 26203 13212
rect 26145 13203 26203 13209
rect 11606 13172 11612 13184
rect 10244 13144 11612 13172
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 11790 13132 11796 13184
rect 11848 13172 11854 13184
rect 11977 13175 12035 13181
rect 11977 13172 11989 13175
rect 11848 13144 11989 13172
rect 11848 13132 11854 13144
rect 11977 13141 11989 13144
rect 12023 13141 12035 13175
rect 15102 13172 15108 13184
rect 15063 13144 15108 13172
rect 11977 13135 12035 13141
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 15378 13132 15384 13184
rect 15436 13172 15442 13184
rect 18690 13172 18696 13184
rect 15436 13144 18696 13172
rect 15436 13132 15442 13144
rect 18690 13132 18696 13144
rect 18748 13132 18754 13184
rect 20533 13175 20591 13181
rect 20533 13141 20545 13175
rect 20579 13172 20591 13175
rect 21266 13172 21272 13184
rect 20579 13144 21272 13172
rect 20579 13141 20591 13144
rect 20533 13135 20591 13141
rect 21266 13132 21272 13144
rect 21324 13132 21330 13184
rect 24854 13132 24860 13184
rect 24912 13172 24918 13184
rect 25314 13172 25320 13184
rect 24912 13144 25320 13172
rect 24912 13132 24918 13144
rect 25314 13132 25320 13144
rect 25372 13172 25378 13184
rect 26068 13172 26096 13203
rect 27890 13200 27896 13212
rect 27948 13200 27954 13252
rect 28644 13240 28672 13271
rect 29086 13268 29092 13280
rect 29144 13268 29150 13320
rect 29546 13308 29552 13320
rect 29507 13280 29552 13308
rect 29546 13268 29552 13280
rect 29604 13268 29610 13320
rect 28552 13212 28672 13240
rect 27798 13172 27804 13184
rect 25372 13144 26096 13172
rect 27759 13144 27804 13172
rect 25372 13132 25378 13144
rect 27798 13132 27804 13144
rect 27856 13132 27862 13184
rect 27982 13132 27988 13184
rect 28040 13172 28046 13184
rect 28552 13172 28580 13212
rect 28810 13172 28816 13184
rect 28040 13144 28816 13172
rect 28040 13132 28046 13144
rect 28810 13132 28816 13144
rect 28868 13132 28874 13184
rect 1104 13082 30820 13104
rect 1104 13030 10880 13082
rect 10932 13030 10944 13082
rect 10996 13030 11008 13082
rect 11060 13030 11072 13082
rect 11124 13030 11136 13082
rect 11188 13030 20811 13082
rect 20863 13030 20875 13082
rect 20927 13030 20939 13082
rect 20991 13030 21003 13082
rect 21055 13030 21067 13082
rect 21119 13030 30820 13082
rect 1104 13008 30820 13030
rect 10042 12968 10048 12980
rect 10003 12940 10048 12968
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 13814 12968 13820 12980
rect 13775 12940 13820 12968
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 14185 12971 14243 12977
rect 14185 12937 14197 12971
rect 14231 12968 14243 12971
rect 15102 12968 15108 12980
rect 14231 12940 15108 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 15562 12968 15568 12980
rect 15523 12940 15568 12968
rect 15562 12928 15568 12940
rect 15620 12928 15626 12980
rect 16574 12968 16580 12980
rect 15856 12940 16580 12968
rect 10594 12900 10600 12912
rect 9416 12872 10600 12900
rect 9416 12841 9444 12872
rect 10594 12860 10600 12872
rect 10652 12900 10658 12912
rect 11422 12900 11428 12912
rect 10652 12872 11428 12900
rect 10652 12860 10658 12872
rect 11422 12860 11428 12872
rect 11480 12860 11486 12912
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 10134 12832 10140 12844
rect 9631 12804 10140 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 10134 12792 10140 12804
rect 10192 12792 10198 12844
rect 10410 12832 10416 12844
rect 10371 12804 10416 12832
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 11698 12832 11704 12844
rect 11659 12804 11704 12832
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12710 12832 12716 12844
rect 12671 12804 12716 12832
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 15856 12841 15884 12940
rect 16574 12928 16580 12940
rect 16632 12968 16638 12980
rect 16761 12971 16819 12977
rect 16761 12968 16773 12971
rect 16632 12940 16773 12968
rect 16632 12928 16638 12940
rect 16761 12937 16773 12940
rect 16807 12937 16819 12971
rect 16761 12931 16819 12937
rect 18322 12928 18328 12980
rect 18380 12968 18386 12980
rect 18380 12940 18552 12968
rect 18380 12928 18386 12940
rect 16206 12860 16212 12912
rect 16264 12900 16270 12912
rect 16264 12872 16712 12900
rect 16264 12860 16270 12872
rect 15749 12835 15807 12841
rect 15749 12801 15761 12835
rect 15795 12801 15807 12835
rect 15749 12795 15807 12801
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12832 16175 12835
rect 16298 12832 16304 12844
rect 16163 12804 16304 12832
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12764 9551 12767
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 9539 12736 10517 12764
rect 9539 12733 9551 12736
rect 9493 12727 9551 12733
rect 10505 12733 10517 12736
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12764 10747 12767
rect 11514 12764 11520 12776
rect 10735 12736 11520 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 11793 12767 11851 12773
rect 11793 12733 11805 12767
rect 11839 12764 11851 12767
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 11839 12736 12817 12764
rect 11839 12733 11851 12736
rect 11793 12727 11851 12733
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 12989 12767 13047 12773
rect 12989 12733 13001 12767
rect 13035 12733 13047 12767
rect 14274 12764 14280 12776
rect 14235 12736 14280 12764
rect 12989 12727 13047 12733
rect 13004 12696 13032 12727
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14461 12767 14519 12773
rect 14461 12733 14473 12767
rect 14507 12764 14519 12767
rect 15010 12764 15016 12776
rect 14507 12736 15016 12764
rect 14507 12733 14519 12736
rect 14461 12727 14519 12733
rect 14476 12696 14504 12727
rect 15010 12724 15016 12736
rect 15068 12724 15074 12776
rect 15764 12764 15792 12795
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 16684 12841 16712 12872
rect 17034 12860 17040 12912
rect 17092 12900 17098 12912
rect 18414 12900 18420 12912
rect 17092 12872 18420 12900
rect 17092 12860 17098 12872
rect 18414 12860 18420 12872
rect 18472 12860 18478 12912
rect 16669 12835 16727 12841
rect 16669 12801 16681 12835
rect 16715 12832 16727 12835
rect 16715 12804 17264 12832
rect 16715 12801 16727 12804
rect 16669 12795 16727 12801
rect 16850 12764 16856 12776
rect 15764 12736 16856 12764
rect 16850 12724 16856 12736
rect 16908 12724 16914 12776
rect 13004 12668 14504 12696
rect 12158 12588 12164 12640
rect 12216 12628 12222 12640
rect 12342 12628 12348 12640
rect 12216 12600 12348 12628
rect 12216 12588 12222 12600
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 16025 12631 16083 12637
rect 16025 12597 16037 12631
rect 16071 12628 16083 12631
rect 16206 12628 16212 12640
rect 16071 12600 16212 12628
rect 16071 12597 16083 12600
rect 16025 12591 16083 12597
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 17236 12628 17264 12804
rect 18046 12792 18052 12844
rect 18104 12832 18110 12844
rect 18141 12835 18199 12841
rect 18141 12832 18153 12835
rect 18104 12804 18153 12832
rect 18104 12792 18110 12804
rect 18141 12801 18153 12804
rect 18187 12801 18199 12835
rect 18141 12795 18199 12801
rect 18230 12792 18236 12844
rect 18288 12832 18294 12844
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 18288 12804 18337 12832
rect 18288 12792 18294 12804
rect 18325 12801 18337 12804
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 18524 12773 18552 12940
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 23569 12971 23627 12977
rect 18748 12940 22094 12968
rect 18748 12928 18754 12940
rect 19536 12872 20576 12900
rect 18690 12832 18696 12844
rect 18651 12804 18696 12832
rect 18690 12792 18696 12804
rect 18748 12792 18754 12844
rect 19536 12841 19564 12872
rect 19521 12835 19579 12841
rect 19521 12801 19533 12835
rect 19567 12801 19579 12835
rect 19521 12795 19579 12801
rect 19702 12792 19708 12844
rect 19760 12792 19766 12844
rect 19797 12835 19855 12841
rect 19797 12801 19809 12835
rect 19843 12832 19855 12835
rect 20070 12832 20076 12844
rect 19843 12804 20076 12832
rect 19843 12801 19855 12804
rect 19797 12795 19855 12801
rect 20070 12792 20076 12804
rect 20128 12792 20134 12844
rect 20548 12841 20576 12872
rect 20622 12860 20628 12912
rect 20680 12900 20686 12912
rect 22066 12900 22094 12940
rect 23569 12937 23581 12971
rect 23615 12968 23627 12971
rect 26234 12968 26240 12980
rect 23615 12940 26240 12968
rect 23615 12937 23627 12940
rect 23569 12931 23627 12937
rect 23477 12903 23535 12909
rect 23477 12900 23489 12903
rect 20680 12872 21864 12900
rect 22066 12872 23489 12900
rect 20680 12860 20686 12872
rect 20533 12835 20591 12841
rect 20533 12801 20545 12835
rect 20579 12832 20591 12835
rect 20809 12835 20867 12841
rect 20579 12804 20760 12832
rect 20579 12801 20591 12804
rect 20533 12795 20591 12801
rect 18417 12767 18475 12773
rect 18417 12733 18429 12767
rect 18463 12733 18475 12767
rect 18417 12727 18475 12733
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12764 18567 12767
rect 19150 12764 19156 12776
rect 18555 12736 19156 12764
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 18432 12696 18460 12727
rect 19150 12724 19156 12736
rect 19208 12724 19214 12776
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12764 19671 12767
rect 19720 12764 19748 12792
rect 20625 12767 20683 12773
rect 20625 12764 20637 12767
rect 19659 12736 20637 12764
rect 19659 12733 19671 12736
rect 19613 12727 19671 12733
rect 20625 12733 20637 12736
rect 20671 12733 20683 12767
rect 20732 12764 20760 12804
rect 20809 12801 20821 12835
rect 20855 12832 20867 12835
rect 21450 12832 21456 12844
rect 20855 12804 21456 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 20898 12764 20904 12776
rect 20732 12736 20904 12764
rect 20625 12727 20683 12733
rect 20898 12724 20904 12736
rect 20956 12724 20962 12776
rect 19337 12699 19395 12705
rect 19337 12696 19349 12699
rect 18432 12668 19349 12696
rect 19337 12665 19349 12668
rect 19383 12665 19395 12699
rect 19337 12659 19395 12665
rect 19705 12699 19763 12705
rect 19705 12665 19717 12699
rect 19751 12696 19763 12699
rect 20717 12699 20775 12705
rect 20717 12696 20729 12699
rect 19751 12668 20729 12696
rect 19751 12665 19763 12668
rect 19705 12659 19763 12665
rect 20640 12640 20668 12668
rect 20717 12665 20729 12668
rect 20763 12665 20775 12699
rect 20717 12659 20775 12665
rect 18690 12628 18696 12640
rect 17236 12600 18696 12628
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 18874 12628 18880 12640
rect 18835 12600 18880 12628
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 19610 12588 19616 12640
rect 19668 12628 19674 12640
rect 20070 12628 20076 12640
rect 19668 12600 20076 12628
rect 19668 12588 19674 12600
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 20346 12628 20352 12640
rect 20307 12600 20352 12628
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 20622 12588 20628 12640
rect 20680 12588 20686 12640
rect 21100 12628 21128 12804
rect 21450 12792 21456 12804
rect 21508 12792 21514 12844
rect 21836 12841 21864 12872
rect 23477 12869 23489 12872
rect 23523 12869 23535 12903
rect 24210 12900 24216 12912
rect 24123 12872 24216 12900
rect 23477 12863 23535 12869
rect 24136 12841 24164 12872
rect 24210 12860 24216 12872
rect 24268 12900 24274 12912
rect 24394 12900 24400 12912
rect 24268 12872 24400 12900
rect 24268 12860 24274 12872
rect 24394 12860 24400 12872
rect 24452 12860 24458 12912
rect 24762 12900 24768 12912
rect 24504 12872 24768 12900
rect 24504 12844 24532 12872
rect 24762 12860 24768 12872
rect 24820 12860 24826 12912
rect 21821 12835 21879 12841
rect 21821 12801 21833 12835
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12801 24179 12835
rect 24121 12795 24179 12801
rect 24305 12835 24363 12841
rect 24305 12801 24317 12835
rect 24351 12801 24363 12835
rect 24305 12795 24363 12801
rect 22097 12767 22155 12773
rect 22097 12733 22109 12767
rect 22143 12764 22155 12767
rect 22186 12764 22192 12776
rect 22143 12736 22192 12764
rect 22143 12733 22155 12736
rect 22097 12727 22155 12733
rect 22186 12724 22192 12736
rect 22244 12724 22250 12776
rect 24320 12764 24348 12795
rect 24486 12792 24492 12844
rect 24544 12832 24550 12844
rect 24673 12835 24731 12841
rect 24544 12804 24637 12832
rect 24544 12792 24550 12804
rect 24673 12801 24685 12835
rect 24719 12832 24731 12835
rect 24854 12832 24860 12844
rect 24719 12804 24860 12832
rect 24719 12801 24731 12804
rect 24673 12795 24731 12801
rect 24854 12792 24860 12804
rect 24912 12792 24918 12844
rect 25332 12832 25360 12940
rect 26234 12928 26240 12940
rect 26292 12928 26298 12980
rect 27614 12928 27620 12980
rect 27672 12968 27678 12980
rect 28537 12971 28595 12977
rect 28537 12968 28549 12971
rect 27672 12940 28549 12968
rect 27672 12928 27678 12940
rect 28537 12937 28549 12940
rect 28583 12968 28595 12971
rect 29546 12968 29552 12980
rect 28583 12940 29552 12968
rect 28583 12937 28595 12940
rect 28537 12931 28595 12937
rect 29546 12928 29552 12940
rect 29604 12928 29610 12980
rect 29730 12968 29736 12980
rect 29691 12940 29736 12968
rect 29730 12928 29736 12940
rect 29788 12928 29794 12980
rect 25406 12860 25412 12912
rect 25464 12900 25470 12912
rect 25961 12903 26019 12909
rect 25961 12900 25973 12903
rect 25464 12872 25973 12900
rect 25464 12860 25470 12872
rect 25961 12869 25973 12872
rect 26007 12869 26019 12903
rect 28718 12900 28724 12912
rect 25961 12863 26019 12869
rect 27172 12872 28724 12900
rect 25590 12832 25596 12844
rect 25332 12804 25596 12832
rect 25590 12792 25596 12804
rect 25648 12792 25654 12844
rect 25777 12835 25835 12841
rect 25777 12801 25789 12835
rect 25823 12801 25835 12835
rect 25777 12795 25835 12801
rect 26145 12835 26203 12841
rect 26145 12801 26157 12835
rect 26191 12801 26203 12835
rect 26145 12795 26203 12801
rect 26421 12835 26479 12841
rect 26421 12801 26433 12835
rect 26467 12832 26479 12835
rect 26786 12832 26792 12844
rect 26467 12804 26792 12832
rect 26467 12801 26479 12804
rect 26421 12795 26479 12801
rect 22296 12736 24348 12764
rect 24397 12767 24455 12773
rect 22296 12708 22324 12736
rect 24397 12733 24409 12767
rect 24443 12764 24455 12767
rect 24443 12736 24716 12764
rect 24443 12733 24455 12736
rect 24397 12727 24455 12733
rect 24688 12708 24716 12736
rect 25406 12724 25412 12776
rect 25464 12764 25470 12776
rect 25792 12764 25820 12795
rect 25464 12736 25820 12764
rect 26160 12764 26188 12795
rect 26786 12792 26792 12804
rect 26844 12792 26850 12844
rect 27172 12841 27200 12872
rect 28718 12860 28724 12872
rect 28776 12860 28782 12912
rect 28810 12860 28816 12912
rect 28868 12900 28874 12912
rect 28868 12872 29408 12900
rect 28868 12860 28874 12872
rect 27157 12835 27215 12841
rect 27157 12801 27169 12835
rect 27203 12801 27215 12835
rect 27157 12795 27215 12801
rect 27424 12835 27482 12841
rect 27424 12801 27436 12835
rect 27470 12832 27482 12835
rect 27798 12832 27804 12844
rect 27470 12804 27804 12832
rect 27470 12801 27482 12804
rect 27424 12795 27482 12801
rect 27798 12792 27804 12804
rect 27856 12792 27862 12844
rect 28258 12792 28264 12844
rect 28316 12832 28322 12844
rect 28997 12835 29055 12841
rect 28997 12832 29009 12835
rect 28316 12804 29009 12832
rect 28316 12792 28322 12804
rect 28997 12801 29009 12804
rect 29043 12801 29055 12835
rect 29178 12832 29184 12844
rect 29139 12804 29184 12832
rect 28997 12795 29055 12801
rect 29178 12792 29184 12804
rect 29236 12792 29242 12844
rect 29380 12841 29408 12872
rect 29365 12835 29423 12841
rect 29365 12801 29377 12835
rect 29411 12801 29423 12835
rect 29365 12795 29423 12801
rect 29549 12835 29607 12841
rect 29549 12801 29561 12835
rect 29595 12832 29607 12835
rect 30098 12832 30104 12844
rect 29595 12804 30104 12832
rect 29595 12801 29607 12804
rect 29549 12795 29607 12801
rect 30098 12792 30104 12804
rect 30156 12792 30162 12844
rect 26160 12736 26280 12764
rect 25464 12724 25470 12736
rect 21450 12656 21456 12708
rect 21508 12696 21514 12708
rect 22278 12696 22284 12708
rect 21508 12668 22284 12696
rect 21508 12656 21514 12668
rect 22278 12656 22284 12668
rect 22336 12656 22342 12708
rect 24670 12656 24676 12708
rect 24728 12656 24734 12708
rect 21910 12628 21916 12640
rect 21100 12600 21916 12628
rect 21910 12588 21916 12600
rect 21968 12588 21974 12640
rect 24854 12628 24860 12640
rect 24815 12600 24860 12628
rect 24854 12588 24860 12600
rect 24912 12588 24918 12640
rect 26252 12628 26280 12736
rect 28534 12724 28540 12776
rect 28592 12764 28598 12776
rect 29273 12767 29331 12773
rect 29273 12764 29285 12767
rect 28592 12736 29285 12764
rect 28592 12724 28598 12736
rect 29273 12733 29285 12736
rect 29319 12733 29331 12767
rect 29273 12727 29331 12733
rect 30006 12628 30012 12640
rect 26252 12600 30012 12628
rect 30006 12588 30012 12600
rect 30064 12588 30070 12640
rect 1104 12538 30820 12560
rect 1104 12486 5915 12538
rect 5967 12486 5979 12538
rect 6031 12486 6043 12538
rect 6095 12486 6107 12538
rect 6159 12486 6171 12538
rect 6223 12486 15846 12538
rect 15898 12486 15910 12538
rect 15962 12486 15974 12538
rect 16026 12486 16038 12538
rect 16090 12486 16102 12538
rect 16154 12486 25776 12538
rect 25828 12486 25840 12538
rect 25892 12486 25904 12538
rect 25956 12486 25968 12538
rect 26020 12486 26032 12538
rect 26084 12486 30820 12538
rect 1104 12464 30820 12486
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10321 12427 10379 12433
rect 10321 12424 10333 12427
rect 10192 12396 10333 12424
rect 10192 12384 10198 12396
rect 10321 12393 10333 12396
rect 10367 12393 10379 12427
rect 10321 12387 10379 12393
rect 11517 12427 11575 12433
rect 11517 12393 11529 12427
rect 11563 12424 11575 12427
rect 12066 12424 12072 12436
rect 11563 12396 12072 12424
rect 11563 12393 11575 12396
rect 11517 12387 11575 12393
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 15654 12424 15660 12436
rect 12400 12396 15660 12424
rect 12400 12384 12406 12396
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 17954 12424 17960 12436
rect 16592 12396 17960 12424
rect 10594 12316 10600 12368
rect 10652 12356 10658 12368
rect 10652 12328 10916 12356
rect 10652 12316 10658 12328
rect 10778 12288 10784 12300
rect 10739 12260 10784 12288
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 10888 12297 10916 12328
rect 11882 12316 11888 12368
rect 11940 12356 11946 12368
rect 14093 12359 14151 12365
rect 14093 12356 14105 12359
rect 11940 12328 14105 12356
rect 11940 12316 11946 12328
rect 14093 12325 14105 12328
rect 14139 12325 14151 12359
rect 14093 12319 14151 12325
rect 16592 12300 16620 12396
rect 17954 12384 17960 12396
rect 18012 12384 18018 12436
rect 18690 12424 18696 12436
rect 18651 12396 18696 12424
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 19610 12384 19616 12436
rect 19668 12424 19674 12436
rect 21818 12424 21824 12436
rect 19668 12396 20668 12424
rect 19668 12384 19674 12396
rect 20640 12368 20668 12396
rect 21192 12396 21824 12424
rect 20622 12316 20628 12368
rect 20680 12356 20686 12368
rect 21192 12365 21220 12396
rect 21818 12384 21824 12396
rect 21876 12384 21882 12436
rect 21177 12359 21235 12365
rect 21177 12356 21189 12359
rect 20680 12328 21189 12356
rect 20680 12316 20686 12328
rect 21177 12325 21189 12328
rect 21223 12325 21235 12359
rect 21542 12356 21548 12368
rect 21177 12319 21235 12325
rect 21376 12328 21548 12356
rect 21376 12300 21404 12328
rect 21542 12316 21548 12328
rect 21600 12316 21606 12368
rect 24394 12316 24400 12368
rect 24452 12356 24458 12368
rect 26510 12356 26516 12368
rect 24452 12328 24532 12356
rect 26471 12328 26516 12356
rect 24452 12316 24458 12328
rect 10873 12291 10931 12297
rect 10873 12257 10885 12291
rect 10919 12257 10931 12291
rect 10873 12251 10931 12257
rect 11514 12248 11520 12300
rect 11572 12288 11578 12300
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 11572 12260 12081 12288
rect 11572 12248 11578 12260
rect 12069 12257 12081 12260
rect 12115 12257 12127 12291
rect 12069 12251 12127 12257
rect 12250 12248 12256 12300
rect 12308 12288 12314 12300
rect 14737 12291 14795 12297
rect 12308 12260 12940 12288
rect 12308 12248 12314 12260
rect 10686 12220 10692 12232
rect 10647 12192 10692 12220
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 11330 12180 11336 12232
rect 11388 12220 11394 12232
rect 12342 12220 12348 12232
rect 11388 12192 12348 12220
rect 11388 12180 11394 12192
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 12912 12229 12940 12260
rect 14737 12257 14749 12291
rect 14783 12288 14795 12291
rect 15010 12288 15016 12300
rect 14783 12260 15016 12288
rect 14783 12257 14795 12260
rect 14737 12251 14795 12257
rect 15010 12248 15016 12260
rect 15068 12248 15074 12300
rect 16574 12288 16580 12300
rect 16487 12260 16580 12288
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 17310 12288 17316 12300
rect 17271 12260 17316 12288
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 20898 12248 20904 12300
rect 20956 12288 20962 12300
rect 21358 12288 21364 12300
rect 20956 12260 21128 12288
rect 21271 12260 21364 12288
rect 20956 12248 20962 12260
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12189 12955 12223
rect 15378 12220 15384 12232
rect 15339 12192 15384 12220
rect 12897 12183 12955 12189
rect 12820 12152 12848 12183
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12189 16267 12223
rect 16209 12183 16267 12189
rect 16357 12223 16415 12229
rect 16357 12189 16369 12223
rect 16403 12220 16415 12223
rect 16592 12220 16620 12248
rect 16403 12192 16620 12220
rect 16715 12223 16773 12229
rect 16403 12189 16415 12192
rect 16357 12183 16415 12189
rect 16715 12189 16727 12223
rect 16761 12220 16773 12223
rect 17580 12223 17638 12229
rect 16761 12192 17540 12220
rect 16761 12189 16773 12192
rect 16715 12183 16773 12189
rect 13906 12152 13912 12164
rect 12820 12124 13912 12152
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 14918 12152 14924 12164
rect 14056 12124 14924 12152
rect 14056 12112 14062 12124
rect 14918 12112 14924 12124
rect 14976 12152 14982 12164
rect 16224 12152 16252 12183
rect 16482 12152 16488 12164
rect 14976 12124 16252 12152
rect 16443 12124 16488 12152
rect 14976 12112 14982 12124
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 16577 12155 16635 12161
rect 16577 12121 16589 12155
rect 16623 12152 16635 12155
rect 17034 12152 17040 12164
rect 16623 12124 17040 12152
rect 16623 12121 16635 12124
rect 16577 12115 16635 12121
rect 17034 12112 17040 12124
rect 17092 12112 17098 12164
rect 11882 12084 11888 12096
rect 11843 12056 11888 12084
rect 11882 12044 11888 12056
rect 11940 12044 11946 12096
rect 11977 12087 12035 12093
rect 11977 12053 11989 12087
rect 12023 12084 12035 12087
rect 12066 12084 12072 12096
rect 12023 12056 12072 12084
rect 12023 12053 12035 12056
rect 11977 12047 12035 12053
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 13078 12084 13084 12096
rect 13039 12056 13084 12084
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 13722 12044 13728 12096
rect 13780 12084 13786 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 13780 12056 14473 12084
rect 13780 12044 13786 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 14461 12047 14519 12053
rect 14553 12087 14611 12093
rect 14553 12053 14565 12087
rect 14599 12084 14611 12087
rect 15102 12084 15108 12096
rect 14599 12056 15108 12084
rect 14599 12053 14611 12056
rect 14553 12047 14611 12053
rect 15102 12044 15108 12056
rect 15160 12044 15166 12096
rect 15654 12084 15660 12096
rect 15615 12056 15660 12084
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 16853 12087 16911 12093
rect 16853 12053 16865 12087
rect 16899 12084 16911 12087
rect 16942 12084 16948 12096
rect 16899 12056 16948 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 17512 12084 17540 12192
rect 17580 12189 17592 12223
rect 17626 12220 17638 12223
rect 18874 12220 18880 12232
rect 17626 12192 18880 12220
rect 17626 12189 17638 12192
rect 17580 12183 17638 12189
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 19334 12220 19340 12232
rect 19291 12192 19340 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 19334 12180 19340 12192
rect 19392 12220 19398 12232
rect 21100 12229 21128 12260
rect 21358 12248 21364 12260
rect 21416 12248 21422 12300
rect 21560 12260 22131 12288
rect 21085 12223 21143 12229
rect 19392 12192 21036 12220
rect 19392 12180 19398 12192
rect 19518 12161 19524 12164
rect 19512 12115 19524 12161
rect 19576 12152 19582 12164
rect 21008 12152 21036 12192
rect 21085 12189 21097 12223
rect 21131 12220 21143 12223
rect 21560 12220 21588 12260
rect 21994 12223 22052 12229
rect 21994 12220 22006 12223
rect 21131 12192 21588 12220
rect 21928 12192 22006 12220
rect 21131 12189 21143 12192
rect 21085 12183 21143 12189
rect 21928 12152 21956 12192
rect 21994 12189 22006 12192
rect 22040 12189 22052 12223
rect 22103 12220 22131 12260
rect 22738 12220 22744 12232
rect 22103 12192 22744 12220
rect 21994 12183 22052 12189
rect 22738 12180 22744 12192
rect 22796 12180 22802 12232
rect 24210 12180 24216 12232
rect 24268 12220 24274 12232
rect 24397 12223 24455 12229
rect 24397 12220 24409 12223
rect 24268 12192 24409 12220
rect 24268 12180 24274 12192
rect 24397 12189 24409 12192
rect 24443 12189 24455 12223
rect 24504 12220 24532 12328
rect 26510 12316 26516 12328
rect 26568 12316 26574 12368
rect 27798 12356 27804 12368
rect 26620 12328 27804 12356
rect 24670 12288 24676 12300
rect 24631 12260 24676 12288
rect 24670 12248 24676 12260
rect 24728 12248 24734 12300
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 24504 12192 24593 12220
rect 24397 12183 24455 12189
rect 24581 12189 24593 12192
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 24949 12223 25007 12229
rect 24949 12189 24961 12223
rect 24995 12189 25007 12223
rect 26234 12220 26240 12232
rect 26195 12192 26240 12220
rect 24949 12183 25007 12189
rect 22094 12152 22100 12164
rect 19576 12124 19612 12152
rect 19720 12124 20760 12152
rect 21008 12124 22100 12152
rect 19518 12112 19524 12115
rect 19576 12112 19582 12124
rect 19720 12084 19748 12124
rect 17512 12056 19748 12084
rect 19794 12044 19800 12096
rect 19852 12084 19858 12096
rect 20625 12087 20683 12093
rect 20625 12084 20637 12087
rect 19852 12056 20637 12084
rect 19852 12044 19858 12056
rect 20625 12053 20637 12056
rect 20671 12053 20683 12087
rect 20732 12084 20760 12124
rect 22094 12112 22100 12124
rect 22152 12112 22158 12164
rect 22278 12161 22284 12164
rect 22272 12115 22284 12161
rect 22336 12152 22342 12164
rect 22336 12124 22372 12152
rect 22278 12112 22284 12115
rect 22336 12112 22342 12124
rect 23750 12112 23756 12164
rect 23808 12152 23814 12164
rect 24486 12152 24492 12164
rect 23808 12124 24492 12152
rect 23808 12112 23814 12124
rect 24486 12112 24492 12124
rect 24544 12152 24550 12164
rect 24780 12152 24808 12183
rect 24544 12124 24808 12152
rect 24964 12152 24992 12183
rect 26234 12180 26240 12192
rect 26292 12180 26298 12232
rect 26620 12229 26648 12328
rect 27798 12316 27804 12328
rect 27856 12316 27862 12368
rect 26329 12223 26387 12229
rect 26329 12189 26341 12223
rect 26375 12189 26387 12223
rect 26329 12183 26387 12189
rect 26605 12223 26663 12229
rect 26605 12189 26617 12223
rect 26651 12189 26663 12223
rect 26786 12220 26792 12232
rect 26747 12192 26792 12220
rect 26605 12183 26663 12189
rect 25682 12152 25688 12164
rect 24964 12124 25688 12152
rect 24544 12112 24550 12124
rect 25682 12112 25688 12124
rect 25740 12152 25746 12164
rect 26344 12152 26372 12183
rect 26786 12180 26792 12192
rect 26844 12180 26850 12232
rect 27525 12223 27583 12229
rect 27525 12189 27537 12223
rect 27571 12189 27583 12223
rect 27525 12183 27583 12189
rect 25740 12124 26372 12152
rect 25740 12112 25746 12124
rect 21361 12087 21419 12093
rect 21361 12084 21373 12087
rect 20732 12056 21373 12084
rect 20625 12047 20683 12053
rect 21361 12053 21373 12056
rect 21407 12053 21419 12087
rect 21361 12047 21419 12053
rect 21450 12044 21456 12096
rect 21508 12084 21514 12096
rect 22370 12084 22376 12096
rect 21508 12056 22376 12084
rect 21508 12044 21514 12056
rect 22370 12044 22376 12056
rect 22428 12084 22434 12096
rect 23385 12087 23443 12093
rect 23385 12084 23397 12087
rect 22428 12056 23397 12084
rect 22428 12044 22434 12056
rect 23385 12053 23397 12056
rect 23431 12053 23443 12087
rect 25130 12084 25136 12096
rect 25091 12056 25136 12084
rect 23385 12047 23443 12053
rect 25130 12044 25136 12056
rect 25188 12044 25194 12096
rect 26142 12044 26148 12096
rect 26200 12084 26206 12096
rect 27540 12084 27568 12183
rect 27706 12180 27712 12232
rect 27764 12220 27770 12232
rect 27801 12223 27859 12229
rect 27801 12220 27813 12223
rect 27764 12192 27813 12220
rect 27764 12180 27770 12192
rect 27801 12189 27813 12192
rect 27847 12220 27859 12223
rect 28258 12220 28264 12232
rect 27847 12192 28264 12220
rect 27847 12189 27859 12192
rect 27801 12183 27859 12189
rect 28258 12180 28264 12192
rect 28316 12180 28322 12232
rect 28997 12223 29055 12229
rect 28997 12189 29009 12223
rect 29043 12220 29055 12223
rect 29178 12220 29184 12232
rect 29043 12192 29184 12220
rect 29043 12189 29055 12192
rect 28997 12183 29055 12189
rect 29178 12180 29184 12192
rect 29236 12180 29242 12232
rect 30101 12223 30159 12229
rect 30101 12189 30113 12223
rect 30147 12220 30159 12223
rect 30190 12220 30196 12232
rect 30147 12192 30196 12220
rect 30147 12189 30159 12192
rect 30101 12183 30159 12189
rect 30190 12180 30196 12192
rect 30248 12180 30254 12232
rect 26200 12056 27568 12084
rect 26200 12044 26206 12056
rect 27706 12044 27712 12096
rect 27764 12084 27770 12096
rect 28813 12087 28871 12093
rect 28813 12084 28825 12087
rect 27764 12056 28825 12084
rect 27764 12044 27770 12056
rect 28813 12053 28825 12056
rect 28859 12053 28871 12087
rect 28813 12047 28871 12053
rect 28902 12044 28908 12096
rect 28960 12084 28966 12096
rect 29917 12087 29975 12093
rect 29917 12084 29929 12087
rect 28960 12056 29929 12084
rect 28960 12044 28966 12056
rect 29917 12053 29929 12056
rect 29963 12053 29975 12087
rect 29917 12047 29975 12053
rect 1104 11994 30820 12016
rect 1104 11942 10880 11994
rect 10932 11942 10944 11994
rect 10996 11942 11008 11994
rect 11060 11942 11072 11994
rect 11124 11942 11136 11994
rect 11188 11942 20811 11994
rect 20863 11942 20875 11994
rect 20927 11942 20939 11994
rect 20991 11942 21003 11994
rect 21055 11942 21067 11994
rect 21119 11942 30820 11994
rect 1104 11920 30820 11942
rect 12066 11880 12072 11892
rect 12027 11852 12072 11880
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 12897 11883 12955 11889
rect 12897 11880 12909 11883
rect 12768 11852 12909 11880
rect 12768 11840 12774 11852
rect 12897 11849 12909 11852
rect 12943 11849 12955 11883
rect 12897 11843 12955 11849
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13541 11883 13599 11889
rect 13541 11880 13553 11883
rect 13412 11852 13553 11880
rect 13412 11840 13418 11852
rect 13541 11849 13553 11852
rect 13587 11849 13599 11883
rect 13541 11843 13599 11849
rect 13722 11840 13728 11892
rect 13780 11880 13786 11892
rect 13909 11883 13967 11889
rect 13909 11880 13921 11883
rect 13780 11852 13921 11880
rect 13780 11840 13786 11852
rect 13909 11849 13921 11852
rect 13955 11849 13967 11883
rect 13909 11843 13967 11849
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 14734 11880 14740 11892
rect 14240 11852 14740 11880
rect 14240 11840 14246 11852
rect 14734 11840 14740 11852
rect 14792 11880 14798 11892
rect 15102 11880 15108 11892
rect 14792 11852 14964 11880
rect 15063 11852 15108 11880
rect 14792 11840 14798 11852
rect 9858 11812 9864 11824
rect 9819 11784 9864 11812
rect 9858 11772 9864 11784
rect 9916 11772 9922 11824
rect 10045 11815 10103 11821
rect 10045 11781 10057 11815
rect 10091 11812 10103 11815
rect 14458 11812 14464 11824
rect 10091 11784 14464 11812
rect 10091 11781 10103 11784
rect 10045 11775 10103 11781
rect 14458 11772 14464 11784
rect 14516 11812 14522 11824
rect 14642 11812 14648 11824
rect 14516 11784 14648 11812
rect 14516 11772 14522 11784
rect 14642 11772 14648 11784
rect 14700 11772 14706 11824
rect 11422 11704 11428 11756
rect 11480 11744 11486 11756
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 11480 11716 11989 11744
rect 11480 11704 11486 11716
rect 11977 11713 11989 11716
rect 12023 11713 12035 11747
rect 12158 11744 12164 11756
rect 12119 11716 12164 11744
rect 11977 11707 12035 11713
rect 12158 11704 12164 11716
rect 12216 11704 12222 11756
rect 13078 11744 13084 11756
rect 13039 11716 13084 11744
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11744 14795 11747
rect 14829 11747 14887 11753
rect 14829 11744 14841 11747
rect 14783 11716 14841 11744
rect 14783 11713 14795 11716
rect 14737 11707 14795 11713
rect 14829 11713 14841 11716
rect 14875 11713 14887 11747
rect 14936 11744 14964 11852
rect 15102 11840 15108 11852
rect 15160 11840 15166 11892
rect 16482 11840 16488 11892
rect 16540 11880 16546 11892
rect 18049 11883 18107 11889
rect 18049 11880 18061 11883
rect 16540 11852 18061 11880
rect 16540 11840 16546 11852
rect 18049 11849 18061 11852
rect 18095 11849 18107 11883
rect 19518 11880 19524 11892
rect 19479 11852 19524 11880
rect 18049 11843 18107 11849
rect 19518 11840 19524 11852
rect 19576 11840 19582 11892
rect 21269 11883 21327 11889
rect 20732 11852 21211 11880
rect 16500 11812 16528 11840
rect 15764 11784 16528 11812
rect 16776 11784 17724 11812
rect 15764 11753 15792 11784
rect 15749 11747 15807 11753
rect 14936 11716 15148 11744
rect 14829 11707 14887 11713
rect 13998 11676 14004 11688
rect 13959 11648 14004 11676
rect 13998 11636 14004 11648
rect 14056 11636 14062 11688
rect 14182 11636 14188 11688
rect 14240 11676 14246 11688
rect 15010 11676 15016 11688
rect 14240 11648 15016 11676
rect 14240 11636 14246 11648
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 15120 11685 15148 11716
rect 15749 11713 15761 11747
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11744 15991 11747
rect 16206 11744 16212 11756
rect 15979 11716 16212 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 16666 11744 16672 11756
rect 16627 11716 16672 11744
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 15105 11679 15163 11685
rect 15105 11645 15117 11679
rect 15151 11645 15163 11679
rect 15105 11639 15163 11645
rect 16025 11679 16083 11685
rect 16025 11645 16037 11679
rect 16071 11676 16083 11679
rect 16298 11676 16304 11688
rect 16071 11648 16304 11676
rect 16071 11645 16083 11648
rect 16025 11639 16083 11645
rect 16298 11636 16304 11648
rect 16356 11676 16362 11688
rect 16776 11676 16804 11784
rect 16942 11753 16948 11756
rect 16936 11744 16948 11753
rect 16903 11716 16948 11744
rect 16936 11707 16948 11716
rect 16942 11704 16948 11707
rect 17000 11704 17006 11756
rect 16356 11648 16804 11676
rect 16356 11636 16362 11648
rect 14921 11611 14979 11617
rect 14921 11577 14933 11611
rect 14967 11608 14979 11611
rect 15565 11611 15623 11617
rect 15565 11608 15577 11611
rect 14967 11580 15577 11608
rect 14967 11577 14979 11580
rect 14921 11571 14979 11577
rect 15565 11577 15577 11580
rect 15611 11577 15623 11611
rect 17696 11608 17724 11784
rect 18230 11772 18236 11824
rect 18288 11812 18294 11824
rect 20346 11812 20352 11824
rect 18288 11784 19012 11812
rect 18288 11772 18294 11784
rect 18046 11704 18052 11756
rect 18104 11744 18110 11756
rect 18782 11744 18788 11756
rect 18104 11716 18788 11744
rect 18104 11704 18110 11716
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 18984 11753 19012 11784
rect 19076 11784 20352 11812
rect 19076 11753 19104 11784
rect 20346 11772 20352 11784
rect 20404 11772 20410 11824
rect 18969 11747 19027 11753
rect 18969 11713 18981 11747
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 19061 11747 19119 11753
rect 19061 11713 19073 11747
rect 19107 11713 19119 11747
rect 19061 11707 19119 11713
rect 19337 11747 19395 11753
rect 19337 11713 19349 11747
rect 19383 11744 19395 11747
rect 19794 11744 19800 11756
rect 19383 11716 19800 11744
rect 19383 11713 19395 11716
rect 19337 11707 19395 11713
rect 19150 11676 19156 11688
rect 19111 11648 19156 11676
rect 19150 11636 19156 11648
rect 19208 11636 19214 11688
rect 19352 11608 19380 11707
rect 19794 11704 19800 11716
rect 19852 11704 19858 11756
rect 20732 11753 20760 11852
rect 21183 11812 21211 11852
rect 21269 11849 21281 11883
rect 21315 11880 21327 11883
rect 22278 11880 22284 11892
rect 21315 11852 22284 11880
rect 21315 11849 21327 11852
rect 21269 11843 21327 11849
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 23477 11883 23535 11889
rect 23477 11849 23489 11883
rect 23523 11849 23535 11883
rect 25314 11880 25320 11892
rect 25275 11852 25320 11880
rect 23477 11843 23535 11849
rect 21818 11812 21824 11824
rect 21183 11784 21824 11812
rect 21818 11772 21824 11784
rect 21876 11772 21882 11824
rect 21910 11772 21916 11824
rect 21968 11812 21974 11824
rect 23492 11812 23520 11843
rect 25314 11840 25320 11852
rect 25372 11840 25378 11892
rect 21968 11784 23520 11812
rect 24204 11815 24262 11821
rect 21968 11772 21974 11784
rect 24204 11781 24216 11815
rect 24250 11812 24262 11815
rect 24854 11812 24860 11824
rect 24250 11784 24860 11812
rect 24250 11781 24262 11784
rect 24204 11775 24262 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 25498 11772 25504 11824
rect 25556 11812 25562 11824
rect 25869 11815 25927 11821
rect 25869 11812 25881 11815
rect 25556 11784 25881 11812
rect 25556 11772 25562 11784
rect 25869 11781 25881 11784
rect 25915 11781 25927 11815
rect 28534 11812 28540 11824
rect 25869 11775 25927 11781
rect 27816 11784 28540 11812
rect 20990 11753 20996 11756
rect 20533 11747 20591 11753
rect 20533 11713 20545 11747
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 20947 11747 20996 11753
rect 20947 11713 20959 11747
rect 20993 11713 20996 11747
rect 20947 11707 20996 11713
rect 17696 11580 19380 11608
rect 20548 11608 20576 11707
rect 20990 11704 20996 11707
rect 21048 11704 21054 11756
rect 21085 11747 21143 11753
rect 21085 11713 21097 11747
rect 21131 11744 21143 11747
rect 21450 11744 21456 11756
rect 21131 11716 21456 11744
rect 21131 11713 21143 11716
rect 21085 11707 21143 11713
rect 21450 11704 21456 11716
rect 21508 11704 21514 11756
rect 22094 11704 22100 11756
rect 22152 11744 22158 11756
rect 22370 11753 22376 11756
rect 22152 11716 22197 11744
rect 22152 11704 22158 11716
rect 22364 11707 22376 11753
rect 22428 11744 22434 11756
rect 23934 11744 23940 11756
rect 22428 11716 22464 11744
rect 23895 11716 23940 11744
rect 22370 11704 22376 11707
rect 22428 11704 22434 11716
rect 23934 11704 23940 11716
rect 23992 11704 23998 11756
rect 27525 11747 27583 11753
rect 27525 11713 27537 11747
rect 27571 11713 27583 11747
rect 27706 11744 27712 11756
rect 27667 11716 27712 11744
rect 27525 11707 27583 11713
rect 20806 11676 20812 11688
rect 20767 11648 20812 11676
rect 20806 11636 20812 11648
rect 20864 11636 20870 11688
rect 27540 11676 27568 11707
rect 27706 11704 27712 11716
rect 27764 11704 27770 11756
rect 27816 11753 27844 11784
rect 28534 11772 28540 11784
rect 28592 11772 28598 11824
rect 27801 11747 27859 11753
rect 27801 11713 27813 11747
rect 27847 11713 27859 11747
rect 28074 11744 28080 11756
rect 28035 11716 28080 11744
rect 27801 11707 27859 11713
rect 28074 11704 28080 11716
rect 28132 11704 28138 11756
rect 28994 11753 29000 11756
rect 28988 11707 29000 11753
rect 29052 11744 29058 11756
rect 29052 11716 29088 11744
rect 28994 11704 29000 11707
rect 29052 11704 29058 11716
rect 27614 11676 27620 11688
rect 27540 11648 27620 11676
rect 27614 11636 27620 11648
rect 27672 11636 27678 11688
rect 27893 11679 27951 11685
rect 27893 11645 27905 11679
rect 27939 11645 27951 11679
rect 28718 11676 28724 11688
rect 28679 11648 28724 11676
rect 27893 11639 27951 11645
rect 21266 11608 21272 11620
rect 20548 11580 21272 11608
rect 15565 11571 15623 11577
rect 21266 11568 21272 11580
rect 21324 11568 21330 11620
rect 26053 11611 26111 11617
rect 22020 11580 22140 11608
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 10229 11543 10287 11549
rect 10229 11540 10241 11543
rect 9640 11512 10241 11540
rect 9640 11500 9646 11512
rect 10229 11509 10241 11512
rect 10275 11509 10287 11543
rect 10229 11503 10287 11509
rect 14737 11543 14795 11549
rect 14737 11509 14749 11543
rect 14783 11540 14795 11543
rect 15286 11540 15292 11552
rect 14783 11512 15292 11540
rect 14783 11509 14795 11512
rect 14737 11503 14795 11509
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 15654 11500 15660 11552
rect 15712 11540 15718 11552
rect 22020 11540 22048 11580
rect 15712 11512 22048 11540
rect 22112 11540 22140 11580
rect 26053 11577 26065 11611
rect 26099 11608 26111 11611
rect 26878 11608 26884 11620
rect 26099 11580 26884 11608
rect 26099 11577 26111 11580
rect 26053 11571 26111 11577
rect 26878 11568 26884 11580
rect 26936 11568 26942 11620
rect 27908 11608 27936 11639
rect 28718 11636 28724 11648
rect 28776 11636 28782 11688
rect 28626 11608 28632 11620
rect 27908 11580 28632 11608
rect 28626 11568 28632 11580
rect 28684 11568 28690 11620
rect 25590 11540 25596 11552
rect 22112 11512 25596 11540
rect 15712 11500 15718 11512
rect 25590 11500 25596 11512
rect 25648 11500 25654 11552
rect 28261 11543 28319 11549
rect 28261 11509 28273 11543
rect 28307 11540 28319 11543
rect 29086 11540 29092 11552
rect 28307 11512 29092 11540
rect 28307 11509 28319 11512
rect 28261 11503 28319 11509
rect 29086 11500 29092 11512
rect 29144 11500 29150 11552
rect 30098 11540 30104 11552
rect 30059 11512 30104 11540
rect 30098 11500 30104 11512
rect 30156 11500 30162 11552
rect 1104 11450 30820 11472
rect 1104 11398 5915 11450
rect 5967 11398 5979 11450
rect 6031 11398 6043 11450
rect 6095 11398 6107 11450
rect 6159 11398 6171 11450
rect 6223 11398 15846 11450
rect 15898 11398 15910 11450
rect 15962 11398 15974 11450
rect 16026 11398 16038 11450
rect 16090 11398 16102 11450
rect 16154 11398 25776 11450
rect 25828 11398 25840 11450
rect 25892 11398 25904 11450
rect 25956 11398 25968 11450
rect 26020 11398 26032 11450
rect 26084 11398 30820 11450
rect 1104 11376 30820 11398
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 10505 11339 10563 11345
rect 10505 11336 10517 11339
rect 10468 11308 10517 11336
rect 10468 11296 10474 11308
rect 10505 11305 10517 11308
rect 10551 11305 10563 11339
rect 11882 11336 11888 11348
rect 11843 11308 11888 11336
rect 10505 11299 10563 11305
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 12526 11336 12532 11348
rect 12406 11308 12532 11336
rect 9401 11271 9459 11277
rect 9401 11268 9413 11271
rect 2148 11240 9413 11268
rect 2148 11141 2176 11240
rect 9401 11237 9413 11240
rect 9447 11237 9459 11271
rect 10597 11271 10655 11277
rect 9401 11231 9459 11237
rect 9508 11240 10548 11268
rect 9508 11200 9536 11240
rect 2746 11172 9536 11200
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1443 11104 2145 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11132 2375 11135
rect 2746 11132 2774 11172
rect 9950 11160 9956 11212
rect 10008 11200 10014 11212
rect 10520 11200 10548 11240
rect 10597 11237 10609 11271
rect 10643 11268 10655 11271
rect 11977 11271 12035 11277
rect 11977 11268 11989 11271
rect 10643 11240 11989 11268
rect 10643 11237 10655 11240
rect 10597 11231 10655 11237
rect 11977 11237 11989 11240
rect 12023 11268 12035 11271
rect 12406 11268 12434 11308
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 16117 11339 16175 11345
rect 16117 11305 16129 11339
rect 16163 11336 16175 11339
rect 16206 11336 16212 11348
rect 16163 11308 16212 11336
rect 16163 11305 16175 11308
rect 16117 11299 16175 11305
rect 16206 11296 16212 11308
rect 16264 11296 16270 11348
rect 16850 11336 16856 11348
rect 16811 11308 16856 11336
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 20809 11339 20867 11345
rect 20809 11305 20821 11339
rect 20855 11336 20867 11339
rect 21358 11336 21364 11348
rect 20855 11308 21364 11336
rect 20855 11305 20867 11308
rect 20809 11299 20867 11305
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 22097 11339 22155 11345
rect 22097 11305 22109 11339
rect 22143 11336 22155 11339
rect 22370 11336 22376 11348
rect 22143 11308 22376 11336
rect 22143 11305 22155 11308
rect 22097 11299 22155 11305
rect 22370 11296 22376 11308
rect 22428 11296 22434 11348
rect 23753 11339 23811 11345
rect 23753 11305 23765 11339
rect 23799 11336 23811 11339
rect 24026 11336 24032 11348
rect 23799 11308 24032 11336
rect 23799 11305 23811 11308
rect 23753 11299 23811 11305
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 25682 11296 25688 11348
rect 25740 11336 25746 11348
rect 25777 11339 25835 11345
rect 25777 11336 25789 11339
rect 25740 11308 25789 11336
rect 25740 11296 25746 11308
rect 25777 11305 25789 11308
rect 25823 11305 25835 11339
rect 25777 11299 25835 11305
rect 26786 11296 26792 11348
rect 26844 11336 26850 11348
rect 26844 11308 28672 11336
rect 26844 11296 26850 11308
rect 12023 11240 12434 11268
rect 12023 11237 12035 11240
rect 11977 11231 12035 11237
rect 19426 11228 19432 11280
rect 19484 11268 19490 11280
rect 20622 11268 20628 11280
rect 19484 11240 20628 11268
rect 19484 11228 19490 11240
rect 20622 11228 20628 11240
rect 20680 11268 20686 11280
rect 21450 11268 21456 11280
rect 20680 11240 21456 11268
rect 20680 11228 20686 11240
rect 21450 11228 21456 11240
rect 21508 11228 21514 11280
rect 26694 11268 26700 11280
rect 26655 11240 26700 11268
rect 26694 11228 26700 11240
rect 26752 11228 26758 11280
rect 27617 11271 27675 11277
rect 27617 11237 27629 11271
rect 27663 11237 27675 11271
rect 28644 11268 28672 11308
rect 28718 11296 28724 11348
rect 28776 11336 28782 11348
rect 29733 11339 29791 11345
rect 29733 11336 29745 11339
rect 28776 11308 29745 11336
rect 28776 11296 28782 11308
rect 29733 11305 29745 11308
rect 29779 11305 29791 11339
rect 29733 11299 29791 11305
rect 28994 11268 29000 11280
rect 28644 11240 28764 11268
rect 28955 11240 29000 11268
rect 27617 11231 27675 11237
rect 11238 11200 11244 11212
rect 10008 11172 10456 11200
rect 10520 11172 11244 11200
rect 10008 11160 10014 11172
rect 9582 11132 9588 11144
rect 2363 11104 2774 11132
rect 9543 11104 9588 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 10134 11132 10140 11144
rect 10095 11104 10140 11132
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10428 11141 10456 11172
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 12986 11200 12992 11212
rect 11716 11172 12992 11200
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11101 10471 11135
rect 10686 11132 10692 11144
rect 10647 11104 10692 11132
rect 10413 11095 10471 11101
rect 2222 11064 2228 11076
rect 2183 11036 2228 11064
rect 2222 11024 2228 11036
rect 2280 11024 2286 11076
rect 10336 11064 10364 11095
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 11514 11132 11520 11144
rect 11475 11104 11520 11132
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11716 11141 11744 11172
rect 12986 11160 12992 11172
rect 13044 11200 13050 11212
rect 14182 11200 14188 11212
rect 13044 11172 14188 11200
rect 13044 11160 13050 11172
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 16482 11200 16488 11212
rect 15948 11172 16488 11200
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 10594 11064 10600 11076
rect 10336 11036 10600 11064
rect 10594 11024 10600 11036
rect 10652 11064 10658 11076
rect 11716 11064 11744 11095
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 12066 11132 12072 11144
rect 11848 11104 11893 11132
rect 12027 11104 12072 11132
rect 11848 11092 11854 11104
rect 12066 11092 12072 11104
rect 12124 11092 12130 11144
rect 15197 11135 15255 11141
rect 15197 11101 15209 11135
rect 15243 11132 15255 11135
rect 15562 11132 15568 11144
rect 15243 11104 15568 11132
rect 15243 11101 15255 11104
rect 15197 11095 15255 11101
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 15948 11141 15976 11172
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 18506 11160 18512 11212
rect 18564 11200 18570 11212
rect 19150 11200 19156 11212
rect 18564 11172 19156 11200
rect 18564 11160 18570 11172
rect 19150 11160 19156 11172
rect 19208 11200 19214 11212
rect 19613 11203 19671 11209
rect 19613 11200 19625 11203
rect 19208 11172 19625 11200
rect 19208 11160 19214 11172
rect 19613 11169 19625 11172
rect 19659 11169 19671 11203
rect 19613 11163 19671 11169
rect 20806 11160 20812 11212
rect 20864 11200 20870 11212
rect 21637 11203 21695 11209
rect 21637 11200 21649 11203
rect 20864 11172 21649 11200
rect 20864 11160 20870 11172
rect 21637 11169 21649 11172
rect 21683 11200 21695 11203
rect 22186 11200 22192 11212
rect 21683 11172 22192 11200
rect 21683 11169 21695 11172
rect 21637 11163 21695 11169
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 23934 11160 23940 11212
rect 23992 11200 23998 11212
rect 24397 11203 24455 11209
rect 24397 11200 24409 11203
rect 23992 11172 24409 11200
rect 23992 11160 23998 11172
rect 24397 11169 24409 11172
rect 24443 11169 24455 11203
rect 24397 11163 24455 11169
rect 26510 11160 26516 11212
rect 26568 11200 26574 11212
rect 27632 11200 27660 11231
rect 26568 11172 27016 11200
rect 27632 11172 28488 11200
rect 26568 11160 26574 11172
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11101 15991 11135
rect 15933 11095 15991 11101
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11132 16175 11135
rect 16298 11132 16304 11144
rect 16163 11104 16304 11132
rect 16163 11101 16175 11104
rect 16117 11095 16175 11101
rect 16298 11092 16304 11104
rect 16356 11132 16362 11144
rect 16761 11135 16819 11141
rect 16761 11132 16773 11135
rect 16356 11104 16773 11132
rect 16356 11092 16362 11104
rect 16761 11101 16773 11104
rect 16807 11101 16819 11135
rect 16761 11095 16819 11101
rect 18782 11092 18788 11144
rect 18840 11132 18846 11144
rect 19242 11132 19248 11144
rect 18840 11104 19248 11132
rect 18840 11092 18846 11104
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 19426 11132 19432 11144
rect 19387 11104 19432 11132
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 10652 11036 11744 11064
rect 10652 11024 10658 11036
rect 14918 11024 14924 11076
rect 14976 11064 14982 11076
rect 18230 11064 18236 11076
rect 14976 11036 18236 11064
rect 14976 11024 14982 11036
rect 18230 11024 18236 11036
rect 18288 11024 18294 11076
rect 18966 11024 18972 11076
rect 19024 11064 19030 11076
rect 19536 11064 19564 11095
rect 19702 11092 19708 11144
rect 19760 11132 19766 11144
rect 19797 11135 19855 11141
rect 19797 11132 19809 11135
rect 19760 11104 19809 11132
rect 19760 11092 19766 11104
rect 19797 11101 19809 11104
rect 19843 11101 19855 11135
rect 20714 11132 20720 11144
rect 20675 11104 20720 11132
rect 19797 11095 19855 11101
rect 20714 11092 20720 11104
rect 20772 11092 20778 11144
rect 21266 11092 21272 11144
rect 21324 11132 21330 11144
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 21324 11104 21373 11132
rect 21324 11092 21330 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21542 11132 21548 11144
rect 21503 11104 21548 11132
rect 21361 11095 21419 11101
rect 21542 11092 21548 11104
rect 21600 11092 21606 11144
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11101 21787 11135
rect 21910 11132 21916 11144
rect 21871 11104 21916 11132
rect 21729 11095 21787 11101
rect 19024 11036 19564 11064
rect 19024 11024 19030 11036
rect 21174 11024 21180 11076
rect 21232 11064 21238 11076
rect 21744 11064 21772 11095
rect 21910 11092 21916 11104
rect 21968 11092 21974 11144
rect 22370 11092 22376 11144
rect 22428 11132 22434 11144
rect 22738 11132 22744 11144
rect 22428 11104 22744 11132
rect 22428 11092 22434 11104
rect 22738 11092 22744 11104
rect 22796 11132 22802 11144
rect 23661 11135 23719 11141
rect 23661 11132 23673 11135
rect 22796 11104 23673 11132
rect 22796 11092 22802 11104
rect 23661 11101 23673 11104
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 24664 11135 24722 11141
rect 24664 11101 24676 11135
rect 24710 11132 24722 11135
rect 25130 11132 25136 11144
rect 24710 11104 25136 11132
rect 24710 11101 24722 11104
rect 24664 11095 24722 11101
rect 25130 11092 25136 11104
rect 25188 11092 25194 11144
rect 25590 11092 25596 11144
rect 25648 11132 25654 11144
rect 26329 11135 26387 11141
rect 26329 11132 26341 11135
rect 25648 11104 26341 11132
rect 25648 11092 25654 11104
rect 26329 11101 26341 11104
rect 26375 11101 26387 11135
rect 26602 11132 26608 11144
rect 26563 11104 26608 11132
rect 26329 11095 26387 11101
rect 26602 11092 26608 11104
rect 26660 11092 26666 11144
rect 26988 11141 27016 11172
rect 26789 11135 26847 11141
rect 26789 11101 26801 11135
rect 26835 11101 26847 11135
rect 26789 11095 26847 11101
rect 26973 11135 27031 11141
rect 26973 11101 26985 11135
rect 27019 11101 27031 11135
rect 27798 11132 27804 11144
rect 27759 11104 27804 11132
rect 26973 11095 27031 11101
rect 21818 11064 21824 11076
rect 21232 11036 21824 11064
rect 21232 11024 21238 11036
rect 21818 11024 21824 11036
rect 21876 11024 21882 11076
rect 1578 10996 1584 11008
rect 1539 10968 1584 10996
rect 1578 10956 1584 10968
rect 1636 10956 1642 11008
rect 15562 10956 15568 11008
rect 15620 10996 15626 11008
rect 16301 10999 16359 11005
rect 16301 10996 16313 10999
rect 15620 10968 16313 10996
rect 15620 10956 15626 10968
rect 16301 10965 16313 10968
rect 16347 10965 16359 10999
rect 16301 10959 16359 10965
rect 19518 10956 19524 11008
rect 19576 10996 19582 11008
rect 19981 10999 20039 11005
rect 19981 10996 19993 10999
rect 19576 10968 19993 10996
rect 19576 10956 19582 10968
rect 19981 10965 19993 10968
rect 20027 10965 20039 10999
rect 26804 10996 26832 11095
rect 27798 11092 27804 11104
rect 27856 11092 27862 11144
rect 28258 11132 28264 11144
rect 28219 11104 28264 11132
rect 28258 11092 28264 11104
rect 28316 11092 28322 11144
rect 28460 11141 28488 11172
rect 28534 11160 28540 11212
rect 28592 11200 28598 11212
rect 28736 11200 28764 11240
rect 28994 11228 29000 11240
rect 29052 11228 29058 11280
rect 30098 11200 30104 11212
rect 28592 11172 28637 11200
rect 28736 11172 30104 11200
rect 28592 11160 28598 11172
rect 28445 11135 28503 11141
rect 28445 11101 28457 11135
rect 28491 11101 28503 11135
rect 28626 11132 28632 11144
rect 28587 11104 28632 11132
rect 28445 11095 28503 11101
rect 28626 11092 28632 11104
rect 28684 11092 28690 11144
rect 28736 11132 28764 11172
rect 30098 11160 30104 11172
rect 30156 11160 30162 11212
rect 28813 11135 28871 11141
rect 28813 11132 28825 11135
rect 28736 11104 28825 11132
rect 28813 11101 28825 11104
rect 28859 11101 28871 11135
rect 28813 11095 28871 11101
rect 26878 11024 26884 11076
rect 26936 11064 26942 11076
rect 29641 11067 29699 11073
rect 29641 11064 29653 11067
rect 26936 11036 29653 11064
rect 26936 11024 26942 11036
rect 29641 11033 29653 11036
rect 29687 11033 29699 11067
rect 29641 11027 29699 11033
rect 28074 10996 28080 11008
rect 26804 10968 28080 10996
rect 19981 10959 20039 10965
rect 28074 10956 28080 10968
rect 28132 10956 28138 11008
rect 1104 10906 30820 10928
rect 1104 10854 10880 10906
rect 10932 10854 10944 10906
rect 10996 10854 11008 10906
rect 11060 10854 11072 10906
rect 11124 10854 11136 10906
rect 11188 10854 20811 10906
rect 20863 10854 20875 10906
rect 20927 10854 20939 10906
rect 20991 10854 21003 10906
rect 21055 10854 21067 10906
rect 21119 10854 30820 10906
rect 1104 10832 30820 10854
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10781 10795 10839 10801
rect 10781 10792 10793 10795
rect 10192 10764 10793 10792
rect 10192 10752 10198 10764
rect 10781 10761 10793 10764
rect 10827 10761 10839 10795
rect 10781 10755 10839 10761
rect 11514 10752 11520 10804
rect 11572 10792 11578 10804
rect 11885 10795 11943 10801
rect 11885 10792 11897 10795
rect 11572 10764 11897 10792
rect 11572 10752 11578 10764
rect 11885 10761 11897 10764
rect 11931 10761 11943 10795
rect 11885 10755 11943 10761
rect 12066 10752 12072 10804
rect 12124 10792 12130 10804
rect 12345 10795 12403 10801
rect 12345 10792 12357 10795
rect 12124 10764 12357 10792
rect 12124 10752 12130 10764
rect 12345 10761 12357 10764
rect 12391 10761 12403 10795
rect 12710 10792 12716 10804
rect 12671 10764 12716 10792
rect 12345 10755 12403 10761
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 21913 10795 21971 10801
rect 21913 10761 21925 10795
rect 21959 10792 21971 10795
rect 22002 10792 22008 10804
rect 21959 10764 22008 10792
rect 21959 10761 21971 10764
rect 21913 10755 21971 10761
rect 22002 10752 22008 10764
rect 22060 10752 22066 10804
rect 26510 10752 26516 10804
rect 26568 10792 26574 10804
rect 26568 10764 27660 10792
rect 26568 10752 26574 10764
rect 10413 10727 10471 10733
rect 10413 10693 10425 10727
rect 10459 10724 10471 10727
rect 10502 10724 10508 10736
rect 10459 10696 10508 10724
rect 10459 10693 10471 10696
rect 10413 10687 10471 10693
rect 10502 10684 10508 10696
rect 10560 10724 10566 10736
rect 19702 10724 19708 10736
rect 10560 10696 11560 10724
rect 10560 10684 10566 10696
rect 10594 10656 10600 10668
rect 10555 10628 10600 10656
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 11532 10665 11560 10696
rect 15764 10696 19708 10724
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10656 11759 10659
rect 12434 10656 12440 10668
rect 11747 10628 12440 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 14918 10656 14924 10668
rect 14879 10628 14924 10656
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 15562 10656 15568 10668
rect 15523 10628 15568 10656
rect 15562 10616 15568 10628
rect 15620 10616 15626 10668
rect 15764 10665 15792 10696
rect 19702 10684 19708 10696
rect 19760 10684 19766 10736
rect 19978 10684 19984 10736
rect 20036 10724 20042 10736
rect 20901 10727 20959 10733
rect 20901 10724 20913 10727
rect 20036 10696 20913 10724
rect 20036 10684 20042 10696
rect 20901 10693 20913 10696
rect 20947 10693 20959 10727
rect 20901 10687 20959 10693
rect 25608 10696 27016 10724
rect 25608 10668 25636 10696
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 12802 10588 12808 10600
rect 12763 10560 12808 10588
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 12986 10588 12992 10600
rect 12947 10560 12992 10588
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 15470 10548 15476 10600
rect 15528 10588 15534 10600
rect 15764 10588 15792 10619
rect 15838 10616 15844 10668
rect 15896 10656 15902 10668
rect 15933 10659 15991 10665
rect 15933 10656 15945 10659
rect 15896 10628 15945 10656
rect 15896 10616 15902 10628
rect 15933 10625 15945 10628
rect 15979 10656 15991 10659
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 15979 10628 16681 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 16942 10616 16948 10668
rect 17000 10656 17006 10668
rect 17589 10659 17647 10665
rect 17589 10656 17601 10659
rect 17000 10628 17601 10656
rect 17000 10616 17006 10628
rect 17589 10625 17601 10628
rect 17635 10625 17647 10659
rect 18506 10656 18512 10668
rect 18467 10628 18512 10656
rect 17589 10619 17647 10625
rect 18506 10616 18512 10628
rect 18564 10616 18570 10668
rect 19242 10616 19248 10668
rect 19300 10656 19306 10668
rect 19797 10659 19855 10665
rect 19797 10656 19809 10659
rect 19300 10628 19809 10656
rect 19300 10616 19306 10628
rect 19797 10625 19809 10628
rect 19843 10625 19855 10659
rect 19797 10619 19855 10625
rect 20622 10616 20628 10668
rect 20680 10656 20686 10668
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 20680 10628 21833 10656
rect 20680 10616 20686 10628
rect 21821 10625 21833 10628
rect 21867 10625 21879 10659
rect 21821 10619 21879 10625
rect 24029 10659 24087 10665
rect 24029 10625 24041 10659
rect 24075 10656 24087 10659
rect 25590 10656 25596 10668
rect 24075 10628 25360 10656
rect 25551 10628 25596 10656
rect 24075 10625 24087 10628
rect 24029 10619 24087 10625
rect 15528 10560 15792 10588
rect 18233 10591 18291 10597
rect 15528 10548 15534 10560
rect 18233 10557 18245 10591
rect 18279 10588 18291 10591
rect 18598 10588 18604 10600
rect 18279 10560 18604 10588
rect 18279 10557 18291 10560
rect 18233 10551 18291 10557
rect 18598 10548 18604 10560
rect 18656 10588 18662 10600
rect 19058 10588 19064 10600
rect 18656 10560 19064 10588
rect 18656 10548 18662 10560
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 19521 10591 19579 10597
rect 19521 10557 19533 10591
rect 19567 10588 19579 10591
rect 20438 10588 20444 10600
rect 19567 10560 20444 10588
rect 19567 10557 19579 10560
rect 19521 10551 19579 10557
rect 20438 10548 20444 10560
rect 20496 10548 20502 10600
rect 21085 10591 21143 10597
rect 21085 10557 21097 10591
rect 21131 10588 21143 10591
rect 21910 10588 21916 10600
rect 21131 10560 21916 10588
rect 21131 10557 21143 10560
rect 21085 10551 21143 10557
rect 21910 10548 21916 10560
rect 21968 10548 21974 10600
rect 17773 10523 17831 10529
rect 17773 10489 17785 10523
rect 17819 10520 17831 10523
rect 18966 10520 18972 10532
rect 17819 10492 18972 10520
rect 17819 10489 17831 10492
rect 17773 10483 17831 10489
rect 18966 10480 18972 10492
rect 19024 10480 19030 10532
rect 20456 10520 20484 10548
rect 24044 10520 24072 10619
rect 24210 10548 24216 10600
rect 24268 10588 24274 10600
rect 24305 10591 24363 10597
rect 24305 10588 24317 10591
rect 24268 10560 24317 10588
rect 24268 10548 24274 10560
rect 24305 10557 24317 10560
rect 24351 10557 24363 10591
rect 25332 10588 25360 10628
rect 25590 10616 25596 10628
rect 25648 10616 25654 10668
rect 25682 10616 25688 10668
rect 25740 10656 25746 10668
rect 25777 10659 25835 10665
rect 25777 10656 25789 10659
rect 25740 10628 25789 10656
rect 25740 10616 25746 10628
rect 25777 10625 25789 10628
rect 25823 10625 25835 10659
rect 25777 10619 25835 10625
rect 26145 10659 26203 10665
rect 26145 10625 26157 10659
rect 26191 10625 26203 10659
rect 26145 10619 26203 10625
rect 26421 10659 26479 10665
rect 26421 10625 26433 10659
rect 26467 10656 26479 10659
rect 26510 10656 26516 10668
rect 26467 10628 26516 10656
rect 26467 10625 26479 10628
rect 26421 10619 26479 10625
rect 26050 10588 26056 10600
rect 25332 10560 26056 10588
rect 24305 10551 24363 10557
rect 26050 10548 26056 10560
rect 26108 10548 26114 10600
rect 26160 10588 26188 10619
rect 26510 10616 26516 10628
rect 26568 10616 26574 10668
rect 26988 10665 27016 10696
rect 26973 10659 27031 10665
rect 26973 10625 26985 10659
rect 27019 10625 27031 10659
rect 27154 10656 27160 10668
rect 27115 10628 27160 10656
rect 26973 10619 27031 10625
rect 27154 10616 27160 10628
rect 27212 10616 27218 10668
rect 27632 10665 27660 10764
rect 28074 10752 28080 10804
rect 28132 10792 28138 10804
rect 30101 10795 30159 10801
rect 30101 10792 30113 10795
rect 28132 10764 30113 10792
rect 28132 10752 28138 10764
rect 30101 10761 30113 10764
rect 30147 10761 30159 10795
rect 30101 10755 30159 10761
rect 28988 10727 29046 10733
rect 28988 10693 29000 10727
rect 29034 10724 29046 10727
rect 29086 10724 29092 10736
rect 29034 10696 29092 10724
rect 29034 10693 29046 10696
rect 28988 10687 29046 10693
rect 29086 10684 29092 10696
rect 29144 10684 29150 10736
rect 27525 10659 27583 10665
rect 27525 10625 27537 10659
rect 27571 10625 27583 10659
rect 27525 10619 27583 10625
rect 27617 10659 27675 10665
rect 27617 10625 27629 10659
rect 27663 10625 27675 10659
rect 27617 10619 27675 10625
rect 26786 10588 26792 10600
rect 26160 10560 26792 10588
rect 26786 10548 26792 10560
rect 26844 10548 26850 10600
rect 27062 10588 27068 10600
rect 27023 10560 27068 10588
rect 27062 10548 27068 10560
rect 27120 10548 27126 10600
rect 27540 10588 27568 10619
rect 28534 10588 28540 10600
rect 27540 10560 28540 10588
rect 28534 10548 28540 10560
rect 28592 10548 28598 10600
rect 28718 10588 28724 10600
rect 28679 10560 28724 10588
rect 28718 10548 28724 10560
rect 28776 10548 28782 10600
rect 20456 10492 24072 10520
rect 24578 10480 24584 10532
rect 24636 10520 24642 10532
rect 25593 10523 25651 10529
rect 25593 10520 25605 10523
rect 24636 10492 25605 10520
rect 24636 10480 24642 10492
rect 25593 10489 25605 10492
rect 25639 10489 25651 10523
rect 25593 10483 25651 10489
rect 15013 10455 15071 10461
rect 15013 10421 15025 10455
rect 15059 10452 15071 10455
rect 15654 10452 15660 10464
rect 15059 10424 15660 10452
rect 15059 10421 15071 10424
rect 15013 10415 15071 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 16206 10412 16212 10464
rect 16264 10452 16270 10464
rect 16761 10455 16819 10461
rect 16761 10452 16773 10455
rect 16264 10424 16773 10452
rect 16264 10412 16270 10424
rect 16761 10421 16773 10424
rect 16807 10421 16819 10455
rect 16761 10415 16819 10421
rect 1104 10362 30820 10384
rect 1104 10310 5915 10362
rect 5967 10310 5979 10362
rect 6031 10310 6043 10362
rect 6095 10310 6107 10362
rect 6159 10310 6171 10362
rect 6223 10310 15846 10362
rect 15898 10310 15910 10362
rect 15962 10310 15974 10362
rect 16026 10310 16038 10362
rect 16090 10310 16102 10362
rect 16154 10310 25776 10362
rect 25828 10310 25840 10362
rect 25892 10310 25904 10362
rect 25956 10310 25968 10362
rect 26020 10310 26032 10362
rect 26084 10310 30820 10362
rect 1104 10288 30820 10310
rect 10597 10251 10655 10257
rect 10597 10217 10609 10251
rect 10643 10248 10655 10251
rect 10686 10248 10692 10260
rect 10643 10220 10692 10248
rect 10643 10217 10655 10220
rect 10597 10211 10655 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 12986 10248 12992 10260
rect 12492 10220 12537 10248
rect 12820 10220 12992 10248
rect 12492 10208 12498 10220
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 10744 10084 11253 10112
rect 10744 10072 10750 10084
rect 11241 10081 11253 10084
rect 11287 10112 11299 10115
rect 12820 10112 12848 10220
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 14093 10251 14151 10257
rect 14093 10217 14105 10251
rect 14139 10248 14151 10251
rect 14274 10248 14280 10260
rect 14139 10220 14280 10248
rect 14139 10217 14151 10220
rect 14093 10211 14151 10217
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 16574 10248 16580 10260
rect 14884 10220 16436 10248
rect 16535 10220 16580 10248
rect 14884 10208 14890 10220
rect 15933 10183 15991 10189
rect 15933 10180 15945 10183
rect 12912 10152 15945 10180
rect 12912 10121 12940 10152
rect 15933 10149 15945 10152
rect 15979 10149 15991 10183
rect 15933 10143 15991 10149
rect 11287 10084 12848 10112
rect 12897 10115 12955 10121
rect 11287 10081 11299 10084
rect 11241 10075 11299 10081
rect 12897 10081 12909 10115
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 12986 10072 12992 10124
rect 13044 10112 13050 10124
rect 14734 10112 14740 10124
rect 13044 10084 13089 10112
rect 14695 10084 14740 10112
rect 13044 10072 13050 10084
rect 14734 10072 14740 10084
rect 14792 10072 14798 10124
rect 16206 10112 16212 10124
rect 15672 10084 16212 10112
rect 10502 10004 10508 10056
rect 10560 10044 10566 10056
rect 10870 10044 10876 10056
rect 10560 10016 10876 10044
rect 10560 10004 10566 10016
rect 10870 10004 10876 10016
rect 10928 10044 10934 10056
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10928 10016 10977 10044
rect 10928 10004 10934 10016
rect 10965 10013 10977 10016
rect 11011 10013 11023 10047
rect 10965 10007 11023 10013
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12768 10016 12817 10044
rect 12768 10004 12774 10016
rect 12805 10013 12817 10016
rect 12851 10013 12863 10047
rect 15286 10044 15292 10056
rect 15247 10016 15292 10044
rect 12805 10007 12863 10013
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 15437 10047 15495 10053
rect 15437 10013 15449 10047
rect 15483 10044 15495 10047
rect 15672 10044 15700 10084
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 15483 10016 15700 10044
rect 15483 10013 15495 10016
rect 15437 10007 15495 10013
rect 15746 10004 15752 10056
rect 15804 10053 15810 10056
rect 15804 10044 15812 10053
rect 16408 10044 16436 10220
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 18414 10248 18420 10260
rect 18375 10220 18420 10248
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 19426 10248 19432 10260
rect 19260 10220 19432 10248
rect 16592 10180 16620 10208
rect 19260 10180 19288 10220
rect 19426 10208 19432 10220
rect 19484 10248 19490 10260
rect 20622 10248 20628 10260
rect 19484 10220 20628 10248
rect 19484 10208 19490 10220
rect 20622 10208 20628 10220
rect 20680 10208 20686 10260
rect 28534 10248 28540 10260
rect 28495 10220 28540 10248
rect 28534 10208 28540 10220
rect 28592 10208 28598 10260
rect 22186 10180 22192 10192
rect 16592 10152 17264 10180
rect 16485 10047 16543 10053
rect 16485 10044 16497 10047
rect 15804 10016 15849 10044
rect 16408 10016 16497 10044
rect 15804 10007 15812 10016
rect 16485 10013 16497 10016
rect 16531 10044 16543 10047
rect 16942 10044 16948 10056
rect 16531 10016 16948 10044
rect 16531 10013 16543 10016
rect 16485 10007 16543 10013
rect 15804 10004 15810 10007
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17126 10044 17132 10056
rect 17087 10016 17132 10044
rect 17126 10004 17132 10016
rect 17184 10004 17190 10056
rect 17236 10053 17264 10152
rect 17328 10152 19288 10180
rect 21652 10152 22192 10180
rect 17222 10047 17280 10053
rect 17222 10013 17234 10047
rect 17268 10013 17280 10047
rect 17222 10007 17280 10013
rect 10778 9936 10784 9988
rect 10836 9976 10842 9988
rect 11057 9979 11115 9985
rect 11057 9976 11069 9979
rect 10836 9948 11069 9976
rect 10836 9936 10842 9948
rect 11057 9945 11069 9948
rect 11103 9945 11115 9979
rect 11057 9939 11115 9945
rect 14461 9979 14519 9985
rect 14461 9945 14473 9979
rect 14507 9976 14519 9979
rect 15194 9976 15200 9988
rect 14507 9948 15200 9976
rect 14507 9945 14519 9948
rect 14461 9939 14519 9945
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 15565 9979 15623 9985
rect 15565 9945 15577 9979
rect 15611 9945 15623 9979
rect 15565 9939 15623 9945
rect 14090 9868 14096 9920
rect 14148 9908 14154 9920
rect 14553 9911 14611 9917
rect 14553 9908 14565 9911
rect 14148 9880 14565 9908
rect 14148 9868 14154 9880
rect 14553 9877 14565 9880
rect 14599 9877 14611 9911
rect 14553 9871 14611 9877
rect 14918 9868 14924 9920
rect 14976 9908 14982 9920
rect 15580 9908 15608 9939
rect 15654 9936 15660 9988
rect 15712 9976 15718 9988
rect 17328 9976 17356 10152
rect 18046 10112 18052 10124
rect 17420 10084 18052 10112
rect 17420 10053 17448 10084
rect 18046 10072 18052 10084
rect 18104 10072 18110 10124
rect 21174 10072 21180 10124
rect 21232 10112 21238 10124
rect 21652 10121 21680 10152
rect 22186 10140 22192 10152
rect 22244 10140 22250 10192
rect 21637 10115 21695 10121
rect 21637 10112 21649 10115
rect 21232 10084 21649 10112
rect 21232 10072 21238 10084
rect 21637 10081 21649 10084
rect 21683 10081 21695 10115
rect 21637 10075 21695 10081
rect 21729 10115 21787 10121
rect 21729 10081 21741 10115
rect 21775 10112 21787 10115
rect 21818 10112 21824 10124
rect 21775 10084 21824 10112
rect 21775 10081 21787 10084
rect 21729 10075 21787 10081
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 24949 10115 25007 10121
rect 24949 10081 24961 10115
rect 24995 10112 25007 10115
rect 26970 10112 26976 10124
rect 24995 10084 26976 10112
rect 24995 10081 25007 10084
rect 24949 10075 25007 10081
rect 26970 10072 26976 10084
rect 27028 10072 27034 10124
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10013 17463 10047
rect 17405 10007 17463 10013
rect 17635 10047 17693 10053
rect 17635 10013 17647 10047
rect 17681 10044 17693 10047
rect 19058 10044 19064 10056
rect 17681 10016 19064 10044
rect 17681 10013 17693 10016
rect 17635 10007 17693 10013
rect 19058 10004 19064 10016
rect 19116 10004 19122 10056
rect 19245 10047 19303 10053
rect 19245 10013 19257 10047
rect 19291 10044 19303 10047
rect 19334 10044 19340 10056
rect 19291 10016 19340 10044
rect 19291 10013 19303 10016
rect 19245 10007 19303 10013
rect 19334 10004 19340 10016
rect 19392 10004 19398 10056
rect 19518 10053 19524 10056
rect 19512 10044 19524 10053
rect 19479 10016 19524 10044
rect 19512 10007 19524 10016
rect 19518 10004 19524 10007
rect 19576 10004 19582 10056
rect 21266 10004 21272 10056
rect 21324 10044 21330 10056
rect 21361 10047 21419 10053
rect 21361 10044 21373 10047
rect 21324 10016 21373 10044
rect 21324 10004 21330 10016
rect 21361 10013 21373 10016
rect 21407 10013 21419 10047
rect 21361 10007 21419 10013
rect 21450 10004 21456 10056
rect 21508 10044 21514 10056
rect 21545 10047 21603 10053
rect 21545 10044 21557 10047
rect 21508 10016 21557 10044
rect 21508 10004 21514 10016
rect 21545 10013 21557 10016
rect 21591 10013 21603 10047
rect 21545 10007 21603 10013
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10013 21971 10047
rect 25222 10044 25228 10056
rect 25183 10016 25228 10044
rect 21913 10007 21971 10013
rect 17497 9979 17555 9985
rect 17497 9976 17509 9979
rect 15712 9948 15757 9976
rect 17328 9948 17509 9976
rect 15712 9936 15718 9948
rect 17497 9945 17509 9948
rect 17543 9945 17555 9979
rect 17954 9976 17960 9988
rect 17497 9939 17555 9945
rect 17604 9948 17960 9976
rect 17604 9908 17632 9948
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 18322 9976 18328 9988
rect 18283 9948 18328 9976
rect 18322 9936 18328 9948
rect 18380 9936 18386 9988
rect 21928 9976 21956 10007
rect 25222 10004 25228 10016
rect 25280 10004 25286 10056
rect 26329 10047 26387 10053
rect 26329 10013 26341 10047
rect 26375 10044 26387 10047
rect 26878 10044 26884 10056
rect 26375 10016 26884 10044
rect 26375 10013 26387 10016
rect 26329 10007 26387 10013
rect 26878 10004 26884 10016
rect 26936 10004 26942 10056
rect 27157 10047 27215 10053
rect 27157 10013 27169 10047
rect 27203 10044 27215 10047
rect 28718 10044 28724 10056
rect 27203 10016 28724 10044
rect 27203 10013 27215 10016
rect 27157 10007 27215 10013
rect 28718 10004 28724 10016
rect 28776 10004 28782 10056
rect 30098 10044 30104 10056
rect 30059 10016 30104 10044
rect 30098 10004 30104 10016
rect 30156 10004 30162 10056
rect 21284 9948 21956 9976
rect 27424 9979 27482 9985
rect 21284 9920 21312 9948
rect 27424 9945 27436 9979
rect 27470 9976 27482 9979
rect 27522 9976 27528 9988
rect 27470 9948 27528 9976
rect 27470 9945 27482 9948
rect 27424 9939 27482 9945
rect 27522 9936 27528 9948
rect 27580 9936 27586 9988
rect 17770 9908 17776 9920
rect 14976 9880 17632 9908
rect 17731 9880 17776 9908
rect 14976 9868 14982 9880
rect 17770 9868 17776 9880
rect 17828 9868 17834 9920
rect 19702 9868 19708 9920
rect 19760 9908 19766 9920
rect 20625 9911 20683 9917
rect 20625 9908 20637 9911
rect 19760 9880 20637 9908
rect 19760 9868 19766 9880
rect 20625 9877 20637 9880
rect 20671 9877 20683 9911
rect 20625 9871 20683 9877
rect 21266 9868 21272 9920
rect 21324 9868 21330 9920
rect 22097 9911 22155 9917
rect 22097 9877 22109 9911
rect 22143 9908 22155 9911
rect 22278 9908 22284 9920
rect 22143 9880 22284 9908
rect 22143 9877 22155 9880
rect 22097 9871 22155 9877
rect 22278 9868 22284 9880
rect 22336 9868 22342 9920
rect 23934 9868 23940 9920
rect 23992 9908 23998 9920
rect 26421 9911 26479 9917
rect 26421 9908 26433 9911
rect 23992 9880 26433 9908
rect 23992 9868 23998 9880
rect 26421 9877 26433 9880
rect 26467 9877 26479 9911
rect 26421 9871 26479 9877
rect 29270 9868 29276 9920
rect 29328 9908 29334 9920
rect 29917 9911 29975 9917
rect 29917 9908 29929 9911
rect 29328 9880 29929 9908
rect 29328 9868 29334 9880
rect 29917 9877 29929 9880
rect 29963 9877 29975 9911
rect 29917 9871 29975 9877
rect 1104 9818 30820 9840
rect 1104 9766 10880 9818
rect 10932 9766 10944 9818
rect 10996 9766 11008 9818
rect 11060 9766 11072 9818
rect 11124 9766 11136 9818
rect 11188 9766 20811 9818
rect 20863 9766 20875 9818
rect 20927 9766 20939 9818
rect 20991 9766 21003 9818
rect 21055 9766 21067 9818
rect 21119 9766 30820 9818
rect 1104 9744 30820 9766
rect 10229 9707 10287 9713
rect 10229 9673 10241 9707
rect 10275 9704 10287 9707
rect 10594 9704 10600 9716
rect 10275 9676 10600 9704
rect 10275 9673 10287 9676
rect 10229 9667 10287 9673
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 12621 9707 12679 9713
rect 12621 9673 12633 9707
rect 12667 9704 12679 9707
rect 12802 9704 12808 9716
rect 12667 9676 12808 9704
rect 12667 9673 12679 9676
rect 12621 9667 12679 9673
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 15194 9664 15200 9716
rect 15252 9704 15258 9716
rect 15841 9707 15899 9713
rect 15841 9704 15853 9707
rect 15252 9676 15853 9704
rect 15252 9664 15258 9676
rect 15841 9673 15853 9676
rect 15887 9673 15899 9707
rect 18046 9704 18052 9716
rect 18007 9676 18052 9704
rect 15841 9667 15899 9673
rect 18046 9664 18052 9676
rect 18104 9664 18110 9716
rect 25317 9707 25375 9713
rect 25317 9673 25329 9707
rect 25363 9704 25375 9707
rect 25363 9676 25397 9704
rect 25363 9673 25375 9676
rect 25317 9667 25375 9673
rect 10686 9596 10692 9648
rect 10744 9636 10750 9648
rect 14369 9639 14427 9645
rect 10744 9608 10824 9636
rect 10744 9596 10750 9608
rect 10502 9528 10508 9580
rect 10560 9568 10566 9580
rect 10597 9571 10655 9577
rect 10597 9568 10609 9571
rect 10560 9540 10609 9568
rect 10560 9528 10566 9540
rect 10597 9537 10609 9540
rect 10643 9537 10655 9571
rect 10597 9531 10655 9537
rect 10796 9509 10824 9608
rect 14369 9605 14381 9639
rect 14415 9636 14427 9639
rect 16936 9639 16994 9645
rect 14415 9608 16068 9636
rect 14415 9605 14427 9608
rect 14369 9599 14427 9605
rect 12158 9568 12164 9580
rect 12119 9540 12164 9568
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12406 9540 13001 9568
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9469 10747 9503
rect 10689 9463 10747 9469
rect 10781 9503 10839 9509
rect 10781 9469 10793 9503
rect 10827 9469 10839 9503
rect 10781 9463 10839 9469
rect 10704 9364 10732 9463
rect 11977 9435 12035 9441
rect 11977 9401 11989 9435
rect 12023 9432 12035 9435
rect 12406 9432 12434 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9568 14059 9571
rect 14090 9568 14096 9580
rect 14047 9540 14096 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 14185 9571 14243 9577
rect 14185 9537 14197 9571
rect 14231 9568 14243 9571
rect 14642 9568 14648 9580
rect 14231 9540 14648 9568
rect 14231 9537 14243 9540
rect 14185 9531 14243 9537
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9568 15163 9571
rect 15194 9568 15200 9580
rect 15151 9540 15200 9568
rect 15151 9537 15163 9540
rect 15105 9531 15163 9537
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15289 9571 15347 9577
rect 15289 9537 15301 9571
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 13081 9503 13139 9509
rect 13081 9500 13093 9503
rect 12768 9472 13093 9500
rect 12768 9460 12774 9472
rect 13081 9469 13093 9472
rect 13127 9469 13139 9503
rect 13081 9463 13139 9469
rect 13262 9460 13268 9512
rect 13320 9500 13326 9512
rect 14734 9500 14740 9512
rect 13320 9472 14740 9500
rect 13320 9460 13326 9472
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 15304 9500 15332 9531
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 16040 9577 16068 9608
rect 16936 9605 16948 9639
rect 16982 9636 16994 9639
rect 17770 9636 17776 9648
rect 16982 9608 17776 9636
rect 16982 9605 16994 9608
rect 16936 9599 16994 9605
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 17954 9596 17960 9648
rect 18012 9636 18018 9648
rect 18012 9608 18828 9636
rect 18012 9596 18018 9608
rect 18800 9580 18828 9608
rect 19904 9608 22048 9636
rect 16025 9571 16083 9577
rect 15436 9540 15481 9568
rect 15436 9528 15442 9540
rect 16025 9537 16037 9571
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 18230 9528 18236 9580
rect 18288 9568 18294 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18288 9540 18521 9568
rect 18288 9528 18294 9540
rect 18509 9537 18521 9540
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 18598 9528 18604 9580
rect 18656 9568 18662 9580
rect 18782 9568 18788 9580
rect 18656 9540 18701 9568
rect 18743 9540 18788 9568
rect 18656 9528 18662 9540
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 19058 9577 19064 9580
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9537 18935 9571
rect 18877 9531 18935 9537
rect 19015 9571 19064 9577
rect 19015 9537 19027 9571
rect 19061 9537 19064 9571
rect 19015 9531 19064 9537
rect 15746 9500 15752 9512
rect 15304 9472 15752 9500
rect 15746 9460 15752 9472
rect 15804 9460 15810 9512
rect 16666 9500 16672 9512
rect 16627 9472 16672 9500
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 14921 9435 14979 9441
rect 14921 9432 14933 9435
rect 12023 9404 12434 9432
rect 13648 9404 14933 9432
rect 12023 9401 12035 9404
rect 11977 9395 12035 9401
rect 13648 9364 13676 9404
rect 14921 9401 14933 9404
rect 14967 9401 14979 9435
rect 18892 9432 18920 9531
rect 19058 9528 19064 9531
rect 19116 9528 19122 9580
rect 19334 9528 19340 9580
rect 19392 9568 19398 9580
rect 19904 9577 19932 9608
rect 19889 9571 19947 9577
rect 19889 9568 19901 9571
rect 19392 9540 19901 9568
rect 19392 9528 19398 9540
rect 19889 9537 19901 9540
rect 19935 9537 19947 9571
rect 19889 9531 19947 9537
rect 20156 9571 20214 9577
rect 20156 9537 20168 9571
rect 20202 9568 20214 9571
rect 21358 9568 21364 9580
rect 20202 9540 21364 9568
rect 20202 9537 20214 9540
rect 20156 9531 20214 9537
rect 21358 9528 21364 9540
rect 21416 9528 21422 9580
rect 22020 9577 22048 9608
rect 22370 9596 22376 9648
rect 22428 9636 22434 9648
rect 25332 9636 25360 9667
rect 22428 9608 25360 9636
rect 26237 9639 26295 9645
rect 22428 9596 22434 9608
rect 26237 9605 26249 9639
rect 26283 9636 26295 9639
rect 26970 9636 26976 9648
rect 26283 9608 26976 9636
rect 26283 9605 26295 9608
rect 26237 9599 26295 9605
rect 26970 9596 26976 9608
rect 27028 9596 27034 9648
rect 22005 9571 22063 9577
rect 22005 9537 22017 9571
rect 22051 9568 22063 9571
rect 22094 9568 22100 9580
rect 22051 9540 22100 9568
rect 22051 9537 22063 9540
rect 22005 9531 22063 9537
rect 22094 9528 22100 9540
rect 22152 9528 22158 9580
rect 22278 9577 22284 9580
rect 22272 9568 22284 9577
rect 22239 9540 22284 9568
rect 22272 9531 22284 9540
rect 22278 9528 22284 9531
rect 22336 9528 22342 9580
rect 23934 9568 23940 9580
rect 23895 9540 23940 9568
rect 23934 9528 23940 9540
rect 23992 9528 23998 9580
rect 24026 9528 24032 9580
rect 24084 9568 24090 9580
rect 24193 9571 24251 9577
rect 24193 9568 24205 9571
rect 24084 9540 24205 9568
rect 24084 9528 24090 9540
rect 24193 9537 24205 9540
rect 24239 9537 24251 9571
rect 24193 9531 24251 9537
rect 26142 9528 26148 9580
rect 26200 9568 26206 9580
rect 27433 9571 27491 9577
rect 27433 9568 27445 9571
rect 26200 9540 27445 9568
rect 26200 9528 26206 9540
rect 27433 9537 27445 9540
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 27614 9528 27620 9580
rect 27672 9568 27678 9580
rect 27709 9571 27767 9577
rect 27709 9568 27721 9571
rect 27672 9540 27721 9568
rect 27672 9528 27678 9540
rect 27709 9537 27721 9540
rect 27755 9537 27767 9571
rect 27709 9531 27767 9537
rect 28988 9571 29046 9577
rect 28988 9537 29000 9571
rect 29034 9568 29046 9571
rect 29546 9568 29552 9580
rect 29034 9540 29552 9568
rect 29034 9537 29046 9540
rect 28988 9531 29046 9537
rect 29546 9528 29552 9540
rect 29604 9528 29610 9580
rect 21266 9460 21272 9512
rect 21324 9500 21330 9512
rect 28718 9500 28724 9512
rect 21324 9472 21404 9500
rect 28679 9472 28724 9500
rect 21324 9460 21330 9472
rect 18892 9404 19932 9432
rect 14921 9395 14979 9401
rect 19150 9364 19156 9376
rect 10704 9336 13676 9364
rect 19111 9336 19156 9364
rect 19150 9324 19156 9336
rect 19208 9324 19214 9376
rect 19904 9364 19932 9404
rect 20622 9364 20628 9376
rect 19904 9336 20628 9364
rect 20622 9324 20628 9336
rect 20680 9324 20686 9376
rect 20806 9324 20812 9376
rect 20864 9364 20870 9376
rect 20990 9364 20996 9376
rect 20864 9336 20996 9364
rect 20864 9324 20870 9336
rect 20990 9324 20996 9336
rect 21048 9364 21054 9376
rect 21269 9367 21327 9373
rect 21269 9364 21281 9367
rect 21048 9336 21281 9364
rect 21048 9324 21054 9336
rect 21269 9333 21281 9336
rect 21315 9333 21327 9367
rect 21376 9364 21404 9472
rect 28718 9460 28724 9472
rect 28776 9460 28782 9512
rect 23198 9392 23204 9444
rect 23256 9432 23262 9444
rect 26421 9435 26479 9441
rect 23256 9404 23980 9432
rect 23256 9392 23262 9404
rect 23385 9367 23443 9373
rect 23385 9364 23397 9367
rect 21376 9336 23397 9364
rect 21269 9327 21327 9333
rect 23385 9333 23397 9336
rect 23431 9333 23443 9367
rect 23952 9364 23980 9404
rect 26421 9401 26433 9435
rect 26467 9432 26479 9435
rect 28074 9432 28080 9444
rect 26467 9404 28080 9432
rect 26467 9401 26479 9404
rect 26421 9395 26479 9401
rect 28074 9392 28080 9404
rect 28132 9392 28138 9444
rect 30006 9392 30012 9444
rect 30064 9432 30070 9444
rect 30101 9435 30159 9441
rect 30101 9432 30113 9435
rect 30064 9404 30113 9432
rect 30064 9392 30070 9404
rect 30101 9401 30113 9404
rect 30147 9401 30159 9435
rect 30101 9395 30159 9401
rect 24210 9364 24216 9376
rect 23952 9336 24216 9364
rect 23385 9327 23443 9333
rect 24210 9324 24216 9336
rect 24268 9324 24274 9376
rect 1104 9274 30820 9296
rect 1104 9222 5915 9274
rect 5967 9222 5979 9274
rect 6031 9222 6043 9274
rect 6095 9222 6107 9274
rect 6159 9222 6171 9274
rect 6223 9222 15846 9274
rect 15898 9222 15910 9274
rect 15962 9222 15974 9274
rect 16026 9222 16038 9274
rect 16090 9222 16102 9274
rect 16154 9222 25776 9274
rect 25828 9222 25840 9274
rect 25892 9222 25904 9274
rect 25956 9222 25968 9274
rect 26020 9222 26032 9274
rect 26084 9222 30820 9274
rect 1104 9200 30820 9222
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 10965 9163 11023 9169
rect 10965 9160 10977 9163
rect 10836 9132 10977 9160
rect 10836 9120 10842 9132
rect 10965 9129 10977 9132
rect 11011 9129 11023 9163
rect 10965 9123 11023 9129
rect 12158 9120 12164 9172
rect 12216 9160 12222 9172
rect 13173 9163 13231 9169
rect 13173 9160 13185 9163
rect 12216 9132 13185 9160
rect 12216 9120 12222 9132
rect 13173 9129 13185 9132
rect 13219 9129 13231 9163
rect 13173 9123 13231 9129
rect 13998 9120 14004 9172
rect 14056 9160 14062 9172
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 14056 9132 14197 9160
rect 14056 9120 14062 9132
rect 14185 9129 14197 9132
rect 14231 9129 14243 9163
rect 14185 9123 14243 9129
rect 15378 9120 15384 9172
rect 15436 9160 15442 9172
rect 15657 9163 15715 9169
rect 15657 9160 15669 9163
rect 15436 9132 15669 9160
rect 15436 9120 15442 9132
rect 15657 9129 15669 9132
rect 15703 9129 15715 9163
rect 15657 9123 15715 9129
rect 16853 9163 16911 9169
rect 16853 9129 16865 9163
rect 16899 9160 16911 9163
rect 18322 9160 18328 9172
rect 16899 9132 18328 9160
rect 16899 9129 16911 9132
rect 16853 9123 16911 9129
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 19058 9120 19064 9172
rect 19116 9160 19122 9172
rect 19797 9163 19855 9169
rect 19797 9160 19809 9163
rect 19116 9132 19809 9160
rect 19116 9120 19122 9132
rect 19797 9129 19809 9132
rect 19843 9129 19855 9163
rect 19797 9123 19855 9129
rect 22186 9120 22192 9172
rect 22244 9120 22250 9172
rect 22557 9163 22615 9169
rect 22557 9129 22569 9163
rect 22603 9160 22615 9163
rect 24026 9160 24032 9172
rect 22603 9132 24032 9160
rect 22603 9129 22615 9132
rect 22557 9123 22615 9129
rect 24026 9120 24032 9132
rect 24084 9120 24090 9172
rect 28166 9120 28172 9172
rect 28224 9160 28230 9172
rect 28629 9163 28687 9169
rect 28629 9160 28641 9163
rect 28224 9132 28641 9160
rect 28224 9120 28230 9132
rect 28629 9129 28641 9132
rect 28675 9129 28687 9163
rect 28629 9123 28687 9129
rect 21358 9052 21364 9104
rect 21416 9092 21422 9104
rect 22204 9092 22232 9120
rect 21416 9064 21461 9092
rect 21928 9064 22232 9092
rect 21416 9052 21422 9064
rect 11609 9027 11667 9033
rect 11609 8993 11621 9027
rect 11655 9024 11667 9027
rect 13262 9024 13268 9036
rect 11655 8996 13268 9024
rect 11655 8993 11667 8996
rect 11609 8987 11667 8993
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 14734 8984 14740 9036
rect 14792 9024 14798 9036
rect 14829 9027 14887 9033
rect 14829 9024 14841 9027
rect 14792 8996 14841 9024
rect 14792 8984 14798 8996
rect 14829 8993 14841 8996
rect 14875 8993 14887 9027
rect 14829 8987 14887 8993
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 2222 8956 2228 8968
rect 1443 8928 2228 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 11756 8928 13001 8956
rect 11756 8916 11762 8928
rect 12989 8925 13001 8928
rect 13035 8956 13047 8959
rect 14642 8956 14648 8968
rect 13035 8928 14648 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 14642 8916 14648 8928
rect 14700 8916 14706 8968
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 12805 8891 12863 8897
rect 12805 8888 12817 8891
rect 12768 8860 12817 8888
rect 12768 8848 12774 8860
rect 12805 8857 12817 8860
rect 12851 8857 12863 8891
rect 14844 8888 14872 8987
rect 15470 8984 15476 9036
rect 15528 9024 15534 9036
rect 15528 8996 15792 9024
rect 15528 8984 15534 8996
rect 15562 8956 15568 8968
rect 15523 8928 15568 8956
rect 15562 8916 15568 8928
rect 15620 8916 15626 8968
rect 15764 8965 15792 8996
rect 16942 8984 16948 9036
rect 17000 9024 17006 9036
rect 17405 9027 17463 9033
rect 17405 9024 17417 9027
rect 17000 8996 17417 9024
rect 17000 8984 17006 8996
rect 17405 8993 17417 8996
rect 17451 8993 17463 9027
rect 17405 8987 17463 8993
rect 17494 8984 17500 9036
rect 17552 9024 17558 9036
rect 17681 9027 17739 9033
rect 17681 9024 17693 9027
rect 17552 8996 17693 9024
rect 17552 8984 17558 8996
rect 17681 8993 17693 8996
rect 17727 9024 17739 9027
rect 18598 9024 18604 9036
rect 17727 8996 18604 9024
rect 17727 8993 17739 8996
rect 17681 8987 17739 8993
rect 18598 8984 18604 8996
rect 18656 8984 18662 9036
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 16761 8959 16819 8965
rect 16761 8925 16773 8959
rect 16807 8956 16819 8959
rect 16960 8956 16988 8984
rect 16807 8928 16988 8956
rect 16807 8925 16819 8928
rect 16761 8919 16819 8925
rect 18322 8916 18328 8968
rect 18380 8956 18386 8968
rect 19242 8956 19248 8968
rect 18380 8928 19248 8956
rect 18380 8916 18386 8928
rect 19242 8916 19248 8928
rect 19300 8956 19306 8968
rect 19705 8959 19763 8965
rect 19705 8956 19717 8959
rect 19300 8928 19717 8956
rect 19300 8916 19306 8928
rect 19705 8925 19717 8928
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 20530 8916 20536 8968
rect 20588 8956 20594 8968
rect 20898 8965 20904 8968
rect 20717 8959 20775 8965
rect 20717 8956 20729 8959
rect 20588 8928 20729 8956
rect 20588 8916 20594 8928
rect 20717 8925 20729 8928
rect 20763 8925 20775 8959
rect 20717 8919 20775 8925
rect 20865 8959 20904 8965
rect 20865 8925 20877 8959
rect 20865 8919 20904 8925
rect 20898 8916 20904 8919
rect 20956 8916 20962 8968
rect 20990 8916 20996 8968
rect 21048 8956 21054 8968
rect 21223 8959 21281 8965
rect 21048 8928 21093 8956
rect 21048 8916 21054 8928
rect 21223 8925 21235 8959
rect 21269 8956 21281 8959
rect 21818 8956 21824 8968
rect 21269 8928 21824 8956
rect 21269 8925 21281 8928
rect 21223 8919 21281 8925
rect 21818 8916 21824 8928
rect 21876 8916 21882 8968
rect 21928 8965 21956 9064
rect 23106 9052 23112 9104
rect 23164 9092 23170 9104
rect 23164 9064 23428 9092
rect 23164 9052 23170 9064
rect 22186 9024 22192 9036
rect 22021 8996 22192 9024
rect 22021 8965 22049 8996
rect 22186 8984 22192 8996
rect 22244 8984 22250 9036
rect 23400 9033 23428 9064
rect 23385 9027 23443 9033
rect 23385 8993 23397 9027
rect 23431 8993 23443 9027
rect 23385 8987 23443 8993
rect 24946 8984 24952 9036
rect 25004 9024 25010 9036
rect 25685 9027 25743 9033
rect 25685 9024 25697 9027
rect 25004 8996 25697 9024
rect 25004 8984 25010 8996
rect 25685 8993 25697 8996
rect 25731 8993 25743 9027
rect 25685 8987 25743 8993
rect 26789 9027 26847 9033
rect 26789 8993 26801 9027
rect 26835 9024 26847 9027
rect 27338 9024 27344 9036
rect 26835 8996 27344 9024
rect 26835 8993 26847 8996
rect 26789 8987 26847 8993
rect 27338 8984 27344 8996
rect 27396 8984 27402 9036
rect 27617 9027 27675 9033
rect 27617 8993 27629 9027
rect 27663 9024 27675 9027
rect 27982 9024 27988 9036
rect 27663 8996 27988 9024
rect 27663 8993 27675 8996
rect 27617 8987 27675 8993
rect 27982 8984 27988 8996
rect 28040 9024 28046 9036
rect 28626 9024 28632 9036
rect 28040 8996 28632 9024
rect 28040 8984 28046 8996
rect 28626 8984 28632 8996
rect 28684 8984 28690 9036
rect 21913 8959 21971 8965
rect 21913 8925 21925 8959
rect 21959 8925 21971 8959
rect 21913 8919 21971 8925
rect 22006 8959 22064 8965
rect 22006 8925 22018 8959
rect 22052 8925 22064 8959
rect 22378 8959 22436 8965
rect 22378 8956 22390 8959
rect 22006 8919 22064 8925
rect 22112 8928 22390 8956
rect 14844 8860 15608 8888
rect 12805 8851 12863 8857
rect 15580 8832 15608 8860
rect 19886 8848 19892 8900
rect 19944 8888 19950 8900
rect 20622 8888 20628 8900
rect 19944 8860 20628 8888
rect 19944 8848 19950 8860
rect 20622 8848 20628 8860
rect 20680 8888 20686 8900
rect 21085 8891 21143 8897
rect 21085 8888 21097 8891
rect 20680 8860 21097 8888
rect 20680 8848 20686 8860
rect 21085 8857 21097 8860
rect 21131 8857 21143 8891
rect 21836 8888 21864 8916
rect 22112 8888 22140 8928
rect 22378 8925 22390 8928
rect 22424 8925 22436 8959
rect 22378 8919 22436 8925
rect 23109 8959 23167 8965
rect 23109 8925 23121 8959
rect 23155 8956 23167 8959
rect 23198 8956 23204 8968
rect 23155 8928 23204 8956
rect 23155 8925 23167 8928
rect 23109 8919 23167 8925
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 23293 8959 23351 8965
rect 23293 8925 23305 8959
rect 23339 8925 23351 8959
rect 23474 8956 23480 8968
rect 23435 8928 23480 8956
rect 23293 8919 23351 8925
rect 21836 8860 22140 8888
rect 22189 8891 22247 8897
rect 21085 8851 21143 8857
rect 22189 8857 22201 8891
rect 22235 8857 22247 8891
rect 22189 8851 22247 8857
rect 22281 8891 22339 8897
rect 22281 8857 22293 8891
rect 22327 8888 22339 8891
rect 22554 8888 22560 8900
rect 22327 8860 22560 8888
rect 22327 8857 22339 8860
rect 22281 8851 22339 8857
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 11333 8823 11391 8829
rect 11333 8820 11345 8823
rect 10836 8792 11345 8820
rect 10836 8780 10842 8792
rect 11333 8789 11345 8792
rect 11379 8789 11391 8823
rect 11333 8783 11391 8789
rect 11422 8780 11428 8832
rect 11480 8820 11486 8832
rect 14550 8820 14556 8832
rect 11480 8792 11525 8820
rect 14511 8792 14556 8820
rect 11480 8780 11486 8792
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 14645 8823 14703 8829
rect 14645 8789 14657 8823
rect 14691 8820 14703 8823
rect 15470 8820 15476 8832
rect 14691 8792 15476 8820
rect 14691 8789 14703 8792
rect 14645 8783 14703 8789
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 15562 8780 15568 8832
rect 15620 8780 15626 8832
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 22204 8820 22232 8851
rect 22554 8848 22560 8860
rect 22612 8888 22618 8900
rect 22738 8888 22744 8900
rect 22612 8860 22744 8888
rect 22612 8848 22618 8860
rect 22738 8848 22744 8860
rect 22796 8888 22802 8900
rect 23308 8888 23336 8919
rect 23474 8916 23480 8928
rect 23532 8916 23538 8968
rect 23661 8959 23719 8965
rect 23661 8925 23673 8959
rect 23707 8956 23719 8959
rect 25314 8956 25320 8968
rect 23707 8928 25320 8956
rect 23707 8925 23719 8928
rect 23661 8919 23719 8925
rect 25314 8916 25320 8928
rect 25372 8916 25378 8968
rect 25409 8959 25467 8965
rect 25409 8925 25421 8959
rect 25455 8956 25467 8959
rect 26142 8956 26148 8968
rect 25455 8928 26148 8956
rect 25455 8925 25467 8928
rect 25409 8919 25467 8925
rect 26142 8916 26148 8928
rect 26200 8916 26206 8968
rect 26697 8959 26755 8965
rect 26697 8925 26709 8959
rect 26743 8956 26755 8959
rect 26970 8956 26976 8968
rect 26743 8928 26976 8956
rect 26743 8925 26755 8928
rect 26697 8919 26755 8925
rect 26970 8916 26976 8928
rect 27028 8916 27034 8968
rect 28810 8956 28816 8968
rect 28771 8928 28816 8956
rect 28810 8916 28816 8928
rect 28868 8916 28874 8968
rect 30098 8956 30104 8968
rect 30059 8928 30104 8956
rect 30098 8916 30104 8928
rect 30156 8916 30162 8968
rect 22796 8860 23336 8888
rect 22796 8848 22802 8860
rect 24118 8848 24124 8900
rect 24176 8888 24182 8900
rect 25130 8888 25136 8900
rect 24176 8860 25136 8888
rect 24176 8848 24182 8860
rect 25130 8848 25136 8860
rect 25188 8848 25194 8900
rect 22370 8820 22376 8832
rect 20772 8792 22376 8820
rect 20772 8780 20778 8792
rect 22370 8780 22376 8792
rect 22428 8780 22434 8832
rect 23845 8823 23903 8829
rect 23845 8789 23857 8823
rect 23891 8820 23903 8823
rect 24210 8820 24216 8832
rect 23891 8792 24216 8820
rect 23891 8789 23903 8792
rect 23845 8783 23903 8789
rect 24210 8780 24216 8792
rect 24268 8780 24274 8832
rect 28810 8780 28816 8832
rect 28868 8820 28874 8832
rect 29917 8823 29975 8829
rect 29917 8820 29929 8823
rect 28868 8792 29929 8820
rect 28868 8780 28874 8792
rect 29917 8789 29929 8792
rect 29963 8789 29975 8823
rect 29917 8783 29975 8789
rect 1104 8730 30820 8752
rect 1104 8678 10880 8730
rect 10932 8678 10944 8730
rect 10996 8678 11008 8730
rect 11060 8678 11072 8730
rect 11124 8678 11136 8730
rect 11188 8678 20811 8730
rect 20863 8678 20875 8730
rect 20927 8678 20939 8730
rect 20991 8678 21003 8730
rect 21055 8678 21067 8730
rect 21119 8678 30820 8730
rect 1104 8656 30820 8678
rect 10778 8616 10784 8628
rect 10739 8588 10784 8616
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 13817 8619 13875 8625
rect 13817 8585 13829 8619
rect 13863 8616 13875 8619
rect 14550 8616 14556 8628
rect 13863 8588 14556 8616
rect 13863 8585 13875 8588
rect 13817 8579 13875 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 15381 8619 15439 8625
rect 15381 8585 15393 8619
rect 15427 8616 15439 8619
rect 16390 8616 16396 8628
rect 15427 8588 16396 8616
rect 15427 8585 15439 8588
rect 15381 8579 15439 8585
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 18782 8576 18788 8628
rect 18840 8616 18846 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 18840 8588 19441 8616
rect 18840 8576 18846 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 19429 8579 19487 8585
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 20128 8588 20545 8616
rect 20128 8576 20134 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 20533 8579 20591 8585
rect 23569 8619 23627 8625
rect 23569 8585 23581 8619
rect 23615 8616 23627 8619
rect 24118 8616 24124 8628
rect 23615 8588 24124 8616
rect 23615 8585 23627 8588
rect 23569 8579 23627 8585
rect 24118 8576 24124 8588
rect 24176 8576 24182 8628
rect 29914 8576 29920 8628
rect 29972 8616 29978 8628
rect 30101 8619 30159 8625
rect 30101 8616 30113 8619
rect 29972 8588 30113 8616
rect 29972 8576 29978 8588
rect 30101 8585 30113 8588
rect 30147 8585 30159 8619
rect 30101 8579 30159 8585
rect 11698 8548 11704 8560
rect 11659 8520 11704 8548
rect 11698 8508 11704 8520
rect 11756 8508 11762 8560
rect 14829 8551 14887 8557
rect 14829 8548 14841 8551
rect 14016 8520 14841 8548
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 10980 8412 11008 8443
rect 11422 8440 11428 8492
rect 11480 8480 11486 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11480 8452 11529 8480
rect 11480 8440 11486 8452
rect 11517 8449 11529 8452
rect 11563 8480 11575 8483
rect 11974 8480 11980 8492
rect 11563 8452 11980 8480
rect 11563 8449 11575 8452
rect 11517 8443 11575 8449
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 12526 8480 12532 8492
rect 12487 8452 12532 8480
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 14016 8489 14044 8520
rect 14829 8517 14841 8520
rect 14875 8517 14887 8551
rect 16853 8551 16911 8557
rect 16853 8548 16865 8551
rect 14829 8511 14887 8517
rect 14936 8520 16865 8548
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 11885 8415 11943 8421
rect 11885 8412 11897 8415
rect 10980 8384 11897 8412
rect 11885 8381 11897 8384
rect 11931 8381 11943 8415
rect 14476 8412 14504 8443
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 14936 8480 14964 8520
rect 16853 8517 16865 8520
rect 16899 8517 16911 8551
rect 16853 8511 16911 8517
rect 18316 8551 18374 8557
rect 18316 8517 18328 8551
rect 18362 8548 18374 8551
rect 19150 8548 19156 8560
rect 18362 8520 19156 8548
rect 18362 8517 18374 8520
rect 18316 8511 18374 8517
rect 19150 8508 19156 8520
rect 19208 8508 19214 8560
rect 19242 8508 19248 8560
rect 19300 8548 19306 8560
rect 20441 8551 20499 8557
rect 20441 8548 20453 8551
rect 19300 8520 20453 8548
rect 19300 8508 19306 8520
rect 20441 8517 20453 8520
rect 20487 8517 20499 8551
rect 20441 8511 20499 8517
rect 22094 8508 22100 8560
rect 22152 8548 22158 8560
rect 22152 8520 22197 8548
rect 22152 8508 22158 8520
rect 22462 8508 22468 8560
rect 22520 8548 22526 8560
rect 22520 8520 23060 8548
rect 22520 8508 22526 8520
rect 23032 8492 23060 8520
rect 24210 8508 24216 8560
rect 24268 8557 24274 8560
rect 24268 8551 24332 8557
rect 24268 8517 24286 8551
rect 24320 8517 24332 8551
rect 27154 8548 27160 8560
rect 24268 8511 24332 8517
rect 25792 8520 27160 8548
rect 24268 8508 24274 8511
rect 15746 8480 15752 8492
rect 14700 8452 14964 8480
rect 15707 8452 15752 8480
rect 14700 8440 14706 8452
rect 15746 8440 15752 8452
rect 15804 8440 15810 8492
rect 15841 8483 15899 8489
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 15887 8452 16681 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 16669 8449 16681 8452
rect 16715 8480 16727 8483
rect 16758 8480 16764 8492
rect 16715 8452 16764 8480
rect 16715 8449 16727 8452
rect 16669 8443 16727 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 21910 8480 21916 8492
rect 21871 8452 21916 8480
rect 21910 8440 21916 8452
rect 21968 8440 21974 8492
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8449 22891 8483
rect 23014 8480 23020 8492
rect 22975 8452 23020 8480
rect 22833 8443 22891 8449
rect 15470 8412 15476 8424
rect 14476 8384 15476 8412
rect 11885 8375 11943 8381
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 15562 8372 15568 8424
rect 15620 8412 15626 8424
rect 15933 8415 15991 8421
rect 15933 8412 15945 8415
rect 15620 8384 15945 8412
rect 15620 8372 15626 8384
rect 15933 8381 15945 8384
rect 15979 8381 15991 8415
rect 18046 8412 18052 8424
rect 15933 8375 15991 8381
rect 16684 8384 18052 8412
rect 16684 8356 16712 8384
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 20622 8372 20628 8424
rect 20680 8412 20686 8424
rect 22462 8412 22468 8424
rect 20680 8384 22468 8412
rect 20680 8372 20686 8384
rect 22462 8372 22468 8384
rect 22520 8372 22526 8424
rect 12345 8347 12403 8353
rect 12345 8313 12357 8347
rect 12391 8344 12403 8347
rect 12434 8344 12440 8356
rect 12391 8316 12440 8344
rect 12391 8313 12403 8316
rect 12345 8307 12403 8313
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 16666 8304 16672 8356
rect 16724 8304 16730 8356
rect 22848 8344 22876 8443
rect 23014 8440 23020 8452
rect 23072 8440 23078 8492
rect 23106 8440 23112 8492
rect 23164 8480 23170 8492
rect 23385 8483 23443 8489
rect 23164 8452 23209 8480
rect 23164 8440 23170 8452
rect 23385 8449 23397 8483
rect 23431 8480 23443 8483
rect 23431 8452 23888 8480
rect 23431 8449 23443 8452
rect 23385 8443 23443 8449
rect 23201 8415 23259 8421
rect 23201 8381 23213 8415
rect 23247 8412 23259 8415
rect 23474 8412 23480 8424
rect 23247 8384 23480 8412
rect 23247 8381 23259 8384
rect 23201 8375 23259 8381
rect 23474 8372 23480 8384
rect 23532 8412 23538 8424
rect 23750 8412 23756 8424
rect 23532 8384 23756 8412
rect 23532 8372 23538 8384
rect 23750 8372 23756 8384
rect 23808 8372 23814 8424
rect 23860 8412 23888 8452
rect 23934 8440 23940 8492
rect 23992 8480 23998 8492
rect 24029 8483 24087 8489
rect 24029 8480 24041 8483
rect 23992 8452 24041 8480
rect 23992 8440 23998 8452
rect 24029 8449 24041 8452
rect 24075 8449 24087 8483
rect 25792 8480 25820 8520
rect 27154 8508 27160 8520
rect 27212 8508 27218 8560
rect 24029 8443 24087 8449
rect 24136 8452 25820 8480
rect 24136 8412 24164 8452
rect 26142 8440 26148 8492
rect 26200 8480 26206 8492
rect 28994 8489 29000 8492
rect 27249 8483 27307 8489
rect 27249 8480 27261 8483
rect 26200 8452 27261 8480
rect 26200 8440 26206 8452
rect 27249 8449 27261 8452
rect 27295 8449 27307 8483
rect 27249 8443 27307 8449
rect 28988 8443 29000 8489
rect 29052 8480 29058 8492
rect 29052 8452 29088 8480
rect 28994 8440 29000 8443
rect 29052 8440 29058 8452
rect 23860 8384 24164 8412
rect 26234 8372 26240 8424
rect 26292 8412 26298 8424
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26292 8384 26985 8412
rect 26292 8372 26298 8384
rect 26973 8381 26985 8384
rect 27019 8412 27031 8415
rect 27338 8412 27344 8424
rect 27019 8384 27344 8412
rect 27019 8381 27031 8384
rect 26973 8375 27031 8381
rect 27338 8372 27344 8384
rect 27396 8372 27402 8424
rect 27706 8372 27712 8424
rect 27764 8412 27770 8424
rect 28718 8412 28724 8424
rect 27764 8384 28724 8412
rect 27764 8372 27770 8384
rect 28718 8372 28724 8384
rect 28776 8372 28782 8424
rect 22848 8316 24072 8344
rect 17034 8276 17040 8288
rect 16995 8248 17040 8276
rect 17034 8236 17040 8248
rect 17092 8236 17098 8288
rect 17954 8236 17960 8288
rect 18012 8276 18018 8288
rect 18230 8276 18236 8288
rect 18012 8248 18236 8276
rect 18012 8236 18018 8248
rect 18230 8236 18236 8248
rect 18288 8236 18294 8288
rect 24044 8276 24072 8316
rect 25314 8304 25320 8356
rect 25372 8344 25378 8356
rect 25409 8347 25467 8353
rect 25409 8344 25421 8347
rect 25372 8316 25421 8344
rect 25372 8304 25378 8316
rect 25409 8313 25421 8316
rect 25455 8313 25467 8347
rect 25409 8307 25467 8313
rect 24946 8276 24952 8288
rect 24044 8248 24952 8276
rect 24946 8236 24952 8248
rect 25004 8236 25010 8288
rect 1104 8186 30820 8208
rect 1104 8134 5915 8186
rect 5967 8134 5979 8186
rect 6031 8134 6043 8186
rect 6095 8134 6107 8186
rect 6159 8134 6171 8186
rect 6223 8134 15846 8186
rect 15898 8134 15910 8186
rect 15962 8134 15974 8186
rect 16026 8134 16038 8186
rect 16090 8134 16102 8186
rect 16154 8134 25776 8186
rect 25828 8134 25840 8186
rect 25892 8134 25904 8186
rect 25956 8134 25968 8186
rect 26020 8134 26032 8186
rect 26084 8134 30820 8186
rect 1104 8112 30820 8134
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 12584 8044 12633 8072
rect 12584 8032 12590 8044
rect 12621 8041 12633 8044
rect 12667 8041 12679 8075
rect 12621 8035 12679 8041
rect 15746 8032 15752 8084
rect 15804 8072 15810 8084
rect 16025 8075 16083 8081
rect 16025 8072 16037 8075
rect 15804 8044 16037 8072
rect 15804 8032 15810 8044
rect 16025 8041 16037 8044
rect 16071 8041 16083 8075
rect 17954 8072 17960 8084
rect 16025 8035 16083 8041
rect 17420 8044 17960 8072
rect 12894 7936 12900 7948
rect 12268 7908 12900 7936
rect 12268 7877 12296 7908
rect 12894 7896 12900 7908
rect 12952 7896 12958 7948
rect 17420 7936 17448 8044
rect 17954 8032 17960 8044
rect 18012 8032 18018 8084
rect 18046 8032 18052 8084
rect 18104 8072 18110 8084
rect 18598 8072 18604 8084
rect 18104 8044 18604 8072
rect 18104 8032 18110 8044
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 19426 8032 19432 8084
rect 19484 8072 19490 8084
rect 19613 8075 19671 8081
rect 19613 8072 19625 8075
rect 19484 8044 19625 8072
rect 19484 8032 19490 8044
rect 19613 8041 19625 8044
rect 19659 8041 19671 8075
rect 19613 8035 19671 8041
rect 19886 8032 19892 8084
rect 19944 8072 19950 8084
rect 20162 8072 20168 8084
rect 19944 8044 20168 8072
rect 19944 8032 19950 8044
rect 20162 8032 20168 8044
rect 20220 8072 20226 8084
rect 20257 8075 20315 8081
rect 20257 8072 20269 8075
rect 20220 8044 20269 8072
rect 20220 8032 20226 8044
rect 20257 8041 20269 8044
rect 20303 8041 20315 8075
rect 21266 8072 21272 8084
rect 20257 8035 20315 8041
rect 21100 8044 21272 8072
rect 19518 8004 19524 8016
rect 17328 7908 17448 7936
rect 17696 7976 19524 8004
rect 17328 7880 17356 7908
rect 12253 7871 12311 7877
rect 12253 7837 12265 7871
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 12526 7828 12532 7880
rect 12584 7868 12590 7880
rect 13081 7871 13139 7877
rect 13081 7868 13093 7871
rect 12584 7840 13093 7868
rect 12584 7828 12590 7840
rect 13081 7837 13093 7840
rect 13127 7837 13139 7871
rect 14274 7868 14280 7880
rect 14235 7840 14280 7868
rect 13081 7831 13139 7837
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 16209 7871 16267 7877
rect 16209 7837 16221 7871
rect 16255 7868 16267 7871
rect 17034 7868 17040 7880
rect 16255 7840 17040 7868
rect 16255 7837 16267 7840
rect 16209 7831 16267 7837
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 17310 7868 17316 7880
rect 17223 7840 17316 7868
rect 17310 7828 17316 7840
rect 17368 7828 17374 7880
rect 17494 7877 17500 7880
rect 17461 7871 17500 7877
rect 17461 7837 17473 7871
rect 17461 7831 17500 7837
rect 17494 7828 17500 7831
rect 17552 7828 17558 7880
rect 17696 7877 17724 7976
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 19886 7936 19892 7948
rect 19444 7908 19892 7936
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7837 17739 7871
rect 17681 7831 17739 7837
rect 17819 7871 17877 7877
rect 17819 7837 17831 7871
rect 17865 7868 17877 7871
rect 18414 7868 18420 7880
rect 17865 7840 18420 7868
rect 17865 7837 17877 7840
rect 17819 7831 17877 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 19444 7877 19472 7908
rect 19886 7896 19892 7908
rect 19944 7896 19950 7948
rect 21100 7945 21128 8044
rect 21266 8032 21272 8044
rect 21324 8072 21330 8084
rect 21324 8044 22416 8072
rect 21324 8032 21330 8044
rect 22278 8004 22284 8016
rect 22066 7976 22284 8004
rect 21085 7939 21143 7945
rect 21085 7905 21097 7939
rect 21131 7905 21143 7939
rect 21085 7899 21143 7905
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 19702 7828 19708 7880
rect 19760 7868 19766 7880
rect 19760 7840 19805 7868
rect 19760 7828 19766 7840
rect 20070 7828 20076 7880
rect 20128 7868 20134 7880
rect 20165 7871 20223 7877
rect 20165 7868 20177 7871
rect 20128 7840 20177 7868
rect 20128 7828 20134 7840
rect 20165 7837 20177 7840
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 22066 7877 22094 7976
rect 22278 7964 22284 7976
rect 22336 7964 22342 8016
rect 22388 7936 22416 8044
rect 23290 8032 23296 8084
rect 23348 8072 23354 8084
rect 23477 8075 23535 8081
rect 23477 8072 23489 8075
rect 23348 8044 23489 8072
rect 23348 8032 23354 8044
rect 23477 8041 23489 8044
rect 23523 8041 23535 8075
rect 23477 8035 23535 8041
rect 24302 8032 24308 8084
rect 24360 8072 24366 8084
rect 24489 8075 24547 8081
rect 24489 8072 24501 8075
rect 24360 8044 24501 8072
rect 24360 8032 24366 8044
rect 24489 8041 24501 8044
rect 24535 8041 24547 8075
rect 24489 8035 24547 8041
rect 26697 8075 26755 8081
rect 26697 8041 26709 8075
rect 26743 8072 26755 8075
rect 27154 8072 27160 8084
rect 26743 8044 27160 8072
rect 26743 8041 26755 8044
rect 26697 8035 26755 8041
rect 27154 8032 27160 8044
rect 27212 8032 27218 8084
rect 27522 8032 27528 8084
rect 27580 8072 27586 8084
rect 28353 8075 28411 8081
rect 28353 8072 28365 8075
rect 27580 8044 28365 8072
rect 27580 8032 27586 8044
rect 28353 8041 28365 8044
rect 28399 8041 28411 8075
rect 28353 8035 28411 8041
rect 23934 7964 23940 8016
rect 23992 8004 23998 8016
rect 23992 7976 25360 8004
rect 23992 7964 23998 7976
rect 22830 7936 22836 7948
rect 22388 7908 22836 7936
rect 20809 7871 20867 7877
rect 20809 7868 20821 7871
rect 20772 7840 20821 7868
rect 20772 7828 20778 7840
rect 20809 7837 20821 7840
rect 20855 7837 20867 7871
rect 22066 7871 22144 7877
rect 22066 7842 22098 7871
rect 20809 7831 20867 7837
rect 22086 7837 22098 7842
rect 22132 7837 22144 7871
rect 22086 7831 22144 7837
rect 22245 7871 22303 7877
rect 22245 7837 22257 7871
rect 22291 7868 22303 7871
rect 22388 7868 22416 7908
rect 22830 7896 22836 7908
rect 22888 7896 22894 7948
rect 25332 7945 25360 7976
rect 27614 7964 27620 8016
rect 27672 8004 27678 8016
rect 28718 8004 28724 8016
rect 27672 7976 28724 8004
rect 27672 7964 27678 7976
rect 28718 7964 28724 7976
rect 28776 7964 28782 8016
rect 25317 7939 25375 7945
rect 25317 7905 25329 7939
rect 25363 7905 25375 7939
rect 28902 7936 28908 7948
rect 25317 7899 25375 7905
rect 27816 7908 28908 7936
rect 22291 7840 22416 7868
rect 22603 7871 22661 7877
rect 22291 7837 22303 7840
rect 22245 7831 22303 7837
rect 22603 7837 22615 7871
rect 22649 7868 22661 7871
rect 23198 7868 23204 7880
rect 22649 7840 23204 7868
rect 22649 7837 22661 7840
rect 22603 7831 22661 7837
rect 23198 7828 23204 7840
rect 23256 7828 23262 7880
rect 23385 7871 23443 7877
rect 23385 7837 23397 7871
rect 23431 7868 23443 7871
rect 23566 7868 23572 7880
rect 23431 7840 23572 7868
rect 23431 7837 23443 7840
rect 23385 7831 23443 7837
rect 23566 7828 23572 7840
rect 23624 7828 23630 7880
rect 24302 7828 24308 7880
rect 24360 7868 24366 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 24360 7840 24409 7868
rect 24360 7828 24366 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 25130 7828 25136 7880
rect 25188 7868 25194 7880
rect 25573 7871 25631 7877
rect 25573 7868 25585 7871
rect 25188 7840 25585 7868
rect 25188 7828 25194 7840
rect 25573 7837 25585 7840
rect 25619 7837 25631 7871
rect 27614 7868 27620 7880
rect 27575 7840 27620 7868
rect 25573 7831 25631 7837
rect 27614 7828 27620 7840
rect 27672 7828 27678 7880
rect 27816 7877 27844 7908
rect 28902 7896 28908 7908
rect 28960 7896 28966 7948
rect 27801 7871 27859 7877
rect 27801 7837 27813 7871
rect 27847 7837 27859 7871
rect 27801 7831 27859 7837
rect 27893 7871 27951 7877
rect 27893 7837 27905 7871
rect 27939 7837 27951 7871
rect 27893 7831 27951 7837
rect 12437 7803 12495 7809
rect 12437 7769 12449 7803
rect 12483 7800 12495 7803
rect 12802 7800 12808 7812
rect 12483 7772 12808 7800
rect 12483 7769 12495 7772
rect 12437 7763 12495 7769
rect 12802 7760 12808 7772
rect 12860 7800 12866 7812
rect 13630 7800 13636 7812
rect 12860 7772 13636 7800
rect 12860 7760 12866 7772
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 17589 7803 17647 7809
rect 17589 7769 17601 7803
rect 17635 7769 17647 7803
rect 17589 7763 17647 7769
rect 18509 7803 18567 7809
rect 18509 7769 18521 7803
rect 18555 7800 18567 7803
rect 21910 7800 21916 7812
rect 18555 7772 21916 7800
rect 18555 7769 18567 7772
rect 18509 7763 18567 7769
rect 12342 7692 12348 7744
rect 12400 7732 12406 7744
rect 13265 7735 13323 7741
rect 13265 7732 13277 7735
rect 12400 7704 13277 7732
rect 12400 7692 12406 7704
rect 13265 7701 13277 7704
rect 13311 7701 13323 7735
rect 13265 7695 13323 7701
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 14277 7735 14335 7741
rect 14277 7732 14289 7735
rect 13412 7704 14289 7732
rect 13412 7692 13418 7704
rect 14277 7701 14289 7704
rect 14323 7701 14335 7735
rect 17604 7732 17632 7763
rect 21910 7760 21916 7772
rect 21968 7760 21974 7812
rect 22370 7800 22376 7812
rect 22066 7772 22376 7800
rect 17678 7732 17684 7744
rect 17604 7704 17684 7732
rect 14277 7695 14335 7701
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 17954 7732 17960 7744
rect 17915 7704 17960 7732
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 19245 7735 19303 7741
rect 19245 7732 19257 7735
rect 18104 7704 19257 7732
rect 18104 7692 18110 7704
rect 19245 7701 19257 7704
rect 19291 7701 19303 7735
rect 19245 7695 19303 7701
rect 19426 7692 19432 7744
rect 19484 7732 19490 7744
rect 22066 7732 22094 7772
rect 22370 7760 22376 7772
rect 22428 7760 22434 7812
rect 22462 7760 22468 7812
rect 22520 7800 22526 7812
rect 23474 7800 23480 7812
rect 22520 7772 23480 7800
rect 22520 7760 22526 7772
rect 23474 7760 23480 7772
rect 23532 7760 23538 7812
rect 27908 7800 27936 7831
rect 27982 7828 27988 7880
rect 28040 7868 28046 7880
rect 28169 7871 28227 7877
rect 28040 7840 28085 7868
rect 28040 7828 28046 7840
rect 28169 7837 28181 7871
rect 28215 7868 28227 7871
rect 28534 7868 28540 7880
rect 28215 7840 28540 7868
rect 28215 7837 28227 7840
rect 28169 7831 28227 7837
rect 28534 7828 28540 7840
rect 28592 7828 28598 7880
rect 30098 7868 30104 7880
rect 30059 7840 30104 7868
rect 30098 7828 30104 7840
rect 30156 7828 30162 7880
rect 28074 7800 28080 7812
rect 27908 7772 28080 7800
rect 28074 7760 28080 7772
rect 28132 7760 28138 7812
rect 19484 7704 22094 7732
rect 19484 7692 19490 7704
rect 22278 7692 22284 7744
rect 22336 7732 22342 7744
rect 22741 7735 22799 7741
rect 22741 7732 22753 7735
rect 22336 7704 22753 7732
rect 22336 7692 22342 7704
rect 22741 7701 22753 7704
rect 22787 7701 22799 7735
rect 22741 7695 22799 7701
rect 27614 7692 27620 7744
rect 27672 7732 27678 7744
rect 29917 7735 29975 7741
rect 29917 7732 29929 7735
rect 27672 7704 29929 7732
rect 27672 7692 27678 7704
rect 29917 7701 29929 7704
rect 29963 7701 29975 7735
rect 29917 7695 29975 7701
rect 1104 7642 30820 7664
rect 1104 7590 10880 7642
rect 10932 7590 10944 7642
rect 10996 7590 11008 7642
rect 11060 7590 11072 7642
rect 11124 7590 11136 7642
rect 11188 7590 20811 7642
rect 20863 7590 20875 7642
rect 20927 7590 20939 7642
rect 20991 7590 21003 7642
rect 21055 7590 21067 7642
rect 21119 7590 30820 7642
rect 1104 7568 30820 7590
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 14274 7528 14280 7540
rect 13412 7500 14280 7528
rect 13412 7488 13418 7500
rect 14274 7488 14280 7500
rect 14332 7528 14338 7540
rect 14645 7531 14703 7537
rect 14645 7528 14657 7531
rect 14332 7500 14657 7528
rect 14332 7488 14338 7500
rect 14645 7497 14657 7500
rect 14691 7497 14703 7531
rect 14645 7491 14703 7497
rect 19518 7488 19524 7540
rect 19576 7528 19582 7540
rect 23014 7528 23020 7540
rect 19576 7500 23020 7528
rect 19576 7488 19582 7500
rect 23014 7488 23020 7500
rect 23072 7528 23078 7540
rect 24121 7531 24179 7537
rect 24121 7528 24133 7531
rect 23072 7500 24133 7528
rect 23072 7488 23078 7500
rect 24121 7497 24133 7500
rect 24167 7528 24179 7531
rect 24302 7528 24308 7540
rect 24167 7500 24308 7528
rect 24167 7497 24179 7500
rect 24121 7491 24179 7497
rect 24302 7488 24308 7500
rect 24360 7488 24366 7540
rect 27890 7488 27896 7540
rect 27948 7528 27954 7540
rect 28353 7531 28411 7537
rect 28353 7528 28365 7531
rect 27948 7500 28365 7528
rect 27948 7488 27954 7500
rect 28353 7497 28365 7500
rect 28399 7497 28411 7531
rect 29546 7528 29552 7540
rect 29507 7500 29552 7528
rect 28353 7491 28411 7497
rect 29546 7488 29552 7500
rect 29604 7488 29610 7540
rect 14090 7420 14096 7472
rect 14148 7460 14154 7472
rect 14185 7463 14243 7469
rect 14185 7460 14197 7463
rect 14148 7432 14197 7460
rect 14148 7420 14154 7432
rect 14185 7429 14197 7432
rect 14231 7429 14243 7463
rect 14185 7423 14243 7429
rect 17028 7463 17086 7469
rect 17028 7429 17040 7463
rect 17074 7460 17086 7463
rect 17954 7460 17960 7472
rect 17074 7432 17960 7460
rect 17074 7429 17086 7432
rect 17028 7423 17086 7429
rect 17954 7420 17960 7432
rect 18012 7420 18018 7472
rect 20162 7420 20168 7472
rect 20220 7460 20226 7472
rect 21542 7460 21548 7472
rect 20220 7432 21548 7460
rect 20220 7420 20226 7432
rect 21542 7420 21548 7432
rect 21600 7420 21606 7472
rect 22922 7460 22928 7472
rect 21836 7432 22928 7460
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7392 1455 7395
rect 1854 7392 1860 7404
rect 1443 7364 1860 7392
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 1854 7352 1860 7364
rect 1912 7352 1918 7404
rect 12342 7392 12348 7404
rect 12303 7364 12348 7392
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 12529 7395 12587 7401
rect 12529 7392 12541 7395
rect 12492 7364 12541 7392
rect 12492 7352 12498 7364
rect 12529 7361 12541 7364
rect 12575 7361 12587 7395
rect 12529 7355 12587 7361
rect 13262 7352 13268 7404
rect 13320 7392 13326 7404
rect 14826 7392 14832 7404
rect 13320 7364 13365 7392
rect 14787 7364 14832 7392
rect 13320 7352 13326 7364
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 16666 7352 16672 7404
rect 16724 7392 16730 7404
rect 16761 7395 16819 7401
rect 16761 7392 16773 7395
rect 16724 7364 16773 7392
rect 16724 7352 16730 7364
rect 16761 7361 16773 7364
rect 16807 7361 16819 7395
rect 16761 7355 16819 7361
rect 18598 7352 18604 7404
rect 18656 7392 18662 7404
rect 19337 7395 19395 7401
rect 19337 7392 19349 7395
rect 18656 7364 19349 7392
rect 18656 7352 18662 7364
rect 19337 7361 19349 7364
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 19604 7395 19662 7401
rect 19604 7361 19616 7395
rect 19650 7392 19662 7395
rect 20438 7392 20444 7404
rect 19650 7364 20444 7392
rect 19650 7361 19662 7364
rect 19604 7355 19662 7361
rect 20438 7352 20444 7364
rect 20496 7352 20502 7404
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 21836 7401 21864 7432
rect 22922 7420 22928 7432
rect 22980 7420 22986 7472
rect 23474 7420 23480 7472
rect 23532 7460 23538 7472
rect 24394 7460 24400 7472
rect 23532 7432 24400 7460
rect 23532 7420 23538 7432
rect 24394 7420 24400 7432
rect 24452 7460 24458 7472
rect 29086 7460 29092 7472
rect 24452 7432 29092 7460
rect 24452 7420 24458 7432
rect 29086 7420 29092 7432
rect 29144 7420 29150 7472
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 20772 7364 21833 7392
rect 20772 7352 20778 7364
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 22094 7352 22100 7404
rect 22152 7392 22158 7404
rect 22741 7395 22799 7401
rect 22741 7392 22753 7395
rect 22152 7364 22753 7392
rect 22152 7352 22158 7364
rect 22741 7361 22753 7364
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 23008 7395 23066 7401
rect 23008 7361 23020 7395
rect 23054 7392 23066 7395
rect 23382 7392 23388 7404
rect 23054 7364 23388 7392
rect 23054 7361 23066 7364
rect 23008 7355 23066 7361
rect 23382 7352 23388 7364
rect 23440 7352 23446 7404
rect 23750 7352 23756 7404
rect 23808 7392 23814 7404
rect 27246 7401 27252 7404
rect 25317 7395 25375 7401
rect 25317 7392 25329 7395
rect 23808 7364 25329 7392
rect 23808 7352 23814 7364
rect 25317 7361 25329 7364
rect 25363 7361 25375 7395
rect 25317 7355 25375 7361
rect 27240 7355 27252 7401
rect 27304 7392 27310 7404
rect 27304 7364 27340 7392
rect 27246 7352 27252 7355
rect 27304 7352 27310 7364
rect 28350 7352 28356 7404
rect 28408 7392 28414 7404
rect 28718 7392 28724 7404
rect 28408 7364 28724 7392
rect 28408 7352 28414 7364
rect 28718 7352 28724 7364
rect 28776 7392 28782 7404
rect 28813 7395 28871 7401
rect 28813 7392 28825 7395
rect 28776 7364 28825 7392
rect 28776 7352 28782 7364
rect 28813 7361 28825 7364
rect 28859 7361 28871 7395
rect 28813 7355 28871 7361
rect 28997 7395 29055 7401
rect 28997 7361 29009 7395
rect 29043 7392 29055 7395
rect 29270 7392 29276 7404
rect 29043 7364 29276 7392
rect 29043 7361 29055 7364
rect 28997 7355 29055 7361
rect 29270 7352 29276 7364
rect 29328 7352 29334 7404
rect 29365 7395 29423 7401
rect 29365 7361 29377 7395
rect 29411 7392 29423 7395
rect 30006 7392 30012 7404
rect 29411 7364 30012 7392
rect 29411 7361 29423 7364
rect 29365 7355 29423 7361
rect 30006 7352 30012 7364
rect 30064 7352 30070 7404
rect 13354 7284 13360 7336
rect 13412 7333 13418 7336
rect 13412 7327 13440 7333
rect 13428 7293 13440 7327
rect 13412 7287 13440 7293
rect 13412 7284 13418 7287
rect 13538 7284 13544 7336
rect 13596 7324 13602 7336
rect 25041 7327 25099 7333
rect 13596 7296 13641 7324
rect 13596 7284 13602 7296
rect 25041 7293 25053 7327
rect 25087 7324 25099 7327
rect 26234 7324 26240 7336
rect 25087 7296 26240 7324
rect 25087 7293 25099 7296
rect 25041 7287 25099 7293
rect 26234 7284 26240 7296
rect 26292 7284 26298 7336
rect 26973 7327 27031 7333
rect 26973 7293 26985 7327
rect 27019 7293 27031 7327
rect 26973 7287 27031 7293
rect 12989 7259 13047 7265
rect 12989 7225 13001 7259
rect 13035 7225 13047 7259
rect 12989 7219 13047 7225
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 13004 7188 13032 7219
rect 15562 7188 15568 7200
rect 13004 7160 15568 7188
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 17678 7188 17684 7200
rect 16632 7160 17684 7188
rect 16632 7148 16638 7160
rect 17678 7148 17684 7160
rect 17736 7188 17742 7200
rect 18141 7191 18199 7197
rect 18141 7188 18153 7191
rect 17736 7160 18153 7188
rect 17736 7148 17742 7160
rect 18141 7157 18153 7160
rect 18187 7157 18199 7191
rect 18141 7151 18199 7157
rect 20070 7148 20076 7200
rect 20128 7188 20134 7200
rect 20717 7191 20775 7197
rect 20717 7188 20729 7191
rect 20128 7160 20729 7188
rect 20128 7148 20134 7160
rect 20717 7157 20729 7160
rect 20763 7157 20775 7191
rect 20717 7151 20775 7157
rect 20806 7148 20812 7200
rect 20864 7188 20870 7200
rect 21913 7191 21971 7197
rect 21913 7188 21925 7191
rect 20864 7160 21925 7188
rect 20864 7148 20870 7160
rect 21913 7157 21925 7160
rect 21959 7157 21971 7191
rect 26988 7188 27016 7287
rect 28074 7284 28080 7336
rect 28132 7324 28138 7336
rect 28626 7324 28632 7336
rect 28132 7296 28632 7324
rect 28132 7284 28138 7296
rect 28626 7284 28632 7296
rect 28684 7324 28690 7336
rect 29089 7327 29147 7333
rect 29089 7324 29101 7327
rect 28684 7296 29101 7324
rect 28684 7284 28690 7296
rect 29089 7293 29101 7296
rect 29135 7293 29147 7327
rect 29089 7287 29147 7293
rect 29181 7327 29239 7333
rect 29181 7293 29193 7327
rect 29227 7293 29239 7327
rect 29181 7287 29239 7293
rect 27982 7216 27988 7268
rect 28040 7256 28046 7268
rect 28718 7256 28724 7268
rect 28040 7228 28724 7256
rect 28040 7216 28046 7228
rect 28718 7216 28724 7228
rect 28776 7256 28782 7268
rect 29196 7256 29224 7287
rect 28776 7228 29224 7256
rect 28776 7216 28782 7228
rect 27706 7188 27712 7200
rect 26988 7160 27712 7188
rect 21913 7151 21971 7157
rect 27706 7148 27712 7160
rect 27764 7148 27770 7200
rect 1104 7098 30820 7120
rect 1104 7046 5915 7098
rect 5967 7046 5979 7098
rect 6031 7046 6043 7098
rect 6095 7046 6107 7098
rect 6159 7046 6171 7098
rect 6223 7046 15846 7098
rect 15898 7046 15910 7098
rect 15962 7046 15974 7098
rect 16026 7046 16038 7098
rect 16090 7046 16102 7098
rect 16154 7046 25776 7098
rect 25828 7046 25840 7098
rect 25892 7046 25904 7098
rect 25956 7046 25968 7098
rect 26020 7046 26032 7098
rect 26084 7046 30820 7098
rect 1104 7024 30820 7046
rect 12158 6984 12164 6996
rect 11256 6956 12164 6984
rect 11256 6925 11284 6956
rect 12158 6944 12164 6956
rect 12216 6984 12222 6996
rect 15470 6984 15476 6996
rect 12216 6956 13124 6984
rect 15431 6956 15476 6984
rect 12216 6944 12222 6956
rect 11241 6919 11299 6925
rect 11241 6885 11253 6919
rect 11287 6885 11299 6919
rect 11241 6879 11299 6885
rect 13096 6916 13124 6956
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 20254 6984 20260 6996
rect 16960 6956 20260 6984
rect 14734 6916 14740 6928
rect 13096 6888 14740 6916
rect 10594 6848 10600 6860
rect 10507 6820 10600 6848
rect 10594 6808 10600 6820
rect 10652 6848 10658 6860
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 10652 6820 11529 6848
rect 10652 6808 10658 6820
rect 11517 6817 11529 6820
rect 11563 6817 11575 6851
rect 11517 6811 11575 6817
rect 11793 6851 11851 6857
rect 11793 6817 11805 6851
rect 11839 6848 11851 6851
rect 12342 6848 12348 6860
rect 11839 6820 12348 6848
rect 11839 6817 11851 6820
rect 11793 6811 11851 6817
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 10778 6780 10784 6792
rect 10739 6752 10784 6780
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 11698 6789 11704 6792
rect 11655 6783 11704 6789
rect 11655 6749 11667 6783
rect 11701 6749 11704 6783
rect 11655 6743 11704 6749
rect 11698 6740 11704 6743
rect 11756 6740 11762 6792
rect 12894 6780 12900 6792
rect 12855 6752 12900 6780
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 13096 6789 13124 6888
rect 14734 6876 14740 6888
rect 14792 6916 14798 6928
rect 16850 6916 16856 6928
rect 14792 6888 16856 6916
rect 14792 6876 14798 6888
rect 16850 6876 16856 6888
rect 16908 6876 16914 6928
rect 13265 6851 13323 6857
rect 13265 6817 13277 6851
rect 13311 6848 13323 6851
rect 14826 6848 14832 6860
rect 13311 6820 14832 6848
rect 13311 6817 13323 6820
rect 13265 6811 13323 6817
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 16117 6851 16175 6857
rect 16117 6817 16129 6851
rect 16163 6848 16175 6851
rect 16574 6848 16580 6860
rect 16163 6820 16580 6848
rect 16163 6817 16175 6820
rect 16117 6811 16175 6817
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 13538 6740 13544 6792
rect 13596 6780 13602 6792
rect 16132 6780 16160 6811
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 16960 6848 16988 6956
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 20438 6984 20444 6996
rect 20399 6956 20444 6984
rect 20438 6944 20444 6956
rect 20496 6944 20502 6996
rect 22281 6987 22339 6993
rect 22281 6953 22293 6987
rect 22327 6984 22339 6987
rect 22370 6984 22376 6996
rect 22327 6956 22376 6984
rect 22327 6953 22339 6956
rect 22281 6947 22339 6953
rect 22370 6944 22376 6956
rect 22428 6944 22434 6996
rect 23382 6984 23388 6996
rect 23343 6956 23388 6984
rect 23382 6944 23388 6956
rect 23440 6944 23446 6996
rect 27157 6987 27215 6993
rect 27157 6953 27169 6987
rect 27203 6984 27215 6987
rect 27246 6984 27252 6996
rect 27203 6956 27252 6984
rect 27203 6953 27215 6956
rect 27157 6947 27215 6953
rect 27246 6944 27252 6956
rect 27304 6944 27310 6996
rect 27890 6984 27896 6996
rect 27632 6956 27896 6984
rect 18414 6916 18420 6928
rect 16684 6820 16988 6848
rect 17052 6888 18420 6916
rect 16684 6789 16712 6820
rect 13596 6752 16160 6780
rect 16669 6783 16727 6789
rect 13596 6740 13602 6752
rect 16669 6749 16681 6783
rect 16715 6749 16727 6783
rect 16669 6743 16727 6749
rect 16853 6783 16911 6789
rect 16853 6749 16865 6783
rect 16899 6749 16911 6783
rect 16853 6743 16911 6749
rect 16945 6783 17003 6789
rect 16945 6749 16957 6783
rect 16991 6780 17003 6783
rect 17052 6780 17080 6888
rect 18414 6876 18420 6888
rect 18472 6876 18478 6928
rect 20714 6916 20720 6928
rect 20548 6888 20720 6916
rect 17129 6851 17187 6857
rect 17129 6817 17141 6851
rect 17175 6848 17187 6851
rect 18046 6848 18052 6860
rect 17175 6820 18052 6848
rect 17175 6817 17187 6820
rect 17129 6811 17187 6817
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 18325 6851 18383 6857
rect 18325 6817 18337 6851
rect 18371 6817 18383 6851
rect 20548 6848 20576 6888
rect 20714 6876 20720 6888
rect 20772 6876 20778 6928
rect 20806 6848 20812 6860
rect 18325 6811 18383 6817
rect 20180 6820 20576 6848
rect 20640 6820 20812 6848
rect 16991 6752 17080 6780
rect 17221 6783 17279 6789
rect 16991 6749 17003 6752
rect 16945 6743 17003 6749
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 17494 6780 17500 6792
rect 17267 6752 17500 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 15746 6672 15752 6724
rect 15804 6712 15810 6724
rect 15933 6715 15991 6721
rect 15933 6712 15945 6715
rect 15804 6684 15945 6712
rect 15804 6672 15810 6684
rect 15933 6681 15945 6684
rect 15979 6681 15991 6715
rect 15933 6675 15991 6681
rect 16482 6672 16488 6724
rect 16540 6712 16546 6724
rect 16868 6712 16896 6743
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 17954 6780 17960 6792
rect 17915 6752 17960 6780
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 18141 6781 18199 6787
rect 18141 6747 18153 6781
rect 18187 6747 18199 6781
rect 18141 6741 18199 6747
rect 18236 6783 18294 6789
rect 18236 6749 18248 6783
rect 18282 6749 18294 6783
rect 18236 6743 18294 6749
rect 16540 6684 16896 6712
rect 17512 6712 17540 6740
rect 18156 6712 18184 6741
rect 17512 6684 18184 6712
rect 16540 6672 16546 6684
rect 18248 6656 18276 6743
rect 18340 6712 18368 6811
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 18874 6780 18880 6792
rect 18555 6752 18880 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 19797 6783 19855 6789
rect 19797 6749 19809 6783
rect 19843 6749 19855 6783
rect 19797 6743 19855 6749
rect 19945 6783 20003 6789
rect 19945 6749 19957 6783
rect 19991 6780 20003 6783
rect 20180 6780 20208 6820
rect 19991 6752 20208 6780
rect 20303 6783 20361 6789
rect 19991 6749 20003 6752
rect 19945 6743 20003 6749
rect 20303 6749 20315 6783
rect 20349 6780 20361 6783
rect 20438 6780 20444 6792
rect 20349 6752 20444 6780
rect 20349 6749 20361 6752
rect 20303 6743 20361 6749
rect 19334 6712 19340 6724
rect 18340 6684 19340 6712
rect 19334 6672 19340 6684
rect 19392 6672 19398 6724
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 15838 6644 15844 6656
rect 12492 6616 12537 6644
rect 15799 6616 15844 6644
rect 12492 6604 12498 6616
rect 15838 6604 15844 6616
rect 15896 6604 15902 6656
rect 16666 6644 16672 6656
rect 16627 6616 16672 6644
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 18230 6604 18236 6656
rect 18288 6604 18294 6656
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 18693 6647 18751 6653
rect 18693 6644 18705 6647
rect 18564 6616 18705 6644
rect 18564 6604 18570 6616
rect 18693 6613 18705 6616
rect 18739 6613 18751 6647
rect 19812 6644 19840 6743
rect 20438 6740 20444 6752
rect 20496 6780 20502 6792
rect 20640 6780 20668 6820
rect 20806 6808 20812 6820
rect 20864 6808 20870 6860
rect 25314 6808 25320 6860
rect 25372 6848 25378 6860
rect 25501 6851 25559 6857
rect 25501 6848 25513 6851
rect 25372 6820 25513 6848
rect 25372 6808 25378 6820
rect 25501 6817 25513 6820
rect 25547 6817 25559 6851
rect 25501 6811 25559 6817
rect 25593 6851 25651 6857
rect 25593 6817 25605 6851
rect 25639 6848 25651 6851
rect 26142 6848 26148 6860
rect 25639 6820 26148 6848
rect 25639 6817 25651 6820
rect 25593 6811 25651 6817
rect 26142 6808 26148 6820
rect 26200 6848 26206 6860
rect 26789 6851 26847 6857
rect 26789 6848 26801 6851
rect 26200 6820 26801 6848
rect 26200 6808 26206 6820
rect 26789 6817 26801 6820
rect 26835 6817 26847 6851
rect 27632 6848 27660 6956
rect 27890 6944 27896 6956
rect 27948 6944 27954 6996
rect 26789 6811 26847 6817
rect 26988 6820 27660 6848
rect 20496 6752 20668 6780
rect 20496 6740 20502 6752
rect 20714 6740 20720 6792
rect 20772 6780 20778 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20772 6752 20913 6780
rect 20772 6740 20778 6752
rect 20901 6749 20913 6752
rect 20947 6780 20959 6783
rect 22094 6780 22100 6792
rect 20947 6752 22100 6780
rect 20947 6749 20959 6752
rect 20901 6743 20959 6749
rect 22094 6740 22100 6752
rect 22152 6740 22158 6792
rect 22186 6740 22192 6792
rect 22244 6780 22250 6792
rect 22741 6783 22799 6789
rect 22741 6780 22753 6783
rect 22244 6752 22753 6780
rect 22244 6740 22250 6752
rect 22741 6749 22753 6752
rect 22787 6749 22799 6783
rect 22741 6743 22799 6749
rect 22830 6740 22836 6792
rect 22888 6780 22894 6792
rect 22888 6752 22933 6780
rect 22888 6740 22894 6752
rect 23014 6740 23020 6792
rect 23072 6780 23078 6792
rect 23072 6752 23117 6780
rect 23072 6740 23078 6752
rect 23198 6740 23204 6792
rect 23256 6789 23262 6792
rect 23256 6780 23264 6789
rect 23256 6752 23301 6780
rect 23256 6743 23264 6752
rect 23256 6740 23262 6743
rect 24946 6740 24952 6792
rect 25004 6780 25010 6792
rect 25225 6783 25283 6789
rect 25225 6780 25237 6783
rect 25004 6752 25237 6780
rect 25004 6740 25010 6752
rect 25225 6749 25237 6752
rect 25271 6749 25283 6783
rect 25406 6780 25412 6792
rect 25367 6752 25412 6780
rect 25225 6743 25283 6749
rect 20070 6712 20076 6724
rect 20031 6684 20076 6712
rect 20070 6672 20076 6684
rect 20128 6672 20134 6724
rect 20162 6672 20168 6724
rect 20220 6712 20226 6724
rect 21168 6715 21226 6721
rect 20220 6684 20265 6712
rect 20220 6672 20226 6684
rect 21168 6681 21180 6715
rect 21214 6712 21226 6715
rect 22278 6712 22284 6724
rect 21214 6684 22284 6712
rect 21214 6681 21226 6684
rect 21168 6675 21226 6681
rect 22278 6672 22284 6684
rect 22336 6672 22342 6724
rect 23106 6712 23112 6724
rect 23067 6684 23112 6712
rect 23106 6672 23112 6684
rect 23164 6672 23170 6724
rect 25240 6712 25268 6743
rect 25406 6740 25412 6752
rect 25464 6740 25470 6792
rect 25777 6783 25835 6789
rect 25777 6749 25789 6783
rect 25823 6780 25835 6783
rect 26326 6780 26332 6792
rect 25823 6752 26332 6780
rect 25823 6749 25835 6752
rect 25777 6743 25835 6749
rect 26326 6740 26332 6752
rect 26384 6740 26390 6792
rect 26421 6783 26479 6789
rect 26421 6749 26433 6783
rect 26467 6749 26479 6783
rect 26421 6743 26479 6749
rect 26605 6783 26663 6789
rect 26605 6749 26617 6783
rect 26651 6749 26663 6783
rect 26605 6743 26663 6749
rect 26436 6712 26464 6743
rect 25240 6684 26464 6712
rect 26620 6712 26648 6743
rect 26694 6740 26700 6792
rect 26752 6780 26758 6792
rect 26988 6789 27016 6820
rect 26973 6783 27031 6789
rect 26752 6752 26797 6780
rect 26752 6740 26758 6752
rect 26973 6749 26985 6783
rect 27019 6749 27031 6783
rect 26973 6743 27031 6749
rect 27617 6783 27675 6789
rect 27617 6749 27629 6783
rect 27663 6780 27675 6783
rect 27706 6780 27712 6792
rect 27663 6752 27712 6780
rect 27663 6749 27675 6752
rect 27617 6743 27675 6749
rect 27706 6740 27712 6752
rect 27764 6740 27770 6792
rect 30098 6780 30104 6792
rect 27816 6752 29960 6780
rect 30059 6752 30104 6780
rect 27816 6712 27844 6752
rect 27890 6721 27896 6724
rect 26620 6684 27844 6712
rect 27884 6675 27896 6721
rect 27948 6712 27954 6724
rect 27948 6684 27984 6712
rect 27890 6672 27896 6675
rect 27948 6672 27954 6684
rect 21910 6644 21916 6656
rect 19812 6616 21916 6644
rect 18693 6607 18751 6613
rect 21910 6604 21916 6616
rect 21968 6644 21974 6656
rect 22186 6644 22192 6656
rect 21968 6616 22192 6644
rect 21968 6604 21974 6616
rect 22186 6604 22192 6616
rect 22244 6604 22250 6656
rect 22738 6604 22744 6656
rect 22796 6644 22802 6656
rect 22922 6644 22928 6656
rect 22796 6616 22928 6644
rect 22796 6604 22802 6616
rect 22922 6604 22928 6616
rect 22980 6604 22986 6656
rect 25961 6647 26019 6653
rect 25961 6613 25973 6647
rect 26007 6644 26019 6647
rect 27338 6644 27344 6656
rect 26007 6616 27344 6644
rect 26007 6613 26019 6616
rect 25961 6607 26019 6613
rect 27338 6604 27344 6616
rect 27396 6604 27402 6656
rect 27798 6604 27804 6656
rect 27856 6644 27862 6656
rect 29932 6653 29960 6752
rect 30098 6740 30104 6752
rect 30156 6740 30162 6792
rect 28997 6647 29055 6653
rect 28997 6644 29009 6647
rect 27856 6616 29009 6644
rect 27856 6604 27862 6616
rect 28997 6613 29009 6616
rect 29043 6613 29055 6647
rect 28997 6607 29055 6613
rect 29917 6647 29975 6653
rect 29917 6613 29929 6647
rect 29963 6613 29975 6647
rect 29917 6607 29975 6613
rect 1104 6554 30820 6576
rect 1104 6502 10880 6554
rect 10932 6502 10944 6554
rect 10996 6502 11008 6554
rect 11060 6502 11072 6554
rect 11124 6502 11136 6554
rect 11188 6502 20811 6554
rect 20863 6502 20875 6554
rect 20927 6502 20939 6554
rect 20991 6502 21003 6554
rect 21055 6502 21067 6554
rect 21119 6502 30820 6554
rect 1104 6480 30820 6502
rect 11974 6440 11980 6452
rect 11935 6412 11980 6440
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 12492 6412 12537 6440
rect 12492 6400 12498 6412
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 13265 6443 13323 6449
rect 13265 6440 13277 6443
rect 12952 6412 13277 6440
rect 12952 6400 12958 6412
rect 13265 6409 13277 6412
rect 13311 6409 13323 6443
rect 13265 6403 13323 6409
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 13872 6412 15792 6440
rect 13872 6400 13878 6412
rect 15764 6372 15792 6412
rect 15838 6400 15844 6452
rect 15896 6440 15902 6452
rect 15933 6443 15991 6449
rect 15933 6440 15945 6443
rect 15896 6412 15945 6440
rect 15896 6400 15902 6412
rect 15933 6409 15945 6412
rect 15979 6409 15991 6443
rect 19150 6440 19156 6452
rect 15933 6403 15991 6409
rect 16040 6412 19156 6440
rect 16040 6372 16068 6412
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 21634 6400 21640 6452
rect 21692 6440 21698 6452
rect 21913 6443 21971 6449
rect 21913 6440 21925 6443
rect 21692 6412 21925 6440
rect 21692 6400 21698 6412
rect 21913 6409 21925 6412
rect 21959 6409 21971 6443
rect 25682 6440 25688 6452
rect 25643 6412 25688 6440
rect 21913 6403 21971 6409
rect 25682 6400 25688 6412
rect 25740 6400 25746 6452
rect 27890 6440 27896 6452
rect 27851 6412 27896 6440
rect 27890 6400 27896 6412
rect 27948 6400 27954 6452
rect 28994 6400 29000 6452
rect 29052 6440 29058 6452
rect 29089 6443 29147 6449
rect 29089 6440 29101 6443
rect 29052 6412 29101 6440
rect 29052 6400 29058 6412
rect 29089 6409 29101 6412
rect 29135 6409 29147 6443
rect 29089 6403 29147 6409
rect 29917 6443 29975 6449
rect 29917 6409 29929 6443
rect 29963 6409 29975 6443
rect 29917 6403 29975 6409
rect 15764 6344 16068 6372
rect 16850 6332 16856 6384
rect 16908 6372 16914 6384
rect 17678 6372 17684 6384
rect 16908 6344 17684 6372
rect 16908 6332 16914 6344
rect 17678 6332 17684 6344
rect 17736 6332 17742 6384
rect 18414 6372 18420 6384
rect 17972 6344 18420 6372
rect 12345 6307 12403 6313
rect 12345 6273 12357 6307
rect 12391 6304 12403 6307
rect 12434 6304 12440 6316
rect 12391 6276 12440 6304
rect 12391 6273 12403 6276
rect 12345 6267 12403 6273
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6304 13231 6307
rect 14182 6304 14188 6316
rect 13219 6276 14188 6304
rect 13219 6273 13231 6276
rect 13173 6267 13231 6273
rect 14182 6264 14188 6276
rect 14240 6264 14246 6316
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 17405 6307 17463 6313
rect 17405 6304 17417 6307
rect 17368 6276 17417 6304
rect 17368 6264 17374 6276
rect 17405 6273 17417 6276
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 17494 6264 17500 6316
rect 17552 6304 17558 6316
rect 17773 6307 17831 6313
rect 17552 6276 17597 6304
rect 17552 6264 17558 6276
rect 17773 6273 17785 6307
rect 17819 6273 17831 6307
rect 17773 6267 17831 6273
rect 17870 6307 17928 6313
rect 17870 6273 17882 6307
rect 17916 6304 17928 6307
rect 17972 6304 18000 6344
rect 18414 6332 18420 6344
rect 18472 6332 18478 6384
rect 19702 6372 19708 6384
rect 18892 6344 19708 6372
rect 17916 6276 18000 6304
rect 17916 6273 17928 6276
rect 17870 6267 17928 6273
rect 12621 6239 12679 6245
rect 12621 6205 12633 6239
rect 12667 6236 12679 6239
rect 13538 6236 13544 6248
rect 12667 6208 13544 6236
rect 12667 6205 12679 6208
rect 12621 6199 12679 6205
rect 13538 6196 13544 6208
rect 13596 6196 13602 6248
rect 14090 6236 14096 6248
rect 14051 6208 14096 6236
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 14274 6236 14280 6248
rect 14235 6208 14280 6236
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 15010 6236 15016 6248
rect 14971 6208 15016 6236
rect 15010 6196 15016 6208
rect 15068 6196 15074 6248
rect 15102 6196 15108 6248
rect 15160 6245 15166 6248
rect 15160 6239 15188 6245
rect 15176 6205 15188 6239
rect 15160 6199 15188 6205
rect 15289 6239 15347 6245
rect 15289 6205 15301 6239
rect 15335 6236 15347 6239
rect 15470 6236 15476 6248
rect 15335 6208 15476 6236
rect 15335 6205 15347 6208
rect 15289 6199 15347 6205
rect 15160 6196 15166 6199
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 11238 6128 11244 6180
rect 11296 6168 11302 6180
rect 11790 6168 11796 6180
rect 11296 6140 11796 6168
rect 11296 6128 11302 6140
rect 11790 6128 11796 6140
rect 11848 6168 11854 6180
rect 12802 6168 12808 6180
rect 11848 6140 12808 6168
rect 11848 6128 11854 6140
rect 12802 6128 12808 6140
rect 12860 6168 12866 6180
rect 14737 6171 14795 6177
rect 14737 6168 14749 6171
rect 12860 6140 14749 6168
rect 12860 6128 12866 6140
rect 14737 6137 14749 6140
rect 14783 6168 14795 6171
rect 14826 6168 14832 6180
rect 14783 6140 14832 6168
rect 14783 6137 14795 6140
rect 14737 6131 14795 6137
rect 14826 6128 14832 6140
rect 14884 6128 14890 6180
rect 17788 6168 17816 6267
rect 18046 6264 18052 6316
rect 18104 6304 18110 6316
rect 18690 6304 18696 6316
rect 18104 6276 18696 6304
rect 18104 6264 18110 6276
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 18892 6313 18920 6344
rect 19702 6332 19708 6344
rect 19760 6332 19766 6384
rect 25406 6332 25412 6384
rect 25464 6372 25470 6384
rect 29932 6372 29960 6403
rect 25464 6344 29960 6372
rect 25464 6332 25470 6344
rect 18877 6307 18935 6313
rect 18877 6273 18889 6307
rect 18923 6273 18935 6307
rect 18877 6267 18935 6273
rect 18966 6264 18972 6316
rect 19024 6304 19030 6316
rect 19024 6276 19069 6304
rect 19024 6264 19030 6276
rect 19150 6264 19156 6316
rect 19208 6304 19214 6316
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 19208 6276 19257 6304
rect 19208 6264 19214 6276
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 20438 6304 20444 6316
rect 20399 6276 20444 6304
rect 19245 6267 19303 6273
rect 20438 6264 20444 6276
rect 20496 6264 20502 6316
rect 21818 6304 21824 6316
rect 21779 6276 21824 6304
rect 21818 6264 21824 6276
rect 21876 6264 21882 6316
rect 22094 6264 22100 6316
rect 22152 6304 22158 6316
rect 22738 6313 22744 6316
rect 22465 6307 22523 6313
rect 22465 6304 22477 6307
rect 22152 6276 22477 6304
rect 22152 6264 22158 6276
rect 22465 6273 22477 6276
rect 22511 6273 22523 6307
rect 22465 6267 22523 6273
rect 22732 6267 22744 6313
rect 22796 6304 22802 6316
rect 22796 6276 22832 6304
rect 22738 6264 22744 6267
rect 22796 6264 22802 6276
rect 23934 6264 23940 6316
rect 23992 6304 23998 6316
rect 24305 6307 24363 6313
rect 24305 6304 24317 6307
rect 23992 6276 24317 6304
rect 23992 6264 23998 6276
rect 24305 6273 24317 6276
rect 24351 6273 24363 6307
rect 24305 6267 24363 6273
rect 24572 6307 24630 6313
rect 24572 6273 24584 6307
rect 24618 6304 24630 6307
rect 25590 6304 25596 6316
rect 24618 6276 25596 6304
rect 24618 6273 24630 6276
rect 24572 6267 24630 6273
rect 25590 6264 25596 6276
rect 25648 6264 25654 6316
rect 27065 6307 27123 6313
rect 27065 6273 27077 6307
rect 27111 6304 27123 6307
rect 27157 6307 27215 6313
rect 27157 6304 27169 6307
rect 27111 6276 27169 6304
rect 27111 6273 27123 6276
rect 27065 6267 27123 6273
rect 27157 6273 27169 6276
rect 27203 6273 27215 6307
rect 27157 6267 27215 6273
rect 27341 6307 27399 6313
rect 27341 6273 27353 6307
rect 27387 6304 27399 6307
rect 27614 6304 27620 6316
rect 27387 6276 27620 6304
rect 27387 6273 27399 6276
rect 27341 6267 27399 6273
rect 27614 6264 27620 6276
rect 27672 6264 27678 6316
rect 27709 6307 27767 6313
rect 27709 6273 27721 6307
rect 27755 6304 27767 6307
rect 27798 6304 27804 6316
rect 27755 6276 27804 6304
rect 27755 6273 27767 6276
rect 27709 6267 27767 6273
rect 27798 6264 27804 6276
rect 27856 6264 27862 6316
rect 28350 6304 28356 6316
rect 28311 6276 28356 6304
rect 28350 6264 28356 6276
rect 28408 6264 28414 6316
rect 28537 6307 28595 6313
rect 28537 6273 28549 6307
rect 28583 6304 28595 6307
rect 28810 6304 28816 6316
rect 28583 6276 28816 6304
rect 28583 6273 28595 6276
rect 28537 6267 28595 6273
rect 28810 6264 28816 6276
rect 28868 6264 28874 6316
rect 28905 6307 28963 6313
rect 28905 6273 28917 6307
rect 28951 6304 28963 6307
rect 29914 6304 29920 6316
rect 28951 6276 29920 6304
rect 28951 6273 28963 6276
rect 28905 6267 28963 6273
rect 29914 6264 29920 6276
rect 29972 6264 29978 6316
rect 30098 6304 30104 6316
rect 30059 6276 30104 6304
rect 30098 6264 30104 6276
rect 30156 6264 30162 6316
rect 19061 6239 19119 6245
rect 19061 6205 19073 6239
rect 19107 6236 19119 6239
rect 19334 6236 19340 6248
rect 19107 6208 19340 6236
rect 19107 6205 19119 6208
rect 19061 6199 19119 6205
rect 19334 6196 19340 6208
rect 19392 6236 19398 6248
rect 19978 6236 19984 6248
rect 19392 6208 19984 6236
rect 19392 6196 19398 6208
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 20717 6239 20775 6245
rect 20717 6205 20729 6239
rect 20763 6236 20775 6239
rect 21174 6236 21180 6248
rect 20763 6208 21180 6236
rect 20763 6205 20775 6208
rect 20717 6199 20775 6205
rect 21174 6196 21180 6208
rect 21232 6196 21238 6248
rect 26694 6196 26700 6248
rect 26752 6236 26758 6248
rect 27430 6236 27436 6248
rect 26752 6208 27436 6236
rect 26752 6196 26758 6208
rect 27430 6196 27436 6208
rect 27488 6196 27494 6248
rect 27525 6239 27583 6245
rect 27525 6205 27537 6239
rect 27571 6205 27583 6239
rect 28626 6236 28632 6248
rect 28587 6208 28632 6236
rect 27525 6199 27583 6205
rect 21358 6168 21364 6180
rect 17788 6140 21364 6168
rect 21358 6128 21364 6140
rect 21416 6128 21422 6180
rect 22278 6128 22284 6180
rect 22336 6168 22342 6180
rect 22336 6140 22508 6168
rect 22336 6128 22342 6140
rect 18046 6100 18052 6112
rect 18007 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 19426 6100 19432 6112
rect 19387 6072 19432 6100
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 22480 6100 22508 6140
rect 26142 6128 26148 6180
rect 26200 6168 26206 6180
rect 27540 6168 27568 6199
rect 28626 6196 28632 6208
rect 28684 6196 28690 6248
rect 28718 6196 28724 6248
rect 28776 6236 28782 6248
rect 28776 6208 28821 6236
rect 28776 6196 28782 6208
rect 26200 6140 27568 6168
rect 26200 6128 26206 6140
rect 27614 6128 27620 6180
rect 27672 6168 27678 6180
rect 28644 6168 28672 6196
rect 27672 6140 28672 6168
rect 27672 6128 27678 6140
rect 23566 6100 23572 6112
rect 22480 6072 23572 6100
rect 23566 6060 23572 6072
rect 23624 6100 23630 6112
rect 23845 6103 23903 6109
rect 23845 6100 23857 6103
rect 23624 6072 23857 6100
rect 23624 6060 23630 6072
rect 23845 6069 23857 6072
rect 23891 6069 23903 6103
rect 23845 6063 23903 6069
rect 27065 6103 27123 6109
rect 27065 6069 27077 6103
rect 27111 6100 27123 6103
rect 28350 6100 28356 6112
rect 27111 6072 28356 6100
rect 27111 6069 27123 6072
rect 27065 6063 27123 6069
rect 28350 6060 28356 6072
rect 28408 6060 28414 6112
rect 1104 6010 30820 6032
rect 1104 5958 5915 6010
rect 5967 5958 5979 6010
rect 6031 5958 6043 6010
rect 6095 5958 6107 6010
rect 6159 5958 6171 6010
rect 6223 5958 15846 6010
rect 15898 5958 15910 6010
rect 15962 5958 15974 6010
rect 16026 5958 16038 6010
rect 16090 5958 16102 6010
rect 16154 5958 25776 6010
rect 25828 5958 25840 6010
rect 25892 5958 25904 6010
rect 25956 5958 25968 6010
rect 26020 5958 26032 6010
rect 26084 5958 30820 6010
rect 1104 5936 30820 5958
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12492 5868 12537 5896
rect 12492 5856 12498 5868
rect 14550 5856 14556 5908
rect 14608 5896 14614 5908
rect 15102 5896 15108 5908
rect 14608 5868 15108 5896
rect 14608 5856 14614 5868
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15746 5856 15752 5908
rect 15804 5896 15810 5908
rect 15933 5899 15991 5905
rect 15933 5896 15945 5899
rect 15804 5868 15945 5896
rect 15804 5856 15810 5868
rect 15933 5865 15945 5868
rect 15979 5865 15991 5899
rect 15933 5859 15991 5865
rect 18230 5856 18236 5908
rect 18288 5896 18294 5908
rect 19429 5899 19487 5905
rect 19429 5896 19441 5899
rect 18288 5868 19441 5896
rect 18288 5856 18294 5868
rect 19429 5865 19441 5868
rect 19475 5865 19487 5899
rect 19429 5859 19487 5865
rect 21174 5856 21180 5908
rect 21232 5896 21238 5908
rect 22649 5899 22707 5905
rect 21232 5868 22600 5896
rect 21232 5856 21238 5868
rect 9953 5831 10011 5837
rect 9953 5797 9965 5831
rect 9999 5797 10011 5831
rect 9953 5791 10011 5797
rect 9968 5760 9996 5791
rect 10594 5788 10600 5840
rect 10652 5828 10658 5840
rect 10652 5800 11376 5828
rect 10652 5788 10658 5800
rect 10778 5760 10784 5772
rect 9968 5732 10784 5760
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 11238 5760 11244 5772
rect 11199 5732 11244 5760
rect 11238 5720 11244 5732
rect 11296 5720 11302 5772
rect 11348 5760 11376 5800
rect 19518 5788 19524 5840
rect 19576 5828 19582 5840
rect 19705 5831 19763 5837
rect 19705 5828 19717 5831
rect 19576 5800 19717 5828
rect 19576 5788 19582 5800
rect 19705 5797 19717 5800
rect 19751 5797 19763 5831
rect 19705 5791 19763 5797
rect 19797 5831 19855 5837
rect 19797 5797 19809 5831
rect 19843 5828 19855 5831
rect 20070 5828 20076 5840
rect 19843 5800 20076 5828
rect 19843 5797 19855 5800
rect 19797 5791 19855 5797
rect 20070 5788 20076 5800
rect 20128 5788 20134 5840
rect 21818 5828 21824 5840
rect 21008 5800 21824 5828
rect 11514 5760 11520 5772
rect 11348 5732 11520 5760
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 11606 5720 11612 5772
rect 11664 5769 11670 5772
rect 11664 5763 11692 5769
rect 11680 5729 11692 5763
rect 11664 5723 11692 5729
rect 11793 5763 11851 5769
rect 11793 5729 11805 5763
rect 11839 5760 11851 5763
rect 12342 5760 12348 5772
rect 11839 5732 12348 5760
rect 11839 5729 11851 5732
rect 11793 5723 11851 5729
rect 11664 5720 11670 5723
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 13541 5763 13599 5769
rect 13541 5729 13553 5763
rect 13587 5760 13599 5763
rect 13814 5760 13820 5772
rect 13587 5732 13820 5760
rect 13587 5729 13599 5732
rect 13541 5723 13599 5729
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 14734 5760 14740 5772
rect 14695 5732 14740 5760
rect 14734 5720 14740 5732
rect 14792 5720 14798 5772
rect 15102 5720 15108 5772
rect 15160 5769 15166 5772
rect 15160 5763 15188 5769
rect 15176 5729 15188 5763
rect 15160 5723 15188 5729
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5760 15347 5763
rect 15470 5760 15476 5772
rect 15335 5732 15476 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 15160 5720 15166 5723
rect 15470 5720 15476 5732
rect 15528 5720 15534 5772
rect 21008 5760 21036 5800
rect 21174 5760 21180 5772
rect 19628 5732 21036 5760
rect 21135 5732 21180 5760
rect 19628 5704 19656 5732
rect 21174 5720 21180 5732
rect 21232 5720 21238 5772
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10594 5692 10600 5704
rect 10555 5664 10600 5692
rect 10137 5655 10195 5661
rect 10152 5556 10180 5655
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 13262 5692 13268 5704
rect 13223 5664 13268 5692
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 13357 5695 13415 5701
rect 13357 5661 13369 5695
rect 13403 5692 13415 5695
rect 13630 5692 13636 5704
rect 13403 5664 13636 5692
rect 13403 5661 13415 5664
rect 13357 5655 13415 5661
rect 13630 5652 13636 5664
rect 13688 5652 13694 5704
rect 14090 5692 14096 5704
rect 14003 5664 14096 5692
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 14274 5692 14280 5704
rect 14235 5664 14280 5692
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 15010 5652 15016 5704
rect 15068 5692 15074 5704
rect 16390 5692 16396 5704
rect 15068 5664 15113 5692
rect 16351 5664 16396 5692
rect 15068 5652 15074 5664
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 19610 5692 19616 5704
rect 19571 5664 19616 5692
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 19794 5652 19800 5704
rect 19852 5692 19858 5704
rect 19889 5695 19947 5701
rect 19889 5692 19901 5695
rect 19852 5664 19901 5692
rect 19852 5652 19858 5664
rect 19889 5661 19901 5664
rect 19935 5661 19947 5695
rect 19889 5655 19947 5661
rect 20809 5695 20867 5701
rect 20809 5661 20821 5695
rect 20855 5661 20867 5695
rect 20978 5692 20984 5704
rect 20939 5664 20984 5692
rect 20809 5655 20867 5661
rect 14108 5624 14136 5652
rect 14108 5596 14228 5624
rect 11882 5556 11888 5568
rect 10152 5528 11888 5556
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 12986 5516 12992 5568
rect 13044 5556 13050 5568
rect 13541 5559 13599 5565
rect 13541 5556 13553 5559
rect 13044 5528 13553 5556
rect 13044 5516 13050 5528
rect 13541 5525 13553 5528
rect 13587 5525 13599 5559
rect 14200 5556 14228 5596
rect 15010 5556 15016 5568
rect 14200 5528 15016 5556
rect 13541 5519 13599 5525
rect 15010 5516 15016 5528
rect 15068 5516 15074 5568
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 16482 5556 16488 5568
rect 15344 5528 16488 5556
rect 15344 5516 15350 5528
rect 16482 5516 16488 5528
rect 16540 5516 16546 5568
rect 20824 5556 20852 5655
rect 20978 5652 20984 5664
rect 21036 5652 21042 5704
rect 21085 5695 21143 5701
rect 21085 5661 21097 5695
rect 21131 5661 21143 5695
rect 21284 5692 21312 5800
rect 21818 5788 21824 5800
rect 21876 5788 21882 5840
rect 22572 5704 22600 5868
rect 22649 5865 22661 5899
rect 22695 5896 22707 5899
rect 22738 5896 22744 5908
rect 22695 5868 22744 5896
rect 22695 5865 22707 5868
rect 22649 5859 22707 5865
rect 22738 5856 22744 5868
rect 22796 5856 22802 5908
rect 26602 5856 26608 5908
rect 26660 5896 26666 5908
rect 26697 5899 26755 5905
rect 26697 5896 26709 5899
rect 26660 5868 26709 5896
rect 26660 5856 26666 5868
rect 26697 5865 26709 5868
rect 26743 5865 26755 5899
rect 28537 5899 28595 5905
rect 28537 5896 28549 5899
rect 26697 5859 26755 5865
rect 26896 5868 28549 5896
rect 26326 5788 26332 5840
rect 26384 5828 26390 5840
rect 26896 5828 26924 5868
rect 28537 5865 28549 5868
rect 28583 5865 28595 5899
rect 28537 5859 28595 5865
rect 26384 5800 26924 5828
rect 26384 5788 26390 5800
rect 23934 5720 23940 5772
rect 23992 5760 23998 5772
rect 25317 5763 25375 5769
rect 25317 5760 25329 5763
rect 23992 5732 25329 5760
rect 23992 5720 23998 5732
rect 25317 5729 25329 5732
rect 25363 5729 25375 5763
rect 25317 5723 25375 5729
rect 21358 5692 21364 5704
rect 21271 5664 21364 5692
rect 21085 5655 21143 5661
rect 21100 5624 21128 5655
rect 21358 5652 21364 5664
rect 21416 5652 21422 5704
rect 21910 5652 21916 5704
rect 21968 5690 21974 5704
rect 22005 5695 22063 5701
rect 22005 5690 22017 5695
rect 21968 5662 22017 5690
rect 21968 5652 21974 5662
rect 22005 5661 22017 5662
rect 22051 5661 22063 5695
rect 22005 5655 22063 5661
rect 22098 5695 22156 5701
rect 22098 5661 22110 5695
rect 22144 5661 22156 5695
rect 22278 5692 22284 5704
rect 22239 5664 22284 5692
rect 22098 5655 22156 5661
rect 21266 5624 21272 5636
rect 21100 5596 21272 5624
rect 21266 5584 21272 5596
rect 21324 5624 21330 5636
rect 22113 5624 22141 5655
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 22554 5701 22560 5704
rect 22509 5695 22560 5701
rect 22509 5661 22521 5695
rect 22555 5661 22560 5695
rect 22509 5655 22560 5661
rect 22554 5652 22560 5655
rect 22612 5692 22618 5704
rect 23198 5692 23204 5704
rect 22612 5664 23204 5692
rect 22612 5652 22618 5664
rect 23198 5652 23204 5664
rect 23256 5652 23262 5704
rect 27157 5695 27215 5701
rect 27157 5661 27169 5695
rect 27203 5692 27215 5695
rect 27706 5692 27712 5704
rect 27203 5664 27712 5692
rect 27203 5661 27215 5664
rect 27157 5655 27215 5661
rect 27706 5652 27712 5664
rect 27764 5652 27770 5704
rect 21324 5596 22141 5624
rect 22373 5627 22431 5633
rect 21324 5584 21330 5596
rect 22112 5568 22140 5596
rect 22373 5593 22385 5627
rect 22419 5624 22431 5627
rect 22922 5624 22928 5636
rect 22419 5596 22928 5624
rect 22419 5593 22431 5596
rect 22373 5587 22431 5593
rect 22922 5584 22928 5596
rect 22980 5624 22986 5636
rect 25584 5627 25642 5633
rect 22980 5596 24164 5624
rect 22980 5584 22986 5596
rect 21174 5556 21180 5568
rect 20824 5528 21180 5556
rect 21174 5516 21180 5528
rect 21232 5516 21238 5568
rect 21542 5556 21548 5568
rect 21503 5528 21548 5556
rect 21542 5516 21548 5528
rect 21600 5516 21606 5568
rect 22094 5516 22100 5568
rect 22152 5516 22158 5568
rect 24136 5556 24164 5596
rect 25584 5593 25596 5627
rect 25630 5624 25642 5627
rect 26142 5624 26148 5636
rect 25630 5596 26148 5624
rect 25630 5593 25642 5596
rect 25584 5587 25642 5593
rect 26142 5584 26148 5596
rect 26200 5584 26206 5636
rect 27338 5584 27344 5636
rect 27396 5633 27402 5636
rect 27396 5627 27460 5633
rect 27396 5593 27414 5627
rect 27448 5593 27460 5627
rect 29914 5624 29920 5636
rect 29875 5596 29920 5624
rect 27396 5587 27460 5593
rect 27396 5584 27402 5587
rect 29914 5584 29920 5596
rect 29972 5584 29978 5636
rect 29178 5556 29184 5568
rect 24136 5528 29184 5556
rect 29178 5516 29184 5528
rect 29236 5516 29242 5568
rect 30006 5556 30012 5568
rect 29967 5528 30012 5556
rect 30006 5516 30012 5528
rect 30064 5516 30070 5568
rect 1104 5466 30820 5488
rect 1104 5414 10880 5466
rect 10932 5414 10944 5466
rect 10996 5414 11008 5466
rect 11060 5414 11072 5466
rect 11124 5414 11136 5466
rect 11188 5414 20811 5466
rect 20863 5414 20875 5466
rect 20927 5414 20939 5466
rect 20991 5414 21003 5466
rect 21055 5414 21067 5466
rect 21119 5414 30820 5466
rect 1104 5392 30820 5414
rect 11882 5352 11888 5364
rect 11843 5324 11888 5352
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 14274 5312 14280 5364
rect 14332 5352 14338 5364
rect 14829 5355 14887 5361
rect 14829 5352 14841 5355
rect 14332 5324 14841 5352
rect 14332 5312 14338 5324
rect 14829 5321 14841 5324
rect 14875 5321 14887 5355
rect 14829 5315 14887 5321
rect 17678 5312 17684 5364
rect 17736 5352 17742 5364
rect 18417 5355 18475 5361
rect 18417 5352 18429 5355
rect 17736 5324 18429 5352
rect 17736 5312 17742 5324
rect 18417 5321 18429 5324
rect 18463 5321 18475 5355
rect 18417 5315 18475 5321
rect 19150 5312 19156 5364
rect 19208 5352 19214 5364
rect 20349 5355 20407 5361
rect 20349 5352 20361 5355
rect 19208 5324 20361 5352
rect 19208 5312 19214 5324
rect 20349 5321 20361 5324
rect 20395 5321 20407 5355
rect 20349 5315 20407 5321
rect 25590 5312 25596 5364
rect 25648 5352 25654 5364
rect 25777 5355 25835 5361
rect 25777 5352 25789 5355
rect 25648 5324 25789 5352
rect 25648 5312 25654 5324
rect 25777 5321 25789 5324
rect 25823 5321 25835 5355
rect 25777 5315 25835 5321
rect 18230 5284 18236 5296
rect 14476 5256 15424 5284
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5216 1455 5219
rect 1486 5216 1492 5228
rect 1443 5188 1492 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 1486 5176 1492 5188
rect 1544 5176 1550 5228
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5216 11759 5219
rect 12986 5216 12992 5228
rect 11747 5188 12992 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 13173 5219 13231 5225
rect 13173 5185 13185 5219
rect 13219 5216 13231 5219
rect 13219 5188 13584 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 11517 5151 11575 5157
rect 11517 5117 11529 5151
rect 11563 5117 11575 5151
rect 11517 5111 11575 5117
rect 11532 5080 11560 5111
rect 12434 5080 12440 5092
rect 11532 5052 12440 5080
rect 12434 5040 12440 5052
rect 12492 5080 12498 5092
rect 12989 5083 13047 5089
rect 12989 5080 13001 5083
rect 12492 5052 13001 5080
rect 12492 5040 12498 5052
rect 12989 5049 13001 5052
rect 13035 5049 13047 5083
rect 13556 5080 13584 5188
rect 13630 5176 13636 5228
rect 13688 5216 13694 5228
rect 14366 5216 14372 5228
rect 13688 5188 14372 5216
rect 13688 5176 13694 5188
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5148 13783 5151
rect 13814 5148 13820 5160
rect 13771 5120 13820 5148
rect 13771 5117 13783 5120
rect 13725 5111 13783 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14001 5083 14059 5089
rect 14001 5080 14013 5083
rect 13556 5052 14013 5080
rect 12989 5043 13047 5049
rect 14001 5049 14013 5052
rect 14047 5049 14059 5083
rect 14476 5080 14504 5256
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5185 15071 5219
rect 15013 5179 15071 5185
rect 15105 5219 15163 5225
rect 15105 5185 15117 5219
rect 15151 5216 15163 5219
rect 15286 5216 15292 5228
rect 15151 5188 15292 5216
rect 15151 5185 15163 5188
rect 15105 5179 15163 5185
rect 15028 5148 15056 5179
rect 15286 5176 15292 5188
rect 15344 5176 15350 5228
rect 15396 5225 15424 5256
rect 17052 5256 18236 5284
rect 17052 5228 17080 5256
rect 18230 5244 18236 5256
rect 18288 5284 18294 5296
rect 18598 5284 18604 5296
rect 18288 5256 18604 5284
rect 18288 5244 18294 5256
rect 18598 5244 18604 5256
rect 18656 5244 18662 5296
rect 19236 5287 19294 5293
rect 19236 5253 19248 5287
rect 19282 5284 19294 5287
rect 19426 5284 19432 5296
rect 19282 5256 19432 5284
rect 19282 5253 19294 5256
rect 19236 5247 19294 5253
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 19794 5244 19800 5296
rect 19852 5284 19858 5296
rect 19852 5256 22416 5284
rect 19852 5244 19858 5256
rect 15381 5219 15439 5225
rect 15381 5185 15393 5219
rect 15427 5216 15439 5219
rect 15470 5216 15476 5228
rect 15427 5188 15476 5216
rect 15427 5185 15439 5188
rect 15381 5179 15439 5185
rect 15470 5176 15476 5188
rect 15528 5216 15534 5228
rect 17034 5216 17040 5228
rect 15528 5188 16528 5216
rect 16947 5188 17040 5216
rect 15528 5176 15534 5188
rect 15028 5120 15424 5148
rect 15396 5092 15424 5120
rect 14001 5043 14059 5049
rect 14292 5052 14504 5080
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 13262 4972 13268 5024
rect 13320 5012 13326 5024
rect 13817 5015 13875 5021
rect 13817 5012 13829 5015
rect 13320 4984 13829 5012
rect 13320 4972 13326 4984
rect 13817 4981 13829 4984
rect 13863 5012 13875 5015
rect 14292 5012 14320 5052
rect 15378 5040 15384 5092
rect 15436 5040 15442 5092
rect 13863 4984 14320 5012
rect 13863 4981 13875 4984
rect 13817 4975 13875 4981
rect 14366 4972 14372 5024
rect 14424 5012 14430 5024
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 14424 4984 15301 5012
rect 14424 4972 14430 4984
rect 15289 4981 15301 4984
rect 15335 5012 15347 5015
rect 16390 5012 16396 5024
rect 15335 4984 16396 5012
rect 15335 4981 15347 4984
rect 15289 4975 15347 4981
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 16500 5012 16528 5188
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 17304 5219 17362 5225
rect 17304 5185 17316 5219
rect 17350 5216 17362 5219
rect 18046 5216 18052 5228
rect 17350 5188 18052 5216
rect 17350 5185 17362 5188
rect 17304 5179 17362 5185
rect 18046 5176 18052 5188
rect 18104 5176 18110 5228
rect 18616 5216 18644 5244
rect 18969 5219 19027 5225
rect 18969 5216 18981 5219
rect 18616 5188 18981 5216
rect 18969 5185 18981 5188
rect 19015 5185 19027 5219
rect 18969 5179 19027 5185
rect 21174 5176 21180 5228
rect 21232 5216 21238 5228
rect 21726 5216 21732 5228
rect 21232 5188 21732 5216
rect 21232 5176 21238 5188
rect 21726 5176 21732 5188
rect 21784 5216 21790 5228
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 21784 5188 21833 5216
rect 21784 5176 21790 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 22002 5216 22008 5228
rect 21963 5188 22008 5216
rect 21821 5179 21879 5185
rect 22002 5176 22008 5188
rect 22060 5176 22066 5228
rect 22094 5176 22100 5228
rect 22152 5216 22158 5228
rect 22388 5225 22416 5256
rect 23842 5244 23848 5296
rect 23900 5284 23906 5296
rect 30006 5284 30012 5296
rect 23900 5256 30012 5284
rect 23900 5244 23906 5256
rect 22373 5219 22431 5225
rect 22152 5188 22197 5216
rect 22152 5176 22158 5188
rect 22373 5185 22385 5219
rect 22419 5216 22431 5219
rect 23198 5216 23204 5228
rect 22419 5188 23204 5216
rect 22419 5185 22431 5188
rect 22373 5179 22431 5185
rect 23198 5176 23204 5188
rect 23256 5176 23262 5228
rect 24946 5176 24952 5228
rect 25004 5216 25010 5228
rect 25240 5225 25268 5256
rect 30006 5244 30012 5256
rect 30064 5244 30070 5296
rect 25041 5219 25099 5225
rect 25041 5216 25053 5219
rect 25004 5188 25053 5216
rect 25004 5176 25010 5188
rect 25041 5185 25053 5188
rect 25087 5185 25099 5219
rect 25041 5179 25099 5185
rect 25225 5219 25283 5225
rect 25225 5185 25237 5219
rect 25271 5185 25283 5219
rect 25225 5179 25283 5185
rect 25593 5219 25651 5225
rect 25593 5185 25605 5219
rect 25639 5216 25651 5219
rect 25682 5216 25688 5228
rect 25639 5188 25688 5216
rect 25639 5185 25651 5188
rect 25593 5179 25651 5185
rect 25682 5176 25688 5188
rect 25740 5176 25746 5228
rect 29914 5216 29920 5228
rect 29875 5188 29920 5216
rect 29914 5176 29920 5188
rect 29972 5176 29978 5228
rect 22020 5080 22048 5176
rect 22189 5151 22247 5157
rect 22189 5117 22201 5151
rect 22235 5148 22247 5151
rect 22554 5148 22560 5160
rect 22235 5120 22560 5148
rect 22235 5117 22247 5120
rect 22189 5111 22247 5117
rect 22554 5108 22560 5120
rect 22612 5108 22618 5160
rect 25314 5148 25320 5160
rect 25275 5120 25320 5148
rect 25314 5108 25320 5120
rect 25372 5108 25378 5160
rect 25409 5151 25467 5157
rect 25409 5117 25421 5151
rect 25455 5148 25467 5151
rect 25774 5148 25780 5160
rect 25455 5120 25780 5148
rect 25455 5117 25467 5120
rect 25409 5111 25467 5117
rect 25774 5108 25780 5120
rect 25832 5148 25838 5160
rect 26050 5148 26056 5160
rect 25832 5120 26056 5148
rect 25832 5108 25838 5120
rect 26050 5108 26056 5120
rect 26108 5108 26114 5160
rect 28994 5080 29000 5092
rect 22020 5052 29000 5080
rect 28994 5040 29000 5052
rect 29052 5040 29058 5092
rect 18138 5012 18144 5024
rect 16500 4984 18144 5012
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 22554 5012 22560 5024
rect 22515 4984 22560 5012
rect 22554 4972 22560 4984
rect 22612 4972 22618 5024
rect 30006 5012 30012 5024
rect 29967 4984 30012 5012
rect 30006 4972 30012 4984
rect 30064 4972 30070 5024
rect 1104 4922 30820 4944
rect 1104 4870 5915 4922
rect 5967 4870 5979 4922
rect 6031 4870 6043 4922
rect 6095 4870 6107 4922
rect 6159 4870 6171 4922
rect 6223 4870 15846 4922
rect 15898 4870 15910 4922
rect 15962 4870 15974 4922
rect 16026 4870 16038 4922
rect 16090 4870 16102 4922
rect 16154 4870 25776 4922
rect 25828 4870 25840 4922
rect 25892 4870 25904 4922
rect 25956 4870 25968 4922
rect 26020 4870 26032 4922
rect 26084 4870 30820 4922
rect 1104 4848 30820 4870
rect 12710 4808 12716 4820
rect 12671 4780 12716 4808
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 17034 4808 17040 4820
rect 16132 4780 17040 4808
rect 11514 4700 11520 4752
rect 11572 4740 11578 4752
rect 14093 4743 14151 4749
rect 14093 4740 14105 4743
rect 11572 4712 14105 4740
rect 11572 4700 11578 4712
rect 14093 4709 14105 4712
rect 14139 4740 14151 4743
rect 14550 4740 14556 4752
rect 14139 4712 14556 4740
rect 14139 4709 14151 4712
rect 14093 4703 14151 4709
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 13357 4675 13415 4681
rect 13357 4641 13369 4675
rect 13403 4672 13415 4675
rect 13538 4672 13544 4684
rect 13403 4644 13544 4672
rect 13403 4641 13415 4644
rect 13357 4635 13415 4641
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 14461 4675 14519 4681
rect 14461 4641 14473 4675
rect 14507 4672 14519 4675
rect 14734 4672 14740 4684
rect 14507 4644 14740 4672
rect 14507 4641 14519 4644
rect 14461 4635 14519 4641
rect 14734 4632 14740 4644
rect 14792 4632 14798 4684
rect 16132 4681 16160 4780
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 21358 4808 21364 4820
rect 21319 4780 21364 4808
rect 21358 4768 21364 4780
rect 21416 4768 21422 4820
rect 22738 4768 22744 4820
rect 22796 4768 22802 4820
rect 23198 4808 23204 4820
rect 23159 4780 23204 4808
rect 23198 4768 23204 4780
rect 23256 4768 23262 4820
rect 26142 4808 26148 4820
rect 26103 4780 26148 4808
rect 26142 4768 26148 4780
rect 26200 4768 26206 4820
rect 22756 4740 22784 4768
rect 30006 4740 30012 4752
rect 22756 4712 30012 4740
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4641 16175 4675
rect 16117 4635 16175 4641
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14553 4607 14611 4613
rect 14553 4573 14565 4607
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4604 15071 4607
rect 15470 4604 15476 4616
rect 15059 4576 15476 4604
rect 15059 4573 15071 4576
rect 15013 4567 15071 4573
rect 14568 4536 14596 4567
rect 15470 4564 15476 4576
rect 15528 4564 15534 4616
rect 16384 4607 16442 4613
rect 16384 4573 16396 4607
rect 16430 4604 16442 4607
rect 16666 4604 16672 4616
rect 16430 4576 16672 4604
rect 16430 4573 16442 4576
rect 16384 4567 16442 4573
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 19981 4607 20039 4613
rect 19981 4573 19993 4607
rect 20027 4604 20039 4607
rect 20714 4604 20720 4616
rect 20027 4576 20720 4604
rect 20027 4573 20039 4576
rect 19981 4567 20039 4573
rect 20714 4564 20720 4576
rect 20772 4604 20778 4616
rect 21821 4607 21879 4613
rect 21821 4604 21833 4607
rect 20772 4576 21833 4604
rect 20772 4564 20778 4576
rect 21821 4573 21833 4576
rect 21867 4573 21879 4607
rect 21821 4567 21879 4573
rect 22088 4607 22146 4613
rect 22088 4573 22100 4607
rect 22134 4604 22146 4607
rect 22554 4604 22560 4616
rect 22134 4576 22560 4604
rect 22134 4573 22146 4576
rect 22088 4567 22146 4573
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 24946 4564 24952 4616
rect 25004 4604 25010 4616
rect 25608 4613 25636 4712
rect 30006 4700 30012 4712
rect 30064 4700 30070 4752
rect 25774 4672 25780 4684
rect 25735 4644 25780 4672
rect 25774 4632 25780 4644
rect 25832 4632 25838 4684
rect 25409 4607 25467 4613
rect 25409 4604 25421 4607
rect 25004 4576 25421 4604
rect 25004 4564 25010 4576
rect 25409 4573 25421 4576
rect 25455 4573 25467 4607
rect 25409 4567 25467 4573
rect 25593 4607 25651 4613
rect 25593 4573 25605 4607
rect 25639 4573 25651 4607
rect 25593 4567 25651 4573
rect 25685 4607 25743 4613
rect 25685 4573 25697 4607
rect 25731 4573 25743 4607
rect 25685 4567 25743 4573
rect 25961 4607 26019 4613
rect 25961 4573 25973 4607
rect 26007 4604 26019 4607
rect 26602 4604 26608 4616
rect 26007 4576 26608 4604
rect 26007 4573 26019 4576
rect 25961 4567 26019 4573
rect 20248 4539 20306 4545
rect 14568 4508 15148 4536
rect 13078 4468 13084 4480
rect 13039 4440 13084 4468
rect 13078 4428 13084 4440
rect 13136 4428 13142 4480
rect 13170 4428 13176 4480
rect 13228 4468 13234 4480
rect 15120 4477 15148 4508
rect 20248 4505 20260 4539
rect 20294 4536 20306 4539
rect 21542 4536 21548 4548
rect 20294 4508 21548 4536
rect 20294 4505 20306 4508
rect 20248 4499 20306 4505
rect 21542 4496 21548 4508
rect 21600 4496 21606 4548
rect 25314 4496 25320 4548
rect 25372 4536 25378 4548
rect 25700 4536 25728 4567
rect 26602 4564 26608 4576
rect 26660 4564 26666 4616
rect 29914 4536 29920 4548
rect 25372 4508 25728 4536
rect 29875 4508 29920 4536
rect 25372 4496 25378 4508
rect 29914 4496 29920 4508
rect 29972 4496 29978 4548
rect 15105 4471 15163 4477
rect 13228 4440 13273 4468
rect 13228 4428 13234 4440
rect 15105 4437 15117 4471
rect 15151 4468 15163 4471
rect 15378 4468 15384 4480
rect 15151 4440 15384 4468
rect 15151 4437 15163 4440
rect 15105 4431 15163 4437
rect 15378 4428 15384 4440
rect 15436 4428 15442 4480
rect 16390 4428 16396 4480
rect 16448 4468 16454 4480
rect 17497 4471 17555 4477
rect 17497 4468 17509 4471
rect 16448 4440 17509 4468
rect 16448 4428 16454 4440
rect 17497 4437 17509 4440
rect 17543 4437 17555 4471
rect 17497 4431 17555 4437
rect 23106 4428 23112 4480
rect 23164 4468 23170 4480
rect 30009 4471 30067 4477
rect 30009 4468 30021 4471
rect 23164 4440 30021 4468
rect 23164 4428 23170 4440
rect 30009 4437 30021 4440
rect 30055 4437 30067 4471
rect 30009 4431 30067 4437
rect 1104 4378 30820 4400
rect 1104 4326 10880 4378
rect 10932 4326 10944 4378
rect 10996 4326 11008 4378
rect 11060 4326 11072 4378
rect 11124 4326 11136 4378
rect 11188 4326 20811 4378
rect 20863 4326 20875 4378
rect 20927 4326 20939 4378
rect 20991 4326 21003 4378
rect 21055 4326 21067 4378
rect 21119 4326 30820 4378
rect 1104 4304 30820 4326
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 10560 4100 11713 4128
rect 10560 4088 10566 4100
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 13262 4128 13268 4140
rect 12575 4100 13268 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 13814 4128 13820 4140
rect 13587 4100 13820 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 14366 4128 14372 4140
rect 14327 4100 14372 4128
rect 14366 4088 14372 4100
rect 14424 4088 14430 4140
rect 15197 4131 15255 4137
rect 15197 4097 15209 4131
rect 15243 4097 15255 4131
rect 15378 4128 15384 4140
rect 15339 4100 15384 4128
rect 15197 4091 15255 4097
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 12360 4032 13001 4060
rect 12250 3952 12256 4004
rect 12308 3992 12314 4004
rect 12360 4001 12388 4032
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 12989 4023 13047 4029
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4029 13691 4063
rect 14182 4060 14188 4072
rect 14143 4032 14188 4060
rect 13633 4023 13691 4029
rect 12345 3995 12403 4001
rect 12345 3992 12357 3995
rect 12308 3964 12357 3992
rect 12308 3952 12314 3964
rect 12345 3961 12357 3964
rect 12391 3961 12403 3995
rect 12345 3955 12403 3961
rect 13265 3995 13323 4001
rect 13265 3961 13277 3995
rect 13311 3961 13323 3995
rect 13648 3992 13676 4023
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 14734 4060 14740 4072
rect 14695 4032 14740 4060
rect 14734 4020 14740 4032
rect 14792 4060 14798 4072
rect 15212 4060 15240 4091
rect 15378 4088 15384 4100
rect 15436 4088 15442 4140
rect 17034 4128 17040 4140
rect 16995 4100 17040 4128
rect 17034 4088 17040 4100
rect 17092 4088 17098 4140
rect 18230 4128 18236 4140
rect 18191 4100 18236 4128
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 18506 4137 18512 4140
rect 18500 4128 18512 4137
rect 18467 4100 18512 4128
rect 18500 4091 18512 4100
rect 18506 4088 18512 4091
rect 18564 4088 18570 4140
rect 29825 4131 29883 4137
rect 29825 4097 29837 4131
rect 29871 4128 29883 4131
rect 30006 4128 30012 4140
rect 29871 4100 30012 4128
rect 29871 4097 29883 4100
rect 29825 4091 29883 4097
rect 30006 4088 30012 4100
rect 30064 4088 30070 4140
rect 14792 4032 15240 4060
rect 14792 4020 14798 4032
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 17126 4060 17132 4072
rect 16632 4032 16896 4060
rect 17087 4032 17132 4060
rect 16632 4020 16638 4032
rect 14645 3995 14703 4001
rect 13648 3964 14320 3992
rect 13265 3955 13323 3961
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11204 3896 11529 3924
rect 11204 3884 11210 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 13280 3924 13308 3955
rect 14292 3936 14320 3964
rect 14645 3961 14657 3995
rect 14691 3992 14703 3995
rect 15010 3992 15016 4004
rect 14691 3964 15016 3992
rect 14691 3961 14703 3964
rect 14645 3955 14703 3961
rect 15010 3952 15016 3964
rect 15068 3992 15074 4004
rect 15378 3992 15384 4004
rect 15068 3964 15384 3992
rect 15068 3952 15074 3964
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 16669 3995 16727 4001
rect 16669 3961 16681 3995
rect 16715 3992 16727 3995
rect 16758 3992 16764 4004
rect 16715 3964 16764 3992
rect 16715 3961 16727 3964
rect 16669 3955 16727 3961
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 16868 3992 16896 4032
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 17221 4063 17279 4069
rect 17221 4029 17233 4063
rect 17267 4029 17279 4063
rect 17221 4023 17279 4029
rect 17236 3992 17264 4023
rect 16868 3964 17264 3992
rect 29178 3952 29184 4004
rect 29236 3992 29242 4004
rect 30009 3995 30067 4001
rect 30009 3992 30021 3995
rect 29236 3964 30021 3992
rect 29236 3952 29242 3964
rect 30009 3961 30021 3964
rect 30055 3961 30067 3995
rect 30009 3955 30067 3961
rect 11664 3896 13308 3924
rect 11664 3884 11670 3896
rect 14274 3884 14280 3936
rect 14332 3924 14338 3936
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 14332 3896 15301 3924
rect 14332 3884 14338 3896
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 15289 3887 15347 3893
rect 18874 3884 18880 3936
rect 18932 3924 18938 3936
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 18932 3896 19625 3924
rect 18932 3884 18938 3896
rect 19613 3893 19625 3896
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 1104 3834 30820 3856
rect 1104 3782 5915 3834
rect 5967 3782 5979 3834
rect 6031 3782 6043 3834
rect 6095 3782 6107 3834
rect 6159 3782 6171 3834
rect 6223 3782 15846 3834
rect 15898 3782 15910 3834
rect 15962 3782 15974 3834
rect 16026 3782 16038 3834
rect 16090 3782 16102 3834
rect 16154 3782 25776 3834
rect 25828 3782 25840 3834
rect 25892 3782 25904 3834
rect 25956 3782 25968 3834
rect 26020 3782 26032 3834
rect 26084 3782 30820 3834
rect 1104 3760 30820 3782
rect 10502 3720 10508 3732
rect 10463 3692 10508 3720
rect 10502 3680 10508 3692
rect 10560 3680 10566 3732
rect 12434 3720 12440 3732
rect 11348 3692 12440 3720
rect 11146 3584 11152 3596
rect 11107 3556 11152 3584
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 11348 3593 11376 3692
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 12989 3723 13047 3729
rect 12989 3689 13001 3723
rect 13035 3720 13047 3723
rect 13078 3720 13084 3732
rect 13035 3692 13084 3720
rect 13035 3689 13047 3692
rect 12989 3683 13047 3689
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 16209 3723 16267 3729
rect 16209 3689 16221 3723
rect 16255 3720 16267 3723
rect 17034 3720 17040 3732
rect 16255 3692 17040 3720
rect 16255 3689 16267 3692
rect 16209 3683 16267 3689
rect 17034 3680 17040 3692
rect 17092 3680 17098 3732
rect 11606 3612 11612 3664
rect 11664 3612 11670 3664
rect 11790 3652 11796 3664
rect 11751 3624 11796 3652
rect 11790 3612 11796 3624
rect 11848 3612 11854 3664
rect 14366 3612 14372 3664
rect 14424 3652 14430 3664
rect 14424 3624 14596 3652
rect 14424 3612 14430 3624
rect 11333 3587 11391 3593
rect 11333 3553 11345 3587
rect 11379 3553 11391 3587
rect 11624 3584 11652 3612
rect 12250 3593 12256 3596
rect 12069 3587 12127 3593
rect 12069 3584 12081 3587
rect 11333 3547 11391 3553
rect 11532 3556 12081 3584
rect 10689 3519 10747 3525
rect 10689 3485 10701 3519
rect 10735 3516 10747 3519
rect 11532 3516 11560 3556
rect 12069 3553 12081 3556
rect 12115 3553 12127 3587
rect 12207 3587 12256 3593
rect 12207 3584 12219 3587
rect 12163 3556 12219 3584
rect 12069 3547 12127 3553
rect 12207 3553 12219 3556
rect 12253 3553 12256 3587
rect 12207 3547 12256 3553
rect 12250 3544 12256 3547
rect 12308 3584 12314 3596
rect 12526 3584 12532 3596
rect 12308 3556 12532 3584
rect 12308 3544 12314 3556
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 14568 3593 14596 3624
rect 14826 3612 14832 3664
rect 14884 3652 14890 3664
rect 15013 3655 15071 3661
rect 15013 3652 15025 3655
rect 14884 3624 15025 3652
rect 14884 3612 14890 3624
rect 15013 3621 15025 3624
rect 15059 3621 15071 3655
rect 15013 3615 15071 3621
rect 14553 3587 14611 3593
rect 14553 3553 14565 3587
rect 14599 3553 14611 3587
rect 15102 3584 15108 3596
rect 14553 3547 14611 3553
rect 14660 3556 15108 3584
rect 12342 3516 12348 3528
rect 10735 3488 11560 3516
rect 12303 3488 12348 3516
rect 10735 3485 10747 3488
rect 10689 3479 10747 3485
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 14182 3476 14188 3528
rect 14240 3516 14246 3528
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 14240 3488 14381 3516
rect 14240 3476 14246 3488
rect 14369 3485 14381 3488
rect 14415 3516 14427 3519
rect 14660 3516 14688 3556
rect 15102 3544 15108 3556
rect 15160 3584 15166 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 15160 3556 15301 3584
rect 15160 3544 15166 3556
rect 15289 3553 15301 3556
rect 15335 3584 15347 3587
rect 18874 3584 18880 3596
rect 15335 3556 18880 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 18874 3544 18880 3556
rect 18932 3544 18938 3596
rect 14415 3488 14688 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 15378 3476 15384 3528
rect 15436 3525 15442 3528
rect 15436 3519 15464 3525
rect 15452 3485 15464 3519
rect 15562 3516 15568 3528
rect 15523 3488 15568 3516
rect 15436 3479 15464 3485
rect 15436 3476 15442 3479
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 29822 3516 29828 3528
rect 29783 3488 29828 3516
rect 29822 3476 29828 3488
rect 29880 3476 29886 3528
rect 12342 3340 12348 3392
rect 12400 3380 12406 3392
rect 12894 3380 12900 3392
rect 12400 3352 12900 3380
rect 12400 3340 12406 3352
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 21450 3340 21456 3392
rect 21508 3380 21514 3392
rect 30009 3383 30067 3389
rect 30009 3380 30021 3383
rect 21508 3352 30021 3380
rect 21508 3340 21514 3352
rect 30009 3349 30021 3352
rect 30055 3349 30067 3383
rect 30009 3343 30067 3349
rect 1104 3290 30820 3312
rect 1104 3238 10880 3290
rect 10932 3238 10944 3290
rect 10996 3238 11008 3290
rect 11060 3238 11072 3290
rect 11124 3238 11136 3290
rect 11188 3238 20811 3290
rect 20863 3238 20875 3290
rect 20927 3238 20939 3290
rect 20991 3238 21003 3290
rect 21055 3238 21067 3290
rect 21119 3238 30820 3290
rect 1104 3216 30820 3238
rect 12434 3176 12440 3188
rect 11716 3148 12440 3176
rect 1397 3043 1455 3049
rect 1397 3009 1409 3043
rect 1443 3040 1455 3043
rect 1670 3040 1676 3052
rect 1443 3012 1676 3040
rect 1443 3009 1455 3012
rect 1397 3003 1455 3009
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 11716 3049 11744 3148
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 13170 3136 13176 3188
rect 13228 3176 13234 3188
rect 13357 3179 13415 3185
rect 13357 3176 13369 3179
rect 13228 3148 13369 3176
rect 13228 3136 13234 3148
rect 13357 3145 13369 3148
rect 13403 3145 13415 3179
rect 15470 3176 15476 3188
rect 13357 3139 13415 3145
rect 13832 3148 15476 3176
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11296 3012 11529 3040
rect 11296 3000 11302 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 12526 3000 12532 3052
rect 12584 3049 12590 3052
rect 12584 3043 12612 3049
rect 12600 3009 12612 3043
rect 12584 3003 12612 3009
rect 12584 3000 12590 3003
rect 11606 2932 11612 2984
rect 11664 2972 11670 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 11664 2944 12449 2972
rect 11664 2932 11670 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12713 2975 12771 2981
rect 12713 2941 12725 2975
rect 12759 2972 12771 2975
rect 12894 2972 12900 2984
rect 12759 2944 12900 2972
rect 12759 2941 12771 2944
rect 12713 2935 12771 2941
rect 12894 2932 12900 2944
rect 12952 2972 12958 2984
rect 13832 2972 13860 3148
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 16117 3179 16175 3185
rect 16117 3145 16129 3179
rect 16163 3176 16175 3179
rect 17126 3176 17132 3188
rect 16163 3148 17132 3176
rect 16163 3145 16175 3148
rect 16117 3139 16175 3145
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 29086 3136 29092 3188
rect 29144 3176 29150 3188
rect 29825 3179 29883 3185
rect 29825 3176 29837 3179
rect 29144 3148 29837 3176
rect 29144 3136 29150 3148
rect 29825 3145 29837 3148
rect 29871 3145 29883 3179
rect 29825 3139 29883 3145
rect 14182 3000 14188 3052
rect 14240 3040 14246 3052
rect 14277 3043 14335 3049
rect 14277 3040 14289 3043
rect 14240 3012 14289 3040
rect 14240 3000 14246 3012
rect 14277 3009 14289 3012
rect 14323 3009 14335 3043
rect 14277 3003 14335 3009
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 14461 3043 14519 3049
rect 14461 3040 14473 3043
rect 14424 3012 14473 3040
rect 14424 3000 14430 3012
rect 14461 3009 14473 3012
rect 14507 3009 14519 3043
rect 14461 3003 14519 3009
rect 15194 3000 15200 3052
rect 15252 3040 15258 3052
rect 15378 3049 15384 3052
rect 15335 3043 15384 3049
rect 15252 3012 15297 3040
rect 15252 3000 15258 3012
rect 15335 3009 15347 3043
rect 15381 3009 15384 3043
rect 15335 3003 15384 3009
rect 15378 3000 15384 3003
rect 15436 3000 15442 3052
rect 29733 3043 29791 3049
rect 29733 3009 29745 3043
rect 29779 3040 29791 3043
rect 29914 3040 29920 3052
rect 29779 3012 29920 3040
rect 29779 3009 29791 3012
rect 29733 3003 29791 3009
rect 29914 3000 29920 3012
rect 29972 3000 29978 3052
rect 12952 2944 13860 2972
rect 12952 2932 12958 2944
rect 15470 2932 15476 2984
rect 15528 2972 15534 2984
rect 15528 2944 15573 2972
rect 15528 2932 15534 2944
rect 1578 2904 1584 2916
rect 1539 2876 1584 2904
rect 1578 2864 1584 2876
rect 1636 2864 1642 2916
rect 12158 2904 12164 2916
rect 12119 2876 12164 2904
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 14921 2907 14979 2913
rect 14921 2873 14933 2907
rect 14967 2873 14979 2907
rect 14921 2867 14979 2873
rect 12176 2836 12204 2864
rect 14936 2836 14964 2867
rect 12176 2808 14964 2836
rect 1104 2746 30820 2768
rect 1104 2694 5915 2746
rect 5967 2694 5979 2746
rect 6031 2694 6043 2746
rect 6095 2694 6107 2746
rect 6159 2694 6171 2746
rect 6223 2694 15846 2746
rect 15898 2694 15910 2746
rect 15962 2694 15974 2746
rect 16026 2694 16038 2746
rect 16090 2694 16102 2746
rect 16154 2694 25776 2746
rect 25828 2694 25840 2746
rect 25892 2694 25904 2746
rect 25956 2694 25968 2746
rect 26020 2694 26032 2746
rect 26084 2694 30820 2746
rect 1104 2672 30820 2694
rect 13262 2632 13268 2644
rect 13223 2604 13268 2632
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 14093 2635 14151 2641
rect 14093 2601 14105 2635
rect 14139 2632 14151 2635
rect 14734 2632 14740 2644
rect 14139 2604 14740 2632
rect 14139 2601 14151 2604
rect 14093 2595 14151 2601
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 20162 2592 20168 2644
rect 20220 2632 20226 2644
rect 28905 2635 28963 2641
rect 28905 2632 28917 2635
rect 20220 2604 28917 2632
rect 20220 2592 20226 2604
rect 28905 2601 28917 2604
rect 28951 2601 28963 2635
rect 28905 2595 28963 2601
rect 28994 2592 29000 2644
rect 29052 2632 29058 2644
rect 29825 2635 29883 2641
rect 29825 2632 29837 2635
rect 29052 2604 29837 2632
rect 29052 2592 29058 2604
rect 29825 2601 29837 2604
rect 29871 2601 29883 2635
rect 29825 2595 29883 2601
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2428 1455 2431
rect 9490 2428 9496 2440
rect 1443 2400 9496 2428
rect 1443 2397 1455 2400
rect 1397 2391 1455 2397
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12492 2400 12909 2428
rect 12492 2388 12498 2400
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2428 13139 2431
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13127 2400 14105 2428
rect 13127 2397 13139 2400
rect 13081 2391 13139 2397
rect 14093 2397 14105 2400
rect 14139 2428 14151 2431
rect 14182 2428 14188 2440
rect 14139 2400 14188 2428
rect 14139 2397 14151 2400
rect 14093 2391 14151 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2428 14335 2431
rect 14366 2428 14372 2440
rect 14323 2400 14372 2428
rect 14323 2397 14335 2400
rect 14277 2391 14335 2397
rect 14366 2388 14372 2400
rect 14424 2388 14430 2440
rect 28718 2428 28724 2440
rect 28679 2400 28724 2428
rect 28718 2388 28724 2400
rect 28776 2388 28782 2440
rect 29730 2360 29736 2372
rect 29691 2332 29736 2360
rect 29730 2320 29736 2332
rect 29788 2320 29794 2372
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 1104 2202 30820 2224
rect 1104 2150 10880 2202
rect 10932 2150 10944 2202
rect 10996 2150 11008 2202
rect 11060 2150 11072 2202
rect 11124 2150 11136 2202
rect 11188 2150 20811 2202
rect 20863 2150 20875 2202
rect 20927 2150 20939 2202
rect 20991 2150 21003 2202
rect 21055 2150 21067 2202
rect 21119 2150 30820 2202
rect 1104 2128 30820 2150
<< via1 >>
rect 14188 45772 14240 45824
rect 15568 45772 15620 45824
rect 23296 45772 23348 45824
rect 27068 45772 27120 45824
rect 10880 45670 10932 45722
rect 10944 45670 10996 45722
rect 11008 45670 11060 45722
rect 11072 45670 11124 45722
rect 11136 45670 11188 45722
rect 20811 45670 20863 45722
rect 20875 45670 20927 45722
rect 20939 45670 20991 45722
rect 21003 45670 21055 45722
rect 21067 45670 21119 45722
rect 16672 45568 16724 45620
rect 17500 45568 17552 45620
rect 23848 45568 23900 45620
rect 30012 45611 30064 45620
rect 30012 45577 30021 45611
rect 30021 45577 30055 45611
rect 30055 45577 30064 45611
rect 30012 45568 30064 45577
rect 1584 45475 1636 45484
rect 1584 45441 1593 45475
rect 1593 45441 1627 45475
rect 1627 45441 1636 45475
rect 1584 45432 1636 45441
rect 2596 45432 2648 45484
rect 3424 45432 3476 45484
rect 4160 45432 4212 45484
rect 5724 45432 5776 45484
rect 6920 45432 6972 45484
rect 2688 45407 2740 45416
rect 2688 45373 2697 45407
rect 2697 45373 2731 45407
rect 2731 45373 2740 45407
rect 2688 45364 2740 45373
rect 5356 45407 5408 45416
rect 5356 45373 5365 45407
rect 5365 45373 5399 45407
rect 5399 45373 5408 45407
rect 5356 45364 5408 45373
rect 7932 45432 7984 45484
rect 8760 45432 8812 45484
rect 8852 45364 8904 45416
rect 8944 45296 8996 45348
rect 9496 45432 9548 45484
rect 11244 45432 11296 45484
rect 13452 45432 13504 45484
rect 13820 45432 13872 45484
rect 16396 45500 16448 45552
rect 15292 45475 15344 45484
rect 15292 45441 15301 45475
rect 15301 45441 15335 45475
rect 15335 45441 15344 45475
rect 15292 45432 15344 45441
rect 20996 45500 21048 45552
rect 16948 45475 17000 45484
rect 16948 45441 16957 45475
rect 16957 45441 16991 45475
rect 16991 45441 17000 45475
rect 16948 45432 17000 45441
rect 18420 45475 18472 45484
rect 16672 45364 16724 45416
rect 17408 45364 17460 45416
rect 1400 45271 1452 45280
rect 1400 45237 1409 45271
rect 1409 45237 1443 45271
rect 1443 45237 1452 45271
rect 1400 45228 1452 45237
rect 7012 45271 7064 45280
rect 7012 45237 7021 45271
rect 7021 45237 7055 45271
rect 7055 45237 7064 45271
rect 7012 45228 7064 45237
rect 9864 45228 9916 45280
rect 11704 45271 11756 45280
rect 11704 45237 11713 45271
rect 11713 45237 11747 45271
rect 11747 45237 11756 45271
rect 11704 45228 11756 45237
rect 16580 45296 16632 45348
rect 18420 45441 18429 45475
rect 18429 45441 18463 45475
rect 18463 45441 18472 45475
rect 18420 45432 18472 45441
rect 18512 45432 18564 45484
rect 20536 45432 20588 45484
rect 21088 45432 21140 45484
rect 21456 45500 21508 45552
rect 21732 45432 21784 45484
rect 23848 45475 23900 45484
rect 23848 45441 23857 45475
rect 23857 45441 23891 45475
rect 23891 45441 23900 45475
rect 26148 45475 26200 45484
rect 23848 45432 23900 45441
rect 26148 45441 26157 45475
rect 26157 45441 26191 45475
rect 26191 45441 26200 45475
rect 26148 45432 26200 45441
rect 27436 45475 27488 45484
rect 27436 45441 27445 45475
rect 27445 45441 27479 45475
rect 27479 45441 27488 45475
rect 27436 45432 27488 45441
rect 27620 45432 27672 45484
rect 19340 45407 19392 45416
rect 19340 45373 19349 45407
rect 19349 45373 19383 45407
rect 19383 45373 19392 45407
rect 19340 45364 19392 45373
rect 20444 45364 20496 45416
rect 23204 45364 23256 45416
rect 27528 45407 27580 45416
rect 14280 45228 14332 45280
rect 14464 45271 14516 45280
rect 14464 45237 14473 45271
rect 14473 45237 14507 45271
rect 14507 45237 14516 45271
rect 14464 45228 14516 45237
rect 15108 45271 15160 45280
rect 15108 45237 15117 45271
rect 15117 45237 15151 45271
rect 15151 45237 15160 45271
rect 15108 45228 15160 45237
rect 15200 45228 15252 45280
rect 15660 45228 15712 45280
rect 27528 45373 27537 45407
rect 27537 45373 27571 45407
rect 27571 45373 27580 45407
rect 27528 45364 27580 45373
rect 17040 45228 17092 45280
rect 17592 45228 17644 45280
rect 19432 45228 19484 45280
rect 19616 45271 19668 45280
rect 19616 45237 19625 45271
rect 19625 45237 19659 45271
rect 19659 45237 19668 45271
rect 19616 45228 19668 45237
rect 20628 45228 20680 45280
rect 20996 45228 21048 45280
rect 27712 45296 27764 45348
rect 28540 45475 28592 45484
rect 28540 45441 28549 45475
rect 28549 45441 28583 45475
rect 28583 45441 28592 45475
rect 28540 45432 28592 45441
rect 29184 45432 29236 45484
rect 27160 45228 27212 45280
rect 27252 45228 27304 45280
rect 27528 45228 27580 45280
rect 5915 45126 5967 45178
rect 5979 45126 6031 45178
rect 6043 45126 6095 45178
rect 6107 45126 6159 45178
rect 6171 45126 6223 45178
rect 15846 45126 15898 45178
rect 15910 45126 15962 45178
rect 15974 45126 16026 45178
rect 16038 45126 16090 45178
rect 16102 45126 16154 45178
rect 25776 45126 25828 45178
rect 25840 45126 25892 45178
rect 25904 45126 25956 45178
rect 25968 45126 26020 45178
rect 26032 45126 26084 45178
rect 8944 45024 8996 45076
rect 9772 44956 9824 45008
rect 1400 44888 1452 44940
rect 11244 44888 11296 44940
rect 13912 45024 13964 45076
rect 14740 45024 14792 45076
rect 15016 45024 15068 45076
rect 16580 45067 16632 45076
rect 16580 45033 16589 45067
rect 16589 45033 16623 45067
rect 16623 45033 16632 45067
rect 16580 45024 16632 45033
rect 16948 45024 17000 45076
rect 20720 45067 20772 45076
rect 20720 45033 20729 45067
rect 20729 45033 20763 45067
rect 20763 45033 20772 45067
rect 20720 45024 20772 45033
rect 21088 45024 21140 45076
rect 14372 44956 14424 45008
rect 14464 44956 14516 45008
rect 1860 44820 1912 44872
rect 4896 44820 4948 44872
rect 7196 44820 7248 44872
rect 10232 44820 10284 44872
rect 11796 44820 11848 44872
rect 12532 44820 12584 44872
rect 13544 44863 13596 44872
rect 13544 44829 13553 44863
rect 13553 44829 13587 44863
rect 13587 44829 13596 44863
rect 13544 44820 13596 44829
rect 14740 44863 14792 44872
rect 14740 44829 14749 44863
rect 14749 44829 14783 44863
rect 14783 44829 14792 44863
rect 14740 44820 14792 44829
rect 14924 44863 14976 44872
rect 14924 44829 14933 44863
rect 14933 44829 14967 44863
rect 14967 44829 14976 44863
rect 14924 44820 14976 44829
rect 16212 44888 16264 44940
rect 15752 44863 15804 44872
rect 2412 44795 2464 44804
rect 2412 44761 2421 44795
rect 2421 44761 2455 44795
rect 2455 44761 2464 44795
rect 2412 44752 2464 44761
rect 5172 44727 5224 44736
rect 5172 44693 5181 44727
rect 5181 44693 5215 44727
rect 5215 44693 5224 44727
rect 5172 44684 5224 44693
rect 10048 44684 10100 44736
rect 14648 44752 14700 44804
rect 13452 44684 13504 44736
rect 14464 44684 14516 44736
rect 14924 44684 14976 44736
rect 15292 44752 15344 44804
rect 15752 44829 15761 44863
rect 15761 44829 15795 44863
rect 15795 44829 15804 44863
rect 15752 44820 15804 44829
rect 19248 44956 19300 45008
rect 22192 44956 22244 45008
rect 22376 45024 22428 45076
rect 27528 45024 27580 45076
rect 28264 45067 28316 45076
rect 28264 45033 28273 45067
rect 28273 45033 28307 45067
rect 28307 45033 28316 45067
rect 28264 45024 28316 45033
rect 17224 44888 17276 44940
rect 18420 44888 18472 44940
rect 19984 44888 20036 44940
rect 16856 44863 16908 44872
rect 16856 44829 16865 44863
rect 16865 44829 16899 44863
rect 16899 44829 16908 44863
rect 16856 44820 16908 44829
rect 17316 44752 17368 44804
rect 17776 44820 17828 44872
rect 18052 44820 18104 44872
rect 19892 44863 19944 44872
rect 19892 44829 19901 44863
rect 19901 44829 19935 44863
rect 19935 44829 19944 44863
rect 19892 44820 19944 44829
rect 21456 44888 21508 44940
rect 20996 44863 21048 44872
rect 20996 44829 21005 44863
rect 21005 44829 21039 44863
rect 21039 44829 21048 44863
rect 20996 44820 21048 44829
rect 21456 44752 21508 44804
rect 21640 44752 21692 44804
rect 22376 44888 22428 44940
rect 22468 44888 22520 44940
rect 23940 44888 23992 44940
rect 21916 44863 21968 44872
rect 21916 44829 21917 44863
rect 21917 44829 21951 44863
rect 21951 44829 21968 44863
rect 22836 44863 22888 44872
rect 21916 44820 21968 44829
rect 22836 44829 22845 44863
rect 22845 44829 22879 44863
rect 22879 44829 22888 44863
rect 22836 44820 22888 44829
rect 22192 44752 22244 44804
rect 25044 44820 25096 44872
rect 27160 44888 27212 44940
rect 28080 44820 28132 44872
rect 26332 44752 26384 44804
rect 16672 44684 16724 44736
rect 17868 44684 17920 44736
rect 19340 44684 19392 44736
rect 20076 44727 20128 44736
rect 20076 44693 20085 44727
rect 20085 44693 20119 44727
rect 20119 44693 20128 44727
rect 20076 44684 20128 44693
rect 21272 44727 21324 44736
rect 21272 44693 21281 44727
rect 21281 44693 21315 44727
rect 21315 44693 21324 44727
rect 21272 44684 21324 44693
rect 22100 44684 22152 44736
rect 25320 44684 25372 44736
rect 26792 44684 26844 44736
rect 27528 44684 27580 44736
rect 30012 44727 30064 44736
rect 30012 44693 30021 44727
rect 30021 44693 30055 44727
rect 30055 44693 30064 44727
rect 30012 44684 30064 44693
rect 10880 44582 10932 44634
rect 10944 44582 10996 44634
rect 11008 44582 11060 44634
rect 11072 44582 11124 44634
rect 11136 44582 11188 44634
rect 20811 44582 20863 44634
rect 20875 44582 20927 44634
rect 20939 44582 20991 44634
rect 21003 44582 21055 44634
rect 21067 44582 21119 44634
rect 5172 44480 5224 44532
rect 12624 44480 12676 44532
rect 2780 44412 2832 44464
rect 2044 44387 2096 44396
rect 2044 44353 2053 44387
rect 2053 44353 2087 44387
rect 2087 44353 2096 44387
rect 2044 44344 2096 44353
rect 2412 44344 2464 44396
rect 2596 44319 2648 44328
rect 2596 44285 2605 44319
rect 2605 44285 2639 44319
rect 2639 44285 2648 44319
rect 2596 44276 2648 44285
rect 2688 44276 2740 44328
rect 15660 44480 15712 44532
rect 14924 44455 14976 44464
rect 14924 44421 14933 44455
rect 14933 44421 14967 44455
rect 14967 44421 14976 44455
rect 14924 44412 14976 44421
rect 17500 44480 17552 44532
rect 17868 44455 17920 44464
rect 17868 44421 17877 44455
rect 17877 44421 17911 44455
rect 17911 44421 17920 44455
rect 17868 44412 17920 44421
rect 18512 44412 18564 44464
rect 18696 44412 18748 44464
rect 14004 44344 14056 44396
rect 14188 44344 14240 44396
rect 16396 44344 16448 44396
rect 16488 44344 16540 44396
rect 15016 44319 15068 44328
rect 15016 44285 15025 44319
rect 15025 44285 15059 44319
rect 15059 44285 15068 44319
rect 15016 44276 15068 44285
rect 15200 44319 15252 44328
rect 15200 44285 15209 44319
rect 15209 44285 15243 44319
rect 15243 44285 15252 44319
rect 15200 44276 15252 44285
rect 16764 44276 16816 44328
rect 16948 44276 17000 44328
rect 19340 44344 19392 44396
rect 19708 44344 19760 44396
rect 19432 44319 19484 44328
rect 10876 44208 10928 44260
rect 18696 44208 18748 44260
rect 19432 44285 19441 44319
rect 19441 44285 19475 44319
rect 19475 44285 19484 44319
rect 19432 44276 19484 44285
rect 19892 44412 19944 44464
rect 20260 44387 20312 44396
rect 20260 44353 20269 44387
rect 20269 44353 20303 44387
rect 20303 44353 20312 44387
rect 20260 44344 20312 44353
rect 20352 44276 20404 44328
rect 21180 44344 21232 44396
rect 21640 44344 21692 44396
rect 22008 44387 22060 44396
rect 22008 44353 22017 44387
rect 22017 44353 22051 44387
rect 22051 44353 22060 44387
rect 22008 44344 22060 44353
rect 22928 44387 22980 44396
rect 22928 44353 22937 44387
rect 22937 44353 22971 44387
rect 22971 44353 22980 44387
rect 22928 44344 22980 44353
rect 20812 44276 20864 44328
rect 21732 44276 21784 44328
rect 22100 44276 22152 44328
rect 23388 44276 23440 44328
rect 23572 44319 23624 44328
rect 23572 44285 23581 44319
rect 23581 44285 23615 44319
rect 23615 44285 23624 44319
rect 23572 44276 23624 44285
rect 24860 44344 24912 44396
rect 25688 44387 25740 44396
rect 25688 44353 25697 44387
rect 25697 44353 25731 44387
rect 25731 44353 25740 44387
rect 25688 44344 25740 44353
rect 27528 44480 27580 44532
rect 28448 44523 28500 44532
rect 28448 44489 28457 44523
rect 28457 44489 28491 44523
rect 28491 44489 28500 44523
rect 28448 44480 28500 44489
rect 28540 44480 28592 44532
rect 27896 44412 27948 44464
rect 29552 44387 29604 44396
rect 29552 44353 29561 44387
rect 29561 44353 29595 44387
rect 29595 44353 29604 44387
rect 29552 44344 29604 44353
rect 29920 44387 29972 44396
rect 29920 44353 29929 44387
rect 29929 44353 29963 44387
rect 29963 44353 29972 44387
rect 29920 44344 29972 44353
rect 25136 44276 25188 44328
rect 14188 44140 14240 44192
rect 14740 44140 14792 44192
rect 16304 44140 16356 44192
rect 17316 44140 17368 44192
rect 17960 44140 18012 44192
rect 18972 44140 19024 44192
rect 20444 44183 20496 44192
rect 20444 44149 20453 44183
rect 20453 44149 20487 44183
rect 20487 44149 20496 44183
rect 20444 44140 20496 44149
rect 20720 44140 20772 44192
rect 21732 44140 21784 44192
rect 22836 44140 22888 44192
rect 23112 44183 23164 44192
rect 23112 44149 23121 44183
rect 23121 44149 23155 44183
rect 23155 44149 23164 44183
rect 23112 44140 23164 44149
rect 28080 44208 28132 44260
rect 24952 44183 25004 44192
rect 24952 44149 24961 44183
rect 24961 44149 24995 44183
rect 24995 44149 25004 44183
rect 24952 44140 25004 44149
rect 25228 44140 25280 44192
rect 29000 44208 29052 44260
rect 28264 44183 28316 44192
rect 28264 44149 28273 44183
rect 28273 44149 28307 44183
rect 28307 44149 28316 44183
rect 28264 44140 28316 44149
rect 29644 44140 29696 44192
rect 31576 44115 31628 44124
rect 5915 44038 5967 44090
rect 5979 44038 6031 44090
rect 6043 44038 6095 44090
rect 6107 44038 6159 44090
rect 6171 44038 6223 44090
rect 15846 44038 15898 44090
rect 15910 44038 15962 44090
rect 15974 44038 16026 44090
rect 16038 44038 16090 44090
rect 16102 44038 16154 44090
rect 25776 44038 25828 44090
rect 25840 44038 25892 44090
rect 25904 44038 25956 44090
rect 25968 44038 26020 44090
rect 26032 44038 26084 44090
rect 31576 44081 31585 44115
rect 31585 44081 31619 44115
rect 31619 44081 31628 44115
rect 31576 44072 31628 44081
rect 2044 43936 2096 43988
rect 13820 43936 13872 43988
rect 18604 43936 18656 43988
rect 19432 43979 19484 43988
rect 19432 43945 19441 43979
rect 19441 43945 19475 43979
rect 19475 43945 19484 43979
rect 19432 43936 19484 43945
rect 20444 43979 20496 43988
rect 20444 43945 20453 43979
rect 20453 43945 20487 43979
rect 20487 43945 20496 43979
rect 20444 43936 20496 43945
rect 23572 43936 23624 43988
rect 23664 43936 23716 43988
rect 28264 43979 28316 43988
rect 10876 43843 10928 43852
rect 10876 43809 10885 43843
rect 10885 43809 10919 43843
rect 10919 43809 10928 43843
rect 10876 43800 10928 43809
rect 11244 43800 11296 43852
rect 22836 43868 22888 43920
rect 25136 43911 25188 43920
rect 14464 43800 14516 43852
rect 15016 43800 15068 43852
rect 15200 43800 15252 43852
rect 388 43732 440 43784
rect 11336 43732 11388 43784
rect 13268 43732 13320 43784
rect 13544 43732 13596 43784
rect 15752 43732 15804 43784
rect 14188 43664 14240 43716
rect 14924 43664 14976 43716
rect 15476 43664 15528 43716
rect 16212 43800 16264 43852
rect 16580 43800 16632 43852
rect 17408 43843 17460 43852
rect 17408 43809 17417 43843
rect 17417 43809 17451 43843
rect 17451 43809 17460 43843
rect 17408 43800 17460 43809
rect 19340 43843 19392 43852
rect 19340 43809 19349 43843
rect 19349 43809 19383 43843
rect 19383 43809 19392 43843
rect 19340 43800 19392 43809
rect 16488 43732 16540 43784
rect 16948 43732 17000 43784
rect 17592 43732 17644 43784
rect 20076 43732 20128 43784
rect 22652 43800 22704 43852
rect 20352 43775 20404 43784
rect 20352 43741 20361 43775
rect 20361 43741 20395 43775
rect 20395 43741 20404 43775
rect 20352 43732 20404 43741
rect 20812 43732 20864 43784
rect 21088 43775 21140 43784
rect 21088 43741 21097 43775
rect 21097 43741 21131 43775
rect 21131 43741 21140 43775
rect 21088 43732 21140 43741
rect 21272 43775 21324 43784
rect 21272 43741 21281 43775
rect 21281 43741 21315 43775
rect 21315 43741 21324 43775
rect 21272 43732 21324 43741
rect 22468 43775 22520 43784
rect 22468 43741 22477 43775
rect 22477 43741 22511 43775
rect 22511 43741 22520 43775
rect 22468 43732 22520 43741
rect 22560 43732 22612 43784
rect 23204 43732 23256 43784
rect 23572 43732 23624 43784
rect 24492 43800 24544 43852
rect 25136 43877 25145 43911
rect 25145 43877 25179 43911
rect 25179 43877 25188 43911
rect 25136 43868 25188 43877
rect 25412 43800 25464 43852
rect 25872 43800 25924 43852
rect 28264 43945 28273 43979
rect 28273 43945 28307 43979
rect 28307 43945 28316 43979
rect 28264 43936 28316 43945
rect 30840 43936 30892 43988
rect 30012 43911 30064 43920
rect 30012 43877 30021 43911
rect 30021 43877 30055 43911
rect 30055 43877 30064 43911
rect 30012 43868 30064 43877
rect 29092 43800 29144 43852
rect 24400 43775 24452 43784
rect 24400 43741 24409 43775
rect 24409 43741 24443 43775
rect 24443 43741 24452 43775
rect 24400 43732 24452 43741
rect 24584 43773 24636 43784
rect 24584 43739 24615 43773
rect 24615 43739 24636 43773
rect 24584 43732 24636 43739
rect 24676 43775 24728 43784
rect 24676 43741 24685 43775
rect 24685 43741 24719 43775
rect 24719 43741 24728 43775
rect 24952 43775 25004 43784
rect 24676 43732 24728 43741
rect 24952 43741 24961 43775
rect 24961 43741 24995 43775
rect 24995 43741 25004 43775
rect 24952 43732 25004 43741
rect 26056 43732 26108 43784
rect 11244 43639 11296 43648
rect 11244 43605 11253 43639
rect 11253 43605 11287 43639
rect 11287 43605 11296 43639
rect 11244 43596 11296 43605
rect 14464 43596 14516 43648
rect 14556 43596 14608 43648
rect 15384 43596 15436 43648
rect 16212 43639 16264 43648
rect 16212 43605 16221 43639
rect 16221 43605 16255 43639
rect 16255 43605 16264 43639
rect 16212 43596 16264 43605
rect 16396 43596 16448 43648
rect 17592 43596 17644 43648
rect 18788 43596 18840 43648
rect 20260 43664 20312 43716
rect 20628 43664 20680 43716
rect 24124 43664 24176 43716
rect 24308 43664 24360 43716
rect 27068 43732 27120 43784
rect 28080 43732 28132 43784
rect 29000 43732 29052 43784
rect 26240 43707 26292 43716
rect 26240 43673 26274 43707
rect 26274 43673 26292 43707
rect 26240 43664 26292 43673
rect 19984 43596 20036 43648
rect 22376 43596 22428 43648
rect 23388 43596 23440 43648
rect 23848 43639 23900 43648
rect 23848 43605 23857 43639
rect 23857 43605 23891 43639
rect 23891 43605 23900 43639
rect 23848 43596 23900 43605
rect 23940 43596 23992 43648
rect 26608 43596 26660 43648
rect 10880 43494 10932 43546
rect 10944 43494 10996 43546
rect 11008 43494 11060 43546
rect 11072 43494 11124 43546
rect 11136 43494 11188 43546
rect 20811 43494 20863 43546
rect 20875 43494 20927 43546
rect 20939 43494 20991 43546
rect 21003 43494 21055 43546
rect 21067 43494 21119 43546
rect 13544 43392 13596 43444
rect 14188 43435 14240 43444
rect 14188 43401 14197 43435
rect 14197 43401 14231 43435
rect 14231 43401 14240 43435
rect 14188 43392 14240 43401
rect 15108 43392 15160 43444
rect 15292 43435 15344 43444
rect 15292 43401 15301 43435
rect 15301 43401 15335 43435
rect 15335 43401 15344 43435
rect 16764 43435 16816 43444
rect 15292 43392 15344 43401
rect 16764 43401 16773 43435
rect 16773 43401 16807 43435
rect 16807 43401 16816 43435
rect 16764 43392 16816 43401
rect 17592 43392 17644 43444
rect 1584 43299 1636 43308
rect 1584 43265 1593 43299
rect 1593 43265 1627 43299
rect 1627 43265 1636 43299
rect 1584 43256 1636 43265
rect 14832 43324 14884 43376
rect 17224 43324 17276 43376
rect 19524 43324 19576 43376
rect 14096 43256 14148 43308
rect 17132 43256 17184 43308
rect 15200 43188 15252 43240
rect 17040 43188 17092 43240
rect 17960 43256 18012 43308
rect 18144 43256 18196 43308
rect 19616 43299 19668 43308
rect 19616 43265 19625 43299
rect 19625 43265 19659 43299
rect 19659 43265 19668 43299
rect 19616 43256 19668 43265
rect 17408 43231 17460 43240
rect 17408 43197 17417 43231
rect 17417 43197 17451 43231
rect 17451 43197 17460 43231
rect 17408 43188 17460 43197
rect 18604 43188 18656 43240
rect 21180 43392 21232 43444
rect 22468 43392 22520 43444
rect 23204 43392 23256 43444
rect 24400 43392 24452 43444
rect 24492 43392 24544 43444
rect 25320 43392 25372 43444
rect 26332 43392 26384 43444
rect 26516 43392 26568 43444
rect 21180 43256 21232 43308
rect 22192 43256 22244 43308
rect 22744 43299 22796 43308
rect 11244 43120 11296 43172
rect 21916 43188 21968 43240
rect 22744 43265 22753 43299
rect 22753 43265 22787 43299
rect 22787 43265 22796 43299
rect 22744 43256 22796 43265
rect 23112 43256 23164 43308
rect 23480 43256 23532 43308
rect 23848 43324 23900 43376
rect 24952 43324 25004 43376
rect 28908 43392 28960 43444
rect 10876 43052 10928 43104
rect 14924 43052 14976 43104
rect 15016 43052 15068 43104
rect 18512 43052 18564 43104
rect 18696 43095 18748 43104
rect 18696 43061 18705 43095
rect 18705 43061 18739 43095
rect 18739 43061 18748 43095
rect 18696 43052 18748 43061
rect 19064 43095 19116 43104
rect 19064 43061 19073 43095
rect 19073 43061 19107 43095
rect 19107 43061 19116 43095
rect 19064 43052 19116 43061
rect 19708 43095 19760 43104
rect 19708 43061 19717 43095
rect 19717 43061 19751 43095
rect 19751 43061 19760 43095
rect 19708 43052 19760 43061
rect 20720 43120 20772 43172
rect 23388 43120 23440 43172
rect 25320 43256 25372 43308
rect 25688 43299 25740 43308
rect 25688 43265 25697 43299
rect 25697 43265 25731 43299
rect 25731 43265 25740 43299
rect 25688 43256 25740 43265
rect 25872 43299 25924 43308
rect 25872 43265 25881 43299
rect 25881 43265 25915 43299
rect 25915 43265 25924 43299
rect 25872 43256 25924 43265
rect 26792 43256 26844 43308
rect 26976 43299 27028 43308
rect 26976 43265 26985 43299
rect 26985 43265 27019 43299
rect 27019 43265 27028 43299
rect 26976 43256 27028 43265
rect 27068 43256 27120 43308
rect 25596 43188 25648 43240
rect 26332 43120 26384 43172
rect 27804 43120 27856 43172
rect 28080 43120 28132 43172
rect 20628 43095 20680 43104
rect 20628 43061 20637 43095
rect 20637 43061 20671 43095
rect 20671 43061 20680 43095
rect 22100 43095 22152 43104
rect 20628 43052 20680 43061
rect 22100 43061 22109 43095
rect 22109 43061 22143 43095
rect 22143 43061 22152 43095
rect 22100 43052 22152 43061
rect 22284 43052 22336 43104
rect 24584 43052 24636 43104
rect 25504 43052 25556 43104
rect 25688 43052 25740 43104
rect 27160 43095 27212 43104
rect 27160 43061 27169 43095
rect 27169 43061 27203 43095
rect 27203 43061 27212 43095
rect 27160 43052 27212 43061
rect 27712 43052 27764 43104
rect 28264 43095 28316 43104
rect 28264 43061 28273 43095
rect 28273 43061 28307 43095
rect 28307 43061 28316 43095
rect 28264 43052 28316 43061
rect 30012 43095 30064 43104
rect 30012 43061 30021 43095
rect 30021 43061 30055 43095
rect 30055 43061 30064 43095
rect 30012 43052 30064 43061
rect 5915 42950 5967 43002
rect 5979 42950 6031 43002
rect 6043 42950 6095 43002
rect 6107 42950 6159 43002
rect 6171 42950 6223 43002
rect 15846 42950 15898 43002
rect 15910 42950 15962 43002
rect 15974 42950 16026 43002
rect 16038 42950 16090 43002
rect 16102 42950 16154 43002
rect 25776 42950 25828 43002
rect 25840 42950 25892 43002
rect 25904 42950 25956 43002
rect 25968 42950 26020 43002
rect 26032 42950 26084 43002
rect 16212 42848 16264 42900
rect 17040 42848 17092 42900
rect 17408 42848 17460 42900
rect 17684 42780 17736 42832
rect 10876 42755 10928 42764
rect 10876 42721 10885 42755
rect 10885 42721 10919 42755
rect 10919 42721 10928 42755
rect 10876 42712 10928 42721
rect 15476 42755 15528 42764
rect 15476 42721 15485 42755
rect 15485 42721 15519 42755
rect 15519 42721 15528 42755
rect 15476 42712 15528 42721
rect 17316 42712 17368 42764
rect 17776 42755 17828 42764
rect 17776 42721 17785 42755
rect 17785 42721 17819 42755
rect 17819 42721 17828 42755
rect 17776 42712 17828 42721
rect 18420 42712 18472 42764
rect 11336 42644 11388 42696
rect 14464 42644 14516 42696
rect 15108 42644 15160 42696
rect 15752 42644 15804 42696
rect 15200 42576 15252 42628
rect 16488 42644 16540 42696
rect 19708 42848 19760 42900
rect 25136 42780 25188 42832
rect 25412 42780 25464 42832
rect 25872 42780 25924 42832
rect 25044 42712 25096 42764
rect 17040 42576 17092 42628
rect 20076 42644 20128 42696
rect 20628 42644 20680 42696
rect 22744 42687 22796 42696
rect 11244 42551 11296 42560
rect 11244 42517 11253 42551
rect 11253 42517 11287 42551
rect 11287 42517 11296 42551
rect 11244 42508 11296 42517
rect 14648 42508 14700 42560
rect 17224 42508 17276 42560
rect 17684 42551 17736 42560
rect 17684 42517 17693 42551
rect 17693 42517 17727 42551
rect 17727 42517 17736 42551
rect 17684 42508 17736 42517
rect 17776 42508 17828 42560
rect 19800 42551 19852 42560
rect 19800 42517 19809 42551
rect 19809 42517 19843 42551
rect 19843 42517 19852 42551
rect 19800 42508 19852 42517
rect 21180 42576 21232 42628
rect 22744 42653 22753 42687
rect 22753 42653 22787 42687
rect 22787 42653 22796 42687
rect 22744 42644 22796 42653
rect 27160 42712 27212 42764
rect 27436 42712 27488 42764
rect 25320 42644 25372 42696
rect 25596 42644 25648 42696
rect 22928 42551 22980 42560
rect 22928 42517 22937 42551
rect 22937 42517 22971 42551
rect 22971 42517 22980 42551
rect 22928 42508 22980 42517
rect 23388 42551 23440 42560
rect 23388 42517 23397 42551
rect 23397 42517 23431 42551
rect 23431 42517 23440 42551
rect 23388 42508 23440 42517
rect 24952 42576 25004 42628
rect 24676 42508 24728 42560
rect 24768 42508 24820 42560
rect 25688 42508 25740 42560
rect 25872 42687 25924 42696
rect 25872 42653 25881 42687
rect 25881 42653 25915 42687
rect 25915 42653 25924 42687
rect 25872 42644 25924 42653
rect 26240 42687 26292 42696
rect 26240 42653 26249 42687
rect 26249 42653 26283 42687
rect 26283 42653 26292 42687
rect 26700 42687 26752 42696
rect 26240 42644 26292 42653
rect 26700 42653 26709 42687
rect 26709 42653 26743 42687
rect 26743 42653 26752 42687
rect 26700 42644 26752 42653
rect 27344 42687 27396 42696
rect 27344 42653 27353 42687
rect 27353 42653 27387 42687
rect 27387 42653 27396 42687
rect 27344 42644 27396 42653
rect 28448 42644 28500 42696
rect 28908 42644 28960 42696
rect 26148 42576 26200 42628
rect 26608 42508 26660 42560
rect 27528 42551 27580 42560
rect 27528 42517 27537 42551
rect 27537 42517 27571 42551
rect 27571 42517 27580 42551
rect 27528 42508 27580 42517
rect 29736 42576 29788 42628
rect 28632 42551 28684 42560
rect 28632 42517 28641 42551
rect 28641 42517 28675 42551
rect 28675 42517 28684 42551
rect 28632 42508 28684 42517
rect 30012 42551 30064 42560
rect 30012 42517 30021 42551
rect 30021 42517 30055 42551
rect 30055 42517 30064 42551
rect 30012 42508 30064 42517
rect 10880 42406 10932 42458
rect 10944 42406 10996 42458
rect 11008 42406 11060 42458
rect 11072 42406 11124 42458
rect 11136 42406 11188 42458
rect 20811 42406 20863 42458
rect 20875 42406 20927 42458
rect 20939 42406 20991 42458
rect 21003 42406 21055 42458
rect 21067 42406 21119 42458
rect 17684 42304 17736 42356
rect 18512 42304 18564 42356
rect 19064 42304 19116 42356
rect 20628 42304 20680 42356
rect 21180 42347 21232 42356
rect 21180 42313 21189 42347
rect 21189 42313 21223 42347
rect 21223 42313 21232 42347
rect 21180 42304 21232 42313
rect 23848 42347 23900 42356
rect 23848 42313 23857 42347
rect 23857 42313 23891 42347
rect 23891 42313 23900 42347
rect 23848 42304 23900 42313
rect 26700 42304 26752 42356
rect 26792 42304 26844 42356
rect 11244 42236 11296 42288
rect 17408 42236 17460 42288
rect 14372 42168 14424 42220
rect 15016 42211 15068 42220
rect 15016 42177 15025 42211
rect 15025 42177 15059 42211
rect 15059 42177 15068 42211
rect 15016 42168 15068 42177
rect 15200 42211 15252 42220
rect 15200 42177 15209 42211
rect 15209 42177 15243 42211
rect 15243 42177 15252 42211
rect 15200 42168 15252 42177
rect 15108 42100 15160 42152
rect 17776 42168 17828 42220
rect 16948 42143 17000 42152
rect 16948 42109 16957 42143
rect 16957 42109 16991 42143
rect 16991 42109 17000 42143
rect 16948 42100 17000 42109
rect 17132 42100 17184 42152
rect 18604 42100 18656 42152
rect 19432 42236 19484 42288
rect 19708 42236 19760 42288
rect 19800 42236 19852 42288
rect 19524 42211 19576 42220
rect 19524 42177 19533 42211
rect 19533 42177 19567 42211
rect 19567 42177 19576 42211
rect 19524 42168 19576 42177
rect 18788 42100 18840 42152
rect 19340 42100 19392 42152
rect 19892 42168 19944 42220
rect 19984 42168 20036 42220
rect 20628 42211 20680 42220
rect 20628 42177 20637 42211
rect 20637 42177 20671 42211
rect 20671 42177 20680 42211
rect 20628 42168 20680 42177
rect 21272 42211 21324 42220
rect 21272 42177 21281 42211
rect 21281 42177 21315 42211
rect 21315 42177 21324 42211
rect 21272 42168 21324 42177
rect 22652 42236 22704 42288
rect 23020 42211 23072 42220
rect 23020 42177 23029 42211
rect 23029 42177 23063 42211
rect 23063 42177 23072 42211
rect 23388 42236 23440 42288
rect 24032 42211 24084 42220
rect 23020 42168 23072 42177
rect 24032 42177 24041 42211
rect 24041 42177 24075 42211
rect 24075 42177 24084 42211
rect 24032 42168 24084 42177
rect 24124 42168 24176 42220
rect 26976 42168 27028 42220
rect 21548 42100 21600 42152
rect 24216 42100 24268 42152
rect 24768 42143 24820 42152
rect 24768 42109 24777 42143
rect 24777 42109 24811 42143
rect 24811 42109 24820 42143
rect 24768 42100 24820 42109
rect 27436 42236 27488 42288
rect 27712 42236 27764 42288
rect 27988 42236 28040 42288
rect 28540 42211 28592 42220
rect 28540 42177 28549 42211
rect 28549 42177 28583 42211
rect 28583 42177 28592 42211
rect 28540 42168 28592 42177
rect 14832 42007 14884 42016
rect 14832 41973 14841 42007
rect 14841 41973 14875 42007
rect 14875 41973 14884 42007
rect 14832 41964 14884 41973
rect 18512 41964 18564 42016
rect 19892 42032 19944 42084
rect 26976 42032 27028 42084
rect 21088 41964 21140 42016
rect 25044 41964 25096 42016
rect 28264 41964 28316 42016
rect 28632 41964 28684 42016
rect 30012 42007 30064 42016
rect 30012 41973 30021 42007
rect 30021 41973 30055 42007
rect 30055 41973 30064 42007
rect 30012 41964 30064 41973
rect 5915 41862 5967 41914
rect 5979 41862 6031 41914
rect 6043 41862 6095 41914
rect 6107 41862 6159 41914
rect 6171 41862 6223 41914
rect 15846 41862 15898 41914
rect 15910 41862 15962 41914
rect 15974 41862 16026 41914
rect 16038 41862 16090 41914
rect 16102 41862 16154 41914
rect 25776 41862 25828 41914
rect 25840 41862 25892 41914
rect 25904 41862 25956 41914
rect 25968 41862 26020 41914
rect 26032 41862 26084 41914
rect 21272 41760 21324 41812
rect 27344 41760 27396 41812
rect 28632 41760 28684 41812
rect 28816 41803 28868 41812
rect 28816 41769 28825 41803
rect 28825 41769 28859 41803
rect 28859 41769 28868 41803
rect 28816 41760 28868 41769
rect 29092 41760 29144 41812
rect 16948 41692 17000 41744
rect 19984 41692 20036 41744
rect 21088 41692 21140 41744
rect 14464 41624 14516 41676
rect 15292 41624 15344 41676
rect 16488 41624 16540 41676
rect 14648 41599 14700 41608
rect 14648 41565 14657 41599
rect 14657 41565 14691 41599
rect 14691 41565 14700 41599
rect 14648 41556 14700 41565
rect 2596 41488 2648 41540
rect 17500 41599 17552 41608
rect 16672 41488 16724 41540
rect 17500 41565 17509 41599
rect 17509 41565 17543 41599
rect 17543 41565 17552 41599
rect 17500 41556 17552 41565
rect 20076 41667 20128 41676
rect 20076 41633 20085 41667
rect 20085 41633 20119 41667
rect 20119 41633 20128 41667
rect 20076 41624 20128 41633
rect 19064 41556 19116 41608
rect 23848 41624 23900 41676
rect 24032 41692 24084 41744
rect 25228 41692 25280 41744
rect 28540 41692 28592 41744
rect 21272 41556 21324 41608
rect 23388 41556 23440 41608
rect 24124 41556 24176 41608
rect 24308 41556 24360 41608
rect 25136 41624 25188 41676
rect 26976 41624 27028 41676
rect 25504 41556 25556 41608
rect 27528 41556 27580 41608
rect 27988 41599 28040 41608
rect 27988 41565 27997 41599
rect 27997 41565 28031 41599
rect 28031 41565 28040 41599
rect 27988 41556 28040 41565
rect 18512 41488 18564 41540
rect 19616 41488 19668 41540
rect 14280 41463 14332 41472
rect 14280 41429 14289 41463
rect 14289 41429 14323 41463
rect 14323 41429 14332 41463
rect 14280 41420 14332 41429
rect 15568 41420 15620 41472
rect 16856 41420 16908 41472
rect 19248 41463 19300 41472
rect 19248 41429 19257 41463
rect 19257 41429 19291 41463
rect 19291 41429 19300 41463
rect 19248 41420 19300 41429
rect 20720 41420 20772 41472
rect 21456 41463 21508 41472
rect 21456 41429 21465 41463
rect 21465 41429 21499 41463
rect 21499 41429 21508 41463
rect 21456 41420 21508 41429
rect 21824 41420 21876 41472
rect 25044 41488 25096 41540
rect 26240 41531 26292 41540
rect 26240 41497 26274 41531
rect 26274 41497 26292 41531
rect 26240 41488 26292 41497
rect 27160 41488 27212 41540
rect 23572 41420 23624 41472
rect 24584 41420 24636 41472
rect 24768 41420 24820 41472
rect 26976 41420 27028 41472
rect 27712 41420 27764 41472
rect 28724 41420 28776 41472
rect 30012 41463 30064 41472
rect 30012 41429 30021 41463
rect 30021 41429 30055 41463
rect 30055 41429 30064 41463
rect 30012 41420 30064 41429
rect 10880 41318 10932 41370
rect 10944 41318 10996 41370
rect 11008 41318 11060 41370
rect 11072 41318 11124 41370
rect 11136 41318 11188 41370
rect 20811 41318 20863 41370
rect 20875 41318 20927 41370
rect 20939 41318 20991 41370
rect 21003 41318 21055 41370
rect 21067 41318 21119 41370
rect 13912 41216 13964 41268
rect 14372 41216 14424 41268
rect 16672 41259 16724 41268
rect 16672 41225 16681 41259
rect 16681 41225 16715 41259
rect 16715 41225 16724 41259
rect 16672 41216 16724 41225
rect 18144 41259 18196 41268
rect 18144 41225 18153 41259
rect 18153 41225 18187 41259
rect 18187 41225 18196 41259
rect 18144 41216 18196 41225
rect 26240 41259 26292 41268
rect 26240 41225 26249 41259
rect 26249 41225 26283 41259
rect 26283 41225 26292 41259
rect 26240 41216 26292 41225
rect 26424 41216 26476 41268
rect 1584 41123 1636 41132
rect 1584 41089 1593 41123
rect 1593 41089 1627 41123
rect 1627 41089 1636 41123
rect 1584 41080 1636 41089
rect 14648 41080 14700 41132
rect 15016 41080 15068 41132
rect 18696 41148 18748 41200
rect 16856 41123 16908 41132
rect 16856 41089 16865 41123
rect 16865 41089 16899 41123
rect 16899 41089 16908 41123
rect 16856 41080 16908 41089
rect 19248 41123 19300 41132
rect 19248 41089 19257 41123
rect 19257 41089 19291 41123
rect 19291 41089 19300 41123
rect 19248 41080 19300 41089
rect 23848 41148 23900 41200
rect 15292 41012 15344 41064
rect 17132 41055 17184 41064
rect 17132 41021 17141 41055
rect 17141 41021 17175 41055
rect 17175 41021 17184 41055
rect 17132 41012 17184 41021
rect 18420 41012 18472 41064
rect 21824 41080 21876 41132
rect 24584 41080 24636 41132
rect 14464 40944 14516 40996
rect 12072 40876 12124 40928
rect 14188 40876 14240 40928
rect 18052 40944 18104 40996
rect 20720 41012 20772 41064
rect 21180 41012 21232 41064
rect 21640 41012 21692 41064
rect 23480 41055 23532 41064
rect 23480 41021 23489 41055
rect 23489 41021 23523 41055
rect 23523 41021 23532 41055
rect 23480 41012 23532 41021
rect 25044 41012 25096 41064
rect 25780 41123 25832 41132
rect 25780 41089 25789 41123
rect 25789 41089 25823 41123
rect 25823 41089 25832 41123
rect 25780 41080 25832 41089
rect 26976 41148 27028 41200
rect 28356 41148 28408 41200
rect 26608 41080 26660 41132
rect 28540 41080 28592 41132
rect 29736 41080 29788 41132
rect 19524 40944 19576 40996
rect 21456 40944 21508 40996
rect 22192 40944 22244 40996
rect 23112 40944 23164 40996
rect 25136 40944 25188 40996
rect 26424 41012 26476 41064
rect 28264 41012 28316 41064
rect 29552 41012 29604 41064
rect 28172 40944 28224 40996
rect 16396 40876 16448 40928
rect 17040 40919 17092 40928
rect 17040 40885 17049 40919
rect 17049 40885 17083 40919
rect 17083 40885 17092 40919
rect 17040 40876 17092 40885
rect 17500 40876 17552 40928
rect 17868 40876 17920 40928
rect 18144 40876 18196 40928
rect 20720 40919 20772 40928
rect 20720 40885 20729 40919
rect 20729 40885 20763 40919
rect 20763 40885 20772 40919
rect 20720 40876 20772 40885
rect 21732 40876 21784 40928
rect 24400 40876 24452 40928
rect 27896 40876 27948 40928
rect 28356 40919 28408 40928
rect 28356 40885 28365 40919
rect 28365 40885 28399 40919
rect 28399 40885 28408 40919
rect 28356 40876 28408 40885
rect 29184 40919 29236 40928
rect 29184 40885 29193 40919
rect 29193 40885 29227 40919
rect 29227 40885 29236 40919
rect 29184 40876 29236 40885
rect 30104 40876 30156 40928
rect 5915 40774 5967 40826
rect 5979 40774 6031 40826
rect 6043 40774 6095 40826
rect 6107 40774 6159 40826
rect 6171 40774 6223 40826
rect 15846 40774 15898 40826
rect 15910 40774 15962 40826
rect 15974 40774 16026 40826
rect 16038 40774 16090 40826
rect 16102 40774 16154 40826
rect 25776 40774 25828 40826
rect 25840 40774 25892 40826
rect 25904 40774 25956 40826
rect 25968 40774 26020 40826
rect 26032 40774 26084 40826
rect 12624 40672 12676 40724
rect 5356 40604 5408 40656
rect 11704 40536 11756 40588
rect 14556 40536 14608 40588
rect 15016 40604 15068 40656
rect 16856 40604 16908 40656
rect 19248 40672 19300 40724
rect 19708 40672 19760 40724
rect 20260 40715 20312 40724
rect 20260 40681 20269 40715
rect 20269 40681 20303 40715
rect 20303 40681 20312 40715
rect 20260 40672 20312 40681
rect 20720 40672 20772 40724
rect 21824 40715 21876 40724
rect 21824 40681 21833 40715
rect 21833 40681 21867 40715
rect 21867 40681 21876 40715
rect 21824 40672 21876 40681
rect 23480 40672 23532 40724
rect 26516 40672 26568 40724
rect 28816 40715 28868 40724
rect 28816 40681 28825 40715
rect 28825 40681 28859 40715
rect 28859 40681 28868 40715
rect 28816 40672 28868 40681
rect 29184 40672 29236 40724
rect 19524 40604 19576 40656
rect 20352 40604 20404 40656
rect 21180 40604 21232 40656
rect 14832 40468 14884 40520
rect 15292 40579 15344 40588
rect 15292 40545 15301 40579
rect 15301 40545 15335 40579
rect 15335 40545 15344 40579
rect 15292 40536 15344 40545
rect 16488 40536 16540 40588
rect 15292 40332 15344 40384
rect 16580 40375 16632 40384
rect 16580 40341 16589 40375
rect 16589 40341 16623 40375
rect 16623 40341 16632 40375
rect 16580 40332 16632 40341
rect 16948 40332 17000 40384
rect 17960 40536 18012 40588
rect 18512 40536 18564 40588
rect 22560 40536 22612 40588
rect 25412 40604 25464 40656
rect 27160 40604 27212 40656
rect 28540 40604 28592 40656
rect 25504 40536 25556 40588
rect 18052 40468 18104 40520
rect 19800 40511 19852 40520
rect 18236 40400 18288 40452
rect 18328 40400 18380 40452
rect 18604 40400 18656 40452
rect 19800 40477 19809 40511
rect 19809 40477 19843 40511
rect 19843 40477 19852 40511
rect 19800 40468 19852 40477
rect 20168 40468 20220 40520
rect 21364 40468 21416 40520
rect 22928 40511 22980 40520
rect 22928 40477 22937 40511
rect 22937 40477 22971 40511
rect 22971 40477 22980 40511
rect 22928 40468 22980 40477
rect 23572 40511 23624 40520
rect 23572 40477 23581 40511
rect 23581 40477 23615 40511
rect 23615 40477 23624 40511
rect 23572 40468 23624 40477
rect 19616 40375 19668 40384
rect 19616 40341 19625 40375
rect 19625 40341 19659 40375
rect 19659 40341 19668 40375
rect 19616 40332 19668 40341
rect 21272 40400 21324 40452
rect 23204 40400 23256 40452
rect 23296 40400 23348 40452
rect 25136 40400 25188 40452
rect 21364 40332 21416 40384
rect 22100 40332 22152 40384
rect 24860 40332 24912 40384
rect 25872 40468 25924 40520
rect 26424 40468 26476 40520
rect 26884 40511 26936 40520
rect 26884 40477 26893 40511
rect 26893 40477 26927 40511
rect 26927 40477 26936 40511
rect 26884 40468 26936 40477
rect 28908 40468 28960 40520
rect 29092 40468 29144 40520
rect 26240 40332 26292 40384
rect 26516 40400 26568 40452
rect 27068 40375 27120 40384
rect 27068 40341 27077 40375
rect 27077 40341 27111 40375
rect 27111 40341 27120 40375
rect 27068 40332 27120 40341
rect 28632 40332 28684 40384
rect 30012 40375 30064 40384
rect 30012 40341 30021 40375
rect 30021 40341 30055 40375
rect 30055 40341 30064 40375
rect 30012 40332 30064 40341
rect 10880 40230 10932 40282
rect 10944 40230 10996 40282
rect 11008 40230 11060 40282
rect 11072 40230 11124 40282
rect 11136 40230 11188 40282
rect 20811 40230 20863 40282
rect 20875 40230 20927 40282
rect 20939 40230 20991 40282
rect 21003 40230 21055 40282
rect 21067 40230 21119 40282
rect 14648 40171 14700 40180
rect 14648 40137 14657 40171
rect 14657 40137 14691 40171
rect 14691 40137 14700 40171
rect 14648 40128 14700 40137
rect 16580 40128 16632 40180
rect 17132 40128 17184 40180
rect 21456 40128 21508 40180
rect 22008 40128 22060 40180
rect 22560 40171 22612 40180
rect 22560 40137 22569 40171
rect 22569 40137 22603 40171
rect 22603 40137 22612 40171
rect 22560 40128 22612 40137
rect 22928 40128 22980 40180
rect 25872 40171 25924 40180
rect 25872 40137 25881 40171
rect 25881 40137 25915 40171
rect 25915 40137 25924 40171
rect 25872 40128 25924 40137
rect 26240 40128 26292 40180
rect 26792 40128 26844 40180
rect 27160 40171 27212 40180
rect 27160 40137 27169 40171
rect 27169 40137 27203 40171
rect 27203 40137 27212 40171
rect 27160 40128 27212 40137
rect 27344 40128 27396 40180
rect 29460 40128 29512 40180
rect 14556 40060 14608 40112
rect 12072 40035 12124 40044
rect 12072 40001 12081 40035
rect 12081 40001 12115 40035
rect 12115 40001 12124 40035
rect 12072 39992 12124 40001
rect 12256 40035 12308 40044
rect 12256 40001 12265 40035
rect 12265 40001 12299 40035
rect 12299 40001 12308 40035
rect 12256 39992 12308 40001
rect 14372 39992 14424 40044
rect 15108 40035 15160 40044
rect 15108 40001 15117 40035
rect 15117 40001 15151 40035
rect 15151 40001 15160 40035
rect 15108 39992 15160 40001
rect 16948 39992 17000 40044
rect 17684 39992 17736 40044
rect 19524 39992 19576 40044
rect 19708 40060 19760 40112
rect 20904 40060 20956 40112
rect 15200 39924 15252 39976
rect 17040 39967 17092 39976
rect 17040 39933 17049 39967
rect 17049 39933 17083 39967
rect 17083 39933 17092 39967
rect 17040 39924 17092 39933
rect 19708 39967 19760 39976
rect 19708 39933 19717 39967
rect 19717 39933 19751 39967
rect 19751 39933 19760 39967
rect 19708 39924 19760 39933
rect 20536 39992 20588 40044
rect 21272 40035 21324 40044
rect 21272 40001 21281 40035
rect 21281 40001 21315 40035
rect 21315 40001 21324 40035
rect 21272 39992 21324 40001
rect 22100 40035 22152 40044
rect 22100 40001 22109 40035
rect 22109 40001 22143 40035
rect 22143 40001 22152 40035
rect 23296 40060 23348 40112
rect 23388 40060 23440 40112
rect 22100 39992 22152 40001
rect 22836 39992 22888 40044
rect 23848 40035 23900 40044
rect 23848 40001 23857 40035
rect 23857 40001 23891 40035
rect 23891 40001 23900 40035
rect 23848 39992 23900 40001
rect 23296 39924 23348 39976
rect 24400 40035 24452 40044
rect 24400 40001 24409 40035
rect 24409 40001 24443 40035
rect 24443 40001 24452 40035
rect 24584 40035 24636 40044
rect 24400 39992 24452 40001
rect 24584 40001 24593 40035
rect 24593 40001 24627 40035
rect 24627 40001 24636 40035
rect 24584 39992 24636 40001
rect 26516 40060 26568 40112
rect 26700 40060 26752 40112
rect 29092 40060 29144 40112
rect 26976 40035 27028 40044
rect 26976 40001 26985 40035
rect 26985 40001 27019 40035
rect 27019 40001 27028 40035
rect 26976 39992 27028 40001
rect 28448 39992 28500 40044
rect 28816 39992 28868 40044
rect 24124 39967 24176 39976
rect 24124 39933 24133 39967
rect 24133 39933 24167 39967
rect 24167 39933 24176 39967
rect 24124 39924 24176 39933
rect 24308 39924 24360 39976
rect 24492 39924 24544 39976
rect 29644 39924 29696 39976
rect 23204 39856 23256 39908
rect 23388 39899 23440 39908
rect 23388 39865 23397 39899
rect 23397 39865 23431 39899
rect 23431 39865 23440 39899
rect 23388 39856 23440 39865
rect 16948 39788 17000 39840
rect 17592 39788 17644 39840
rect 20168 39831 20220 39840
rect 20168 39797 20177 39831
rect 20177 39797 20211 39831
rect 20211 39797 20220 39831
rect 20168 39788 20220 39797
rect 20904 39788 20956 39840
rect 21272 39788 21324 39840
rect 23664 39788 23716 39840
rect 24768 39788 24820 39840
rect 25320 39788 25372 39840
rect 26240 39788 26292 39840
rect 27252 39788 27304 39840
rect 28172 39831 28224 39840
rect 28172 39797 28181 39831
rect 28181 39797 28215 39831
rect 28215 39797 28224 39831
rect 28172 39788 28224 39797
rect 29368 39788 29420 39840
rect 30104 39788 30156 39840
rect 5915 39686 5967 39738
rect 5979 39686 6031 39738
rect 6043 39686 6095 39738
rect 6107 39686 6159 39738
rect 6171 39686 6223 39738
rect 15846 39686 15898 39738
rect 15910 39686 15962 39738
rect 15974 39686 16026 39738
rect 16038 39686 16090 39738
rect 16102 39686 16154 39738
rect 25776 39686 25828 39738
rect 25840 39686 25892 39738
rect 25904 39686 25956 39738
rect 25968 39686 26020 39738
rect 26032 39686 26084 39738
rect 19616 39627 19668 39636
rect 19616 39593 19625 39627
rect 19625 39593 19659 39627
rect 19659 39593 19668 39627
rect 19616 39584 19668 39593
rect 22744 39584 22796 39636
rect 23204 39584 23256 39636
rect 24860 39584 24912 39636
rect 25136 39627 25188 39636
rect 25136 39593 25145 39627
rect 25145 39593 25179 39627
rect 25179 39593 25188 39627
rect 25136 39584 25188 39593
rect 1584 39423 1636 39432
rect 1584 39389 1593 39423
rect 1593 39389 1627 39423
rect 1627 39389 1636 39423
rect 1584 39380 1636 39389
rect 16580 39448 16632 39500
rect 17776 39448 17828 39500
rect 19708 39516 19760 39568
rect 27620 39584 27672 39636
rect 29184 39584 29236 39636
rect 25320 39516 25372 39568
rect 25964 39516 26016 39568
rect 18512 39448 18564 39500
rect 21456 39448 21508 39500
rect 21640 39448 21692 39500
rect 15384 39423 15436 39432
rect 15384 39389 15393 39423
rect 15393 39389 15427 39423
rect 15427 39389 15436 39423
rect 15384 39380 15436 39389
rect 15476 39423 15528 39432
rect 15476 39389 15485 39423
rect 15485 39389 15519 39423
rect 15519 39389 15528 39423
rect 15476 39380 15528 39389
rect 15660 39380 15712 39432
rect 16028 39380 16080 39432
rect 17684 39423 17736 39432
rect 17684 39389 17693 39423
rect 17693 39389 17727 39423
rect 17727 39389 17736 39423
rect 17684 39380 17736 39389
rect 17868 39423 17920 39432
rect 17868 39389 17877 39423
rect 17877 39389 17911 39423
rect 17911 39389 17920 39423
rect 17868 39380 17920 39389
rect 18236 39423 18288 39432
rect 18236 39389 18245 39423
rect 18245 39389 18279 39423
rect 18279 39389 18288 39423
rect 18236 39380 18288 39389
rect 23480 39448 23532 39500
rect 24768 39491 24820 39500
rect 24768 39457 24777 39491
rect 24777 39457 24811 39491
rect 24811 39457 24820 39491
rect 24768 39448 24820 39457
rect 25596 39448 25648 39500
rect 22284 39423 22336 39432
rect 22284 39389 22293 39423
rect 22293 39389 22327 39423
rect 22327 39389 22336 39423
rect 22284 39380 22336 39389
rect 22836 39380 22888 39432
rect 18788 39312 18840 39364
rect 20720 39312 20772 39364
rect 23572 39312 23624 39364
rect 23848 39380 23900 39432
rect 24308 39380 24360 39432
rect 24492 39380 24544 39432
rect 24216 39312 24268 39364
rect 25412 39380 25464 39432
rect 24860 39312 24912 39364
rect 25504 39312 25556 39364
rect 25688 39312 25740 39364
rect 25964 39380 26016 39432
rect 26148 39423 26200 39432
rect 26148 39389 26157 39423
rect 26157 39389 26191 39423
rect 26191 39389 26200 39423
rect 26792 39448 26844 39500
rect 27528 39516 27580 39568
rect 28540 39516 28592 39568
rect 26148 39380 26200 39389
rect 26608 39423 26660 39432
rect 26608 39389 26617 39423
rect 26617 39389 26651 39423
rect 26651 39389 26660 39423
rect 26608 39380 26660 39389
rect 27252 39423 27304 39432
rect 27252 39389 27261 39423
rect 27261 39389 27295 39423
rect 27295 39389 27304 39423
rect 27252 39380 27304 39389
rect 12072 39244 12124 39296
rect 15936 39287 15988 39296
rect 15936 39253 15945 39287
rect 15945 39253 15979 39287
rect 15979 39253 15988 39287
rect 15936 39244 15988 39253
rect 18420 39287 18472 39296
rect 18420 39253 18429 39287
rect 18429 39253 18463 39287
rect 18463 39253 18472 39287
rect 18420 39244 18472 39253
rect 19156 39244 19208 39296
rect 20352 39244 20404 39296
rect 21640 39287 21692 39296
rect 21640 39253 21649 39287
rect 21649 39253 21683 39287
rect 21683 39253 21692 39287
rect 21640 39244 21692 39253
rect 22100 39244 22152 39296
rect 26056 39244 26108 39296
rect 26148 39244 26200 39296
rect 28540 39380 28592 39432
rect 28724 39423 28776 39432
rect 28724 39389 28733 39423
rect 28733 39389 28767 39423
rect 28767 39389 28776 39423
rect 28724 39380 28776 39389
rect 29092 39380 29144 39432
rect 28356 39312 28408 39364
rect 27804 39287 27856 39296
rect 27804 39253 27813 39287
rect 27813 39253 27847 39287
rect 27847 39253 27856 39287
rect 27804 39244 27856 39253
rect 28908 39287 28960 39296
rect 28908 39253 28917 39287
rect 28917 39253 28951 39287
rect 28951 39253 28960 39287
rect 28908 39244 28960 39253
rect 10880 39142 10932 39194
rect 10944 39142 10996 39194
rect 11008 39142 11060 39194
rect 11072 39142 11124 39194
rect 11136 39142 11188 39194
rect 20811 39142 20863 39194
rect 20875 39142 20927 39194
rect 20939 39142 20991 39194
rect 21003 39142 21055 39194
rect 21067 39142 21119 39194
rect 15752 39040 15804 39092
rect 16028 39083 16080 39092
rect 16028 39049 16037 39083
rect 16037 39049 16071 39083
rect 16071 39049 16080 39083
rect 16028 39040 16080 39049
rect 20720 39040 20772 39092
rect 22100 39083 22152 39092
rect 22100 39049 22109 39083
rect 22109 39049 22143 39083
rect 22143 39049 22152 39083
rect 23020 39083 23072 39092
rect 22100 39040 22152 39049
rect 23020 39049 23029 39083
rect 23029 39049 23063 39083
rect 23063 39049 23072 39083
rect 23020 39040 23072 39049
rect 23664 39083 23716 39092
rect 23664 39049 23673 39083
rect 23673 39049 23707 39083
rect 23707 39049 23716 39083
rect 23664 39040 23716 39049
rect 23756 39040 23808 39092
rect 28540 39083 28592 39092
rect 12072 38947 12124 38956
rect 12072 38913 12081 38947
rect 12081 38913 12115 38947
rect 12115 38913 12124 38947
rect 12072 38904 12124 38913
rect 12256 38947 12308 38956
rect 12256 38913 12265 38947
rect 12265 38913 12299 38947
rect 12299 38913 12308 38947
rect 12256 38904 12308 38913
rect 14096 38836 14148 38888
rect 18420 38972 18472 39024
rect 15936 38904 15988 38956
rect 16672 38947 16724 38956
rect 16672 38913 16681 38947
rect 16681 38913 16715 38947
rect 16715 38913 16724 38947
rect 16672 38904 16724 38913
rect 16948 38947 17000 38956
rect 16948 38913 16982 38947
rect 16982 38913 17000 38947
rect 18512 38947 18564 38956
rect 16948 38904 17000 38913
rect 18512 38913 18521 38947
rect 18521 38913 18555 38947
rect 18555 38913 18564 38947
rect 18512 38904 18564 38913
rect 19156 38904 19208 38956
rect 19524 38904 19576 38956
rect 19984 38904 20036 38956
rect 21180 38972 21232 39024
rect 21640 38904 21692 38956
rect 26332 38972 26384 39024
rect 27804 38972 27856 39024
rect 28540 39049 28549 39083
rect 28549 39049 28583 39083
rect 28583 39049 28592 39083
rect 28540 39040 28592 39049
rect 23756 38904 23808 38956
rect 24308 38947 24360 38956
rect 19708 38836 19760 38888
rect 20536 38768 20588 38820
rect 24308 38913 24317 38947
rect 24317 38913 24351 38947
rect 24351 38913 24360 38947
rect 24308 38904 24360 38913
rect 24400 38904 24452 38956
rect 24676 38947 24728 38956
rect 24676 38913 24685 38947
rect 24685 38913 24719 38947
rect 24719 38913 24728 38947
rect 24676 38904 24728 38913
rect 25504 38904 25556 38956
rect 25688 38947 25740 38956
rect 25688 38913 25697 38947
rect 25697 38913 25731 38947
rect 25731 38913 25740 38947
rect 25688 38904 25740 38913
rect 25780 38904 25832 38956
rect 26148 38904 26200 38956
rect 24216 38836 24268 38888
rect 25596 38836 25648 38888
rect 27068 38904 27120 38956
rect 28356 38904 28408 38956
rect 25412 38768 25464 38820
rect 25780 38768 25832 38820
rect 26332 38768 26384 38820
rect 29092 38768 29144 38820
rect 18052 38743 18104 38752
rect 18052 38709 18061 38743
rect 18061 38709 18095 38743
rect 18095 38709 18104 38743
rect 18052 38700 18104 38709
rect 18236 38700 18288 38752
rect 24952 38700 25004 38752
rect 27068 38700 27120 38752
rect 29368 38743 29420 38752
rect 29368 38709 29377 38743
rect 29377 38709 29411 38743
rect 29411 38709 29420 38743
rect 29368 38700 29420 38709
rect 5915 38598 5967 38650
rect 5979 38598 6031 38650
rect 6043 38598 6095 38650
rect 6107 38598 6159 38650
rect 6171 38598 6223 38650
rect 15846 38598 15898 38650
rect 15910 38598 15962 38650
rect 15974 38598 16026 38650
rect 16038 38598 16090 38650
rect 16102 38598 16154 38650
rect 25776 38598 25828 38650
rect 25840 38598 25892 38650
rect 25904 38598 25956 38650
rect 25968 38598 26020 38650
rect 26032 38598 26084 38650
rect 16948 38496 17000 38548
rect 15660 38428 15712 38480
rect 15200 38360 15252 38412
rect 15476 38360 15528 38412
rect 10140 38335 10192 38344
rect 10140 38301 10149 38335
rect 10149 38301 10183 38335
rect 10183 38301 10192 38335
rect 10140 38292 10192 38301
rect 14096 38335 14148 38344
rect 14096 38301 14105 38335
rect 14105 38301 14139 38335
rect 14139 38301 14148 38335
rect 14096 38292 14148 38301
rect 16304 38335 16356 38344
rect 10600 38224 10652 38276
rect 15384 38224 15436 38276
rect 16304 38301 16313 38335
rect 16313 38301 16347 38335
rect 16347 38301 16356 38335
rect 16304 38292 16356 38301
rect 18052 38360 18104 38412
rect 17684 38292 17736 38344
rect 18144 38335 18196 38344
rect 18144 38301 18153 38335
rect 18153 38301 18187 38335
rect 18187 38301 18196 38335
rect 18144 38292 18196 38301
rect 19616 38428 19668 38480
rect 20076 38496 20128 38548
rect 16580 38224 16632 38276
rect 17776 38224 17828 38276
rect 18052 38224 18104 38276
rect 20536 38292 20588 38344
rect 21640 38335 21692 38344
rect 21640 38301 21649 38335
rect 21649 38301 21683 38335
rect 21683 38301 21692 38335
rect 21640 38292 21692 38301
rect 22100 38292 22152 38344
rect 24492 38292 24544 38344
rect 24676 38335 24728 38344
rect 24676 38301 24685 38335
rect 24685 38301 24719 38335
rect 24719 38301 24728 38335
rect 24676 38292 24728 38301
rect 24952 38335 25004 38344
rect 24952 38301 24986 38335
rect 24986 38301 25004 38335
rect 24952 38292 25004 38301
rect 25504 38292 25556 38344
rect 26424 38496 26476 38548
rect 26976 38496 27028 38548
rect 28356 38496 28408 38548
rect 27160 38403 27212 38412
rect 27160 38369 27169 38403
rect 27169 38369 27203 38403
rect 27203 38369 27212 38403
rect 27160 38360 27212 38369
rect 26516 38335 26568 38344
rect 26516 38301 26525 38335
rect 26525 38301 26559 38335
rect 26559 38301 26568 38335
rect 26516 38292 26568 38301
rect 27068 38292 27120 38344
rect 28632 38292 28684 38344
rect 20168 38224 20220 38276
rect 11244 38156 11296 38208
rect 16028 38156 16080 38208
rect 17500 38156 17552 38208
rect 18696 38199 18748 38208
rect 18696 38165 18705 38199
rect 18705 38165 18739 38199
rect 18739 38165 18748 38199
rect 18696 38156 18748 38165
rect 21272 38156 21324 38208
rect 21364 38156 21416 38208
rect 21640 38156 21692 38208
rect 21916 38156 21968 38208
rect 22560 38156 22612 38208
rect 23480 38199 23532 38208
rect 23480 38165 23489 38199
rect 23489 38165 23523 38199
rect 23523 38165 23532 38199
rect 23480 38156 23532 38165
rect 30012 38199 30064 38208
rect 30012 38165 30021 38199
rect 30021 38165 30055 38199
rect 30055 38165 30064 38199
rect 30012 38156 30064 38165
rect 10880 38054 10932 38106
rect 10944 38054 10996 38106
rect 11008 38054 11060 38106
rect 11072 38054 11124 38106
rect 11136 38054 11188 38106
rect 20811 38054 20863 38106
rect 20875 38054 20927 38106
rect 20939 38054 20991 38106
rect 21003 38054 21055 38106
rect 21067 38054 21119 38106
rect 7012 37884 7064 37936
rect 9956 37816 10008 37868
rect 10784 37816 10836 37868
rect 14096 37884 14148 37936
rect 13084 37816 13136 37868
rect 14924 37859 14976 37868
rect 10324 37791 10376 37800
rect 10324 37757 10333 37791
rect 10333 37757 10367 37791
rect 10367 37757 10376 37791
rect 10324 37748 10376 37757
rect 10508 37748 10560 37800
rect 14924 37825 14933 37859
rect 14933 37825 14967 37859
rect 14967 37825 14976 37859
rect 14924 37816 14976 37825
rect 15108 37884 15160 37936
rect 15660 37952 15712 38004
rect 18512 37952 18564 38004
rect 22100 37995 22152 38004
rect 22100 37961 22109 37995
rect 22109 37961 22143 37995
rect 22143 37961 22152 37995
rect 22100 37952 22152 37961
rect 22744 37952 22796 38004
rect 26884 37952 26936 38004
rect 15752 37816 15804 37868
rect 16028 37816 16080 37868
rect 18144 37816 18196 37868
rect 18696 37884 18748 37936
rect 20444 37884 20496 37936
rect 19984 37816 20036 37868
rect 25412 37884 25464 37936
rect 28264 37884 28316 37936
rect 20628 37859 20680 37868
rect 20628 37825 20637 37859
rect 20637 37825 20671 37859
rect 20671 37825 20680 37859
rect 20628 37816 20680 37825
rect 22100 37816 22152 37868
rect 22560 37859 22612 37868
rect 22560 37825 22569 37859
rect 22569 37825 22603 37859
rect 22603 37825 22612 37859
rect 22560 37816 22612 37825
rect 23756 37816 23808 37868
rect 24768 37859 24820 37868
rect 24768 37825 24777 37859
rect 24777 37825 24811 37859
rect 24811 37825 24820 37859
rect 24768 37816 24820 37825
rect 25688 37816 25740 37868
rect 26516 37816 26568 37868
rect 27896 37859 27948 37868
rect 27896 37825 27905 37859
rect 27905 37825 27939 37859
rect 27939 37825 27948 37859
rect 27896 37816 27948 37825
rect 28540 37859 28592 37868
rect 28540 37825 28549 37859
rect 28549 37825 28583 37859
rect 28583 37825 28592 37859
rect 28540 37816 28592 37825
rect 15384 37748 15436 37800
rect 20352 37791 20404 37800
rect 20352 37757 20361 37791
rect 20361 37757 20395 37791
rect 20395 37757 20404 37791
rect 20352 37748 20404 37757
rect 20444 37791 20496 37800
rect 20444 37757 20453 37791
rect 20453 37757 20487 37791
rect 20487 37757 20496 37791
rect 20444 37748 20496 37757
rect 16580 37680 16632 37732
rect 17132 37680 17184 37732
rect 10692 37612 10744 37664
rect 13636 37655 13688 37664
rect 13636 37621 13645 37655
rect 13645 37621 13679 37655
rect 13679 37621 13688 37655
rect 13636 37612 13688 37621
rect 16488 37612 16540 37664
rect 16948 37612 17000 37664
rect 18420 37612 18472 37664
rect 19616 37655 19668 37664
rect 19616 37621 19625 37655
rect 19625 37621 19659 37655
rect 19659 37621 19668 37655
rect 19616 37612 19668 37621
rect 20536 37612 20588 37664
rect 21180 37612 21232 37664
rect 22928 37612 22980 37664
rect 23940 37655 23992 37664
rect 23940 37621 23949 37655
rect 23949 37621 23983 37655
rect 23983 37621 23992 37655
rect 23940 37612 23992 37621
rect 29092 37748 29144 37800
rect 28724 37612 28776 37664
rect 29276 37612 29328 37664
rect 29368 37655 29420 37664
rect 29368 37621 29377 37655
rect 29377 37621 29411 37655
rect 29411 37621 29420 37655
rect 29368 37612 29420 37621
rect 5915 37510 5967 37562
rect 5979 37510 6031 37562
rect 6043 37510 6095 37562
rect 6107 37510 6159 37562
rect 6171 37510 6223 37562
rect 15846 37510 15898 37562
rect 15910 37510 15962 37562
rect 15974 37510 16026 37562
rect 16038 37510 16090 37562
rect 16102 37510 16154 37562
rect 25776 37510 25828 37562
rect 25840 37510 25892 37562
rect 25904 37510 25956 37562
rect 25968 37510 26020 37562
rect 26032 37510 26084 37562
rect 13084 37408 13136 37460
rect 15108 37408 15160 37460
rect 21272 37408 21324 37460
rect 23756 37451 23808 37460
rect 23756 37417 23765 37451
rect 23765 37417 23799 37451
rect 23799 37417 23808 37451
rect 23756 37408 23808 37417
rect 24492 37408 24544 37460
rect 12624 37340 12676 37392
rect 1584 37247 1636 37256
rect 1584 37213 1593 37247
rect 1593 37213 1627 37247
rect 1627 37213 1636 37247
rect 1584 37204 1636 37213
rect 10140 37204 10192 37256
rect 10416 37247 10468 37256
rect 10416 37213 10425 37247
rect 10425 37213 10459 37247
rect 10459 37213 10468 37247
rect 10416 37204 10468 37213
rect 10692 37247 10744 37256
rect 10692 37213 10726 37247
rect 10726 37213 10744 37247
rect 10692 37204 10744 37213
rect 13268 37272 13320 37324
rect 18788 37340 18840 37392
rect 23204 37340 23256 37392
rect 28264 37408 28316 37460
rect 29368 37408 29420 37460
rect 15200 37315 15252 37324
rect 15200 37281 15209 37315
rect 15209 37281 15243 37315
rect 15243 37281 15252 37315
rect 15200 37272 15252 37281
rect 15660 37315 15712 37324
rect 15660 37281 15669 37315
rect 15669 37281 15703 37315
rect 15703 37281 15712 37315
rect 15660 37272 15712 37281
rect 19984 37272 20036 37324
rect 20076 37272 20128 37324
rect 9956 37136 10008 37188
rect 12532 37136 12584 37188
rect 10692 37068 10744 37120
rect 10784 37068 10836 37120
rect 12164 37068 12216 37120
rect 12900 37204 12952 37256
rect 13636 37204 13688 37256
rect 15016 37204 15068 37256
rect 14740 37136 14792 37188
rect 15384 37204 15436 37256
rect 16580 37204 16632 37256
rect 16764 37136 16816 37188
rect 18696 37136 18748 37188
rect 19248 37247 19300 37256
rect 19248 37213 19257 37247
rect 19257 37213 19291 37247
rect 19291 37213 19300 37247
rect 19248 37204 19300 37213
rect 22192 37204 22244 37256
rect 22928 37204 22980 37256
rect 23020 37247 23072 37256
rect 23020 37213 23029 37247
rect 23029 37213 23063 37247
rect 23063 37213 23072 37247
rect 23296 37315 23348 37324
rect 23296 37281 23305 37315
rect 23305 37281 23339 37315
rect 23339 37281 23348 37315
rect 23296 37272 23348 37281
rect 23020 37204 23072 37213
rect 23388 37247 23440 37256
rect 23388 37213 23397 37247
rect 23397 37213 23431 37247
rect 23431 37213 23440 37247
rect 23940 37272 23992 37324
rect 23388 37204 23440 37213
rect 20628 37136 20680 37188
rect 20904 37179 20956 37188
rect 20904 37145 20938 37179
rect 20938 37145 20956 37179
rect 20904 37136 20956 37145
rect 22100 37136 22152 37188
rect 24492 37204 24544 37256
rect 24952 37204 25004 37256
rect 26148 37272 26200 37324
rect 25780 37204 25832 37256
rect 26700 37204 26752 37256
rect 27988 37340 28040 37392
rect 27344 37204 27396 37256
rect 27804 37247 27856 37256
rect 27804 37213 27813 37247
rect 27813 37213 27847 37247
rect 27847 37213 27856 37247
rect 27804 37204 27856 37213
rect 29092 37272 29144 37324
rect 17040 37068 17092 37120
rect 21364 37068 21416 37120
rect 22928 37068 22980 37120
rect 23296 37068 23348 37120
rect 25780 37068 25832 37120
rect 27344 37111 27396 37120
rect 27344 37077 27353 37111
rect 27353 37077 27387 37111
rect 27387 37077 27396 37111
rect 27344 37068 27396 37077
rect 27988 37111 28040 37120
rect 27988 37077 27997 37111
rect 27997 37077 28031 37111
rect 28031 37077 28040 37111
rect 27988 37068 28040 37077
rect 28816 37111 28868 37120
rect 28816 37077 28825 37111
rect 28825 37077 28859 37111
rect 28859 37077 28868 37111
rect 28816 37068 28868 37077
rect 28908 37068 28960 37120
rect 10880 36966 10932 37018
rect 10944 36966 10996 37018
rect 11008 36966 11060 37018
rect 11072 36966 11124 37018
rect 11136 36966 11188 37018
rect 20811 36966 20863 37018
rect 20875 36966 20927 37018
rect 20939 36966 20991 37018
rect 21003 36966 21055 37018
rect 21067 36966 21119 37018
rect 10600 36907 10652 36916
rect 10600 36873 10609 36907
rect 10609 36873 10643 36907
rect 10643 36873 10652 36907
rect 10600 36864 10652 36873
rect 10692 36864 10744 36916
rect 12072 36864 12124 36916
rect 8852 36771 8904 36780
rect 8852 36737 8861 36771
rect 8861 36737 8895 36771
rect 8895 36737 8904 36771
rect 8852 36728 8904 36737
rect 9680 36728 9732 36780
rect 9956 36796 10008 36848
rect 19432 36864 19484 36916
rect 10048 36771 10100 36780
rect 10048 36737 10057 36771
rect 10057 36737 10091 36771
rect 10091 36737 10100 36771
rect 10048 36728 10100 36737
rect 10324 36728 10376 36780
rect 11244 36728 11296 36780
rect 13176 36728 13228 36780
rect 12164 36660 12216 36712
rect 9312 36524 9364 36576
rect 10416 36592 10468 36644
rect 10508 36524 10560 36576
rect 11796 36567 11848 36576
rect 11796 36533 11805 36567
rect 11805 36533 11839 36567
rect 11839 36533 11848 36567
rect 11796 36524 11848 36533
rect 12624 36703 12676 36712
rect 12624 36669 12633 36703
rect 12633 36669 12667 36703
rect 12667 36669 12676 36703
rect 12624 36660 12676 36669
rect 15200 36771 15252 36780
rect 15200 36737 15209 36771
rect 15209 36737 15243 36771
rect 15243 36737 15252 36771
rect 15200 36728 15252 36737
rect 15384 36728 15436 36780
rect 17224 36771 17276 36780
rect 17224 36737 17233 36771
rect 17233 36737 17267 36771
rect 17267 36737 17276 36771
rect 17224 36728 17276 36737
rect 17684 36728 17736 36780
rect 19248 36796 19300 36848
rect 17224 36592 17276 36644
rect 18052 36660 18104 36712
rect 22100 36728 22152 36780
rect 22652 36771 22704 36780
rect 22652 36737 22661 36771
rect 22661 36737 22695 36771
rect 22695 36737 22704 36771
rect 22652 36728 22704 36737
rect 18788 36592 18840 36644
rect 19432 36660 19484 36712
rect 22376 36660 22428 36712
rect 22928 36771 22980 36780
rect 22928 36737 22937 36771
rect 22937 36737 22971 36771
rect 22971 36737 22980 36771
rect 22928 36728 22980 36737
rect 23296 36864 23348 36916
rect 24492 36864 24544 36916
rect 24860 36796 24912 36848
rect 19524 36592 19576 36644
rect 17132 36524 17184 36576
rect 22744 36524 22796 36576
rect 23480 36728 23532 36780
rect 25688 36771 25740 36780
rect 25688 36737 25697 36771
rect 25697 36737 25731 36771
rect 25731 36737 25740 36771
rect 25688 36728 25740 36737
rect 26056 36796 26108 36848
rect 26148 36728 26200 36780
rect 28816 36864 28868 36916
rect 28448 36796 28500 36848
rect 25780 36660 25832 36712
rect 26976 36703 27028 36712
rect 26976 36669 26985 36703
rect 26985 36669 27019 36703
rect 27019 36669 27028 36703
rect 26976 36660 27028 36669
rect 29092 36635 29144 36644
rect 29092 36601 29101 36635
rect 29101 36601 29135 36635
rect 29135 36601 29144 36635
rect 29092 36592 29144 36601
rect 29368 36524 29420 36576
rect 5915 36422 5967 36474
rect 5979 36422 6031 36474
rect 6043 36422 6095 36474
rect 6107 36422 6159 36474
rect 6171 36422 6223 36474
rect 15846 36422 15898 36474
rect 15910 36422 15962 36474
rect 15974 36422 16026 36474
rect 16038 36422 16090 36474
rect 16102 36422 16154 36474
rect 25776 36422 25828 36474
rect 25840 36422 25892 36474
rect 25904 36422 25956 36474
rect 25968 36422 26020 36474
rect 26032 36422 26084 36474
rect 13268 36320 13320 36372
rect 19156 36320 19208 36372
rect 19800 36320 19852 36372
rect 22376 36320 22428 36372
rect 24584 36320 24636 36372
rect 28264 36363 28316 36372
rect 28264 36329 28273 36363
rect 28273 36329 28307 36363
rect 28307 36329 28316 36363
rect 28264 36320 28316 36329
rect 28908 36363 28960 36372
rect 28908 36329 28917 36363
rect 28917 36329 28951 36363
rect 28951 36329 28960 36363
rect 28908 36320 28960 36329
rect 13820 36252 13872 36304
rect 22652 36252 22704 36304
rect 23020 36252 23072 36304
rect 23296 36252 23348 36304
rect 25044 36252 25096 36304
rect 26700 36252 26752 36304
rect 11244 36116 11296 36168
rect 10784 36091 10836 36100
rect 10784 36057 10793 36091
rect 10793 36057 10827 36091
rect 10827 36057 10836 36091
rect 10784 36048 10836 36057
rect 11612 36116 11664 36168
rect 12624 36116 12676 36168
rect 9680 35980 9732 36032
rect 12900 36048 12952 36100
rect 11980 35980 12032 36032
rect 12164 35980 12216 36032
rect 13268 36116 13320 36168
rect 13544 36116 13596 36168
rect 16672 36184 16724 36236
rect 19616 36184 19668 36236
rect 20076 36184 20128 36236
rect 22928 36184 22980 36236
rect 24860 36184 24912 36236
rect 25688 36227 25740 36236
rect 25688 36193 25697 36227
rect 25697 36193 25731 36227
rect 25731 36193 25740 36227
rect 25688 36184 25740 36193
rect 17132 36159 17184 36168
rect 13912 36048 13964 36100
rect 15844 36048 15896 36100
rect 17132 36125 17166 36159
rect 17166 36125 17184 36159
rect 17132 36116 17184 36125
rect 18604 36116 18656 36168
rect 19064 36116 19116 36168
rect 13268 35980 13320 36032
rect 15200 35980 15252 36032
rect 15752 35980 15804 36032
rect 17684 35980 17736 36032
rect 18696 35980 18748 36032
rect 19064 35980 19116 36032
rect 21272 36048 21324 36100
rect 22100 36159 22152 36168
rect 22100 36125 22109 36159
rect 22109 36125 22143 36159
rect 22143 36125 22152 36159
rect 22100 36116 22152 36125
rect 22744 36116 22796 36168
rect 24492 36116 24544 36168
rect 27988 36116 28040 36168
rect 28172 36116 28224 36168
rect 29276 36116 29328 36168
rect 21364 35980 21416 36032
rect 23112 36048 23164 36100
rect 23020 36023 23072 36032
rect 23020 35989 23029 36023
rect 23029 35989 23063 36023
rect 23063 35989 23072 36023
rect 23020 35980 23072 35989
rect 23756 36023 23808 36032
rect 23756 35989 23765 36023
rect 23765 35989 23799 36023
rect 23799 35989 23808 36023
rect 23756 35980 23808 35989
rect 27344 36048 27396 36100
rect 27712 35980 27764 36032
rect 30012 36023 30064 36032
rect 30012 35989 30021 36023
rect 30021 35989 30055 36023
rect 30055 35989 30064 36023
rect 30012 35980 30064 35989
rect 10880 35878 10932 35930
rect 10944 35878 10996 35930
rect 11008 35878 11060 35930
rect 11072 35878 11124 35930
rect 11136 35878 11188 35930
rect 20811 35878 20863 35930
rect 20875 35878 20927 35930
rect 20939 35878 20991 35930
rect 21003 35878 21055 35930
rect 21067 35878 21119 35930
rect 10416 35708 10468 35760
rect 11796 35708 11848 35760
rect 9312 35683 9364 35692
rect 9312 35649 9346 35683
rect 9346 35649 9364 35683
rect 9312 35640 9364 35649
rect 12072 35683 12124 35692
rect 12072 35649 12081 35683
rect 12081 35649 12115 35683
rect 12115 35649 12124 35683
rect 12072 35640 12124 35649
rect 12256 35683 12308 35692
rect 12256 35649 12265 35683
rect 12265 35649 12299 35683
rect 12299 35649 12308 35683
rect 12256 35640 12308 35649
rect 13544 35640 13596 35692
rect 13268 35615 13320 35624
rect 13268 35581 13277 35615
rect 13277 35581 13311 35615
rect 13311 35581 13320 35615
rect 13268 35572 13320 35581
rect 14464 35572 14516 35624
rect 15384 35683 15436 35692
rect 15384 35649 15393 35683
rect 15393 35649 15427 35683
rect 15427 35649 15436 35683
rect 15384 35640 15436 35649
rect 15476 35615 15528 35624
rect 15476 35581 15485 35615
rect 15485 35581 15519 35615
rect 15519 35581 15528 35615
rect 15476 35572 15528 35581
rect 15752 35708 15804 35760
rect 19984 35708 20036 35760
rect 20628 35776 20680 35828
rect 20812 35708 20864 35760
rect 22928 35776 22980 35828
rect 23204 35776 23256 35828
rect 26516 35776 26568 35828
rect 27804 35819 27856 35828
rect 27804 35785 27813 35819
rect 27813 35785 27847 35819
rect 27847 35785 27856 35819
rect 27804 35776 27856 35785
rect 27896 35776 27948 35828
rect 17132 35640 17184 35692
rect 17960 35683 18012 35692
rect 17960 35649 17969 35683
rect 17969 35649 18003 35683
rect 18003 35649 18012 35683
rect 17960 35640 18012 35649
rect 18328 35640 18380 35692
rect 19432 35640 19484 35692
rect 19616 35640 19668 35692
rect 22652 35708 22704 35760
rect 15844 35615 15896 35624
rect 15844 35581 15853 35615
rect 15853 35581 15887 35615
rect 15887 35581 15896 35615
rect 15844 35572 15896 35581
rect 16580 35572 16632 35624
rect 18880 35615 18932 35624
rect 18880 35581 18889 35615
rect 18889 35581 18923 35615
rect 18923 35581 18932 35615
rect 18880 35572 18932 35581
rect 19708 35572 19760 35624
rect 22100 35572 22152 35624
rect 23388 35640 23440 35692
rect 23756 35640 23808 35692
rect 25136 35640 25188 35692
rect 27712 35640 27764 35692
rect 28632 35683 28684 35692
rect 28632 35649 28641 35683
rect 28641 35649 28675 35683
rect 28675 35649 28684 35683
rect 28632 35640 28684 35649
rect 29092 35683 29144 35692
rect 29092 35649 29101 35683
rect 29101 35649 29135 35683
rect 29135 35649 29144 35683
rect 29092 35640 29144 35649
rect 23848 35572 23900 35624
rect 9680 35436 9732 35488
rect 13912 35436 13964 35488
rect 14464 35436 14516 35488
rect 19800 35504 19852 35556
rect 24952 35504 25004 35556
rect 18052 35436 18104 35488
rect 20260 35436 20312 35488
rect 22836 35436 22888 35488
rect 23572 35436 23624 35488
rect 26424 35436 26476 35488
rect 29920 35436 29972 35488
rect 5915 35334 5967 35386
rect 5979 35334 6031 35386
rect 6043 35334 6095 35386
rect 6107 35334 6159 35386
rect 6171 35334 6223 35386
rect 15846 35334 15898 35386
rect 15910 35334 15962 35386
rect 15974 35334 16026 35386
rect 16038 35334 16090 35386
rect 16102 35334 16154 35386
rect 25776 35334 25828 35386
rect 25840 35334 25892 35386
rect 25904 35334 25956 35386
rect 25968 35334 26020 35386
rect 26032 35334 26084 35386
rect 14464 35232 14516 35284
rect 16672 35232 16724 35284
rect 16764 35232 16816 35284
rect 17960 35232 18012 35284
rect 18512 35232 18564 35284
rect 19616 35232 19668 35284
rect 23388 35275 23440 35284
rect 18144 35164 18196 35216
rect 18880 35164 18932 35216
rect 21272 35207 21324 35216
rect 21272 35173 21281 35207
rect 21281 35173 21315 35207
rect 21315 35173 21324 35207
rect 21272 35164 21324 35173
rect 1584 35071 1636 35080
rect 1584 35037 1593 35071
rect 1593 35037 1627 35071
rect 1627 35037 1636 35071
rect 1584 35028 1636 35037
rect 10140 35028 10192 35080
rect 12256 35071 12308 35080
rect 12256 35037 12265 35071
rect 12265 35037 12299 35071
rect 12299 35037 12308 35071
rect 12256 35028 12308 35037
rect 15200 35028 15252 35080
rect 15384 35071 15436 35080
rect 15384 35037 15393 35071
rect 15393 35037 15427 35071
rect 15427 35037 15436 35071
rect 15384 35028 15436 35037
rect 19708 35096 19760 35148
rect 19800 35096 19852 35148
rect 20352 35096 20404 35148
rect 16764 35028 16816 35080
rect 17776 35028 17828 35080
rect 19064 35028 19116 35080
rect 20444 35028 20496 35080
rect 13176 34960 13228 35012
rect 15660 34960 15712 35012
rect 20168 34960 20220 35012
rect 11244 34892 11296 34944
rect 14924 34892 14976 34944
rect 17040 34892 17092 34944
rect 17408 34892 17460 34944
rect 19524 34892 19576 34944
rect 20904 35071 20956 35080
rect 20904 35037 20913 35071
rect 20913 35037 20947 35071
rect 20947 35037 20956 35071
rect 20904 35028 20956 35037
rect 21364 35028 21416 35080
rect 23388 35241 23397 35275
rect 23397 35241 23431 35275
rect 23431 35241 23440 35275
rect 23388 35232 23440 35241
rect 25136 35275 25188 35284
rect 25136 35241 25145 35275
rect 25145 35241 25179 35275
rect 25179 35241 25188 35275
rect 25136 35232 25188 35241
rect 26976 35232 27028 35284
rect 24400 35164 24452 35216
rect 28356 35232 28408 35284
rect 28540 35232 28592 35284
rect 29920 35275 29972 35284
rect 29092 35164 29144 35216
rect 29920 35241 29929 35275
rect 29929 35241 29963 35275
rect 29963 35241 29972 35275
rect 29920 35232 29972 35241
rect 23480 35028 23532 35080
rect 24860 35096 24912 35148
rect 24952 35071 25004 35080
rect 21824 35003 21876 35012
rect 21824 34969 21833 35003
rect 21833 34969 21867 35003
rect 21867 34969 21876 35003
rect 21824 34960 21876 34969
rect 24124 34960 24176 35012
rect 24492 34960 24544 35012
rect 24952 35037 24961 35071
rect 24961 35037 24995 35071
rect 24995 35037 25004 35071
rect 24952 35028 25004 35037
rect 26424 35071 26476 35080
rect 26424 35037 26433 35071
rect 26433 35037 26467 35071
rect 26467 35037 26476 35071
rect 26424 35028 26476 35037
rect 30104 35096 30156 35148
rect 28264 35071 28316 35080
rect 28264 35037 28273 35071
rect 28273 35037 28307 35071
rect 28307 35037 28316 35071
rect 28264 35028 28316 35037
rect 28724 35071 28776 35080
rect 28724 35037 28733 35071
rect 28733 35037 28767 35071
rect 28767 35037 28776 35071
rect 28724 35028 28776 35037
rect 29460 34960 29512 35012
rect 22008 34892 22060 34944
rect 22376 34892 22428 34944
rect 27988 34892 28040 34944
rect 28908 34935 28960 34944
rect 28908 34901 28917 34935
rect 28917 34901 28951 34935
rect 28951 34901 28960 34935
rect 28908 34892 28960 34901
rect 29000 34892 29052 34944
rect 10880 34790 10932 34842
rect 10944 34790 10996 34842
rect 11008 34790 11060 34842
rect 11072 34790 11124 34842
rect 11136 34790 11188 34842
rect 20811 34790 20863 34842
rect 20875 34790 20927 34842
rect 20939 34790 20991 34842
rect 21003 34790 21055 34842
rect 21067 34790 21119 34842
rect 10692 34731 10744 34740
rect 10692 34697 10701 34731
rect 10701 34697 10735 34731
rect 10735 34697 10744 34731
rect 10692 34688 10744 34697
rect 11336 34688 11388 34740
rect 17224 34731 17276 34740
rect 10048 34552 10100 34604
rect 12164 34552 12216 34604
rect 13544 34552 13596 34604
rect 14280 34552 14332 34604
rect 11520 34527 11572 34536
rect 11520 34493 11529 34527
rect 11529 34493 11563 34527
rect 11563 34493 11572 34527
rect 11520 34484 11572 34493
rect 15016 34552 15068 34604
rect 17224 34697 17233 34731
rect 17233 34697 17267 34731
rect 17267 34697 17276 34731
rect 17224 34688 17276 34697
rect 17316 34688 17368 34740
rect 18788 34620 18840 34672
rect 19248 34620 19300 34672
rect 18512 34595 18564 34604
rect 15476 34416 15528 34468
rect 16212 34484 16264 34536
rect 18512 34561 18521 34595
rect 18521 34561 18555 34595
rect 18555 34561 18564 34595
rect 18512 34552 18564 34561
rect 18880 34595 18932 34604
rect 18880 34561 18889 34595
rect 18889 34561 18923 34595
rect 18923 34561 18932 34595
rect 18880 34552 18932 34561
rect 19340 34552 19392 34604
rect 19616 34620 19668 34672
rect 20168 34688 20220 34740
rect 21824 34688 21876 34740
rect 22652 34688 22704 34740
rect 24676 34731 24728 34740
rect 24676 34697 24685 34731
rect 24685 34697 24719 34731
rect 24719 34697 24728 34731
rect 24676 34688 24728 34697
rect 19524 34595 19576 34604
rect 19524 34561 19533 34595
rect 19533 34561 19567 34595
rect 19567 34561 19576 34595
rect 19524 34552 19576 34561
rect 19800 34595 19852 34604
rect 19800 34561 19809 34595
rect 19809 34561 19843 34595
rect 19843 34561 19852 34595
rect 19800 34552 19852 34561
rect 20444 34620 20496 34672
rect 20536 34620 20588 34672
rect 17868 34416 17920 34468
rect 19156 34484 19208 34536
rect 12900 34391 12952 34400
rect 12900 34357 12909 34391
rect 12909 34357 12943 34391
rect 12943 34357 12952 34391
rect 12900 34348 12952 34357
rect 18144 34348 18196 34400
rect 19248 34416 19300 34468
rect 20168 34484 20220 34536
rect 21180 34552 21232 34604
rect 22376 34595 22428 34604
rect 22376 34561 22385 34595
rect 22385 34561 22419 34595
rect 22419 34561 22428 34595
rect 22376 34552 22428 34561
rect 23848 34595 23900 34604
rect 23848 34561 23857 34595
rect 23857 34561 23891 34595
rect 23891 34561 23900 34595
rect 23848 34552 23900 34561
rect 24032 34552 24084 34604
rect 24492 34595 24544 34604
rect 24492 34561 24501 34595
rect 24501 34561 24535 34595
rect 24535 34561 24544 34595
rect 24492 34552 24544 34561
rect 24860 34552 24912 34604
rect 26608 34688 26660 34740
rect 28448 34731 28500 34740
rect 28448 34697 28457 34731
rect 28457 34697 28491 34731
rect 28491 34697 28500 34731
rect 28448 34688 28500 34697
rect 29000 34688 29052 34740
rect 29460 34688 29512 34740
rect 28724 34620 28776 34672
rect 26976 34595 27028 34604
rect 26976 34561 26985 34595
rect 26985 34561 27019 34595
rect 27019 34561 27028 34595
rect 26976 34552 27028 34561
rect 28172 34552 28224 34604
rect 28356 34552 28408 34604
rect 29092 34552 29144 34604
rect 24308 34416 24360 34468
rect 24676 34416 24728 34468
rect 29828 34484 29880 34536
rect 19524 34348 19576 34400
rect 21456 34348 21508 34400
rect 25228 34348 25280 34400
rect 27160 34391 27212 34400
rect 27160 34357 27169 34391
rect 27169 34357 27203 34391
rect 27203 34357 27212 34391
rect 27160 34348 27212 34357
rect 29276 34348 29328 34400
rect 5915 34246 5967 34298
rect 5979 34246 6031 34298
rect 6043 34246 6095 34298
rect 6107 34246 6159 34298
rect 6171 34246 6223 34298
rect 15846 34246 15898 34298
rect 15910 34246 15962 34298
rect 15974 34246 16026 34298
rect 16038 34246 16090 34298
rect 16102 34246 16154 34298
rect 25776 34246 25828 34298
rect 25840 34246 25892 34298
rect 25904 34246 25956 34298
rect 25968 34246 26020 34298
rect 26032 34246 26084 34298
rect 1400 34144 1452 34196
rect 11520 34144 11572 34196
rect 13176 34187 13228 34196
rect 13176 34153 13185 34187
rect 13185 34153 13219 34187
rect 13219 34153 13228 34187
rect 13176 34144 13228 34153
rect 17776 34144 17828 34196
rect 12256 34076 12308 34128
rect 16672 34076 16724 34128
rect 23664 34144 23716 34196
rect 24492 34144 24544 34196
rect 26608 34187 26660 34196
rect 26608 34153 26617 34187
rect 26617 34153 26651 34187
rect 26651 34153 26660 34187
rect 26608 34144 26660 34153
rect 29276 34144 29328 34196
rect 29920 34187 29972 34196
rect 29920 34153 29929 34187
rect 29929 34153 29963 34187
rect 29963 34153 29972 34187
rect 29920 34144 29972 34153
rect 30104 34187 30156 34196
rect 30104 34153 30113 34187
rect 30113 34153 30147 34187
rect 30147 34153 30156 34187
rect 30104 34144 30156 34153
rect 19156 34076 19208 34128
rect 15384 34051 15436 34060
rect 10232 33940 10284 33992
rect 10600 33940 10652 33992
rect 11244 33940 11296 33992
rect 12256 33983 12308 33992
rect 10048 33872 10100 33924
rect 12256 33949 12265 33983
rect 12265 33949 12299 33983
rect 12299 33949 12308 33983
rect 12256 33940 12308 33949
rect 15108 33940 15160 33992
rect 15384 34017 15393 34051
rect 15393 34017 15427 34051
rect 15427 34017 15436 34051
rect 15384 34008 15436 34017
rect 17776 34008 17828 34060
rect 18236 34051 18288 34060
rect 12716 33872 12768 33924
rect 15844 33872 15896 33924
rect 10232 33847 10284 33856
rect 10232 33813 10241 33847
rect 10241 33813 10275 33847
rect 10275 33813 10284 33847
rect 10232 33804 10284 33813
rect 11520 33804 11572 33856
rect 16672 33872 16724 33924
rect 17684 33940 17736 33992
rect 17868 33940 17920 33992
rect 18236 34017 18245 34051
rect 18245 34017 18279 34051
rect 18279 34017 18288 34051
rect 18236 34008 18288 34017
rect 29092 34076 29144 34128
rect 25228 34051 25280 34060
rect 25228 34017 25237 34051
rect 25237 34017 25271 34051
rect 25271 34017 25280 34051
rect 25228 34008 25280 34017
rect 26884 34008 26936 34060
rect 18328 33940 18380 33992
rect 19248 33940 19300 33992
rect 19524 33983 19576 33992
rect 19524 33949 19533 33983
rect 19533 33949 19567 33983
rect 19567 33949 19576 33983
rect 19524 33940 19576 33949
rect 19800 33940 19852 33992
rect 20444 33940 20496 33992
rect 21272 33940 21324 33992
rect 22284 33940 22336 33992
rect 24860 33940 24912 33992
rect 27068 33983 27120 33992
rect 27068 33949 27077 33983
rect 27077 33949 27111 33983
rect 27111 33949 27120 33983
rect 27068 33940 27120 33949
rect 16764 33847 16816 33856
rect 16764 33813 16773 33847
rect 16773 33813 16807 33847
rect 16807 33813 16816 33847
rect 16764 33804 16816 33813
rect 17592 33804 17644 33856
rect 18512 33804 18564 33856
rect 19248 33847 19300 33856
rect 19248 33813 19257 33847
rect 19257 33813 19291 33847
rect 19291 33813 19300 33847
rect 19248 33804 19300 33813
rect 19340 33804 19392 33856
rect 19616 33804 19668 33856
rect 20076 33847 20128 33856
rect 20076 33813 20085 33847
rect 20085 33813 20119 33847
rect 20119 33813 20128 33847
rect 20076 33804 20128 33813
rect 21456 33915 21508 33924
rect 21456 33881 21490 33915
rect 21490 33881 21508 33915
rect 21456 33872 21508 33881
rect 24400 33872 24452 33924
rect 24952 33872 25004 33924
rect 26148 33872 26200 33924
rect 26332 33872 26384 33924
rect 27436 33872 27488 33924
rect 22560 33847 22612 33856
rect 22560 33813 22569 33847
rect 22569 33813 22603 33847
rect 22603 33813 22612 33847
rect 22560 33804 22612 33813
rect 22744 33804 22796 33856
rect 27620 33804 27672 33856
rect 27988 33940 28040 33992
rect 28632 33872 28684 33924
rect 28724 33804 28776 33856
rect 28908 33847 28960 33856
rect 28908 33813 28917 33847
rect 28917 33813 28951 33847
rect 28951 33813 28960 33847
rect 28908 33804 28960 33813
rect 10880 33702 10932 33754
rect 10944 33702 10996 33754
rect 11008 33702 11060 33754
rect 11072 33702 11124 33754
rect 11136 33702 11188 33754
rect 20811 33702 20863 33754
rect 20875 33702 20927 33754
rect 20939 33702 20991 33754
rect 21003 33702 21055 33754
rect 21067 33702 21119 33754
rect 1400 33643 1452 33652
rect 1400 33609 1409 33643
rect 1409 33609 1443 33643
rect 1443 33609 1452 33643
rect 1400 33600 1452 33609
rect 11428 33600 11480 33652
rect 11888 33643 11940 33652
rect 11888 33609 11897 33643
rect 11897 33609 11931 33643
rect 11931 33609 11940 33643
rect 12716 33643 12768 33652
rect 11888 33600 11940 33609
rect 12716 33609 12725 33643
rect 12725 33609 12759 33643
rect 12759 33609 12768 33643
rect 12716 33600 12768 33609
rect 11520 33575 11572 33584
rect 11520 33541 11529 33575
rect 11529 33541 11563 33575
rect 11563 33541 11572 33575
rect 11520 33532 11572 33541
rect 1584 33507 1636 33516
rect 1584 33473 1593 33507
rect 1593 33473 1627 33507
rect 1627 33473 1636 33507
rect 1584 33464 1636 33473
rect 12072 33507 12124 33516
rect 9956 33396 10008 33448
rect 10324 33396 10376 33448
rect 12072 33473 12081 33507
rect 12081 33473 12115 33507
rect 12115 33473 12124 33507
rect 12072 33464 12124 33473
rect 14004 33600 14056 33652
rect 14556 33600 14608 33652
rect 17776 33600 17828 33652
rect 19708 33600 19760 33652
rect 20260 33600 20312 33652
rect 21456 33600 21508 33652
rect 22284 33643 22336 33652
rect 22284 33609 22293 33643
rect 22293 33609 22327 33643
rect 22327 33609 22336 33643
rect 22284 33600 22336 33609
rect 26148 33643 26200 33652
rect 26148 33609 26157 33643
rect 26157 33609 26191 33643
rect 26191 33609 26200 33643
rect 26148 33600 26200 33609
rect 15108 33532 15160 33584
rect 15292 33532 15344 33584
rect 10692 33328 10744 33380
rect 13360 33328 13412 33380
rect 15016 33507 15068 33516
rect 15016 33473 15025 33507
rect 15025 33473 15059 33507
rect 15059 33473 15068 33507
rect 15016 33464 15068 33473
rect 15476 33464 15528 33516
rect 16764 33532 16816 33584
rect 15844 33464 15896 33516
rect 16856 33507 16908 33516
rect 14464 33328 14516 33380
rect 15292 33439 15344 33448
rect 15292 33405 15301 33439
rect 15301 33405 15335 33439
rect 15335 33405 15344 33439
rect 15292 33396 15344 33405
rect 16856 33473 16865 33507
rect 16865 33473 16899 33507
rect 16899 33473 16908 33507
rect 16856 33464 16908 33473
rect 17776 33464 17828 33516
rect 17960 33507 18012 33516
rect 17960 33473 17969 33507
rect 17969 33473 18003 33507
rect 18003 33473 18012 33507
rect 17960 33464 18012 33473
rect 18512 33464 18564 33516
rect 19708 33464 19760 33516
rect 20720 33507 20772 33516
rect 20720 33473 20729 33507
rect 20729 33473 20763 33507
rect 20763 33473 20772 33507
rect 20720 33464 20772 33473
rect 20812 33507 20864 33516
rect 20812 33473 20821 33507
rect 20821 33473 20855 33507
rect 20855 33473 20864 33507
rect 22192 33532 22244 33584
rect 22560 33532 22612 33584
rect 27436 33600 27488 33652
rect 20812 33464 20864 33473
rect 22100 33507 22152 33516
rect 22100 33473 22109 33507
rect 22109 33473 22143 33507
rect 22143 33473 22152 33507
rect 22744 33507 22796 33516
rect 22100 33464 22152 33473
rect 22744 33473 22753 33507
rect 22753 33473 22787 33507
rect 22787 33473 22796 33507
rect 22744 33464 22796 33473
rect 22836 33464 22888 33516
rect 23572 33464 23624 33516
rect 24676 33464 24728 33516
rect 25504 33464 25556 33516
rect 26608 33464 26660 33516
rect 17684 33396 17736 33448
rect 22560 33396 22612 33448
rect 26884 33396 26936 33448
rect 9680 33303 9732 33312
rect 9680 33269 9689 33303
rect 9689 33269 9723 33303
rect 9723 33269 9732 33303
rect 9680 33260 9732 33269
rect 12256 33260 12308 33312
rect 12716 33260 12768 33312
rect 13268 33260 13320 33312
rect 15292 33260 15344 33312
rect 16212 33260 16264 33312
rect 17868 33328 17920 33380
rect 17408 33303 17460 33312
rect 17408 33269 17417 33303
rect 17417 33269 17451 33303
rect 17451 33269 17460 33303
rect 17408 33260 17460 33269
rect 24400 33260 24452 33312
rect 24860 33260 24912 33312
rect 25596 33260 25648 33312
rect 27712 33600 27764 33652
rect 28632 33643 28684 33652
rect 28632 33609 28641 33643
rect 28641 33609 28675 33643
rect 28675 33609 28684 33643
rect 28632 33600 28684 33609
rect 27804 33464 27856 33516
rect 29828 33507 29880 33516
rect 29828 33473 29837 33507
rect 29837 33473 29871 33507
rect 29871 33473 29880 33507
rect 29828 33464 29880 33473
rect 30012 33303 30064 33312
rect 30012 33269 30021 33303
rect 30021 33269 30055 33303
rect 30055 33269 30064 33303
rect 30012 33260 30064 33269
rect 5915 33158 5967 33210
rect 5979 33158 6031 33210
rect 6043 33158 6095 33210
rect 6107 33158 6159 33210
rect 6171 33158 6223 33210
rect 15846 33158 15898 33210
rect 15910 33158 15962 33210
rect 15974 33158 16026 33210
rect 16038 33158 16090 33210
rect 16102 33158 16154 33210
rect 25776 33158 25828 33210
rect 25840 33158 25892 33210
rect 25904 33158 25956 33210
rect 25968 33158 26020 33210
rect 26032 33158 26084 33210
rect 9956 33099 10008 33108
rect 9956 33065 9965 33099
rect 9965 33065 9999 33099
rect 9999 33065 10008 33099
rect 9956 33056 10008 33065
rect 10324 32988 10376 33040
rect 16304 33056 16356 33108
rect 16672 33056 16724 33108
rect 17132 33056 17184 33108
rect 17776 33099 17828 33108
rect 17776 33065 17785 33099
rect 17785 33065 17819 33099
rect 17819 33065 17828 33099
rect 17776 33056 17828 33065
rect 17960 32920 18012 32972
rect 19248 32920 19300 32972
rect 26976 33056 27028 33108
rect 24768 32988 24820 33040
rect 28264 33056 28316 33108
rect 28448 33056 28500 33108
rect 28724 33056 28776 33108
rect 25136 32920 25188 32972
rect 26240 32920 26292 32972
rect 26516 32920 26568 32972
rect 27160 32920 27212 32972
rect 9956 32852 10008 32904
rect 10232 32852 10284 32904
rect 10416 32895 10468 32904
rect 10416 32861 10425 32895
rect 10425 32861 10459 32895
rect 10459 32861 10468 32895
rect 10416 32852 10468 32861
rect 11244 32852 11296 32904
rect 11704 32895 11756 32904
rect 11704 32861 11713 32895
rect 11713 32861 11747 32895
rect 11747 32861 11756 32895
rect 11704 32852 11756 32861
rect 12072 32852 12124 32904
rect 13268 32852 13320 32904
rect 14188 32895 14240 32904
rect 14188 32861 14197 32895
rect 14197 32861 14231 32895
rect 14231 32861 14240 32895
rect 14188 32852 14240 32861
rect 11336 32827 11388 32836
rect 11336 32793 11345 32827
rect 11345 32793 11379 32827
rect 11379 32793 11388 32827
rect 11336 32784 11388 32793
rect 12992 32784 13044 32836
rect 15200 32784 15252 32836
rect 17408 32784 17460 32836
rect 19616 32852 19668 32904
rect 23480 32852 23532 32904
rect 24860 32852 24912 32904
rect 26148 32852 26200 32904
rect 28264 32852 28316 32904
rect 10600 32716 10652 32768
rect 11428 32759 11480 32768
rect 11428 32725 11437 32759
rect 11437 32725 11471 32759
rect 11471 32725 11480 32759
rect 11428 32716 11480 32725
rect 11888 32716 11940 32768
rect 12808 32716 12860 32768
rect 15016 32716 15068 32768
rect 16764 32716 16816 32768
rect 20720 32784 20772 32836
rect 21364 32784 21416 32836
rect 23112 32784 23164 32836
rect 27620 32784 27672 32836
rect 17960 32716 18012 32768
rect 18880 32716 18932 32768
rect 23388 32716 23440 32768
rect 25228 32716 25280 32768
rect 30104 32716 30156 32768
rect 10880 32614 10932 32666
rect 10944 32614 10996 32666
rect 11008 32614 11060 32666
rect 11072 32614 11124 32666
rect 11136 32614 11188 32666
rect 20811 32614 20863 32666
rect 20875 32614 20927 32666
rect 20939 32614 20991 32666
rect 21003 32614 21055 32666
rect 21067 32614 21119 32666
rect 11704 32555 11756 32564
rect 11704 32521 11713 32555
rect 11713 32521 11747 32555
rect 11747 32521 11756 32555
rect 11704 32512 11756 32521
rect 12992 32555 13044 32564
rect 12992 32521 13001 32555
rect 13001 32521 13035 32555
rect 13035 32521 13044 32555
rect 12992 32512 13044 32521
rect 15108 32512 15160 32564
rect 20720 32512 20772 32564
rect 21272 32555 21324 32564
rect 21272 32521 21281 32555
rect 21281 32521 21315 32555
rect 21315 32521 21324 32555
rect 21272 32512 21324 32521
rect 22100 32512 22152 32564
rect 22836 32555 22888 32564
rect 22836 32521 22845 32555
rect 22845 32521 22879 32555
rect 22879 32521 22888 32555
rect 22836 32512 22888 32521
rect 23480 32555 23532 32564
rect 23480 32521 23489 32555
rect 23489 32521 23523 32555
rect 23523 32521 23532 32555
rect 23480 32512 23532 32521
rect 27804 32512 27856 32564
rect 28172 32512 28224 32564
rect 13452 32444 13504 32496
rect 14004 32444 14056 32496
rect 11796 32376 11848 32428
rect 12348 32376 12400 32428
rect 12440 32419 12492 32428
rect 12440 32385 12449 32419
rect 12449 32385 12483 32419
rect 12483 32385 12492 32419
rect 12440 32376 12492 32385
rect 12808 32419 12860 32428
rect 10324 32351 10376 32360
rect 10324 32317 10333 32351
rect 10333 32317 10367 32351
rect 10367 32317 10376 32351
rect 10324 32308 10376 32317
rect 10692 32308 10744 32360
rect 11520 32308 11572 32360
rect 12808 32385 12817 32419
rect 12817 32385 12851 32419
rect 12851 32385 12860 32419
rect 12808 32376 12860 32385
rect 13360 32376 13412 32428
rect 14464 32419 14516 32428
rect 12624 32240 12676 32292
rect 14464 32385 14473 32419
rect 14473 32385 14507 32419
rect 14507 32385 14516 32419
rect 14464 32376 14516 32385
rect 15016 32419 15068 32428
rect 14280 32308 14332 32360
rect 15016 32385 15025 32419
rect 15025 32385 15059 32419
rect 15059 32385 15068 32419
rect 15016 32376 15068 32385
rect 15200 32419 15252 32428
rect 15200 32385 15209 32419
rect 15209 32385 15243 32419
rect 15243 32385 15252 32419
rect 15200 32376 15252 32385
rect 16212 32376 16264 32428
rect 17132 32419 17184 32428
rect 17132 32385 17141 32419
rect 17141 32385 17175 32419
rect 17175 32385 17184 32419
rect 17132 32376 17184 32385
rect 17776 32419 17828 32428
rect 17776 32385 17785 32419
rect 17785 32385 17819 32419
rect 17819 32385 17828 32419
rect 17776 32376 17828 32385
rect 19248 32419 19300 32428
rect 19248 32385 19257 32419
rect 19257 32385 19291 32419
rect 19291 32385 19300 32419
rect 19248 32376 19300 32385
rect 20076 32376 20128 32428
rect 23204 32444 23256 32496
rect 22100 32419 22152 32428
rect 14556 32240 14608 32292
rect 15476 32308 15528 32360
rect 22100 32385 22109 32419
rect 22109 32385 22143 32419
rect 22143 32385 22152 32419
rect 26884 32444 26936 32496
rect 27252 32444 27304 32496
rect 27712 32487 27764 32496
rect 22100 32376 22152 32385
rect 15292 32240 15344 32292
rect 15660 32240 15712 32292
rect 9588 32172 9640 32224
rect 13452 32172 13504 32224
rect 16856 32172 16908 32224
rect 19616 32172 19668 32224
rect 21364 32308 21416 32360
rect 20444 32240 20496 32292
rect 22560 32308 22612 32360
rect 23388 32376 23440 32428
rect 25596 32419 25648 32428
rect 25596 32385 25605 32419
rect 25605 32385 25639 32419
rect 25639 32385 25648 32419
rect 25596 32376 25648 32385
rect 26148 32376 26200 32428
rect 26424 32376 26476 32428
rect 27068 32376 27120 32428
rect 27160 32419 27212 32428
rect 27160 32385 27169 32419
rect 27169 32385 27203 32419
rect 27203 32385 27212 32419
rect 27712 32453 27721 32487
rect 27721 32453 27755 32487
rect 27755 32453 27764 32487
rect 27712 32444 27764 32453
rect 27160 32376 27212 32385
rect 28632 32444 28684 32496
rect 28724 32444 28776 32496
rect 28448 32419 28500 32428
rect 28448 32385 28457 32419
rect 28457 32385 28491 32419
rect 28491 32385 28500 32419
rect 28448 32376 28500 32385
rect 29184 32376 29236 32428
rect 24400 32308 24452 32360
rect 25504 32308 25556 32360
rect 26240 32240 26292 32292
rect 26884 32240 26936 32292
rect 27436 32308 27488 32360
rect 28908 32283 28960 32292
rect 28908 32249 28917 32283
rect 28917 32249 28951 32283
rect 28951 32249 28960 32283
rect 28908 32240 28960 32249
rect 24768 32215 24820 32224
rect 24768 32181 24777 32215
rect 24777 32181 24811 32215
rect 24811 32181 24820 32215
rect 24768 32172 24820 32181
rect 25688 32172 25740 32224
rect 26792 32172 26844 32224
rect 27160 32172 27212 32224
rect 29276 32215 29328 32224
rect 29276 32181 29285 32215
rect 29285 32181 29319 32215
rect 29319 32181 29328 32215
rect 29276 32172 29328 32181
rect 29828 32172 29880 32224
rect 5915 32070 5967 32122
rect 5979 32070 6031 32122
rect 6043 32070 6095 32122
rect 6107 32070 6159 32122
rect 6171 32070 6223 32122
rect 15846 32070 15898 32122
rect 15910 32070 15962 32122
rect 15974 32070 16026 32122
rect 16038 32070 16090 32122
rect 16102 32070 16154 32122
rect 25776 32070 25828 32122
rect 25840 32070 25892 32122
rect 25904 32070 25956 32122
rect 25968 32070 26020 32122
rect 26032 32070 26084 32122
rect 10324 31968 10376 32020
rect 11796 32011 11848 32020
rect 11796 31977 11805 32011
rect 11805 31977 11839 32011
rect 11839 31977 11848 32011
rect 11796 31968 11848 31977
rect 12348 31968 12400 32020
rect 15660 31968 15712 32020
rect 16304 31968 16356 32020
rect 23112 32011 23164 32020
rect 23112 31977 23121 32011
rect 23121 31977 23155 32011
rect 23155 31977 23164 32011
rect 23112 31968 23164 31977
rect 24676 32011 24728 32020
rect 24676 31977 24685 32011
rect 24685 31977 24719 32011
rect 24719 31977 24728 32011
rect 24676 31968 24728 31977
rect 24860 32011 24912 32020
rect 24860 31977 24869 32011
rect 24869 31977 24903 32011
rect 24903 31977 24912 32011
rect 24860 31968 24912 31977
rect 26148 31968 26200 32020
rect 26884 31968 26936 32020
rect 10232 31900 10284 31952
rect 10692 31832 10744 31884
rect 11888 31832 11940 31884
rect 12624 31832 12676 31884
rect 10416 31764 10468 31816
rect 10784 31764 10836 31816
rect 11244 31764 11296 31816
rect 11796 31764 11848 31816
rect 15016 31764 15068 31816
rect 15936 31764 15988 31816
rect 16672 31900 16724 31952
rect 18236 31900 18288 31952
rect 16948 31807 17000 31816
rect 12532 31696 12584 31748
rect 16948 31773 16957 31807
rect 16957 31773 16991 31807
rect 16991 31773 17000 31807
rect 16948 31764 17000 31773
rect 16764 31696 16816 31748
rect 18512 31832 18564 31884
rect 18328 31764 18380 31816
rect 21456 31900 21508 31952
rect 22928 31900 22980 31952
rect 26792 31900 26844 31952
rect 21364 31875 21416 31884
rect 21364 31841 21373 31875
rect 21373 31841 21407 31875
rect 21407 31841 21416 31875
rect 21364 31832 21416 31841
rect 22008 31832 22060 31884
rect 21272 31764 21324 31816
rect 22100 31764 22152 31816
rect 26332 31832 26384 31884
rect 26884 31832 26936 31884
rect 18604 31696 18656 31748
rect 19248 31696 19300 31748
rect 10508 31628 10560 31680
rect 15384 31628 15436 31680
rect 16948 31628 17000 31680
rect 17408 31628 17460 31680
rect 17868 31628 17920 31680
rect 22560 31628 22612 31680
rect 23388 31764 23440 31816
rect 23664 31807 23716 31816
rect 23664 31773 23673 31807
rect 23673 31773 23707 31807
rect 23707 31773 23716 31807
rect 23664 31764 23716 31773
rect 24400 31807 24452 31816
rect 24400 31773 24409 31807
rect 24409 31773 24443 31807
rect 24443 31773 24452 31807
rect 24400 31764 24452 31773
rect 25688 31764 25740 31816
rect 26424 31807 26476 31816
rect 26424 31773 26433 31807
rect 26433 31773 26467 31807
rect 26467 31773 26476 31807
rect 26424 31764 26476 31773
rect 26516 31696 26568 31748
rect 26792 31807 26844 31816
rect 26792 31773 26801 31807
rect 26801 31773 26835 31807
rect 26835 31773 26844 31807
rect 28264 31968 28316 32020
rect 28724 31900 28776 31952
rect 26792 31764 26844 31773
rect 27252 31764 27304 31816
rect 29000 31807 29052 31816
rect 29000 31773 29009 31807
rect 29009 31773 29043 31807
rect 29043 31773 29052 31807
rect 29000 31764 29052 31773
rect 30104 31696 30156 31748
rect 27436 31628 27488 31680
rect 30012 31671 30064 31680
rect 30012 31637 30021 31671
rect 30021 31637 30055 31671
rect 30055 31637 30064 31671
rect 30012 31628 30064 31637
rect 10880 31526 10932 31578
rect 10944 31526 10996 31578
rect 11008 31526 11060 31578
rect 11072 31526 11124 31578
rect 11136 31526 11188 31578
rect 20811 31526 20863 31578
rect 20875 31526 20927 31578
rect 20939 31526 20991 31578
rect 21003 31526 21055 31578
rect 21067 31526 21119 31578
rect 10416 31424 10468 31476
rect 10692 31424 10744 31476
rect 11336 31424 11388 31476
rect 12808 31467 12860 31476
rect 12808 31433 12817 31467
rect 12817 31433 12851 31467
rect 12851 31433 12860 31467
rect 12808 31424 12860 31433
rect 15936 31424 15988 31476
rect 23204 31467 23256 31476
rect 23204 31433 23213 31467
rect 23213 31433 23247 31467
rect 23247 31433 23256 31467
rect 23204 31424 23256 31433
rect 26148 31424 26200 31476
rect 12440 31356 12492 31408
rect 8208 31288 8260 31340
rect 8852 31331 8904 31340
rect 8852 31297 8886 31331
rect 8886 31297 8904 31331
rect 8852 31288 8904 31297
rect 10416 31288 10468 31340
rect 11520 31288 11572 31340
rect 11704 31288 11756 31340
rect 11796 31331 11848 31340
rect 11796 31297 11805 31331
rect 11805 31297 11839 31331
rect 11839 31297 11848 31331
rect 12900 31331 12952 31340
rect 11796 31288 11848 31297
rect 12900 31297 12909 31331
rect 12909 31297 12943 31331
rect 12943 31297 12952 31331
rect 12900 31288 12952 31297
rect 1400 31263 1452 31272
rect 1400 31229 1409 31263
rect 1409 31229 1443 31263
rect 1443 31229 1452 31263
rect 1400 31220 1452 31229
rect 9956 31195 10008 31204
rect 9956 31161 9965 31195
rect 9965 31161 9999 31195
rect 9999 31161 10008 31195
rect 9956 31152 10008 31161
rect 10508 31152 10560 31204
rect 10784 31220 10836 31272
rect 11888 31220 11940 31272
rect 13452 31356 13504 31408
rect 17684 31356 17736 31408
rect 15292 31288 15344 31340
rect 17960 31331 18012 31340
rect 13084 31220 13136 31272
rect 17960 31297 17969 31331
rect 17969 31297 18003 31331
rect 18003 31297 18012 31331
rect 17960 31288 18012 31297
rect 18236 31356 18288 31408
rect 20168 31356 20220 31408
rect 20720 31356 20772 31408
rect 21732 31356 21784 31408
rect 21916 31356 21968 31408
rect 18420 31288 18472 31340
rect 19064 31288 19116 31340
rect 19340 31331 19392 31340
rect 19340 31297 19354 31331
rect 19354 31297 19388 31331
rect 19388 31297 19392 31331
rect 19340 31288 19392 31297
rect 19708 31288 19760 31340
rect 22008 31331 22060 31340
rect 18144 31263 18196 31272
rect 11428 31152 11480 31204
rect 18144 31229 18153 31263
rect 18153 31229 18187 31263
rect 18187 31229 18196 31263
rect 18144 31220 18196 31229
rect 18512 31220 18564 31272
rect 22008 31297 22017 31331
rect 22017 31297 22051 31331
rect 22051 31297 22060 31331
rect 22008 31288 22060 31297
rect 26700 31356 26752 31408
rect 27068 31356 27120 31408
rect 27436 31399 27488 31408
rect 27436 31365 27470 31399
rect 27470 31365 27488 31399
rect 27436 31356 27488 31365
rect 28724 31424 28776 31476
rect 29000 31424 29052 31476
rect 22836 31288 22888 31340
rect 23572 31288 23624 31340
rect 27160 31331 27212 31340
rect 27160 31297 27169 31331
rect 27169 31297 27203 31331
rect 27203 31297 27212 31331
rect 27160 31288 27212 31297
rect 21916 31220 21968 31272
rect 22560 31220 22612 31272
rect 24032 31220 24084 31272
rect 24216 31263 24268 31272
rect 24216 31229 24225 31263
rect 24225 31229 24259 31263
rect 24259 31229 24268 31263
rect 24216 31220 24268 31229
rect 24860 31220 24912 31272
rect 25688 31263 25740 31272
rect 25688 31229 25697 31263
rect 25697 31229 25731 31263
rect 25731 31229 25740 31263
rect 25688 31220 25740 31229
rect 26056 31220 26108 31272
rect 28632 31152 28684 31204
rect 28908 31152 28960 31204
rect 10600 31127 10652 31136
rect 10600 31093 10609 31127
rect 10609 31093 10643 31127
rect 10643 31093 10652 31127
rect 10600 31084 10652 31093
rect 11888 31084 11940 31136
rect 16764 31084 16816 31136
rect 17960 31084 18012 31136
rect 18604 31084 18656 31136
rect 20352 31084 20404 31136
rect 21180 31127 21232 31136
rect 21180 31093 21189 31127
rect 21189 31093 21223 31127
rect 21223 31093 21232 31127
rect 21180 31084 21232 31093
rect 21364 31084 21416 31136
rect 23020 31084 23072 31136
rect 29092 31084 29144 31136
rect 29920 31084 29972 31136
rect 5915 30982 5967 31034
rect 5979 30982 6031 31034
rect 6043 30982 6095 31034
rect 6107 30982 6159 31034
rect 6171 30982 6223 31034
rect 15846 30982 15898 31034
rect 15910 30982 15962 31034
rect 15974 30982 16026 31034
rect 16038 30982 16090 31034
rect 16102 30982 16154 31034
rect 25776 30982 25828 31034
rect 25840 30982 25892 31034
rect 25904 30982 25956 31034
rect 25968 30982 26020 31034
rect 26032 30982 26084 31034
rect 10600 30880 10652 30932
rect 11980 30812 12032 30864
rect 12348 30812 12400 30864
rect 12716 30744 12768 30796
rect 14004 30744 14056 30796
rect 23664 30880 23716 30932
rect 17960 30812 18012 30864
rect 22836 30812 22888 30864
rect 11428 30719 11480 30728
rect 10048 30608 10100 30660
rect 11428 30685 11437 30719
rect 11437 30685 11471 30719
rect 11471 30685 11480 30719
rect 11428 30676 11480 30685
rect 11980 30676 12032 30728
rect 12256 30719 12308 30728
rect 12256 30685 12265 30719
rect 12265 30685 12299 30719
rect 12299 30685 12308 30719
rect 12256 30676 12308 30685
rect 13084 30719 13136 30728
rect 13084 30685 13093 30719
rect 13093 30685 13127 30719
rect 13127 30685 13136 30719
rect 13084 30676 13136 30685
rect 14372 30719 14424 30728
rect 14372 30685 14381 30719
rect 14381 30685 14415 30719
rect 14415 30685 14424 30719
rect 14372 30676 14424 30685
rect 12072 30608 12124 30660
rect 12440 30651 12492 30660
rect 12440 30617 12449 30651
rect 12449 30617 12483 30651
rect 12483 30617 12492 30651
rect 12440 30608 12492 30617
rect 9496 30540 9548 30592
rect 9772 30540 9824 30592
rect 10232 30540 10284 30592
rect 10416 30540 10468 30592
rect 11796 30540 11848 30592
rect 12992 30540 13044 30592
rect 16212 30608 16264 30660
rect 16856 30608 16908 30660
rect 17684 30744 17736 30796
rect 18144 30744 18196 30796
rect 20352 30787 20404 30796
rect 20352 30753 20361 30787
rect 20361 30753 20395 30787
rect 20395 30753 20404 30787
rect 20352 30744 20404 30753
rect 22008 30744 22060 30796
rect 17500 30608 17552 30660
rect 19340 30676 19392 30728
rect 21364 30676 21416 30728
rect 21456 30676 21508 30728
rect 21916 30676 21968 30728
rect 22560 30719 22612 30728
rect 22560 30685 22569 30719
rect 22569 30685 22603 30719
rect 22603 30685 22612 30719
rect 22560 30676 22612 30685
rect 23572 30719 23624 30728
rect 15200 30540 15252 30592
rect 17316 30540 17368 30592
rect 17960 30608 18012 30660
rect 18236 30651 18288 30660
rect 18236 30617 18245 30651
rect 18245 30617 18279 30651
rect 18279 30617 18288 30651
rect 18236 30608 18288 30617
rect 18420 30651 18472 30660
rect 18420 30617 18429 30651
rect 18429 30617 18463 30651
rect 18463 30617 18472 30651
rect 18420 30608 18472 30617
rect 18880 30608 18932 30660
rect 17776 30583 17828 30592
rect 17776 30549 17785 30583
rect 17785 30549 17819 30583
rect 17819 30549 17828 30583
rect 17776 30540 17828 30549
rect 20444 30608 20496 30660
rect 23572 30685 23581 30719
rect 23581 30685 23615 30719
rect 23615 30685 23624 30719
rect 23572 30676 23624 30685
rect 24584 30719 24636 30728
rect 24584 30685 24593 30719
rect 24593 30685 24627 30719
rect 24627 30685 24636 30719
rect 24584 30676 24636 30685
rect 26148 30880 26200 30932
rect 29920 30923 29972 30932
rect 29920 30889 29929 30923
rect 29929 30889 29963 30923
rect 29963 30889 29972 30923
rect 29920 30880 29972 30889
rect 30104 30923 30156 30932
rect 30104 30889 30113 30923
rect 30113 30889 30147 30923
rect 30147 30889 30156 30923
rect 30104 30880 30156 30889
rect 23480 30608 23532 30660
rect 25136 30608 25188 30660
rect 28356 30676 28408 30728
rect 28632 30676 28684 30728
rect 26516 30608 26568 30660
rect 27712 30608 27764 30660
rect 19892 30540 19944 30592
rect 22376 30540 22428 30592
rect 28172 30540 28224 30592
rect 28448 30583 28500 30592
rect 28448 30549 28457 30583
rect 28457 30549 28491 30583
rect 28491 30549 28500 30583
rect 28448 30540 28500 30549
rect 10880 30438 10932 30490
rect 10944 30438 10996 30490
rect 11008 30438 11060 30490
rect 11072 30438 11124 30490
rect 11136 30438 11188 30490
rect 20811 30438 20863 30490
rect 20875 30438 20927 30490
rect 20939 30438 20991 30490
rect 21003 30438 21055 30490
rect 21067 30438 21119 30490
rect 8852 30336 8904 30388
rect 10324 30336 10376 30388
rect 11244 30336 11296 30388
rect 12716 30379 12768 30388
rect 9772 30268 9824 30320
rect 8852 30243 8904 30252
rect 8852 30209 8861 30243
rect 8861 30209 8895 30243
rect 8895 30209 8904 30243
rect 8852 30200 8904 30209
rect 9312 30200 9364 30252
rect 10232 30200 10284 30252
rect 10324 30243 10376 30252
rect 10324 30209 10333 30243
rect 10333 30209 10367 30243
rect 10367 30209 10376 30243
rect 10324 30200 10376 30209
rect 10508 30200 10560 30252
rect 10600 30064 10652 30116
rect 12716 30345 12725 30379
rect 12725 30345 12759 30379
rect 12759 30345 12768 30379
rect 12716 30336 12768 30345
rect 12808 30336 12860 30388
rect 25136 30379 25188 30388
rect 12164 30268 12216 30320
rect 12624 30268 12676 30320
rect 16856 30268 16908 30320
rect 16948 30268 17000 30320
rect 11888 30243 11940 30252
rect 11888 30209 11897 30243
rect 11897 30209 11931 30243
rect 11931 30209 11940 30243
rect 11888 30200 11940 30209
rect 12072 30243 12124 30252
rect 12072 30209 12081 30243
rect 12081 30209 12115 30243
rect 12115 30209 12124 30243
rect 12072 30200 12124 30209
rect 14188 30200 14240 30252
rect 14740 30243 14792 30252
rect 14740 30209 14774 30243
rect 14774 30209 14792 30243
rect 14740 30200 14792 30209
rect 18144 30268 18196 30320
rect 25136 30345 25145 30379
rect 25145 30345 25179 30379
rect 25179 30345 25188 30379
rect 25136 30336 25188 30345
rect 28356 30379 28408 30388
rect 28356 30345 28365 30379
rect 28365 30345 28399 30379
rect 28399 30345 28408 30379
rect 28356 30336 28408 30345
rect 17316 30243 17368 30252
rect 17316 30209 17325 30243
rect 17325 30209 17359 30243
rect 17359 30209 17368 30243
rect 17592 30243 17644 30252
rect 17316 30200 17368 30209
rect 17592 30209 17601 30243
rect 17601 30209 17635 30243
rect 17635 30209 17644 30243
rect 17592 30200 17644 30209
rect 18236 30243 18288 30252
rect 18236 30209 18245 30243
rect 18245 30209 18279 30243
rect 18279 30209 18288 30243
rect 18236 30200 18288 30209
rect 18696 30200 18748 30252
rect 18788 30243 18840 30252
rect 18788 30209 18797 30243
rect 18797 30209 18831 30243
rect 18831 30209 18840 30243
rect 18788 30200 18840 30209
rect 19524 30200 19576 30252
rect 19800 30200 19852 30252
rect 20720 30243 20772 30252
rect 20720 30209 20729 30243
rect 20729 30209 20763 30243
rect 20763 30209 20772 30243
rect 20720 30200 20772 30209
rect 21364 30268 21416 30320
rect 21732 30268 21784 30320
rect 22376 30311 22428 30320
rect 22376 30277 22410 30311
rect 22410 30277 22428 30311
rect 22376 30268 22428 30277
rect 23756 30268 23808 30320
rect 24124 30200 24176 30252
rect 24216 30200 24268 30252
rect 25688 30268 25740 30320
rect 27712 30311 27764 30320
rect 13268 30132 13320 30184
rect 13636 30132 13688 30184
rect 16764 30132 16816 30184
rect 12716 30064 12768 30116
rect 19248 30132 19300 30184
rect 20168 30132 20220 30184
rect 20260 30132 20312 30184
rect 19432 30064 19484 30116
rect 20444 30064 20496 30116
rect 24860 30200 24912 30252
rect 26148 30200 26200 30252
rect 26424 30200 26476 30252
rect 27068 30200 27120 30252
rect 27712 30277 27721 30311
rect 27721 30277 27755 30311
rect 27755 30277 27764 30311
rect 27712 30268 27764 30277
rect 28448 30268 28500 30320
rect 28172 30243 28224 30252
rect 28172 30209 28181 30243
rect 28181 30209 28215 30243
rect 28215 30209 28224 30243
rect 28172 30200 28224 30209
rect 29000 30200 29052 30252
rect 24768 30175 24820 30184
rect 24768 30141 24777 30175
rect 24777 30141 24811 30175
rect 24811 30141 24820 30175
rect 24768 30132 24820 30141
rect 26792 30132 26844 30184
rect 26424 30064 26476 30116
rect 11980 29996 12032 30048
rect 13544 29996 13596 30048
rect 15200 29996 15252 30048
rect 15476 29996 15528 30048
rect 16948 29996 17000 30048
rect 17868 29996 17920 30048
rect 18512 29996 18564 30048
rect 20076 29996 20128 30048
rect 23480 30039 23532 30048
rect 23480 30005 23489 30039
rect 23489 30005 23523 30039
rect 23523 30005 23532 30039
rect 23480 29996 23532 30005
rect 23848 29996 23900 30048
rect 28080 29996 28132 30048
rect 30012 30039 30064 30048
rect 30012 30005 30021 30039
rect 30021 30005 30055 30039
rect 30055 30005 30064 30039
rect 30012 29996 30064 30005
rect 5915 29894 5967 29946
rect 5979 29894 6031 29946
rect 6043 29894 6095 29946
rect 6107 29894 6159 29946
rect 6171 29894 6223 29946
rect 15846 29894 15898 29946
rect 15910 29894 15962 29946
rect 15974 29894 16026 29946
rect 16038 29894 16090 29946
rect 16102 29894 16154 29946
rect 25776 29894 25828 29946
rect 25840 29894 25892 29946
rect 25904 29894 25956 29946
rect 25968 29894 26020 29946
rect 26032 29894 26084 29946
rect 8852 29792 8904 29844
rect 10232 29656 10284 29708
rect 10692 29656 10744 29708
rect 9312 29588 9364 29640
rect 9588 29631 9640 29640
rect 9588 29597 9594 29631
rect 9594 29597 9628 29631
rect 9628 29597 9640 29631
rect 10048 29631 10100 29640
rect 9588 29588 9640 29597
rect 10048 29597 10057 29631
rect 10057 29597 10091 29631
rect 10091 29597 10100 29631
rect 10048 29588 10100 29597
rect 10600 29588 10652 29640
rect 11520 29792 11572 29844
rect 14372 29792 14424 29844
rect 14740 29792 14792 29844
rect 15384 29792 15436 29844
rect 16488 29792 16540 29844
rect 18788 29792 18840 29844
rect 19708 29835 19760 29844
rect 19708 29801 19717 29835
rect 19717 29801 19751 29835
rect 19751 29801 19760 29835
rect 19708 29792 19760 29801
rect 22560 29792 22612 29844
rect 24584 29792 24636 29844
rect 11428 29724 11480 29776
rect 12808 29724 12860 29776
rect 11336 29631 11388 29640
rect 11336 29597 11344 29631
rect 11344 29597 11378 29631
rect 11378 29597 11388 29631
rect 11336 29588 11388 29597
rect 9864 29520 9916 29572
rect 12072 29588 12124 29640
rect 11980 29520 12032 29572
rect 8392 29452 8444 29504
rect 9772 29452 9824 29504
rect 10784 29452 10836 29504
rect 11428 29452 11480 29504
rect 12992 29631 13044 29640
rect 12992 29597 13002 29631
rect 13002 29597 13036 29631
rect 13036 29597 13044 29631
rect 12992 29588 13044 29597
rect 13176 29631 13228 29640
rect 13176 29597 13185 29631
rect 13185 29597 13219 29631
rect 13219 29597 13228 29631
rect 15476 29656 15528 29708
rect 13176 29588 13228 29597
rect 13544 29520 13596 29572
rect 15568 29588 15620 29640
rect 15660 29588 15712 29640
rect 16028 29631 16080 29640
rect 16028 29597 16037 29631
rect 16037 29597 16071 29631
rect 16071 29597 16080 29631
rect 16028 29588 16080 29597
rect 16120 29588 16172 29640
rect 17868 29656 17920 29708
rect 16764 29631 16816 29640
rect 16764 29597 16773 29631
rect 16773 29597 16807 29631
rect 16807 29597 16816 29631
rect 16764 29588 16816 29597
rect 14924 29520 14976 29572
rect 14096 29452 14148 29504
rect 15200 29452 15252 29504
rect 16856 29452 16908 29504
rect 18144 29588 18196 29640
rect 17224 29452 17276 29504
rect 19156 29724 19208 29776
rect 24768 29724 24820 29776
rect 24860 29724 24912 29776
rect 23848 29699 23900 29708
rect 23848 29665 23857 29699
rect 23857 29665 23891 29699
rect 23891 29665 23900 29699
rect 23848 29656 23900 29665
rect 24952 29656 25004 29708
rect 19432 29588 19484 29640
rect 20352 29588 20404 29640
rect 21272 29588 21324 29640
rect 22928 29631 22980 29640
rect 21364 29520 21416 29572
rect 19524 29452 19576 29504
rect 20720 29452 20772 29504
rect 22928 29597 22937 29631
rect 22937 29597 22971 29631
rect 22971 29597 22980 29631
rect 22928 29588 22980 29597
rect 24676 29588 24728 29640
rect 27344 29792 27396 29844
rect 29000 29835 29052 29844
rect 29000 29801 29009 29835
rect 29009 29801 29043 29835
rect 29043 29801 29052 29835
rect 29000 29792 29052 29801
rect 30104 29792 30156 29844
rect 29092 29724 29144 29776
rect 24952 29520 25004 29572
rect 27160 29588 27212 29640
rect 28632 29588 28684 29640
rect 29828 29631 29880 29640
rect 29828 29597 29837 29631
rect 29837 29597 29871 29631
rect 29871 29597 29880 29631
rect 29828 29588 29880 29597
rect 25504 29520 25556 29572
rect 27344 29520 27396 29572
rect 21732 29452 21784 29504
rect 22744 29452 22796 29504
rect 23756 29452 23808 29504
rect 25044 29452 25096 29504
rect 26424 29452 26476 29504
rect 27436 29495 27488 29504
rect 27436 29461 27445 29495
rect 27445 29461 27479 29495
rect 27479 29461 27488 29495
rect 27436 29452 27488 29461
rect 10880 29350 10932 29402
rect 10944 29350 10996 29402
rect 11008 29350 11060 29402
rect 11072 29350 11124 29402
rect 11136 29350 11188 29402
rect 20811 29350 20863 29402
rect 20875 29350 20927 29402
rect 20939 29350 20991 29402
rect 21003 29350 21055 29402
rect 21067 29350 21119 29402
rect 9772 29248 9824 29300
rect 11244 29248 11296 29300
rect 12256 29248 12308 29300
rect 13176 29248 13228 29300
rect 16120 29291 16172 29300
rect 16120 29257 16129 29291
rect 16129 29257 16163 29291
rect 16163 29257 16172 29291
rect 16120 29248 16172 29257
rect 16764 29248 16816 29300
rect 20260 29291 20312 29300
rect 2320 29112 2372 29164
rect 7840 29180 7892 29232
rect 10140 29180 10192 29232
rect 12440 29180 12492 29232
rect 14188 29223 14240 29232
rect 14188 29189 14197 29223
rect 14197 29189 14231 29223
rect 14231 29189 14240 29223
rect 14188 29180 14240 29189
rect 18236 29180 18288 29232
rect 20260 29257 20269 29291
rect 20269 29257 20303 29291
rect 20303 29257 20312 29291
rect 20260 29248 20312 29257
rect 25504 29291 25556 29300
rect 25504 29257 25513 29291
rect 25513 29257 25547 29291
rect 25547 29257 25556 29291
rect 25504 29248 25556 29257
rect 27160 29291 27212 29300
rect 8392 29112 8444 29164
rect 9680 29112 9732 29164
rect 10692 29155 10744 29164
rect 10692 29121 10701 29155
rect 10701 29121 10735 29155
rect 10735 29121 10744 29155
rect 10692 29112 10744 29121
rect 10784 29155 10836 29164
rect 10784 29121 10793 29155
rect 10793 29121 10827 29155
rect 10827 29121 10836 29155
rect 11520 29155 11572 29164
rect 10784 29112 10836 29121
rect 11520 29121 11529 29155
rect 11529 29121 11563 29155
rect 11563 29121 11572 29155
rect 11520 29112 11572 29121
rect 8300 29087 8352 29096
rect 8300 29053 8309 29087
rect 8309 29053 8343 29087
rect 8343 29053 8352 29087
rect 8300 29044 8352 29053
rect 9312 29044 9364 29096
rect 11152 29044 11204 29096
rect 11336 29044 11388 29096
rect 11796 29155 11848 29164
rect 11796 29121 11805 29155
rect 11805 29121 11839 29155
rect 11839 29121 11848 29155
rect 12072 29155 12124 29164
rect 11796 29112 11848 29121
rect 12072 29121 12081 29155
rect 12081 29121 12115 29155
rect 12115 29121 12124 29155
rect 12072 29112 12124 29121
rect 12624 29112 12676 29164
rect 11888 29087 11940 29096
rect 11888 29053 11897 29087
rect 11897 29053 11931 29087
rect 11931 29053 11940 29087
rect 11888 29044 11940 29053
rect 13268 29044 13320 29096
rect 13636 29044 13688 29096
rect 1584 29019 1636 29028
rect 1584 28985 1593 29019
rect 1593 28985 1627 29019
rect 1627 28985 1636 29019
rect 1584 28976 1636 28985
rect 9864 28976 9916 29028
rect 11796 28976 11848 29028
rect 11980 28976 12032 29028
rect 12808 28976 12860 29028
rect 14924 29112 14976 29164
rect 15476 29112 15528 29164
rect 16856 29112 16908 29164
rect 17224 29112 17276 29164
rect 18052 29112 18104 29164
rect 19432 29155 19484 29164
rect 16764 29044 16816 29096
rect 19432 29121 19441 29155
rect 19441 29121 19475 29155
rect 19475 29121 19484 29155
rect 19432 29112 19484 29121
rect 20076 29155 20128 29164
rect 20076 29121 20085 29155
rect 20085 29121 20119 29155
rect 20119 29121 20128 29155
rect 20076 29112 20128 29121
rect 21180 29112 21232 29164
rect 23664 29180 23716 29232
rect 24492 29180 24544 29232
rect 22100 29112 22152 29164
rect 16488 28976 16540 29028
rect 19156 28976 19208 29028
rect 24216 29112 24268 29164
rect 24676 29112 24728 29164
rect 24860 29044 24912 29096
rect 21180 28976 21232 29028
rect 23388 29019 23440 29028
rect 23388 28985 23397 29019
rect 23397 28985 23431 29019
rect 23431 28985 23440 29019
rect 23388 28976 23440 28985
rect 7932 28908 7984 28960
rect 10600 28908 10652 28960
rect 15384 28908 15436 28960
rect 16672 28908 16724 28960
rect 19984 28908 20036 28960
rect 22284 28908 22336 28960
rect 23848 28908 23900 28960
rect 24584 28976 24636 29028
rect 24768 28976 24820 29028
rect 27160 29257 27169 29291
rect 27169 29257 27203 29291
rect 27203 29257 27212 29291
rect 27160 29248 27212 29257
rect 27436 29248 27488 29300
rect 29184 29291 29236 29300
rect 29184 29257 29193 29291
rect 29193 29257 29227 29291
rect 29227 29257 29236 29291
rect 29184 29248 29236 29257
rect 27068 29112 27120 29164
rect 28632 29155 28684 29164
rect 28632 29121 28641 29155
rect 28641 29121 28675 29155
rect 28675 29121 28684 29155
rect 28632 29112 28684 29121
rect 27436 29044 27488 29096
rect 27528 29044 27580 29096
rect 26516 28976 26568 29028
rect 30012 29019 30064 29028
rect 30012 28985 30021 29019
rect 30021 28985 30055 29019
rect 30055 28985 30064 29019
rect 30012 28976 30064 28985
rect 29092 28908 29144 28960
rect 5915 28806 5967 28858
rect 5979 28806 6031 28858
rect 6043 28806 6095 28858
rect 6107 28806 6159 28858
rect 6171 28806 6223 28858
rect 15846 28806 15898 28858
rect 15910 28806 15962 28858
rect 15974 28806 16026 28858
rect 16038 28806 16090 28858
rect 16102 28806 16154 28858
rect 25776 28806 25828 28858
rect 25840 28806 25892 28858
rect 25904 28806 25956 28858
rect 25968 28806 26020 28858
rect 26032 28806 26084 28858
rect 8300 28704 8352 28756
rect 10324 28704 10376 28756
rect 11428 28704 11480 28756
rect 12256 28704 12308 28756
rect 22928 28747 22980 28756
rect 11520 28636 11572 28688
rect 14096 28636 14148 28688
rect 8208 28568 8260 28620
rect 18420 28636 18472 28688
rect 22928 28713 22937 28747
rect 22937 28713 22971 28747
rect 22971 28713 22980 28747
rect 22928 28704 22980 28713
rect 24860 28747 24912 28756
rect 24860 28713 24869 28747
rect 24869 28713 24903 28747
rect 24903 28713 24912 28747
rect 24860 28704 24912 28713
rect 27344 28747 27396 28756
rect 27344 28713 27353 28747
rect 27353 28713 27387 28747
rect 27387 28713 27396 28747
rect 27344 28704 27396 28713
rect 18880 28568 18932 28620
rect 21272 28568 21324 28620
rect 21732 28611 21784 28620
rect 7932 28543 7984 28552
rect 7932 28509 7941 28543
rect 7941 28509 7975 28543
rect 7975 28509 7984 28543
rect 7932 28500 7984 28509
rect 9864 28543 9916 28552
rect 9864 28509 9873 28543
rect 9873 28509 9907 28543
rect 9907 28509 9916 28543
rect 9864 28500 9916 28509
rect 11796 28500 11848 28552
rect 12164 28500 12216 28552
rect 13912 28500 13964 28552
rect 10600 28432 10652 28484
rect 12440 28432 12492 28484
rect 14740 28500 14792 28552
rect 15568 28543 15620 28552
rect 15108 28432 15160 28484
rect 15568 28509 15577 28543
rect 15577 28509 15611 28543
rect 15611 28509 15620 28543
rect 15568 28500 15620 28509
rect 16672 28500 16724 28552
rect 16856 28543 16908 28552
rect 16856 28509 16865 28543
rect 16865 28509 16899 28543
rect 16899 28509 16908 28543
rect 16856 28500 16908 28509
rect 17868 28432 17920 28484
rect 18236 28500 18288 28552
rect 19064 28500 19116 28552
rect 19156 28500 19208 28552
rect 19340 28500 19392 28552
rect 21456 28500 21508 28552
rect 21732 28577 21741 28611
rect 21741 28577 21775 28611
rect 21775 28577 21784 28611
rect 21732 28568 21784 28577
rect 21640 28543 21692 28552
rect 21640 28509 21649 28543
rect 21649 28509 21683 28543
rect 21683 28509 21692 28543
rect 21640 28500 21692 28509
rect 23388 28568 23440 28620
rect 22192 28500 22244 28552
rect 23664 28543 23716 28552
rect 23664 28509 23673 28543
rect 23673 28509 23707 28543
rect 23707 28509 23716 28543
rect 23664 28500 23716 28509
rect 24768 28543 24820 28552
rect 24768 28509 24777 28543
rect 24777 28509 24811 28543
rect 24811 28509 24820 28543
rect 24768 28500 24820 28509
rect 26516 28500 26568 28552
rect 29828 28543 29880 28552
rect 29828 28509 29837 28543
rect 29837 28509 29871 28543
rect 29871 28509 29880 28543
rect 29828 28500 29880 28509
rect 10048 28364 10100 28416
rect 10692 28407 10744 28416
rect 10692 28373 10717 28407
rect 10717 28373 10744 28407
rect 11520 28407 11572 28416
rect 10692 28364 10744 28373
rect 11520 28373 11529 28407
rect 11529 28373 11563 28407
rect 11563 28373 11572 28407
rect 11520 28364 11572 28373
rect 11704 28364 11756 28416
rect 12256 28407 12308 28416
rect 12256 28373 12265 28407
rect 12265 28373 12299 28407
rect 12299 28373 12308 28407
rect 12256 28364 12308 28373
rect 14832 28364 14884 28416
rect 17316 28364 17368 28416
rect 18788 28364 18840 28416
rect 19515 28475 19567 28484
rect 19515 28441 19524 28475
rect 19524 28441 19558 28475
rect 19558 28441 19567 28475
rect 19515 28432 19567 28441
rect 26424 28432 26476 28484
rect 19340 28364 19392 28416
rect 19892 28364 19944 28416
rect 22100 28407 22152 28416
rect 22100 28373 22109 28407
rect 22109 28373 22143 28407
rect 22143 28373 22152 28407
rect 22100 28364 22152 28373
rect 23848 28364 23900 28416
rect 24124 28364 24176 28416
rect 25044 28364 25096 28416
rect 30012 28407 30064 28416
rect 30012 28373 30021 28407
rect 30021 28373 30055 28407
rect 30055 28373 30064 28407
rect 30012 28364 30064 28373
rect 10880 28262 10932 28314
rect 10944 28262 10996 28314
rect 11008 28262 11060 28314
rect 11072 28262 11124 28314
rect 11136 28262 11188 28314
rect 20811 28262 20863 28314
rect 20875 28262 20927 28314
rect 20939 28262 20991 28314
rect 21003 28262 21055 28314
rect 21067 28262 21119 28314
rect 9956 28160 10008 28212
rect 16672 28160 16724 28212
rect 17316 28160 17368 28212
rect 17868 28203 17920 28212
rect 11888 28092 11940 28144
rect 7840 28024 7892 28076
rect 10508 28024 10560 28076
rect 15200 28092 15252 28144
rect 15752 28092 15804 28144
rect 17868 28169 17877 28203
rect 17877 28169 17911 28203
rect 17911 28169 17920 28203
rect 17868 28160 17920 28169
rect 19248 28160 19300 28212
rect 13268 28024 13320 28076
rect 14188 28024 14240 28076
rect 10140 27999 10192 28008
rect 10140 27965 10149 27999
rect 10149 27965 10183 27999
rect 10183 27965 10192 27999
rect 10140 27956 10192 27965
rect 10600 27956 10652 28008
rect 17592 28024 17644 28076
rect 18420 28024 18472 28076
rect 17868 27956 17920 28008
rect 17316 27888 17368 27940
rect 18972 28092 19024 28144
rect 19524 28160 19576 28212
rect 21640 28160 21692 28212
rect 24124 28160 24176 28212
rect 19064 28067 19116 28076
rect 19064 28033 19073 28067
rect 19073 28033 19107 28067
rect 19107 28033 19116 28067
rect 19064 28024 19116 28033
rect 19892 28024 19944 28076
rect 20812 28092 20864 28144
rect 21272 28092 21324 28144
rect 20352 27999 20404 28008
rect 20352 27965 20361 27999
rect 20361 27965 20395 27999
rect 20395 27965 20404 27999
rect 20352 27956 20404 27965
rect 20720 28024 20772 28076
rect 21456 28024 21508 28076
rect 22284 28024 22336 28076
rect 22560 28024 22612 28076
rect 23480 28024 23532 28076
rect 24952 28160 25004 28212
rect 27068 28160 27120 28212
rect 24492 28092 24544 28144
rect 24860 28067 24912 28076
rect 21732 27956 21784 28008
rect 21916 27956 21968 28008
rect 23572 27956 23624 28008
rect 24860 28033 24869 28067
rect 24869 28033 24903 28067
rect 24903 28033 24912 28067
rect 24860 28024 24912 28033
rect 19340 27888 19392 27940
rect 22284 27888 22336 27940
rect 8024 27820 8076 27872
rect 9772 27820 9824 27872
rect 11796 27820 11848 27872
rect 14280 27820 14332 27872
rect 15292 27820 15344 27872
rect 19064 27820 19116 27872
rect 19800 27820 19852 27872
rect 22468 27820 22520 27872
rect 22652 27820 22704 27872
rect 22928 27820 22980 27872
rect 23940 27820 23992 27872
rect 30012 27863 30064 27872
rect 30012 27829 30021 27863
rect 30021 27829 30055 27863
rect 30055 27829 30064 27863
rect 30012 27820 30064 27829
rect 5915 27718 5967 27770
rect 5979 27718 6031 27770
rect 6043 27718 6095 27770
rect 6107 27718 6159 27770
rect 6171 27718 6223 27770
rect 15846 27718 15898 27770
rect 15910 27718 15962 27770
rect 15974 27718 16026 27770
rect 16038 27718 16090 27770
rect 16102 27718 16154 27770
rect 25776 27718 25828 27770
rect 25840 27718 25892 27770
rect 25904 27718 25956 27770
rect 25968 27718 26020 27770
rect 26032 27718 26084 27770
rect 12072 27616 12124 27668
rect 14740 27616 14792 27668
rect 15568 27616 15620 27668
rect 16672 27616 16724 27668
rect 18420 27616 18472 27668
rect 9956 27548 10008 27600
rect 11428 27548 11480 27600
rect 10048 27480 10100 27532
rect 11244 27480 11296 27532
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 8024 27455 8076 27464
rect 8024 27421 8033 27455
rect 8033 27421 8067 27455
rect 8067 27421 8076 27455
rect 8024 27412 8076 27421
rect 10140 27412 10192 27464
rect 11888 27548 11940 27600
rect 14280 27548 14332 27600
rect 15200 27591 15252 27600
rect 15200 27557 15209 27591
rect 15209 27557 15243 27591
rect 15243 27557 15252 27591
rect 15200 27548 15252 27557
rect 15660 27548 15712 27600
rect 17684 27548 17736 27600
rect 20352 27616 20404 27668
rect 12256 27480 12308 27532
rect 14372 27480 14424 27532
rect 15292 27523 15344 27532
rect 9588 27387 9640 27396
rect 9588 27353 9597 27387
rect 9597 27353 9631 27387
rect 9631 27353 9640 27387
rect 9588 27344 9640 27353
rect 9864 27344 9916 27396
rect 10232 27344 10284 27396
rect 11428 27387 11480 27396
rect 11428 27353 11437 27387
rect 11437 27353 11471 27387
rect 11471 27353 11480 27387
rect 11428 27344 11480 27353
rect 12992 27412 13044 27464
rect 14740 27412 14792 27464
rect 12624 27344 12676 27396
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 7748 27276 7800 27328
rect 10508 27319 10560 27328
rect 10508 27285 10517 27319
rect 10517 27285 10551 27319
rect 10551 27285 10560 27319
rect 10508 27276 10560 27285
rect 10692 27276 10744 27328
rect 12072 27276 12124 27328
rect 13084 27319 13136 27328
rect 13084 27285 13093 27319
rect 13093 27285 13127 27319
rect 13127 27285 13136 27319
rect 13084 27276 13136 27285
rect 14464 27344 14516 27396
rect 15292 27489 15301 27523
rect 15301 27489 15335 27523
rect 15335 27489 15344 27523
rect 15292 27480 15344 27489
rect 16120 27455 16172 27464
rect 16120 27421 16129 27455
rect 16129 27421 16163 27455
rect 16163 27421 16172 27455
rect 16120 27412 16172 27421
rect 17868 27523 17920 27532
rect 17868 27489 17877 27523
rect 17877 27489 17911 27523
rect 17911 27489 17920 27523
rect 18236 27523 18288 27532
rect 17868 27480 17920 27489
rect 18236 27489 18245 27523
rect 18245 27489 18279 27523
rect 18279 27489 18288 27523
rect 18236 27480 18288 27489
rect 20076 27480 20128 27532
rect 20536 27480 20588 27532
rect 21456 27616 21508 27668
rect 22560 27659 22612 27668
rect 22560 27625 22569 27659
rect 22569 27625 22603 27659
rect 22603 27625 22612 27659
rect 22560 27616 22612 27625
rect 27528 27548 27580 27600
rect 17316 27412 17368 27464
rect 17684 27455 17736 27464
rect 17684 27421 17693 27455
rect 17693 27421 17727 27455
rect 17727 27421 17736 27455
rect 17684 27412 17736 27421
rect 18328 27412 18380 27464
rect 19432 27412 19484 27464
rect 19892 27455 19944 27464
rect 19892 27421 19901 27455
rect 19901 27421 19935 27455
rect 19935 27421 19944 27455
rect 19892 27412 19944 27421
rect 24860 27480 24912 27532
rect 23848 27455 23900 27464
rect 19708 27344 19760 27396
rect 20628 27344 20680 27396
rect 21272 27344 21324 27396
rect 22284 27344 22336 27396
rect 23848 27421 23857 27455
rect 23857 27421 23891 27455
rect 23891 27421 23900 27455
rect 23848 27412 23900 27421
rect 23940 27412 23992 27464
rect 25044 27455 25096 27464
rect 25044 27421 25053 27455
rect 25053 27421 25087 27455
rect 25087 27421 25096 27455
rect 25044 27412 25096 27421
rect 29828 27480 29880 27532
rect 25688 27455 25740 27464
rect 25688 27421 25697 27455
rect 25697 27421 25731 27455
rect 25731 27421 25740 27455
rect 25688 27412 25740 27421
rect 26332 27455 26384 27464
rect 15568 27319 15620 27328
rect 15568 27285 15577 27319
rect 15577 27285 15611 27319
rect 15611 27285 15620 27319
rect 15568 27276 15620 27285
rect 15752 27276 15804 27328
rect 16212 27276 16264 27328
rect 19064 27276 19116 27328
rect 25320 27344 25372 27396
rect 26332 27421 26341 27455
rect 26341 27421 26375 27455
rect 26375 27421 26384 27455
rect 26332 27412 26384 27421
rect 23940 27276 23992 27328
rect 24400 27319 24452 27328
rect 24400 27285 24409 27319
rect 24409 27285 24443 27319
rect 24443 27285 24452 27319
rect 24400 27276 24452 27285
rect 25136 27319 25188 27328
rect 25136 27285 25145 27319
rect 25145 27285 25179 27319
rect 25179 27285 25188 27319
rect 25136 27276 25188 27285
rect 10880 27174 10932 27226
rect 10944 27174 10996 27226
rect 11008 27174 11060 27226
rect 11072 27174 11124 27226
rect 11136 27174 11188 27226
rect 20811 27174 20863 27226
rect 20875 27174 20927 27226
rect 20939 27174 20991 27226
rect 21003 27174 21055 27226
rect 21067 27174 21119 27226
rect 10508 27072 10560 27124
rect 12992 27072 13044 27124
rect 13268 27115 13320 27124
rect 13268 27081 13277 27115
rect 13277 27081 13311 27115
rect 13311 27081 13320 27115
rect 13268 27072 13320 27081
rect 15016 27115 15068 27124
rect 9312 26979 9364 26988
rect 9312 26945 9321 26979
rect 9321 26945 9355 26979
rect 9355 26945 9364 26979
rect 9312 26936 9364 26945
rect 9956 26936 10008 26988
rect 10048 26936 10100 26988
rect 10692 26936 10744 26988
rect 10784 26936 10836 26988
rect 12440 26936 12492 26988
rect 14464 27004 14516 27056
rect 12808 26936 12860 26988
rect 13268 26936 13320 26988
rect 14280 26979 14332 26988
rect 8852 26868 8904 26920
rect 10508 26911 10560 26920
rect 10508 26877 10517 26911
rect 10517 26877 10551 26911
rect 10551 26877 10560 26911
rect 10508 26868 10560 26877
rect 1676 26800 1728 26852
rect 13084 26868 13136 26920
rect 12624 26843 12676 26852
rect 8944 26775 8996 26784
rect 8944 26741 8953 26775
rect 8953 26741 8987 26775
rect 8987 26741 8996 26775
rect 8944 26732 8996 26741
rect 10232 26732 10284 26784
rect 12624 26809 12633 26843
rect 12633 26809 12667 26843
rect 12667 26809 12676 26843
rect 12624 26800 12676 26809
rect 13728 26732 13780 26784
rect 13912 26775 13964 26784
rect 13912 26741 13921 26775
rect 13921 26741 13955 26775
rect 13955 26741 13964 26775
rect 13912 26732 13964 26741
rect 14280 26945 14289 26979
rect 14289 26945 14323 26979
rect 14323 26945 14332 26979
rect 14280 26936 14332 26945
rect 15016 27081 15025 27115
rect 15025 27081 15059 27115
rect 15059 27081 15068 27115
rect 15016 27072 15068 27081
rect 16120 27072 16172 27124
rect 17684 27072 17736 27124
rect 19156 27115 19208 27124
rect 19156 27081 19165 27115
rect 19165 27081 19199 27115
rect 19199 27081 19208 27115
rect 19156 27072 19208 27081
rect 21916 27072 21968 27124
rect 22100 27072 22152 27124
rect 22376 27115 22428 27124
rect 22376 27081 22385 27115
rect 22385 27081 22419 27115
rect 22419 27081 22428 27115
rect 22376 27072 22428 27081
rect 23572 27115 23624 27124
rect 23572 27081 23581 27115
rect 23581 27081 23615 27115
rect 23615 27081 23624 27115
rect 23572 27072 23624 27081
rect 23940 27115 23992 27124
rect 23940 27081 23949 27115
rect 23949 27081 23983 27115
rect 23983 27081 23992 27115
rect 23940 27072 23992 27081
rect 16856 26936 16908 26988
rect 18236 27004 18288 27056
rect 19892 27004 19944 27056
rect 20904 27004 20956 27056
rect 18880 26936 18932 26988
rect 20536 26979 20588 26988
rect 18236 26868 18288 26920
rect 18696 26868 18748 26920
rect 20536 26945 20545 26979
rect 20545 26945 20579 26979
rect 20579 26945 20588 26979
rect 20536 26936 20588 26945
rect 20628 26936 20680 26988
rect 23756 27004 23808 27056
rect 25136 27004 25188 27056
rect 20904 26911 20956 26920
rect 15200 26800 15252 26852
rect 18328 26843 18380 26852
rect 18328 26809 18337 26843
rect 18337 26809 18371 26843
rect 18371 26809 18380 26843
rect 18328 26800 18380 26809
rect 18880 26800 18932 26852
rect 20904 26877 20913 26911
rect 20913 26877 20947 26911
rect 20947 26877 20956 26911
rect 20904 26868 20956 26877
rect 21180 26936 21232 26988
rect 22468 26936 22520 26988
rect 24308 26936 24360 26988
rect 26240 26936 26292 26988
rect 21916 26868 21968 26920
rect 25412 26911 25464 26920
rect 20536 26800 20588 26852
rect 25412 26877 25421 26911
rect 25421 26877 25455 26911
rect 25455 26877 25464 26911
rect 25412 26868 25464 26877
rect 25504 26911 25556 26920
rect 25504 26877 25513 26911
rect 25513 26877 25547 26911
rect 25547 26877 25556 26911
rect 25504 26868 25556 26877
rect 24676 26800 24728 26852
rect 30012 26843 30064 26852
rect 30012 26809 30021 26843
rect 30021 26809 30055 26843
rect 30055 26809 30064 26843
rect 30012 26800 30064 26809
rect 14648 26732 14700 26784
rect 15292 26732 15344 26784
rect 15476 26732 15528 26784
rect 16304 26732 16356 26784
rect 21272 26775 21324 26784
rect 21272 26741 21281 26775
rect 21281 26741 21315 26775
rect 21315 26741 21324 26775
rect 21272 26732 21324 26741
rect 25688 26732 25740 26784
rect 5915 26630 5967 26682
rect 5979 26630 6031 26682
rect 6043 26630 6095 26682
rect 6107 26630 6159 26682
rect 6171 26630 6223 26682
rect 15846 26630 15898 26682
rect 15910 26630 15962 26682
rect 15974 26630 16026 26682
rect 16038 26630 16090 26682
rect 16102 26630 16154 26682
rect 25776 26630 25828 26682
rect 25840 26630 25892 26682
rect 25904 26630 25956 26682
rect 25968 26630 26020 26682
rect 26032 26630 26084 26682
rect 9588 26528 9640 26580
rect 11336 26528 11388 26580
rect 12808 26571 12860 26580
rect 12808 26537 12817 26571
rect 12817 26537 12851 26571
rect 12851 26537 12860 26571
rect 12808 26528 12860 26537
rect 9680 26460 9732 26512
rect 13912 26460 13964 26512
rect 15200 26528 15252 26580
rect 16856 26528 16908 26580
rect 17316 26528 17368 26580
rect 20076 26528 20128 26580
rect 21916 26571 21968 26580
rect 8944 26392 8996 26444
rect 13820 26392 13872 26444
rect 14280 26392 14332 26444
rect 9036 26367 9088 26376
rect 9036 26333 9045 26367
rect 9045 26333 9079 26367
rect 9079 26333 9088 26367
rect 9036 26324 9088 26333
rect 9128 26324 9180 26376
rect 11244 26324 11296 26376
rect 12164 26367 12216 26376
rect 12164 26333 12173 26367
rect 12173 26333 12207 26367
rect 12207 26333 12216 26367
rect 12164 26324 12216 26333
rect 12992 26367 13044 26376
rect 12992 26333 13001 26367
rect 13001 26333 13035 26367
rect 13035 26333 13044 26367
rect 12992 26324 13044 26333
rect 13176 26367 13228 26376
rect 13176 26333 13185 26367
rect 13185 26333 13219 26367
rect 13219 26333 13228 26367
rect 13176 26324 13228 26333
rect 15016 26392 15068 26444
rect 16028 26460 16080 26512
rect 21916 26537 21925 26571
rect 21925 26537 21959 26571
rect 21959 26537 21968 26571
rect 21916 26528 21968 26537
rect 22652 26571 22704 26580
rect 22652 26537 22661 26571
rect 22661 26537 22695 26571
rect 22695 26537 22704 26571
rect 22652 26528 22704 26537
rect 26332 26528 26384 26580
rect 14648 26367 14700 26376
rect 14648 26333 14657 26367
rect 14657 26333 14691 26367
rect 14691 26333 14700 26367
rect 15476 26367 15528 26376
rect 14648 26324 14700 26333
rect 15476 26333 15485 26367
rect 15485 26333 15519 26367
rect 15519 26333 15528 26367
rect 15476 26324 15528 26333
rect 18880 26392 18932 26444
rect 20536 26435 20588 26444
rect 20536 26401 20545 26435
rect 20545 26401 20579 26435
rect 20579 26401 20588 26435
rect 20536 26392 20588 26401
rect 23664 26392 23716 26444
rect 25504 26435 25556 26444
rect 25504 26401 25513 26435
rect 25513 26401 25547 26435
rect 25547 26401 25556 26435
rect 25504 26392 25556 26401
rect 17960 26324 18012 26376
rect 18420 26324 18472 26376
rect 19156 26324 19208 26376
rect 21180 26324 21232 26376
rect 22560 26324 22612 26376
rect 23572 26367 23624 26376
rect 23572 26333 23581 26367
rect 23581 26333 23615 26367
rect 23615 26333 23624 26367
rect 23572 26324 23624 26333
rect 25228 26367 25280 26376
rect 25228 26333 25237 26367
rect 25237 26333 25271 26367
rect 25271 26333 25280 26367
rect 25228 26324 25280 26333
rect 26792 26324 26844 26376
rect 29828 26367 29880 26376
rect 29828 26333 29837 26367
rect 29837 26333 29871 26367
rect 29871 26333 29880 26367
rect 29828 26324 29880 26333
rect 2228 26188 2280 26240
rect 10508 26231 10560 26240
rect 10508 26197 10517 26231
rect 10517 26197 10551 26231
rect 10551 26197 10560 26231
rect 13360 26256 13412 26308
rect 13728 26256 13780 26308
rect 15200 26256 15252 26308
rect 16488 26256 16540 26308
rect 16672 26256 16724 26308
rect 19524 26256 19576 26308
rect 20260 26256 20312 26308
rect 21272 26256 21324 26308
rect 24492 26256 24544 26308
rect 10508 26188 10560 26197
rect 15936 26188 15988 26240
rect 23480 26188 23532 26240
rect 30012 26231 30064 26240
rect 30012 26197 30021 26231
rect 30021 26197 30055 26231
rect 30055 26197 30064 26231
rect 30012 26188 30064 26197
rect 10880 26086 10932 26138
rect 10944 26086 10996 26138
rect 11008 26086 11060 26138
rect 11072 26086 11124 26138
rect 11136 26086 11188 26138
rect 20811 26086 20863 26138
rect 20875 26086 20927 26138
rect 20939 26086 20991 26138
rect 21003 26086 21055 26138
rect 21067 26086 21119 26138
rect 1400 25984 1452 26036
rect 2320 26027 2372 26036
rect 2320 25993 2329 26027
rect 2329 25993 2363 26027
rect 2363 25993 2372 26027
rect 2320 25984 2372 25993
rect 5264 25916 5316 25968
rect 1768 25891 1820 25900
rect 1768 25857 1777 25891
rect 1777 25857 1811 25891
rect 1811 25857 1820 25891
rect 1768 25848 1820 25857
rect 2228 25891 2280 25900
rect 2228 25857 2237 25891
rect 2237 25857 2271 25891
rect 2271 25857 2280 25891
rect 2228 25848 2280 25857
rect 9128 25891 9180 25900
rect 9128 25857 9137 25891
rect 9137 25857 9171 25891
rect 9171 25857 9180 25891
rect 9128 25848 9180 25857
rect 9220 25848 9272 25900
rect 13820 25984 13872 26036
rect 15936 25984 15988 26036
rect 18052 25984 18104 26036
rect 11152 25780 11204 25832
rect 11980 25823 12032 25832
rect 11980 25789 11989 25823
rect 11989 25789 12023 25823
rect 12023 25789 12032 25823
rect 11980 25780 12032 25789
rect 12992 25916 13044 25968
rect 15568 25916 15620 25968
rect 13084 25848 13136 25900
rect 13360 25848 13412 25900
rect 13728 25891 13780 25900
rect 12716 25780 12768 25832
rect 13728 25857 13737 25891
rect 13737 25857 13771 25891
rect 13771 25857 13780 25891
rect 13728 25848 13780 25857
rect 13820 25848 13872 25900
rect 14556 25848 14608 25900
rect 14924 25848 14976 25900
rect 15660 25780 15712 25832
rect 10600 25712 10652 25764
rect 12440 25712 12492 25764
rect 12900 25712 12952 25764
rect 13268 25712 13320 25764
rect 13912 25712 13964 25764
rect 15108 25712 15160 25764
rect 15476 25712 15528 25764
rect 16396 25780 16448 25832
rect 16856 25780 16908 25832
rect 17500 25848 17552 25900
rect 17868 25848 17920 25900
rect 18052 25891 18104 25900
rect 18052 25857 18061 25891
rect 18061 25857 18095 25891
rect 18095 25857 18104 25891
rect 18052 25848 18104 25857
rect 18972 25916 19024 25968
rect 18328 25780 18380 25832
rect 19156 25891 19208 25900
rect 19156 25857 19165 25891
rect 19165 25857 19199 25891
rect 19199 25857 19208 25891
rect 20076 25891 20128 25900
rect 19156 25848 19208 25857
rect 20076 25857 20085 25891
rect 20085 25857 20119 25891
rect 20119 25857 20128 25891
rect 20076 25848 20128 25857
rect 20628 25984 20680 26036
rect 20720 25984 20772 26036
rect 23572 25984 23624 26036
rect 24400 25984 24452 26036
rect 29828 25984 29880 26036
rect 20260 25959 20312 25968
rect 20260 25925 20269 25959
rect 20269 25925 20303 25959
rect 20303 25925 20312 25959
rect 20260 25916 20312 25925
rect 21916 25848 21968 25900
rect 22836 25848 22888 25900
rect 26700 25916 26752 25968
rect 23112 25848 23164 25900
rect 25320 25891 25372 25900
rect 25320 25857 25329 25891
rect 25329 25857 25363 25891
rect 25363 25857 25372 25891
rect 25320 25848 25372 25857
rect 24400 25823 24452 25832
rect 24400 25789 24409 25823
rect 24409 25789 24443 25823
rect 24443 25789 24452 25823
rect 24400 25780 24452 25789
rect 24676 25780 24728 25832
rect 26332 25780 26384 25832
rect 17592 25712 17644 25764
rect 17684 25712 17736 25764
rect 1308 25644 1360 25696
rect 9496 25644 9548 25696
rect 14004 25644 14056 25696
rect 16396 25644 16448 25696
rect 17500 25687 17552 25696
rect 17500 25653 17509 25687
rect 17509 25653 17543 25687
rect 17543 25653 17552 25687
rect 17500 25644 17552 25653
rect 18880 25687 18932 25696
rect 18880 25653 18889 25687
rect 18889 25653 18923 25687
rect 18923 25653 18932 25687
rect 18880 25644 18932 25653
rect 20352 25644 20404 25696
rect 20628 25712 20680 25764
rect 22192 25712 22244 25764
rect 21456 25644 21508 25696
rect 22652 25712 22704 25764
rect 22468 25687 22520 25696
rect 22468 25653 22477 25687
rect 22477 25653 22511 25687
rect 22511 25653 22520 25687
rect 22468 25644 22520 25653
rect 25044 25712 25096 25764
rect 27620 25755 27672 25764
rect 27620 25721 27629 25755
rect 27629 25721 27663 25755
rect 27663 25721 27672 25755
rect 27620 25712 27672 25721
rect 30012 25687 30064 25696
rect 30012 25653 30021 25687
rect 30021 25653 30055 25687
rect 30055 25653 30064 25687
rect 30012 25644 30064 25653
rect 5915 25542 5967 25594
rect 5979 25542 6031 25594
rect 6043 25542 6095 25594
rect 6107 25542 6159 25594
rect 6171 25542 6223 25594
rect 15846 25542 15898 25594
rect 15910 25542 15962 25594
rect 15974 25542 16026 25594
rect 16038 25542 16090 25594
rect 16102 25542 16154 25594
rect 25776 25542 25828 25594
rect 25840 25542 25892 25594
rect 25904 25542 25956 25594
rect 25968 25542 26020 25594
rect 26032 25542 26084 25594
rect 9036 25440 9088 25492
rect 13084 25440 13136 25492
rect 13728 25440 13780 25492
rect 19064 25440 19116 25492
rect 20720 25440 20772 25492
rect 23112 25483 23164 25492
rect 23112 25449 23121 25483
rect 23121 25449 23155 25483
rect 23155 25449 23164 25483
rect 23112 25440 23164 25449
rect 5264 25372 5316 25424
rect 10692 25304 10744 25356
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 11152 25279 11204 25288
rect 11152 25245 11161 25279
rect 11161 25245 11195 25279
rect 11195 25245 11204 25279
rect 11152 25236 11204 25245
rect 8852 25168 8904 25220
rect 9312 25168 9364 25220
rect 10048 25168 10100 25220
rect 10600 25168 10652 25220
rect 11980 25211 12032 25220
rect 11980 25177 11989 25211
rect 11989 25177 12023 25211
rect 12023 25177 12032 25211
rect 11980 25168 12032 25177
rect 13912 25372 13964 25424
rect 16856 25372 16908 25424
rect 18328 25372 18380 25424
rect 19156 25372 19208 25424
rect 13820 25304 13872 25356
rect 16396 25347 16448 25356
rect 16396 25313 16405 25347
rect 16405 25313 16439 25347
rect 16439 25313 16448 25347
rect 16396 25304 16448 25313
rect 13084 25279 13136 25288
rect 13084 25245 13093 25279
rect 13093 25245 13127 25279
rect 13127 25245 13136 25279
rect 13084 25236 13136 25245
rect 13912 25236 13964 25288
rect 14188 25236 14240 25288
rect 14740 25236 14792 25288
rect 16672 25304 16724 25356
rect 17776 25304 17828 25356
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 9956 25100 10008 25152
rect 10324 25100 10376 25152
rect 13084 25100 13136 25152
rect 14004 25168 14056 25220
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 17868 25236 17920 25288
rect 18880 25304 18932 25356
rect 18972 25236 19024 25288
rect 19524 25279 19576 25288
rect 19524 25245 19533 25279
rect 19533 25245 19567 25279
rect 19567 25245 19576 25279
rect 19524 25236 19576 25245
rect 17592 25168 17644 25220
rect 15476 25143 15528 25152
rect 15476 25109 15485 25143
rect 15485 25109 15519 25143
rect 15519 25109 15528 25143
rect 15476 25100 15528 25109
rect 15752 25100 15804 25152
rect 16304 25143 16356 25152
rect 16304 25109 16313 25143
rect 16313 25109 16347 25143
rect 16347 25109 16356 25143
rect 16304 25100 16356 25109
rect 16580 25100 16632 25152
rect 19432 25168 19484 25220
rect 20076 25168 20128 25220
rect 21456 25372 21508 25424
rect 25136 25372 25188 25424
rect 27528 25372 27580 25424
rect 21548 25304 21600 25356
rect 23296 25304 23348 25356
rect 24676 25304 24728 25356
rect 19340 25100 19392 25152
rect 19708 25143 19760 25152
rect 19708 25109 19717 25143
rect 19717 25109 19751 25143
rect 19751 25109 19760 25143
rect 19708 25100 19760 25109
rect 20352 25100 20404 25152
rect 23480 25279 23532 25288
rect 23480 25245 23489 25279
rect 23489 25245 23523 25279
rect 23523 25245 23532 25279
rect 23480 25236 23532 25245
rect 23756 25236 23808 25288
rect 21640 25168 21692 25220
rect 23112 25168 23164 25220
rect 25320 25236 25372 25288
rect 28908 25236 28960 25288
rect 25688 25168 25740 25220
rect 26240 25211 26292 25220
rect 26240 25177 26249 25211
rect 26249 25177 26283 25211
rect 26283 25177 26292 25211
rect 26240 25168 26292 25177
rect 26792 25211 26844 25220
rect 26792 25177 26801 25211
rect 26801 25177 26835 25211
rect 26835 25177 26844 25211
rect 26792 25168 26844 25177
rect 27620 25168 27672 25220
rect 28632 25168 28684 25220
rect 23572 25143 23624 25152
rect 23572 25109 23581 25143
rect 23581 25109 23615 25143
rect 23615 25109 23624 25143
rect 23572 25100 23624 25109
rect 25964 25100 26016 25152
rect 26884 25143 26936 25152
rect 26884 25109 26893 25143
rect 26893 25109 26927 25143
rect 26927 25109 26936 25143
rect 26884 25100 26936 25109
rect 28816 25143 28868 25152
rect 28816 25109 28825 25143
rect 28825 25109 28859 25143
rect 28859 25109 28868 25143
rect 28816 25100 28868 25109
rect 10880 24998 10932 25050
rect 10944 24998 10996 25050
rect 11008 24998 11060 25050
rect 11072 24998 11124 25050
rect 11136 24998 11188 25050
rect 20811 24998 20863 25050
rect 20875 24998 20927 25050
rect 20939 24998 20991 25050
rect 21003 24998 21055 25050
rect 21067 24998 21119 25050
rect 1400 24896 1452 24948
rect 9220 24896 9272 24948
rect 11980 24896 12032 24948
rect 13268 24896 13320 24948
rect 16856 24896 16908 24948
rect 18052 24896 18104 24948
rect 18880 24896 18932 24948
rect 19432 24939 19484 24948
rect 8852 24828 8904 24880
rect 9036 24828 9088 24880
rect 9312 24828 9364 24880
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 1768 24803 1820 24812
rect 1768 24769 1777 24803
rect 1777 24769 1811 24803
rect 1811 24769 1820 24803
rect 1768 24760 1820 24769
rect 2320 24760 2372 24812
rect 8668 24760 8720 24812
rect 9128 24803 9180 24812
rect 9128 24769 9137 24803
rect 9137 24769 9171 24803
rect 9171 24769 9180 24803
rect 9128 24760 9180 24769
rect 9772 24803 9824 24812
rect 9772 24769 9781 24803
rect 9781 24769 9815 24803
rect 9815 24769 9824 24803
rect 9772 24760 9824 24769
rect 10048 24828 10100 24880
rect 10416 24760 10468 24812
rect 10600 24803 10652 24812
rect 10600 24769 10609 24803
rect 10609 24769 10643 24803
rect 10643 24769 10652 24803
rect 10600 24760 10652 24769
rect 11244 24828 11296 24880
rect 11888 24828 11940 24880
rect 13728 24871 13780 24880
rect 13728 24837 13737 24871
rect 13737 24837 13771 24871
rect 13771 24837 13780 24871
rect 13728 24828 13780 24837
rect 14924 24828 14976 24880
rect 10048 24624 10100 24676
rect 13084 24760 13136 24812
rect 14464 24803 14516 24812
rect 10140 24599 10192 24608
rect 10140 24565 10149 24599
rect 10149 24565 10183 24599
rect 10183 24565 10192 24599
rect 10140 24556 10192 24565
rect 10784 24556 10836 24608
rect 13176 24624 13228 24676
rect 11796 24599 11848 24608
rect 11796 24565 11805 24599
rect 11805 24565 11839 24599
rect 11839 24565 11848 24599
rect 11796 24556 11848 24565
rect 12164 24556 12216 24608
rect 13452 24556 13504 24608
rect 14464 24769 14473 24803
rect 14473 24769 14507 24803
rect 14507 24769 14516 24803
rect 14464 24760 14516 24769
rect 17500 24828 17552 24880
rect 19432 24905 19441 24939
rect 19441 24905 19475 24939
rect 19475 24905 19484 24939
rect 19432 24896 19484 24905
rect 25228 24896 25280 24948
rect 25320 24828 25372 24880
rect 14832 24624 14884 24676
rect 18236 24803 18288 24812
rect 15568 24624 15620 24676
rect 18236 24769 18245 24803
rect 18245 24769 18279 24803
rect 18279 24769 18288 24803
rect 18236 24760 18288 24769
rect 18972 24760 19024 24812
rect 19156 24803 19208 24812
rect 19156 24769 19165 24803
rect 19165 24769 19199 24803
rect 19199 24769 19208 24803
rect 19156 24760 19208 24769
rect 19708 24760 19760 24812
rect 20444 24803 20496 24812
rect 20444 24769 20453 24803
rect 20453 24769 20487 24803
rect 20487 24769 20496 24803
rect 20444 24760 20496 24769
rect 22652 24803 22704 24812
rect 22652 24769 22661 24803
rect 22661 24769 22695 24803
rect 22695 24769 22704 24803
rect 22652 24760 22704 24769
rect 23664 24803 23716 24812
rect 23664 24769 23673 24803
rect 23673 24769 23707 24803
rect 23707 24769 23716 24803
rect 23664 24760 23716 24769
rect 24676 24803 24728 24812
rect 24676 24769 24685 24803
rect 24685 24769 24719 24803
rect 24719 24769 24728 24803
rect 24676 24760 24728 24769
rect 28356 24803 28408 24812
rect 17592 24692 17644 24744
rect 18052 24692 18104 24744
rect 19616 24692 19668 24744
rect 20720 24735 20772 24744
rect 20720 24701 20729 24735
rect 20729 24701 20763 24735
rect 20763 24701 20772 24735
rect 20720 24692 20772 24701
rect 22376 24692 22428 24744
rect 23296 24692 23348 24744
rect 23388 24692 23440 24744
rect 24860 24735 24912 24744
rect 24860 24701 24869 24735
rect 24869 24701 24903 24735
rect 24903 24701 24912 24735
rect 24860 24692 24912 24701
rect 15936 24624 15988 24676
rect 16488 24624 16540 24676
rect 19156 24624 19208 24676
rect 19432 24624 19484 24676
rect 24216 24624 24268 24676
rect 28356 24769 28365 24803
rect 28365 24769 28399 24803
rect 28399 24769 28408 24803
rect 28356 24760 28408 24769
rect 28540 24760 28592 24812
rect 25964 24692 26016 24744
rect 29828 24624 29880 24676
rect 30012 24667 30064 24676
rect 30012 24633 30021 24667
rect 30021 24633 30055 24667
rect 30055 24633 30064 24667
rect 30012 24624 30064 24633
rect 17500 24556 17552 24608
rect 19064 24599 19116 24608
rect 19064 24565 19073 24599
rect 19073 24565 19107 24599
rect 19107 24565 19116 24599
rect 19064 24556 19116 24565
rect 22928 24556 22980 24608
rect 23480 24599 23532 24608
rect 23480 24565 23489 24599
rect 23489 24565 23523 24599
rect 23523 24565 23532 24599
rect 23480 24556 23532 24565
rect 25044 24556 25096 24608
rect 28724 24556 28776 24608
rect 5915 24454 5967 24506
rect 5979 24454 6031 24506
rect 6043 24454 6095 24506
rect 6107 24454 6159 24506
rect 6171 24454 6223 24506
rect 15846 24454 15898 24506
rect 15910 24454 15962 24506
rect 15974 24454 16026 24506
rect 16038 24454 16090 24506
rect 16102 24454 16154 24506
rect 25776 24454 25828 24506
rect 25840 24454 25892 24506
rect 25904 24454 25956 24506
rect 25968 24454 26020 24506
rect 26032 24454 26084 24506
rect 8300 24352 8352 24404
rect 9128 24352 9180 24404
rect 9588 24352 9640 24404
rect 12164 24352 12216 24404
rect 13176 24352 13228 24404
rect 15660 24352 15712 24404
rect 16304 24352 16356 24404
rect 22284 24352 22336 24404
rect 22652 24352 22704 24404
rect 23756 24352 23808 24404
rect 24676 24352 24728 24404
rect 1584 24284 1636 24336
rect 11336 24216 11388 24268
rect 8944 24191 8996 24200
rect 8944 24157 8953 24191
rect 8953 24157 8987 24191
rect 8987 24157 8996 24191
rect 8944 24148 8996 24157
rect 9036 24148 9088 24200
rect 9220 24191 9272 24200
rect 9220 24157 9229 24191
rect 9229 24157 9263 24191
rect 9263 24157 9272 24191
rect 9220 24148 9272 24157
rect 8852 24080 8904 24132
rect 9772 24148 9824 24200
rect 10692 24191 10744 24200
rect 10692 24157 10701 24191
rect 10701 24157 10735 24191
rect 10735 24157 10744 24191
rect 10692 24148 10744 24157
rect 11244 24148 11296 24200
rect 9864 24080 9916 24132
rect 11888 24216 11940 24268
rect 11980 24148 12032 24200
rect 12440 24148 12492 24200
rect 17224 24284 17276 24336
rect 13912 24216 13964 24268
rect 14924 24216 14976 24268
rect 12716 24148 12768 24200
rect 13084 24148 13136 24200
rect 15476 24148 15528 24200
rect 16212 24191 16264 24200
rect 16212 24157 16221 24191
rect 16221 24157 16255 24191
rect 16255 24157 16264 24191
rect 16212 24148 16264 24157
rect 17224 24191 17276 24200
rect 17224 24157 17233 24191
rect 17233 24157 17267 24191
rect 17267 24157 17276 24191
rect 17224 24148 17276 24157
rect 17408 24284 17460 24336
rect 19800 24284 19852 24336
rect 26240 24352 26292 24404
rect 26608 24352 26660 24404
rect 17868 24148 17920 24200
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 20444 24148 20496 24200
rect 21272 24148 21324 24200
rect 21824 24148 21876 24200
rect 18236 24080 18288 24132
rect 19892 24080 19944 24132
rect 20076 24080 20128 24132
rect 22284 24216 22336 24268
rect 23204 24216 23256 24268
rect 23296 24216 23348 24268
rect 22468 24148 22520 24200
rect 23480 24191 23532 24200
rect 23480 24157 23489 24191
rect 23489 24157 23523 24191
rect 23523 24157 23532 24191
rect 23480 24148 23532 24157
rect 24584 24191 24636 24200
rect 24584 24157 24593 24191
rect 24593 24157 24627 24191
rect 24627 24157 24636 24191
rect 24584 24148 24636 24157
rect 25136 24284 25188 24336
rect 25320 24259 25372 24268
rect 25320 24225 25329 24259
rect 25329 24225 25363 24259
rect 25363 24225 25372 24259
rect 25320 24216 25372 24225
rect 25136 24148 25188 24200
rect 25596 24191 25648 24200
rect 25596 24157 25605 24191
rect 25605 24157 25639 24191
rect 25639 24157 25648 24191
rect 26608 24191 26660 24200
rect 25596 24148 25648 24157
rect 26608 24157 26617 24191
rect 26617 24157 26651 24191
rect 26651 24157 26660 24191
rect 26608 24148 26660 24157
rect 28816 24284 28868 24336
rect 28080 24216 28132 24268
rect 26884 24191 26936 24200
rect 26884 24157 26893 24191
rect 26893 24157 26927 24191
rect 26927 24157 26936 24191
rect 27160 24191 27212 24200
rect 26884 24148 26936 24157
rect 27160 24157 27169 24191
rect 27169 24157 27203 24191
rect 27203 24157 27212 24191
rect 27160 24148 27212 24157
rect 27804 24191 27856 24200
rect 27804 24157 27813 24191
rect 27813 24157 27847 24191
rect 27847 24157 27856 24191
rect 27804 24148 27856 24157
rect 28264 24148 28316 24200
rect 29828 24191 29880 24200
rect 29828 24157 29837 24191
rect 29837 24157 29871 24191
rect 29871 24157 29880 24191
rect 29828 24148 29880 24157
rect 7564 24012 7616 24064
rect 11336 24012 11388 24064
rect 11704 24055 11756 24064
rect 11704 24021 11713 24055
rect 11713 24021 11747 24055
rect 11747 24021 11756 24055
rect 11704 24012 11756 24021
rect 15292 24012 15344 24064
rect 16856 24012 16908 24064
rect 19432 24012 19484 24064
rect 22284 24012 22336 24064
rect 23480 24012 23532 24064
rect 25780 24055 25832 24064
rect 25780 24021 25789 24055
rect 25789 24021 25823 24055
rect 25823 24021 25832 24055
rect 25780 24012 25832 24021
rect 27068 24012 27120 24064
rect 27344 24055 27396 24064
rect 27344 24021 27353 24055
rect 27353 24021 27387 24055
rect 27387 24021 27396 24055
rect 27344 24012 27396 24021
rect 27436 24012 27488 24064
rect 28172 24012 28224 24064
rect 30012 24055 30064 24064
rect 30012 24021 30021 24055
rect 30021 24021 30055 24055
rect 30055 24021 30064 24055
rect 30012 24012 30064 24021
rect 10880 23910 10932 23962
rect 10944 23910 10996 23962
rect 11008 23910 11060 23962
rect 11072 23910 11124 23962
rect 11136 23910 11188 23962
rect 20811 23910 20863 23962
rect 20875 23910 20927 23962
rect 20939 23910 20991 23962
rect 21003 23910 21055 23962
rect 21067 23910 21119 23962
rect 9036 23808 9088 23860
rect 7564 23715 7616 23724
rect 7564 23681 7598 23715
rect 7598 23681 7616 23715
rect 7564 23672 7616 23681
rect 8852 23740 8904 23792
rect 14280 23808 14332 23860
rect 14464 23808 14516 23860
rect 14924 23808 14976 23860
rect 11428 23740 11480 23792
rect 11704 23740 11756 23792
rect 9680 23672 9732 23724
rect 10600 23672 10652 23724
rect 10968 23672 11020 23724
rect 14740 23740 14792 23792
rect 7288 23647 7340 23656
rect 7288 23613 7297 23647
rect 7297 23613 7331 23647
rect 7331 23613 7340 23647
rect 7288 23604 7340 23613
rect 12440 23604 12492 23656
rect 10876 23536 10928 23588
rect 13360 23672 13412 23724
rect 15016 23715 15068 23724
rect 15016 23681 15025 23715
rect 15025 23681 15059 23715
rect 15059 23681 15068 23715
rect 15016 23672 15068 23681
rect 15476 23740 15528 23792
rect 16672 23740 16724 23792
rect 12992 23647 13044 23656
rect 12992 23613 13001 23647
rect 13001 23613 13035 23647
rect 13035 23613 13044 23647
rect 12992 23604 13044 23613
rect 14464 23604 14516 23656
rect 15108 23647 15160 23656
rect 15108 23613 15117 23647
rect 15117 23613 15151 23647
rect 15151 23613 15160 23647
rect 15108 23604 15160 23613
rect 17500 23715 17552 23724
rect 17500 23681 17509 23715
rect 17509 23681 17543 23715
rect 17543 23681 17552 23715
rect 17500 23672 17552 23681
rect 18328 23740 18380 23792
rect 17960 23715 18012 23724
rect 17960 23681 17969 23715
rect 17969 23681 18003 23715
rect 18003 23681 18012 23715
rect 17960 23672 18012 23681
rect 19064 23672 19116 23724
rect 19340 23672 19392 23724
rect 24492 23808 24544 23860
rect 22192 23740 22244 23792
rect 26332 23808 26384 23860
rect 27712 23808 27764 23860
rect 22928 23715 22980 23724
rect 14832 23536 14884 23588
rect 17040 23536 17092 23588
rect 10416 23468 10468 23520
rect 11980 23511 12032 23520
rect 11980 23477 11989 23511
rect 11989 23477 12023 23511
rect 12023 23477 12032 23511
rect 11980 23468 12032 23477
rect 13084 23468 13136 23520
rect 13544 23468 13596 23520
rect 14648 23511 14700 23520
rect 14648 23477 14657 23511
rect 14657 23477 14691 23511
rect 14691 23477 14700 23511
rect 14648 23468 14700 23477
rect 16304 23468 16356 23520
rect 16948 23511 17000 23520
rect 16948 23477 16957 23511
rect 16957 23477 16991 23511
rect 16991 23477 17000 23511
rect 16948 23468 17000 23477
rect 17224 23468 17276 23520
rect 17592 23468 17644 23520
rect 19616 23511 19668 23520
rect 19616 23477 19625 23511
rect 19625 23477 19659 23511
rect 19659 23477 19668 23511
rect 19616 23468 19668 23477
rect 22928 23681 22937 23715
rect 22937 23681 22971 23715
rect 22971 23681 22980 23715
rect 22928 23672 22980 23681
rect 23112 23715 23164 23724
rect 23112 23681 23121 23715
rect 23121 23681 23155 23715
rect 23155 23681 23164 23715
rect 23112 23672 23164 23681
rect 24860 23672 24912 23724
rect 25780 23672 25832 23724
rect 28448 23740 28500 23792
rect 27988 23672 28040 23724
rect 28816 23672 28868 23724
rect 30104 23715 30156 23724
rect 30104 23681 30113 23715
rect 30113 23681 30147 23715
rect 30147 23681 30156 23715
rect 30104 23672 30156 23681
rect 20444 23604 20496 23656
rect 22836 23604 22888 23656
rect 19892 23536 19944 23588
rect 25320 23468 25372 23520
rect 25596 23468 25648 23520
rect 27804 23468 27856 23520
rect 29828 23468 29880 23520
rect 5915 23366 5967 23418
rect 5979 23366 6031 23418
rect 6043 23366 6095 23418
rect 6107 23366 6159 23418
rect 6171 23366 6223 23418
rect 15846 23366 15898 23418
rect 15910 23366 15962 23418
rect 15974 23366 16026 23418
rect 16038 23366 16090 23418
rect 16102 23366 16154 23418
rect 25776 23366 25828 23418
rect 25840 23366 25892 23418
rect 25904 23366 25956 23418
rect 25968 23366 26020 23418
rect 26032 23366 26084 23418
rect 8300 23307 8352 23316
rect 8300 23273 8309 23307
rect 8309 23273 8343 23307
rect 8343 23273 8352 23307
rect 8300 23264 8352 23273
rect 9680 23307 9732 23316
rect 9680 23273 9689 23307
rect 9689 23273 9723 23307
rect 9723 23273 9732 23307
rect 9680 23264 9732 23273
rect 11888 23307 11940 23316
rect 11888 23273 11897 23307
rect 11897 23273 11931 23307
rect 11931 23273 11940 23307
rect 11888 23264 11940 23273
rect 12624 23264 12676 23316
rect 12992 23264 13044 23316
rect 16948 23264 17000 23316
rect 17040 23264 17092 23316
rect 18328 23264 18380 23316
rect 18880 23264 18932 23316
rect 14096 23196 14148 23248
rect 8300 23128 8352 23180
rect 9220 23171 9272 23180
rect 9220 23137 9229 23171
rect 9229 23137 9263 23171
rect 9263 23137 9272 23171
rect 9220 23128 9272 23137
rect 2320 23103 2372 23112
rect 2320 23069 2329 23103
rect 2329 23069 2363 23103
rect 2363 23069 2372 23103
rect 2320 23060 2372 23069
rect 8944 23103 8996 23112
rect 8944 23069 8953 23103
rect 8953 23069 8987 23103
rect 8987 23069 8996 23103
rect 8944 23060 8996 23069
rect 9404 23060 9456 23112
rect 9864 23060 9916 23112
rect 10140 23128 10192 23180
rect 10416 23128 10468 23180
rect 10600 23171 10652 23180
rect 10600 23137 10609 23171
rect 10609 23137 10643 23171
rect 10643 23137 10652 23171
rect 10600 23128 10652 23137
rect 10968 23128 11020 23180
rect 10876 23060 10928 23112
rect 11336 23060 11388 23112
rect 12716 23128 12768 23180
rect 12440 23060 12492 23112
rect 12900 23060 12952 23112
rect 13176 23060 13228 23112
rect 14648 23196 14700 23248
rect 15936 23239 15988 23248
rect 15936 23205 15945 23239
rect 15945 23205 15979 23239
rect 15979 23205 15988 23239
rect 15936 23196 15988 23205
rect 19616 23264 19668 23316
rect 21916 23264 21968 23316
rect 23388 23264 23440 23316
rect 23756 23264 23808 23316
rect 24860 23307 24912 23316
rect 24860 23273 24869 23307
rect 24869 23273 24903 23307
rect 24903 23273 24912 23307
rect 24860 23264 24912 23273
rect 25412 23264 25464 23316
rect 14366 23171 14418 23180
rect 14366 23137 14375 23171
rect 14375 23137 14409 23171
rect 14409 23137 14418 23171
rect 14366 23128 14418 23137
rect 10324 22992 10376 23044
rect 12072 22992 12124 23044
rect 13268 23035 13320 23044
rect 13268 23001 13277 23035
rect 13277 23001 13311 23035
rect 13311 23001 13320 23035
rect 13268 22992 13320 23001
rect 13544 22992 13596 23044
rect 14372 22992 14424 23044
rect 15200 23060 15252 23112
rect 16212 23128 16264 23180
rect 17316 23171 17368 23180
rect 17316 23137 17325 23171
rect 17325 23137 17359 23171
rect 17359 23137 17368 23171
rect 17316 23128 17368 23137
rect 16304 23103 16356 23112
rect 16304 23069 16313 23103
rect 16313 23069 16347 23103
rect 16347 23069 16356 23103
rect 16304 23060 16356 23069
rect 18328 23060 18380 23112
rect 19340 23060 19392 23112
rect 20720 23128 20772 23180
rect 22836 23196 22888 23248
rect 21640 23171 21692 23180
rect 21640 23137 21649 23171
rect 21649 23137 21683 23171
rect 21683 23137 21692 23171
rect 21640 23128 21692 23137
rect 20352 23060 20404 23112
rect 14924 22992 14976 23044
rect 15016 22992 15068 23044
rect 1584 22967 1636 22976
rect 1584 22933 1593 22967
rect 1593 22933 1627 22967
rect 1627 22933 1636 22967
rect 1584 22924 1636 22933
rect 15200 22924 15252 22976
rect 17408 22992 17460 23044
rect 18604 22992 18656 23044
rect 21732 23060 21784 23112
rect 22468 23103 22520 23112
rect 22468 23069 22477 23103
rect 22477 23069 22511 23103
rect 22511 23069 22520 23103
rect 22468 23060 22520 23069
rect 25596 23196 25648 23248
rect 27160 23196 27212 23248
rect 24492 23128 24544 23180
rect 28080 23128 28132 23180
rect 25044 23060 25096 23112
rect 25504 23103 25556 23112
rect 25504 23069 25513 23103
rect 25513 23069 25547 23103
rect 25547 23069 25556 23103
rect 25504 23060 25556 23069
rect 27344 23060 27396 23112
rect 23388 22992 23440 23044
rect 28356 22992 28408 23044
rect 16948 22924 17000 22976
rect 17040 22924 17092 22976
rect 18880 22924 18932 22976
rect 19248 22924 19300 22976
rect 23664 22924 23716 22976
rect 24676 22924 24728 22976
rect 26516 22924 26568 22976
rect 10880 22822 10932 22874
rect 10944 22822 10996 22874
rect 11008 22822 11060 22874
rect 11072 22822 11124 22874
rect 11136 22822 11188 22874
rect 20811 22822 20863 22874
rect 20875 22822 20927 22874
rect 20939 22822 20991 22874
rect 21003 22822 21055 22874
rect 21067 22822 21119 22874
rect 8300 22720 8352 22772
rect 9772 22720 9824 22772
rect 11980 22720 12032 22772
rect 13268 22720 13320 22772
rect 17040 22720 17092 22772
rect 17132 22720 17184 22772
rect 19708 22763 19760 22772
rect 19708 22729 19717 22763
rect 19717 22729 19751 22763
rect 19751 22729 19760 22763
rect 19708 22720 19760 22729
rect 22008 22720 22060 22772
rect 23388 22720 23440 22772
rect 23664 22720 23716 22772
rect 25136 22720 25188 22772
rect 27988 22763 28040 22772
rect 27988 22729 27997 22763
rect 27997 22729 28031 22763
rect 28031 22729 28040 22763
rect 27988 22720 28040 22729
rect 9496 22652 9548 22704
rect 22192 22652 22244 22704
rect 23756 22695 23808 22704
rect 23756 22661 23765 22695
rect 23765 22661 23799 22695
rect 23799 22661 23808 22695
rect 23756 22652 23808 22661
rect 8392 22584 8444 22636
rect 8944 22627 8996 22636
rect 8944 22593 8953 22627
rect 8953 22593 8987 22627
rect 8987 22593 8996 22627
rect 8944 22584 8996 22593
rect 9128 22584 9180 22636
rect 9772 22584 9824 22636
rect 11244 22584 11296 22636
rect 11888 22584 11940 22636
rect 12716 22584 12768 22636
rect 8576 22448 8628 22500
rect 9680 22516 9732 22568
rect 11336 22516 11388 22568
rect 13544 22584 13596 22636
rect 15200 22627 15252 22636
rect 15200 22593 15209 22627
rect 15209 22593 15243 22627
rect 15243 22593 15252 22627
rect 15200 22584 15252 22593
rect 15292 22584 15344 22636
rect 9956 22448 10008 22500
rect 12164 22448 12216 22500
rect 14740 22516 14792 22568
rect 15200 22448 15252 22500
rect 15476 22627 15528 22636
rect 15476 22593 15485 22627
rect 15485 22593 15519 22627
rect 15519 22593 15528 22627
rect 15752 22627 15804 22636
rect 15476 22584 15528 22593
rect 15752 22593 15761 22627
rect 15761 22593 15795 22627
rect 15795 22593 15804 22627
rect 15752 22584 15804 22593
rect 16580 22584 16632 22636
rect 16948 22584 17000 22636
rect 17408 22584 17460 22636
rect 20812 22627 20864 22636
rect 20812 22593 20821 22627
rect 20821 22593 20855 22627
rect 20855 22593 20864 22627
rect 20812 22584 20864 22593
rect 21272 22584 21324 22636
rect 15752 22448 15804 22500
rect 17500 22516 17552 22568
rect 19156 22516 19208 22568
rect 20628 22516 20680 22568
rect 21640 22584 21692 22636
rect 21916 22584 21968 22636
rect 22560 22584 22612 22636
rect 24768 22652 24820 22704
rect 24584 22584 24636 22636
rect 18420 22448 18472 22500
rect 8484 22423 8536 22432
rect 8484 22389 8493 22423
rect 8493 22389 8527 22423
rect 8527 22389 8536 22423
rect 8484 22380 8536 22389
rect 9864 22380 9916 22432
rect 12532 22380 12584 22432
rect 13084 22380 13136 22432
rect 14372 22380 14424 22432
rect 15384 22380 15436 22432
rect 16948 22380 17000 22432
rect 17684 22380 17736 22432
rect 21364 22380 21416 22432
rect 24860 22516 24912 22568
rect 25596 22516 25648 22568
rect 23112 22448 23164 22500
rect 27344 22584 27396 22636
rect 27528 22652 27580 22704
rect 27804 22627 27856 22636
rect 27804 22593 27813 22627
rect 27813 22593 27847 22627
rect 27847 22593 27856 22627
rect 27804 22584 27856 22593
rect 28448 22627 28500 22636
rect 28448 22593 28457 22627
rect 28457 22593 28491 22627
rect 28491 22593 28500 22627
rect 28448 22584 28500 22593
rect 29000 22584 29052 22636
rect 26884 22516 26936 22568
rect 28080 22516 28132 22568
rect 27988 22448 28040 22500
rect 23020 22380 23072 22432
rect 26332 22423 26384 22432
rect 26332 22389 26341 22423
rect 26341 22389 26375 22423
rect 26375 22389 26384 22423
rect 26332 22380 26384 22389
rect 27620 22380 27672 22432
rect 27804 22380 27856 22432
rect 29552 22380 29604 22432
rect 5915 22278 5967 22330
rect 5979 22278 6031 22330
rect 6043 22278 6095 22330
rect 6107 22278 6159 22330
rect 6171 22278 6223 22330
rect 15846 22278 15898 22330
rect 15910 22278 15962 22330
rect 15974 22278 16026 22330
rect 16038 22278 16090 22330
rect 16102 22278 16154 22330
rect 25776 22278 25828 22330
rect 25840 22278 25892 22330
rect 25904 22278 25956 22330
rect 25968 22278 26020 22330
rect 26032 22278 26084 22330
rect 8300 22219 8352 22228
rect 8300 22185 8309 22219
rect 8309 22185 8343 22219
rect 8343 22185 8352 22219
rect 8300 22176 8352 22185
rect 8944 22176 8996 22228
rect 9772 22176 9824 22228
rect 10784 22176 10836 22228
rect 9864 22151 9916 22160
rect 9864 22117 9873 22151
rect 9873 22117 9907 22151
rect 9907 22117 9916 22151
rect 9864 22108 9916 22117
rect 2136 22040 2188 22092
rect 9588 22040 9640 22092
rect 8576 21972 8628 22024
rect 8668 21972 8720 22024
rect 10048 21972 10100 22024
rect 10048 21836 10100 21888
rect 10692 21972 10744 22024
rect 11152 21972 11204 22024
rect 12532 22176 12584 22228
rect 16580 22176 16632 22228
rect 17224 22176 17276 22228
rect 20720 22176 20772 22228
rect 12992 22108 13044 22160
rect 15568 22083 15620 22092
rect 12440 21972 12492 22024
rect 12624 22015 12676 22024
rect 12624 21981 12633 22015
rect 12633 21981 12667 22015
rect 12667 21981 12676 22015
rect 12624 21972 12676 21981
rect 15568 22049 15577 22083
rect 15577 22049 15611 22083
rect 15611 22049 15620 22083
rect 15568 22040 15620 22049
rect 15384 22015 15436 22024
rect 15384 21981 15393 22015
rect 15393 21981 15427 22015
rect 15427 21981 15436 22015
rect 15384 21972 15436 21981
rect 15476 21972 15528 22024
rect 15844 22040 15896 22092
rect 17040 22108 17092 22160
rect 16856 22083 16908 22092
rect 16856 22049 16865 22083
rect 16865 22049 16899 22083
rect 16899 22049 16908 22083
rect 16856 22040 16908 22049
rect 17224 22040 17276 22092
rect 17500 22040 17552 22092
rect 15752 21972 15804 22024
rect 17316 21972 17368 22024
rect 21456 22108 21508 22160
rect 22468 22108 22520 22160
rect 23112 22176 23164 22228
rect 25504 22176 25556 22228
rect 27620 22176 27672 22228
rect 28356 22176 28408 22228
rect 28632 22176 28684 22228
rect 28908 22176 28960 22228
rect 23756 22108 23808 22160
rect 25596 22108 25648 22160
rect 18144 22015 18196 22024
rect 18144 21981 18153 22015
rect 18153 21981 18187 22015
rect 18187 21981 18196 22015
rect 18144 21972 18196 21981
rect 13820 21904 13872 21956
rect 14188 21904 14240 21956
rect 11520 21836 11572 21888
rect 11704 21879 11756 21888
rect 11704 21845 11713 21879
rect 11713 21845 11747 21879
rect 11747 21845 11756 21879
rect 11704 21836 11756 21845
rect 14832 21836 14884 21888
rect 15016 21879 15068 21888
rect 15016 21845 15025 21879
rect 15025 21845 15059 21879
rect 15059 21845 15068 21879
rect 15016 21836 15068 21845
rect 16580 21879 16632 21888
rect 16580 21845 16589 21879
rect 16589 21845 16623 21879
rect 16623 21845 16632 21879
rect 16580 21836 16632 21845
rect 18420 21972 18472 22024
rect 18788 21972 18840 22024
rect 18604 21904 18656 21956
rect 21916 22040 21968 22092
rect 25688 22083 25740 22092
rect 25688 22049 25697 22083
rect 25697 22049 25731 22083
rect 25731 22049 25740 22083
rect 25688 22040 25740 22049
rect 19064 21836 19116 21888
rect 19800 21879 19852 21888
rect 19800 21845 19809 21879
rect 19809 21845 19843 21879
rect 19843 21845 19852 21879
rect 19800 21836 19852 21845
rect 22008 21972 22060 22024
rect 23388 21972 23440 22024
rect 24216 21972 24268 22024
rect 25412 22015 25464 22024
rect 25412 21981 25421 22015
rect 25421 21981 25455 22015
rect 25455 21981 25464 22015
rect 25412 21972 25464 21981
rect 25596 22015 25648 22024
rect 25596 21981 25605 22015
rect 25605 21981 25639 22015
rect 25639 21981 25648 22015
rect 25596 21972 25648 21981
rect 27436 22040 27488 22092
rect 21272 21904 21324 21956
rect 19984 21836 20036 21888
rect 23940 21904 23992 21956
rect 25320 21904 25372 21956
rect 22100 21836 22152 21888
rect 22744 21836 22796 21888
rect 22928 21836 22980 21888
rect 26792 21904 26844 21956
rect 27160 21972 27212 22024
rect 28080 21972 28132 22024
rect 28724 22040 28776 22092
rect 29000 22083 29052 22092
rect 29000 22049 29009 22083
rect 29009 22049 29043 22083
rect 29043 22049 29052 22083
rect 29000 22040 29052 22049
rect 27344 21904 27396 21956
rect 28356 21904 28408 21956
rect 28632 22015 28684 22024
rect 28632 21981 28641 22015
rect 28641 21981 28675 22015
rect 28675 21981 28684 22015
rect 28632 21972 28684 21981
rect 29552 22015 29604 22024
rect 29552 21981 29561 22015
rect 29561 21981 29595 22015
rect 29595 21981 29604 22015
rect 29552 21972 29604 21981
rect 27068 21836 27120 21888
rect 27252 21836 27304 21888
rect 10880 21734 10932 21786
rect 10944 21734 10996 21786
rect 11008 21734 11060 21786
rect 11072 21734 11124 21786
rect 11136 21734 11188 21786
rect 20811 21734 20863 21786
rect 20875 21734 20927 21786
rect 20939 21734 20991 21786
rect 21003 21734 21055 21786
rect 21067 21734 21119 21786
rect 8668 21632 8720 21684
rect 10692 21632 10744 21684
rect 11244 21632 11296 21684
rect 12164 21632 12216 21684
rect 13452 21632 13504 21684
rect 16580 21632 16632 21684
rect 8484 21564 8536 21616
rect 2136 21539 2188 21548
rect 2136 21505 2145 21539
rect 2145 21505 2179 21539
rect 2179 21505 2188 21539
rect 2136 21496 2188 21505
rect 2320 21539 2372 21548
rect 2320 21505 2329 21539
rect 2329 21505 2363 21539
rect 2363 21505 2372 21539
rect 2320 21496 2372 21505
rect 7288 21496 7340 21548
rect 10416 21496 10468 21548
rect 11428 21496 11480 21548
rect 12992 21564 13044 21616
rect 14832 21607 14884 21616
rect 14832 21573 14841 21607
rect 14841 21573 14875 21607
rect 14875 21573 14884 21607
rect 14832 21564 14884 21573
rect 13820 21496 13872 21548
rect 19432 21564 19484 21616
rect 20536 21632 20588 21684
rect 22008 21632 22060 21684
rect 22468 21632 22520 21684
rect 23388 21632 23440 21684
rect 24952 21632 25004 21684
rect 25688 21632 25740 21684
rect 19984 21564 20036 21616
rect 20260 21607 20312 21616
rect 20260 21573 20269 21607
rect 20269 21573 20303 21607
rect 20303 21573 20312 21607
rect 20260 21564 20312 21573
rect 20352 21564 20404 21616
rect 21916 21564 21968 21616
rect 26148 21607 26200 21616
rect 16304 21496 16356 21548
rect 17592 21496 17644 21548
rect 17868 21496 17920 21548
rect 17960 21496 18012 21548
rect 18604 21496 18656 21548
rect 18788 21539 18840 21548
rect 18788 21505 18797 21539
rect 18797 21505 18831 21539
rect 18831 21505 18840 21539
rect 18788 21496 18840 21505
rect 19156 21496 19208 21548
rect 20168 21496 20220 21548
rect 26148 21573 26157 21607
rect 26157 21573 26191 21607
rect 26191 21573 26200 21607
rect 26148 21564 26200 21573
rect 27160 21564 27212 21616
rect 12072 21471 12124 21480
rect 9956 21403 10008 21412
rect 9956 21369 9965 21403
rect 9965 21369 9999 21403
rect 9999 21369 10008 21403
rect 9956 21360 10008 21369
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 10968 21360 11020 21412
rect 11428 21292 11480 21344
rect 11704 21360 11756 21412
rect 12072 21437 12081 21471
rect 12081 21437 12115 21471
rect 12115 21437 12124 21471
rect 12072 21428 12124 21437
rect 12256 21428 12308 21480
rect 18972 21471 19024 21480
rect 18972 21437 18981 21471
rect 18981 21437 19015 21471
rect 19015 21437 19024 21471
rect 18972 21428 19024 21437
rect 20720 21428 20772 21480
rect 22192 21471 22244 21480
rect 22192 21437 22201 21471
rect 22201 21437 22235 21471
rect 22235 21437 22244 21471
rect 22192 21428 22244 21437
rect 27252 21496 27304 21548
rect 28172 21564 28224 21616
rect 27896 21539 27948 21548
rect 27896 21505 27905 21539
rect 27905 21505 27939 21539
rect 27939 21505 27948 21539
rect 27896 21496 27948 21505
rect 27988 21496 28040 21548
rect 24768 21471 24820 21480
rect 24768 21437 24777 21471
rect 24777 21437 24811 21471
rect 24811 21437 24820 21471
rect 24768 21428 24820 21437
rect 28172 21428 28224 21480
rect 12992 21360 13044 21412
rect 16856 21360 16908 21412
rect 18144 21360 18196 21412
rect 12716 21292 12768 21344
rect 14648 21292 14700 21344
rect 14832 21292 14884 21344
rect 16580 21292 16632 21344
rect 19616 21292 19668 21344
rect 19800 21360 19852 21412
rect 22100 21360 22152 21412
rect 22652 21360 22704 21412
rect 21456 21292 21508 21344
rect 21732 21292 21784 21344
rect 24216 21292 24268 21344
rect 28448 21496 28500 21548
rect 5915 21190 5967 21242
rect 5979 21190 6031 21242
rect 6043 21190 6095 21242
rect 6107 21190 6159 21242
rect 6171 21190 6223 21242
rect 15846 21190 15898 21242
rect 15910 21190 15962 21242
rect 15974 21190 16026 21242
rect 16038 21190 16090 21242
rect 16102 21190 16154 21242
rect 25776 21190 25828 21242
rect 25840 21190 25892 21242
rect 25904 21190 25956 21242
rect 25968 21190 26020 21242
rect 26032 21190 26084 21242
rect 10508 21088 10560 21140
rect 12164 21131 12216 21140
rect 2412 21020 2464 21072
rect 11060 21020 11112 21072
rect 10324 20952 10376 21004
rect 12164 21097 12173 21131
rect 12173 21097 12207 21131
rect 12207 21097 12216 21131
rect 12164 21088 12216 21097
rect 9956 20927 10008 20936
rect 9956 20893 9965 20927
rect 9965 20893 9999 20927
rect 9999 20893 10008 20927
rect 9956 20884 10008 20893
rect 10416 20884 10468 20936
rect 10600 20927 10652 20936
rect 10600 20893 10609 20927
rect 10609 20893 10643 20927
rect 10643 20893 10652 20927
rect 10600 20884 10652 20893
rect 10692 20884 10744 20936
rect 13452 21088 13504 21140
rect 14188 21088 14240 21140
rect 15292 21088 15344 21140
rect 12532 21020 12584 21072
rect 13728 21020 13780 21072
rect 17040 21088 17092 21140
rect 22468 21088 22520 21140
rect 22652 21131 22704 21140
rect 22652 21097 22661 21131
rect 22661 21097 22695 21131
rect 22695 21097 22704 21131
rect 22652 21088 22704 21097
rect 24400 21088 24452 21140
rect 24584 21088 24636 21140
rect 24768 21088 24820 21140
rect 18236 21020 18288 21072
rect 18788 21020 18840 21072
rect 10324 20816 10376 20868
rect 11612 20927 11664 20936
rect 11612 20893 11621 20927
rect 11621 20893 11655 20927
rect 11655 20893 11664 20927
rect 11612 20884 11664 20893
rect 15016 20952 15068 21004
rect 12716 20927 12768 20936
rect 12716 20893 12725 20927
rect 12725 20893 12759 20927
rect 12759 20893 12768 20927
rect 12716 20884 12768 20893
rect 14372 20927 14424 20936
rect 14372 20893 14381 20927
rect 14381 20893 14415 20927
rect 14415 20893 14424 20927
rect 14372 20884 14424 20893
rect 10968 20859 11020 20868
rect 10968 20825 10977 20859
rect 10977 20825 11011 20859
rect 11011 20825 11020 20859
rect 10968 20816 11020 20825
rect 9128 20791 9180 20800
rect 9128 20757 9137 20791
rect 9137 20757 9171 20791
rect 9171 20757 9180 20791
rect 9128 20748 9180 20757
rect 10048 20791 10100 20800
rect 10048 20757 10057 20791
rect 10057 20757 10091 20791
rect 10091 20757 10100 20791
rect 10048 20748 10100 20757
rect 10140 20748 10192 20800
rect 10416 20748 10468 20800
rect 10692 20748 10744 20800
rect 12900 20816 12952 20868
rect 13452 20816 13504 20868
rect 13912 20816 13964 20868
rect 15108 20884 15160 20936
rect 15384 20816 15436 20868
rect 18052 20952 18104 21004
rect 17960 20884 18012 20936
rect 19984 20952 20036 21004
rect 21548 20952 21600 21004
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 20720 20927 20772 20936
rect 20720 20893 20729 20927
rect 20729 20893 20763 20927
rect 20763 20893 20772 20927
rect 20720 20884 20772 20893
rect 22284 20952 22336 21004
rect 23204 20952 23256 21004
rect 23756 20952 23808 21004
rect 24860 20995 24912 21004
rect 24860 20961 24869 20995
rect 24869 20961 24903 20995
rect 24903 20961 24912 20995
rect 24860 20952 24912 20961
rect 27344 21020 27396 21072
rect 16672 20859 16724 20868
rect 16672 20825 16681 20859
rect 16681 20825 16715 20859
rect 16715 20825 16724 20859
rect 16672 20816 16724 20825
rect 17224 20816 17276 20868
rect 18604 20816 18656 20868
rect 18788 20816 18840 20868
rect 18236 20748 18288 20800
rect 20168 20816 20220 20868
rect 20628 20816 20680 20868
rect 22100 20884 22152 20936
rect 22468 20927 22520 20936
rect 22468 20893 22482 20927
rect 22482 20893 22516 20927
rect 22516 20893 22520 20927
rect 22468 20884 22520 20893
rect 22928 20884 22980 20936
rect 23296 20927 23348 20936
rect 23296 20893 23305 20927
rect 23305 20893 23339 20927
rect 23339 20893 23348 20927
rect 23296 20884 23348 20893
rect 20076 20748 20128 20800
rect 20260 20748 20312 20800
rect 20444 20748 20496 20800
rect 21732 20816 21784 20868
rect 22652 20816 22704 20868
rect 22744 20816 22796 20868
rect 24032 20884 24084 20936
rect 24400 20884 24452 20936
rect 21180 20748 21232 20800
rect 22192 20748 22244 20800
rect 22928 20748 22980 20800
rect 24952 20884 25004 20936
rect 25136 20884 25188 20936
rect 25320 20884 25372 20936
rect 25136 20748 25188 20800
rect 25964 20995 26016 21004
rect 25964 20961 25973 20995
rect 25973 20961 26007 20995
rect 26007 20961 26016 20995
rect 25964 20952 26016 20961
rect 26792 20952 26844 21004
rect 27804 20952 27856 21004
rect 27620 20884 27672 20936
rect 28172 20884 28224 20936
rect 28356 20884 28408 20936
rect 29092 20884 29144 20936
rect 26332 20748 26384 20800
rect 27436 20791 27488 20800
rect 27436 20757 27445 20791
rect 27445 20757 27479 20791
rect 27479 20757 27488 20791
rect 27436 20748 27488 20757
rect 10880 20646 10932 20698
rect 10944 20646 10996 20698
rect 11008 20646 11060 20698
rect 11072 20646 11124 20698
rect 11136 20646 11188 20698
rect 20811 20646 20863 20698
rect 20875 20646 20927 20698
rect 20939 20646 20991 20698
rect 21003 20646 21055 20698
rect 21067 20646 21119 20698
rect 9680 20544 9732 20596
rect 12716 20544 12768 20596
rect 13820 20544 13872 20596
rect 14096 20544 14148 20596
rect 9956 20476 10008 20528
rect 10048 20476 10100 20528
rect 10508 20476 10560 20528
rect 11612 20476 11664 20528
rect 11796 20476 11848 20528
rect 12440 20476 12492 20528
rect 15016 20519 15068 20528
rect 8392 20408 8444 20460
rect 9128 20408 9180 20460
rect 12164 20408 12216 20460
rect 13820 20451 13872 20460
rect 13820 20417 13829 20451
rect 13829 20417 13863 20451
rect 13863 20417 13872 20451
rect 13820 20408 13872 20417
rect 14188 20451 14240 20460
rect 14188 20417 14197 20451
rect 14197 20417 14231 20451
rect 14231 20417 14240 20451
rect 14188 20408 14240 20417
rect 15016 20485 15025 20519
rect 15025 20485 15059 20519
rect 15059 20485 15068 20519
rect 15016 20476 15068 20485
rect 19524 20544 19576 20596
rect 19800 20544 19852 20596
rect 20168 20544 20220 20596
rect 24768 20544 24820 20596
rect 25228 20587 25280 20596
rect 25228 20553 25237 20587
rect 25237 20553 25271 20587
rect 25271 20553 25280 20587
rect 25228 20544 25280 20553
rect 20076 20476 20128 20528
rect 20444 20476 20496 20528
rect 14556 20408 14608 20460
rect 15476 20451 15528 20460
rect 15476 20417 15485 20451
rect 15485 20417 15519 20451
rect 15519 20417 15528 20451
rect 15476 20408 15528 20417
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 18328 20451 18380 20460
rect 18328 20417 18337 20451
rect 18337 20417 18371 20451
rect 18371 20417 18380 20451
rect 18328 20408 18380 20417
rect 19984 20408 20036 20460
rect 20628 20408 20680 20460
rect 21180 20476 21232 20528
rect 21272 20519 21324 20528
rect 21272 20485 21281 20519
rect 21281 20485 21315 20519
rect 21315 20485 21324 20519
rect 21272 20476 21324 20485
rect 21916 20476 21968 20528
rect 1584 20340 1636 20392
rect 16580 20340 16632 20392
rect 16856 20340 16908 20392
rect 20076 20340 20128 20392
rect 20444 20340 20496 20392
rect 9128 20272 9180 20324
rect 9956 20204 10008 20256
rect 10324 20204 10376 20256
rect 11244 20272 11296 20324
rect 11704 20272 11756 20324
rect 12348 20272 12400 20324
rect 17408 20272 17460 20324
rect 19432 20272 19484 20324
rect 20168 20272 20220 20324
rect 16488 20204 16540 20256
rect 16672 20247 16724 20256
rect 16672 20213 16681 20247
rect 16681 20213 16715 20247
rect 16715 20213 16724 20247
rect 16672 20204 16724 20213
rect 17132 20204 17184 20256
rect 19524 20204 19576 20256
rect 21456 20340 21508 20392
rect 21916 20340 21968 20392
rect 21640 20204 21692 20256
rect 22100 20451 22152 20460
rect 22100 20417 22109 20451
rect 22109 20417 22143 20451
rect 22143 20417 22152 20451
rect 22100 20408 22152 20417
rect 22284 20408 22336 20460
rect 23020 20408 23072 20460
rect 23204 20408 23256 20460
rect 24676 20451 24728 20460
rect 22468 20340 22520 20392
rect 24676 20417 24685 20451
rect 24685 20417 24719 20451
rect 24719 20417 24728 20451
rect 24676 20408 24728 20417
rect 24768 20451 24820 20460
rect 24768 20417 24777 20451
rect 24777 20417 24811 20451
rect 24811 20417 24820 20451
rect 25044 20451 25096 20460
rect 24768 20408 24820 20417
rect 25044 20417 25053 20451
rect 25053 20417 25087 20451
rect 25087 20417 25096 20451
rect 25044 20408 25096 20417
rect 26148 20544 26200 20596
rect 26240 20544 26292 20596
rect 27620 20544 27672 20596
rect 27436 20476 27488 20528
rect 24584 20340 24636 20392
rect 26240 20451 26292 20460
rect 26240 20417 26249 20451
rect 26249 20417 26283 20451
rect 26283 20417 26292 20451
rect 26240 20408 26292 20417
rect 27252 20408 27304 20460
rect 27896 20451 27948 20460
rect 25964 20383 26016 20392
rect 22560 20315 22612 20324
rect 22560 20281 22569 20315
rect 22569 20281 22603 20315
rect 22603 20281 22612 20315
rect 22560 20272 22612 20281
rect 22744 20272 22796 20324
rect 22836 20204 22888 20256
rect 23756 20204 23808 20256
rect 25964 20349 25973 20383
rect 25973 20349 26007 20383
rect 26007 20349 26016 20383
rect 25964 20340 26016 20349
rect 26148 20340 26200 20392
rect 27896 20417 27905 20451
rect 27905 20417 27939 20451
rect 27939 20417 27948 20451
rect 27896 20408 27948 20417
rect 28448 20408 28500 20460
rect 28172 20340 28224 20392
rect 27712 20272 27764 20324
rect 26608 20204 26660 20256
rect 27528 20204 27580 20256
rect 5915 20102 5967 20154
rect 5979 20102 6031 20154
rect 6043 20102 6095 20154
rect 6107 20102 6159 20154
rect 6171 20102 6223 20154
rect 15846 20102 15898 20154
rect 15910 20102 15962 20154
rect 15974 20102 16026 20154
rect 16038 20102 16090 20154
rect 16102 20102 16154 20154
rect 25776 20102 25828 20154
rect 25840 20102 25892 20154
rect 25904 20102 25956 20154
rect 25968 20102 26020 20154
rect 26032 20102 26084 20154
rect 12164 20043 12216 20052
rect 12164 20009 12173 20043
rect 12173 20009 12207 20043
rect 12207 20009 12216 20043
rect 12164 20000 12216 20009
rect 13544 20000 13596 20052
rect 14096 20000 14148 20052
rect 15476 20000 15528 20052
rect 16580 20000 16632 20052
rect 17316 20000 17368 20052
rect 17408 20000 17460 20052
rect 19432 20000 19484 20052
rect 19984 20043 20036 20052
rect 19984 20009 19993 20043
rect 19993 20009 20027 20043
rect 20027 20009 20036 20043
rect 19984 20000 20036 20009
rect 20628 20000 20680 20052
rect 23112 20000 23164 20052
rect 23388 20000 23440 20052
rect 14924 19932 14976 19984
rect 10784 19864 10836 19916
rect 13820 19864 13872 19916
rect 14096 19864 14148 19916
rect 16672 19932 16724 19984
rect 15568 19907 15620 19916
rect 15568 19873 15577 19907
rect 15577 19873 15611 19907
rect 15611 19873 15620 19907
rect 15568 19864 15620 19873
rect 16304 19864 16356 19916
rect 17500 19864 17552 19916
rect 19156 19864 19208 19916
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 1768 19839 1820 19848
rect 1768 19805 1777 19839
rect 1777 19805 1811 19839
rect 1811 19805 1820 19839
rect 1768 19796 1820 19805
rect 2320 19796 2372 19848
rect 9220 19771 9272 19780
rect 9220 19737 9254 19771
rect 9254 19737 9272 19771
rect 9220 19728 9272 19737
rect 9312 19728 9364 19780
rect 12348 19796 12400 19848
rect 13360 19839 13412 19848
rect 12440 19728 12492 19780
rect 13084 19728 13136 19780
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 16212 19796 16264 19848
rect 16488 19796 16540 19848
rect 17132 19796 17184 19848
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 17960 19839 18012 19848
rect 14188 19728 14240 19780
rect 15568 19728 15620 19780
rect 16764 19728 16816 19780
rect 17960 19805 17969 19839
rect 17969 19805 18003 19839
rect 18003 19805 18012 19839
rect 17960 19796 18012 19805
rect 18788 19796 18840 19848
rect 19340 19796 19392 19848
rect 22284 19932 22336 19984
rect 20168 19864 20220 19916
rect 21180 19864 21232 19916
rect 18880 19728 18932 19780
rect 19616 19839 19668 19848
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 19800 19839 19852 19848
rect 19616 19796 19668 19805
rect 19800 19805 19809 19839
rect 19809 19805 19843 19839
rect 19843 19805 19852 19839
rect 19800 19796 19852 19805
rect 19984 19796 20036 19848
rect 20352 19796 20404 19848
rect 20536 19839 20588 19848
rect 20536 19805 20545 19839
rect 20545 19805 20579 19839
rect 20579 19805 20588 19839
rect 20536 19796 20588 19805
rect 20996 19796 21048 19848
rect 21272 19796 21324 19848
rect 22100 19864 22152 19916
rect 22560 19864 22612 19916
rect 21732 19839 21784 19848
rect 21732 19805 21741 19839
rect 21741 19805 21775 19839
rect 21775 19805 21784 19839
rect 21732 19796 21784 19805
rect 22468 19796 22520 19848
rect 23112 19839 23164 19848
rect 23112 19805 23121 19839
rect 23121 19805 23155 19839
rect 23155 19805 23164 19839
rect 23112 19796 23164 19805
rect 23756 19864 23808 19916
rect 23388 19839 23440 19848
rect 23388 19805 23397 19839
rect 23397 19805 23431 19839
rect 23431 19805 23440 19839
rect 23388 19796 23440 19805
rect 26148 20000 26200 20052
rect 25596 19932 25648 19984
rect 26056 19932 26108 19984
rect 23940 19796 23992 19848
rect 24492 19796 24544 19848
rect 26700 19932 26752 19984
rect 26976 19932 27028 19984
rect 26516 19796 26568 19848
rect 27436 19932 27488 19984
rect 28080 20000 28132 20052
rect 27252 19796 27304 19848
rect 27712 19796 27764 19848
rect 27988 19839 28040 19848
rect 27988 19805 27997 19839
rect 27997 19805 28031 19839
rect 28031 19805 28040 19839
rect 27988 19796 28040 19805
rect 20812 19728 20864 19780
rect 1400 19660 1452 19712
rect 10048 19660 10100 19712
rect 12072 19660 12124 19712
rect 12624 19660 12676 19712
rect 14372 19660 14424 19712
rect 14740 19660 14792 19712
rect 15016 19703 15068 19712
rect 15016 19669 15025 19703
rect 15025 19669 15059 19703
rect 15059 19669 15068 19703
rect 15016 19660 15068 19669
rect 15384 19703 15436 19712
rect 15384 19669 15393 19703
rect 15393 19669 15427 19703
rect 15427 19669 15436 19703
rect 15384 19660 15436 19669
rect 16212 19703 16264 19712
rect 16212 19669 16221 19703
rect 16221 19669 16255 19703
rect 16255 19669 16264 19703
rect 16212 19660 16264 19669
rect 16856 19660 16908 19712
rect 17776 19660 17828 19712
rect 19432 19660 19484 19712
rect 20352 19660 20404 19712
rect 24768 19728 24820 19780
rect 29460 19796 29512 19848
rect 28540 19728 28592 19780
rect 22100 19703 22152 19712
rect 22100 19669 22109 19703
rect 22109 19669 22143 19703
rect 22143 19669 22152 19703
rect 22100 19660 22152 19669
rect 25596 19660 25648 19712
rect 26976 19660 27028 19712
rect 28356 19703 28408 19712
rect 28356 19669 28365 19703
rect 28365 19669 28399 19703
rect 28399 19669 28408 19703
rect 28356 19660 28408 19669
rect 10880 19558 10932 19610
rect 10944 19558 10996 19610
rect 11008 19558 11060 19610
rect 11072 19558 11124 19610
rect 11136 19558 11188 19610
rect 20811 19558 20863 19610
rect 20875 19558 20927 19610
rect 20939 19558 20991 19610
rect 21003 19558 21055 19610
rect 21067 19558 21119 19610
rect 9220 19456 9272 19508
rect 12532 19456 12584 19508
rect 13544 19456 13596 19508
rect 14188 19456 14240 19508
rect 22008 19456 22060 19508
rect 22284 19456 22336 19508
rect 22744 19456 22796 19508
rect 24952 19456 25004 19508
rect 26240 19456 26292 19508
rect 28172 19456 28224 19508
rect 29184 19456 29236 19508
rect 15016 19388 15068 19440
rect 15568 19431 15620 19440
rect 15568 19397 15577 19431
rect 15577 19397 15611 19431
rect 15611 19397 15620 19431
rect 15568 19388 15620 19397
rect 17040 19388 17092 19440
rect 21180 19388 21232 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 9680 19363 9732 19372
rect 9680 19329 9689 19363
rect 9689 19329 9723 19363
rect 9723 19329 9732 19363
rect 9680 19320 9732 19329
rect 9864 19363 9916 19372
rect 9864 19329 9871 19363
rect 9871 19329 9916 19363
rect 9864 19320 9916 19329
rect 10048 19363 10100 19372
rect 10048 19329 10057 19363
rect 10057 19329 10091 19363
rect 10091 19329 10100 19363
rect 10048 19320 10100 19329
rect 10140 19363 10192 19372
rect 10140 19329 10154 19363
rect 10154 19329 10188 19363
rect 10188 19329 10192 19363
rect 10140 19320 10192 19329
rect 11888 19252 11940 19304
rect 10048 19184 10100 19236
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 11612 19116 11664 19168
rect 11888 19116 11940 19168
rect 13084 19363 13136 19372
rect 13084 19329 13093 19363
rect 13093 19329 13127 19363
rect 13127 19329 13136 19363
rect 13084 19320 13136 19329
rect 13912 19363 13964 19372
rect 13912 19329 13921 19363
rect 13921 19329 13955 19363
rect 13955 19329 13964 19363
rect 13912 19320 13964 19329
rect 14188 19320 14240 19372
rect 14740 19363 14792 19372
rect 14372 19294 14424 19346
rect 14740 19329 14749 19363
rect 14749 19329 14783 19363
rect 14783 19329 14792 19363
rect 14740 19320 14792 19329
rect 14924 19363 14976 19372
rect 14924 19329 14933 19363
rect 14933 19329 14967 19363
rect 14967 19329 14976 19363
rect 14924 19320 14976 19329
rect 16212 19320 16264 19372
rect 17316 19320 17368 19372
rect 17776 19363 17828 19372
rect 17776 19329 17783 19363
rect 17783 19329 17828 19363
rect 17776 19320 17828 19329
rect 15016 19252 15068 19304
rect 18052 19363 18104 19372
rect 18052 19329 18066 19363
rect 18066 19329 18100 19363
rect 18100 19329 18104 19363
rect 18052 19320 18104 19329
rect 20536 19320 20588 19372
rect 20720 19320 20772 19372
rect 23664 19388 23716 19440
rect 21916 19320 21968 19372
rect 22100 19363 22152 19372
rect 22100 19329 22134 19363
rect 22134 19329 22152 19363
rect 22100 19320 22152 19329
rect 24216 19363 24268 19372
rect 24216 19329 24250 19363
rect 24250 19329 24268 19363
rect 26240 19363 26292 19372
rect 24216 19320 24268 19329
rect 26240 19329 26249 19363
rect 26249 19329 26283 19363
rect 26283 19329 26292 19363
rect 26240 19320 26292 19329
rect 23664 19252 23716 19304
rect 23940 19295 23992 19304
rect 23940 19261 23949 19295
rect 23949 19261 23983 19295
rect 23983 19261 23992 19295
rect 23940 19252 23992 19261
rect 25688 19252 25740 19304
rect 28448 19320 28500 19372
rect 29000 19363 29052 19372
rect 29000 19329 29034 19363
rect 29034 19329 29052 19363
rect 29000 19320 29052 19329
rect 27528 19252 27580 19304
rect 17684 19184 17736 19236
rect 19156 19184 19208 19236
rect 20904 19184 20956 19236
rect 12532 19116 12584 19168
rect 13176 19116 13228 19168
rect 13820 19116 13872 19168
rect 17960 19116 18012 19168
rect 19524 19116 19576 19168
rect 21732 19116 21784 19168
rect 22008 19116 22060 19168
rect 23664 19116 23716 19168
rect 26332 19184 26384 19236
rect 28448 19184 28500 19236
rect 28724 19184 28776 19236
rect 5915 19014 5967 19066
rect 5979 19014 6031 19066
rect 6043 19014 6095 19066
rect 6107 19014 6159 19066
rect 6171 19014 6223 19066
rect 15846 19014 15898 19066
rect 15910 19014 15962 19066
rect 15974 19014 16026 19066
rect 16038 19014 16090 19066
rect 16102 19014 16154 19066
rect 25776 19014 25828 19066
rect 25840 19014 25892 19066
rect 25904 19014 25956 19066
rect 25968 19014 26020 19066
rect 26032 19014 26084 19066
rect 10140 18912 10192 18964
rect 10508 18912 10560 18964
rect 11796 18912 11848 18964
rect 11888 18912 11940 18964
rect 15384 18955 15436 18964
rect 13360 18844 13412 18896
rect 14188 18844 14240 18896
rect 14464 18844 14516 18896
rect 15384 18921 15393 18955
rect 15393 18921 15427 18955
rect 15427 18921 15436 18955
rect 15384 18912 15436 18921
rect 21732 18912 21784 18964
rect 25044 18912 25096 18964
rect 25320 18912 25372 18964
rect 25504 18912 25556 18964
rect 26516 18912 26568 18964
rect 16396 18844 16448 18896
rect 20720 18844 20772 18896
rect 13084 18776 13136 18828
rect 14556 18776 14608 18828
rect 15384 18776 15436 18828
rect 16028 18776 16080 18828
rect 17500 18776 17552 18828
rect 9312 18708 9364 18760
rect 11612 18708 11664 18760
rect 11888 18708 11940 18760
rect 12256 18708 12308 18760
rect 12716 18708 12768 18760
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 14096 18751 14148 18760
rect 14096 18717 14105 18751
rect 14105 18717 14139 18751
rect 14139 18717 14148 18751
rect 14096 18708 14148 18717
rect 14740 18708 14792 18760
rect 15476 18751 15528 18760
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 15568 18751 15620 18760
rect 15568 18717 15577 18751
rect 15577 18717 15611 18751
rect 15611 18717 15620 18751
rect 15568 18708 15620 18717
rect 16120 18708 16172 18760
rect 17316 18708 17368 18760
rect 17776 18751 17828 18760
rect 17776 18717 17783 18751
rect 17783 18717 17828 18751
rect 17776 18708 17828 18717
rect 18052 18708 18104 18760
rect 18696 18708 18748 18760
rect 19800 18708 19852 18760
rect 12256 18572 12308 18624
rect 17132 18640 17184 18692
rect 17868 18683 17920 18692
rect 17868 18649 17877 18683
rect 17877 18649 17911 18683
rect 17911 18649 17920 18683
rect 17868 18640 17920 18649
rect 20444 18640 20496 18692
rect 20904 18776 20956 18828
rect 22192 18776 22244 18828
rect 23204 18776 23256 18828
rect 23388 18776 23440 18828
rect 25504 18819 25556 18828
rect 25504 18785 25513 18819
rect 25513 18785 25547 18819
rect 25547 18785 25556 18819
rect 25504 18776 25556 18785
rect 21272 18708 21324 18760
rect 23664 18751 23716 18760
rect 23664 18717 23673 18751
rect 23673 18717 23707 18751
rect 23707 18717 23716 18751
rect 23664 18708 23716 18717
rect 24860 18708 24912 18760
rect 25136 18751 25188 18760
rect 25136 18717 25145 18751
rect 25145 18717 25179 18751
rect 25179 18717 25188 18751
rect 25136 18708 25188 18717
rect 25320 18751 25372 18760
rect 25320 18717 25329 18751
rect 25329 18717 25363 18751
rect 25363 18717 25372 18751
rect 25320 18708 25372 18717
rect 25596 18708 25648 18760
rect 26424 18776 26476 18828
rect 29000 18776 29052 18828
rect 29368 18776 29420 18828
rect 25872 18708 25924 18760
rect 27160 18708 27212 18760
rect 27620 18751 27672 18760
rect 27620 18717 27629 18751
rect 27629 18717 27663 18751
rect 27663 18717 27672 18751
rect 27620 18708 27672 18717
rect 28448 18708 28500 18760
rect 28632 18708 28684 18760
rect 26240 18640 26292 18692
rect 29736 18640 29788 18692
rect 14280 18572 14332 18624
rect 15200 18572 15252 18624
rect 17684 18572 17736 18624
rect 18236 18615 18288 18624
rect 18236 18581 18245 18615
rect 18245 18581 18279 18615
rect 18279 18581 18288 18615
rect 18236 18572 18288 18581
rect 19340 18615 19392 18624
rect 19340 18581 19349 18615
rect 19349 18581 19383 18615
rect 19383 18581 19392 18615
rect 19340 18572 19392 18581
rect 20628 18572 20680 18624
rect 22744 18572 22796 18624
rect 23020 18572 23072 18624
rect 23940 18572 23992 18624
rect 24860 18572 24912 18624
rect 29460 18572 29512 18624
rect 10880 18470 10932 18522
rect 10944 18470 10996 18522
rect 11008 18470 11060 18522
rect 11072 18470 11124 18522
rect 11136 18470 11188 18522
rect 20811 18470 20863 18522
rect 20875 18470 20927 18522
rect 20939 18470 20991 18522
rect 21003 18470 21055 18522
rect 21067 18470 21119 18522
rect 10692 18368 10744 18420
rect 12256 18368 12308 18420
rect 2688 18300 2740 18352
rect 13084 18300 13136 18352
rect 15108 18300 15160 18352
rect 7748 18275 7800 18284
rect 7748 18241 7757 18275
rect 7757 18241 7791 18275
rect 7791 18241 7800 18275
rect 7748 18232 7800 18241
rect 8024 18275 8076 18284
rect 8024 18241 8058 18275
rect 8058 18241 8076 18275
rect 11704 18275 11756 18284
rect 8024 18232 8076 18241
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 13176 18275 13228 18284
rect 10784 18164 10836 18216
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 15292 18275 15344 18284
rect 9772 18096 9824 18148
rect 13544 18096 13596 18148
rect 15292 18241 15301 18275
rect 15301 18241 15335 18275
rect 15335 18241 15344 18275
rect 15292 18232 15344 18241
rect 15568 18368 15620 18420
rect 17132 18368 17184 18420
rect 17684 18368 17736 18420
rect 20444 18368 20496 18420
rect 22008 18368 22060 18420
rect 24216 18368 24268 18420
rect 29736 18411 29788 18420
rect 16672 18343 16724 18352
rect 16672 18309 16681 18343
rect 16681 18309 16715 18343
rect 16715 18309 16724 18343
rect 16672 18300 16724 18309
rect 16120 18232 16172 18284
rect 15108 18207 15160 18216
rect 15108 18173 15117 18207
rect 15117 18173 15151 18207
rect 15151 18173 15160 18207
rect 15108 18164 15160 18173
rect 16028 18164 16080 18216
rect 16488 18164 16540 18216
rect 16948 18275 17000 18284
rect 16948 18241 16957 18275
rect 16957 18241 16991 18275
rect 16991 18241 17000 18275
rect 16948 18232 17000 18241
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 18328 18300 18380 18352
rect 19340 18300 19392 18352
rect 17224 18232 17276 18241
rect 17960 18275 18012 18284
rect 17960 18241 17994 18275
rect 17994 18241 18012 18275
rect 17960 18232 18012 18241
rect 20812 18232 20864 18284
rect 22468 18232 22520 18284
rect 23112 18232 23164 18284
rect 23388 18275 23440 18284
rect 23388 18241 23397 18275
rect 23397 18241 23431 18275
rect 23431 18241 23440 18275
rect 23388 18232 23440 18241
rect 23848 18232 23900 18284
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 24952 18232 25004 18284
rect 27620 18300 27672 18352
rect 27988 18300 28040 18352
rect 29092 18300 29144 18352
rect 29736 18377 29745 18411
rect 29745 18377 29779 18411
rect 29779 18377 29788 18411
rect 29736 18368 29788 18377
rect 27252 18232 27304 18284
rect 28356 18232 28408 18284
rect 28724 18232 28776 18284
rect 29460 18232 29512 18284
rect 16764 18164 16816 18216
rect 19340 18164 19392 18216
rect 23204 18164 23256 18216
rect 23756 18207 23808 18216
rect 23756 18173 23765 18207
rect 23765 18173 23799 18207
rect 23799 18173 23808 18207
rect 23756 18164 23808 18173
rect 8392 18028 8444 18080
rect 11520 18071 11572 18080
rect 11520 18037 11529 18071
rect 11529 18037 11563 18071
rect 11563 18037 11572 18071
rect 11520 18028 11572 18037
rect 11796 18028 11848 18080
rect 12256 18028 12308 18080
rect 12440 18071 12492 18080
rect 12440 18037 12449 18071
rect 12449 18037 12483 18071
rect 12483 18037 12492 18071
rect 15752 18096 15804 18148
rect 15844 18096 15896 18148
rect 12440 18028 12492 18037
rect 15108 18028 15160 18080
rect 15660 18028 15712 18080
rect 19432 18096 19484 18148
rect 23020 18096 23072 18148
rect 21180 18028 21232 18080
rect 21456 18028 21508 18080
rect 22192 18028 22244 18080
rect 24860 18028 24912 18080
rect 28264 18164 28316 18216
rect 26332 18096 26384 18148
rect 28540 18139 28592 18148
rect 28540 18105 28549 18139
rect 28549 18105 28583 18139
rect 28583 18105 28592 18139
rect 28540 18096 28592 18105
rect 29092 18096 29144 18148
rect 28080 18028 28132 18080
rect 5915 17926 5967 17978
rect 5979 17926 6031 17978
rect 6043 17926 6095 17978
rect 6107 17926 6159 17978
rect 6171 17926 6223 17978
rect 15846 17926 15898 17978
rect 15910 17926 15962 17978
rect 15974 17926 16026 17978
rect 16038 17926 16090 17978
rect 16102 17926 16154 17978
rect 25776 17926 25828 17978
rect 25840 17926 25892 17978
rect 25904 17926 25956 17978
rect 25968 17926 26020 17978
rect 26032 17926 26084 17978
rect 8024 17824 8076 17876
rect 12716 17867 12768 17876
rect 12716 17833 12725 17867
rect 12725 17833 12759 17867
rect 12759 17833 12768 17867
rect 12716 17824 12768 17833
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 15752 17824 15804 17876
rect 19524 17799 19576 17808
rect 19524 17765 19533 17799
rect 19533 17765 19567 17799
rect 19567 17765 19576 17799
rect 19524 17756 19576 17765
rect 20168 17824 20220 17876
rect 20628 17824 20680 17876
rect 20812 17867 20864 17876
rect 20812 17833 20821 17867
rect 20821 17833 20855 17867
rect 20855 17833 20864 17867
rect 20812 17824 20864 17833
rect 21732 17824 21784 17876
rect 22376 17867 22428 17876
rect 22376 17833 22385 17867
rect 22385 17833 22419 17867
rect 22419 17833 22428 17867
rect 22376 17824 22428 17833
rect 21088 17756 21140 17808
rect 21180 17756 21232 17808
rect 21548 17756 21600 17808
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 1768 17663 1820 17672
rect 1768 17629 1777 17663
rect 1777 17629 1811 17663
rect 1811 17629 1820 17663
rect 1768 17620 1820 17629
rect 11428 17688 11480 17740
rect 11796 17731 11848 17740
rect 11796 17697 11805 17731
rect 11805 17697 11839 17731
rect 11839 17697 11848 17731
rect 11796 17688 11848 17697
rect 11888 17688 11940 17740
rect 13360 17731 13412 17740
rect 13360 17697 13369 17731
rect 13369 17697 13403 17731
rect 13403 17697 13412 17731
rect 13360 17688 13412 17697
rect 10232 17620 10284 17672
rect 9680 17595 9732 17604
rect 9680 17561 9689 17595
rect 9689 17561 9723 17595
rect 9723 17561 9732 17595
rect 9680 17552 9732 17561
rect 10600 17552 10652 17604
rect 11244 17620 11296 17672
rect 11520 17620 11572 17672
rect 13452 17620 13504 17672
rect 14648 17688 14700 17740
rect 16396 17731 16448 17740
rect 16396 17697 16405 17731
rect 16405 17697 16439 17731
rect 16439 17697 16448 17731
rect 16396 17688 16448 17697
rect 19248 17688 19300 17740
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 14556 17663 14608 17672
rect 14556 17629 14565 17663
rect 14565 17629 14599 17663
rect 14599 17629 14608 17663
rect 15200 17663 15252 17672
rect 14556 17620 14608 17629
rect 15200 17629 15209 17663
rect 15209 17629 15243 17663
rect 15243 17629 15252 17663
rect 15200 17620 15252 17629
rect 16212 17663 16264 17672
rect 16212 17629 16221 17663
rect 16221 17629 16255 17663
rect 16255 17629 16264 17663
rect 16212 17620 16264 17629
rect 18328 17620 18380 17672
rect 20352 17688 20404 17740
rect 21456 17688 21508 17740
rect 22008 17756 22060 17808
rect 22744 17824 22796 17876
rect 23572 17867 23624 17876
rect 22836 17756 22888 17808
rect 23572 17833 23581 17867
rect 23581 17833 23615 17867
rect 23615 17833 23624 17867
rect 23572 17824 23624 17833
rect 25320 17824 25372 17876
rect 25688 17824 25740 17876
rect 23572 17688 23624 17740
rect 25596 17688 25648 17740
rect 27620 17756 27672 17808
rect 29460 17756 29512 17808
rect 1400 17484 1452 17536
rect 9772 17527 9824 17536
rect 9772 17493 9781 17527
rect 9781 17493 9815 17527
rect 9815 17493 9824 17527
rect 9772 17484 9824 17493
rect 11336 17484 11388 17536
rect 11520 17484 11572 17536
rect 13728 17484 13780 17536
rect 18236 17552 18288 17604
rect 17132 17484 17184 17536
rect 17868 17484 17920 17536
rect 20076 17552 20128 17604
rect 20628 17663 20680 17672
rect 20628 17629 20661 17663
rect 20661 17629 20680 17663
rect 21640 17663 21692 17672
rect 20628 17620 20680 17629
rect 21640 17629 21649 17663
rect 21649 17629 21683 17663
rect 21683 17629 21692 17663
rect 21640 17620 21692 17629
rect 21732 17620 21784 17672
rect 22008 17663 22060 17672
rect 20812 17552 20864 17604
rect 21548 17552 21600 17604
rect 22008 17629 22017 17663
rect 22017 17629 22051 17663
rect 22051 17629 22060 17663
rect 22008 17620 22060 17629
rect 22192 17663 22244 17672
rect 22192 17629 22201 17663
rect 22201 17629 22235 17663
rect 22235 17629 22244 17663
rect 22836 17663 22888 17672
rect 22192 17620 22244 17629
rect 22836 17629 22845 17663
rect 22845 17629 22879 17663
rect 22879 17629 22888 17663
rect 22836 17620 22888 17629
rect 24216 17620 24268 17672
rect 23664 17552 23716 17604
rect 26056 17620 26108 17672
rect 21272 17484 21324 17536
rect 23112 17484 23164 17536
rect 25044 17552 25096 17604
rect 24952 17484 25004 17536
rect 26976 17688 27028 17740
rect 27528 17731 27580 17740
rect 27528 17697 27537 17731
rect 27537 17697 27571 17731
rect 27571 17697 27580 17731
rect 27528 17688 27580 17697
rect 27988 17688 28040 17740
rect 28816 17688 28868 17740
rect 27620 17620 27672 17672
rect 28540 17620 28592 17672
rect 28356 17552 28408 17604
rect 26332 17484 26384 17536
rect 26424 17484 26476 17536
rect 27896 17484 27948 17536
rect 10880 17382 10932 17434
rect 10944 17382 10996 17434
rect 11008 17382 11060 17434
rect 11072 17382 11124 17434
rect 11136 17382 11188 17434
rect 20811 17382 20863 17434
rect 20875 17382 20927 17434
rect 20939 17382 20991 17434
rect 21003 17382 21055 17434
rect 21067 17382 21119 17434
rect 1584 17280 1636 17332
rect 1400 17187 1452 17196
rect 1400 17153 1409 17187
rect 1409 17153 1443 17187
rect 1443 17153 1452 17187
rect 1400 17144 1452 17153
rect 1492 17144 1544 17196
rect 8392 17144 8444 17196
rect 9312 17144 9364 17196
rect 10416 17076 10468 17128
rect 11704 17280 11756 17332
rect 12440 17323 12492 17332
rect 12440 17289 12449 17323
rect 12449 17289 12483 17323
rect 12483 17289 12492 17323
rect 13728 17323 13780 17332
rect 12440 17280 12492 17289
rect 13728 17289 13737 17323
rect 13737 17289 13771 17323
rect 13771 17289 13780 17323
rect 13728 17280 13780 17289
rect 15384 17280 15436 17332
rect 15476 17280 15528 17332
rect 17132 17323 17184 17332
rect 17132 17289 17141 17323
rect 17141 17289 17175 17323
rect 17175 17289 17184 17323
rect 17132 17280 17184 17289
rect 21640 17280 21692 17332
rect 21732 17280 21784 17332
rect 11796 17212 11848 17264
rect 13452 17144 13504 17196
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 1860 16940 1912 16992
rect 9772 16940 9824 16992
rect 9864 16940 9916 16992
rect 10508 16940 10560 16992
rect 11612 16940 11664 16992
rect 12624 17076 12676 17128
rect 14372 17144 14424 17196
rect 15752 17187 15804 17196
rect 15752 17153 15761 17187
rect 15761 17153 15795 17187
rect 15795 17153 15804 17187
rect 15752 17144 15804 17153
rect 16764 17212 16816 17264
rect 17040 17255 17092 17264
rect 17040 17221 17049 17255
rect 17049 17221 17083 17255
rect 17083 17221 17092 17255
rect 17040 17212 17092 17221
rect 16672 17144 16724 17196
rect 17868 17187 17920 17196
rect 17868 17153 17877 17187
rect 17877 17153 17911 17187
rect 17911 17153 17920 17187
rect 17868 17144 17920 17153
rect 19432 17187 19484 17196
rect 19432 17153 19441 17187
rect 19441 17153 19475 17187
rect 19475 17153 19484 17187
rect 19432 17144 19484 17153
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 20996 17187 21048 17196
rect 20996 17153 21005 17187
rect 21005 17153 21039 17187
rect 21039 17153 21048 17187
rect 20996 17144 21048 17153
rect 21456 17144 21508 17196
rect 22376 17144 22428 17196
rect 23204 17212 23256 17264
rect 25044 17280 25096 17332
rect 26240 17280 26292 17332
rect 27252 17280 27304 17332
rect 23112 17187 23164 17196
rect 12716 17008 12768 17060
rect 16856 17076 16908 17128
rect 17500 17076 17552 17128
rect 19984 17076 20036 17128
rect 21180 17119 21232 17128
rect 21180 17085 21189 17119
rect 21189 17085 21223 17119
rect 21223 17085 21232 17119
rect 21180 17076 21232 17085
rect 22468 17076 22520 17128
rect 23112 17153 23121 17187
rect 23121 17153 23155 17187
rect 23155 17153 23164 17187
rect 23112 17144 23164 17153
rect 25504 17144 25556 17196
rect 27160 17144 27212 17196
rect 28080 17144 28132 17196
rect 28448 17144 28500 17196
rect 28724 17144 28776 17196
rect 23020 17076 23072 17128
rect 23756 17119 23808 17128
rect 23756 17085 23765 17119
rect 23765 17085 23799 17119
rect 23799 17085 23808 17119
rect 23756 17076 23808 17085
rect 27436 17076 27488 17128
rect 27988 17076 28040 17128
rect 15936 17008 15988 17060
rect 21640 17008 21692 17060
rect 22376 17008 22428 17060
rect 23388 17008 23440 17060
rect 15016 16983 15068 16992
rect 15016 16949 15025 16983
rect 15025 16949 15059 16983
rect 15059 16949 15068 16983
rect 15016 16940 15068 16949
rect 15660 16940 15712 16992
rect 20352 16940 20404 16992
rect 20904 16940 20956 16992
rect 21732 16940 21784 16992
rect 25688 16940 25740 16992
rect 29276 16940 29328 16992
rect 29552 16940 29604 16992
rect 5915 16838 5967 16890
rect 5979 16838 6031 16890
rect 6043 16838 6095 16890
rect 6107 16838 6159 16890
rect 6171 16838 6223 16890
rect 15846 16838 15898 16890
rect 15910 16838 15962 16890
rect 15974 16838 16026 16890
rect 16038 16838 16090 16890
rect 16102 16838 16154 16890
rect 25776 16838 25828 16890
rect 25840 16838 25892 16890
rect 25904 16838 25956 16890
rect 25968 16838 26020 16890
rect 26032 16838 26084 16890
rect 9864 16736 9916 16788
rect 10416 16779 10468 16788
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 10416 16745 10425 16779
rect 10425 16745 10459 16779
rect 10459 16745 10468 16779
rect 10416 16736 10468 16745
rect 10692 16736 10744 16788
rect 11796 16736 11848 16788
rect 13452 16779 13504 16788
rect 13452 16745 13461 16779
rect 13461 16745 13495 16779
rect 13495 16745 13504 16779
rect 13452 16736 13504 16745
rect 14740 16736 14792 16788
rect 11612 16668 11664 16720
rect 12716 16668 12768 16720
rect 10784 16600 10836 16652
rect 11336 16643 11388 16652
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 9864 16575 9916 16584
rect 9864 16541 9873 16575
rect 9873 16541 9907 16575
rect 9907 16541 9916 16575
rect 9864 16532 9916 16541
rect 10140 16532 10192 16584
rect 10508 16464 10560 16516
rect 11336 16609 11345 16643
rect 11345 16609 11379 16643
rect 11379 16609 11388 16643
rect 11336 16600 11388 16609
rect 11888 16600 11940 16652
rect 12440 16600 12492 16652
rect 12624 16643 12676 16652
rect 12624 16609 12633 16643
rect 12633 16609 12667 16643
rect 12667 16609 12676 16643
rect 12624 16600 12676 16609
rect 14096 16600 14148 16652
rect 15384 16668 15436 16720
rect 23112 16736 23164 16788
rect 23480 16736 23532 16788
rect 24308 16736 24360 16788
rect 27528 16736 27580 16788
rect 28724 16736 28776 16788
rect 29368 16736 29420 16788
rect 16580 16600 16632 16652
rect 20352 16600 20404 16652
rect 11244 16575 11296 16584
rect 11244 16541 11253 16575
rect 11253 16541 11287 16575
rect 11287 16541 11296 16575
rect 11244 16532 11296 16541
rect 15292 16575 15344 16584
rect 12440 16396 12492 16448
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15292 16532 15344 16541
rect 15936 16532 15988 16584
rect 16488 16532 16540 16584
rect 19340 16532 19392 16584
rect 19892 16532 19944 16584
rect 15384 16464 15436 16516
rect 19524 16507 19576 16516
rect 19524 16473 19558 16507
rect 19558 16473 19576 16507
rect 19524 16464 19576 16473
rect 20996 16600 21048 16652
rect 21272 16575 21324 16584
rect 21272 16541 21281 16575
rect 21281 16541 21315 16575
rect 21315 16541 21324 16575
rect 21272 16532 21324 16541
rect 21456 16600 21508 16652
rect 21640 16575 21692 16584
rect 14096 16439 14148 16448
rect 14096 16405 14105 16439
rect 14105 16405 14139 16439
rect 14139 16405 14148 16439
rect 14096 16396 14148 16405
rect 15016 16396 15068 16448
rect 18512 16396 18564 16448
rect 20352 16396 20404 16448
rect 21180 16464 21232 16516
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 22744 16668 22796 16720
rect 23388 16668 23440 16720
rect 22744 16575 22796 16584
rect 22744 16541 22753 16575
rect 22753 16541 22787 16575
rect 22787 16541 22796 16575
rect 22744 16532 22796 16541
rect 23112 16575 23164 16584
rect 23112 16541 23121 16575
rect 23121 16541 23155 16575
rect 23155 16541 23164 16575
rect 23112 16532 23164 16541
rect 22284 16464 22336 16516
rect 23388 16464 23440 16516
rect 23572 16600 23624 16652
rect 24308 16600 24360 16652
rect 27436 16668 27488 16720
rect 27620 16668 27672 16720
rect 28080 16668 28132 16720
rect 28264 16668 28316 16720
rect 24952 16575 25004 16584
rect 24952 16541 24961 16575
rect 24961 16541 24995 16575
rect 24995 16541 25004 16575
rect 24952 16532 25004 16541
rect 25688 16575 25740 16584
rect 25688 16541 25697 16575
rect 25697 16541 25731 16575
rect 25731 16541 25740 16575
rect 25688 16532 25740 16541
rect 26424 16464 26476 16516
rect 24124 16396 24176 16448
rect 27160 16532 27212 16584
rect 27252 16575 27304 16584
rect 27252 16541 27261 16575
rect 27261 16541 27295 16575
rect 27295 16541 27304 16575
rect 27988 16600 28040 16652
rect 27252 16532 27304 16541
rect 28264 16575 28316 16584
rect 27344 16396 27396 16448
rect 28264 16541 28273 16575
rect 28273 16541 28307 16575
rect 28307 16541 28316 16575
rect 28264 16532 28316 16541
rect 29000 16600 29052 16652
rect 29184 16532 29236 16584
rect 29828 16464 29880 16516
rect 29552 16396 29604 16448
rect 29644 16439 29696 16448
rect 29644 16405 29653 16439
rect 29653 16405 29687 16439
rect 29687 16405 29696 16439
rect 29644 16396 29696 16405
rect 10880 16294 10932 16346
rect 10944 16294 10996 16346
rect 11008 16294 11060 16346
rect 11072 16294 11124 16346
rect 11136 16294 11188 16346
rect 20811 16294 20863 16346
rect 20875 16294 20927 16346
rect 20939 16294 20991 16346
rect 21003 16294 21055 16346
rect 21067 16294 21119 16346
rect 11336 16192 11388 16244
rect 11980 16192 12032 16244
rect 10324 15988 10376 16040
rect 11704 16056 11756 16108
rect 15108 16192 15160 16244
rect 15384 16235 15436 16244
rect 15384 16201 15393 16235
rect 15393 16201 15427 16235
rect 15427 16201 15436 16235
rect 15384 16192 15436 16201
rect 17040 16235 17092 16244
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 19524 16235 19576 16244
rect 19524 16201 19533 16235
rect 19533 16201 19567 16235
rect 19567 16201 19576 16235
rect 19524 16192 19576 16201
rect 13728 16124 13780 16176
rect 18052 16124 18104 16176
rect 20352 16192 20404 16244
rect 22836 16192 22888 16244
rect 23112 16235 23164 16244
rect 23112 16201 23121 16235
rect 23121 16201 23155 16235
rect 23155 16201 23164 16235
rect 23112 16192 23164 16201
rect 24124 16192 24176 16244
rect 27160 16192 27212 16244
rect 28264 16192 28316 16244
rect 11888 15988 11940 16040
rect 13360 15988 13412 16040
rect 13820 16099 13872 16108
rect 13820 16065 13829 16099
rect 13829 16065 13863 16099
rect 13863 16065 13872 16099
rect 13820 16056 13872 16065
rect 14188 16099 14240 16108
rect 13728 15988 13780 16040
rect 14188 16065 14197 16099
rect 14197 16065 14231 16099
rect 14231 16065 14240 16099
rect 14188 16056 14240 16065
rect 16948 16056 17000 16108
rect 18512 16056 18564 16108
rect 18788 16099 18840 16108
rect 18788 16065 18797 16099
rect 18797 16065 18831 16099
rect 18831 16065 18840 16099
rect 18788 16056 18840 16065
rect 11704 15920 11756 15972
rect 12532 15920 12584 15972
rect 15936 15988 15988 16040
rect 14556 15920 14608 15972
rect 10508 15852 10560 15904
rect 12992 15852 13044 15904
rect 14924 15852 14976 15904
rect 16396 15988 16448 16040
rect 16672 15963 16724 15972
rect 16672 15929 16681 15963
rect 16681 15929 16715 15963
rect 16715 15929 16724 15963
rect 16672 15920 16724 15929
rect 16580 15852 16632 15904
rect 17500 15988 17552 16040
rect 19064 16099 19116 16108
rect 19064 16065 19073 16099
rect 19073 16065 19107 16099
rect 19107 16065 19116 16099
rect 19708 16124 19760 16176
rect 21180 16124 21232 16176
rect 19064 16056 19116 16065
rect 20352 16099 20404 16108
rect 20352 16065 20361 16099
rect 20361 16065 20395 16099
rect 20395 16065 20404 16099
rect 20352 16056 20404 16065
rect 21640 16056 21692 16108
rect 22192 16056 22244 16108
rect 23388 16056 23440 16108
rect 27344 16124 27396 16176
rect 27620 16124 27672 16176
rect 29644 16124 29696 16176
rect 25136 16099 25188 16108
rect 25136 16065 25170 16099
rect 25170 16065 25188 16099
rect 25136 16056 25188 16065
rect 27528 16056 27580 16108
rect 19616 15988 19668 16040
rect 20444 15988 20496 16040
rect 21364 15988 21416 16040
rect 21456 15988 21508 16040
rect 23756 15988 23808 16040
rect 24860 16031 24912 16040
rect 24860 15997 24869 16031
rect 24869 15997 24903 16031
rect 24903 15997 24912 16031
rect 24860 15988 24912 15997
rect 26148 15988 26200 16040
rect 27988 15988 28040 16040
rect 28448 16056 28500 16108
rect 19524 15920 19576 15972
rect 19984 15920 20036 15972
rect 28080 15920 28132 15972
rect 28264 15920 28316 15972
rect 19892 15852 19944 15904
rect 21180 15895 21232 15904
rect 21180 15861 21189 15895
rect 21189 15861 21223 15895
rect 21223 15861 21232 15895
rect 21180 15852 21232 15861
rect 22376 15852 22428 15904
rect 22836 15852 22888 15904
rect 26148 15852 26200 15904
rect 27252 15852 27304 15904
rect 5915 15750 5967 15802
rect 5979 15750 6031 15802
rect 6043 15750 6095 15802
rect 6107 15750 6159 15802
rect 6171 15750 6223 15802
rect 15846 15750 15898 15802
rect 15910 15750 15962 15802
rect 15974 15750 16026 15802
rect 16038 15750 16090 15802
rect 16102 15750 16154 15802
rect 25776 15750 25828 15802
rect 25840 15750 25892 15802
rect 25904 15750 25956 15802
rect 25968 15750 26020 15802
rect 26032 15750 26084 15802
rect 11520 15648 11572 15700
rect 11980 15648 12032 15700
rect 14188 15691 14240 15700
rect 14188 15657 14197 15691
rect 14197 15657 14231 15691
rect 14231 15657 14240 15691
rect 14188 15648 14240 15657
rect 18512 15691 18564 15700
rect 18512 15657 18521 15691
rect 18521 15657 18555 15691
rect 18555 15657 18564 15691
rect 18512 15648 18564 15657
rect 19064 15648 19116 15700
rect 10600 15580 10652 15632
rect 2688 15512 2740 15564
rect 12440 15580 12492 15632
rect 13268 15580 13320 15632
rect 13360 15580 13412 15632
rect 13912 15512 13964 15564
rect 16304 15580 16356 15632
rect 16580 15512 16632 15564
rect 18236 15512 18288 15564
rect 19156 15512 19208 15564
rect 23756 15648 23808 15700
rect 25136 15648 25188 15700
rect 28172 15648 28224 15700
rect 23020 15580 23072 15632
rect 28080 15623 28132 15632
rect 22284 15512 22336 15564
rect 28080 15589 28089 15623
rect 28089 15589 28123 15623
rect 28123 15589 28132 15623
rect 28080 15580 28132 15589
rect 28908 15580 28960 15632
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 9864 15444 9916 15496
rect 10048 15444 10100 15496
rect 11428 15487 11480 15496
rect 11428 15453 11437 15487
rect 11437 15453 11471 15487
rect 11471 15453 11480 15487
rect 11428 15444 11480 15453
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 11980 15444 12032 15496
rect 12808 15487 12860 15496
rect 12808 15453 12817 15487
rect 12817 15453 12851 15487
rect 12851 15453 12860 15487
rect 12808 15444 12860 15453
rect 12992 15487 13044 15496
rect 12992 15453 13001 15487
rect 13001 15453 13035 15487
rect 13035 15453 13044 15487
rect 12992 15444 13044 15453
rect 13360 15487 13412 15496
rect 13360 15453 13369 15487
rect 13369 15453 13403 15487
rect 13403 15453 13412 15487
rect 13360 15444 13412 15453
rect 14096 15444 14148 15496
rect 15660 15444 15712 15496
rect 17132 15487 17184 15496
rect 17132 15453 17141 15487
rect 17141 15453 17175 15487
rect 17175 15453 17184 15487
rect 17132 15444 17184 15453
rect 18788 15444 18840 15496
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 19708 15444 19760 15496
rect 22100 15444 22152 15496
rect 24124 15512 24176 15564
rect 23204 15444 23256 15496
rect 23388 15444 23440 15496
rect 23480 15444 23532 15496
rect 24400 15444 24452 15496
rect 1400 15308 1452 15360
rect 9956 15308 10008 15360
rect 11428 15308 11480 15360
rect 15016 15376 15068 15428
rect 19156 15376 19208 15428
rect 15200 15308 15252 15360
rect 15384 15351 15436 15360
rect 15384 15317 15393 15351
rect 15393 15317 15427 15351
rect 15427 15317 15436 15351
rect 15384 15308 15436 15317
rect 16580 15308 16632 15360
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 21824 15376 21876 15428
rect 23940 15376 23992 15428
rect 24860 15487 24912 15496
rect 24860 15453 24869 15487
rect 24869 15453 24903 15487
rect 24903 15453 24912 15487
rect 26148 15512 26200 15564
rect 24860 15444 24912 15453
rect 25320 15376 25372 15428
rect 22008 15308 22060 15360
rect 23020 15308 23072 15360
rect 23572 15308 23624 15360
rect 28448 15444 28500 15496
rect 28172 15376 28224 15428
rect 28908 15444 28960 15496
rect 29092 15376 29144 15428
rect 27252 15308 27304 15360
rect 29184 15308 29236 15360
rect 10880 15206 10932 15258
rect 10944 15206 10996 15258
rect 11008 15206 11060 15258
rect 11072 15206 11124 15258
rect 11136 15206 11188 15258
rect 20811 15206 20863 15258
rect 20875 15206 20927 15258
rect 20939 15206 20991 15258
rect 21003 15206 21055 15258
rect 21067 15206 21119 15258
rect 12992 15104 13044 15156
rect 13728 15104 13780 15156
rect 18144 15104 18196 15156
rect 18880 15104 18932 15156
rect 19156 15104 19208 15156
rect 19524 15104 19576 15156
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 13176 15036 13228 15088
rect 12072 15011 12124 15020
rect 12072 14977 12081 15011
rect 12081 14977 12115 15011
rect 12115 14977 12124 15011
rect 12072 14968 12124 14977
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 13728 14968 13780 15020
rect 14740 14968 14792 15020
rect 15384 15036 15436 15088
rect 20352 15036 20404 15088
rect 20904 15036 20956 15088
rect 15292 14968 15344 15020
rect 18512 14968 18564 15020
rect 9312 14900 9364 14952
rect 1584 14875 1636 14884
rect 1584 14841 1593 14875
rect 1593 14841 1627 14875
rect 1627 14841 1636 14875
rect 1584 14832 1636 14841
rect 11612 14900 11664 14952
rect 11428 14832 11480 14884
rect 10140 14764 10192 14816
rect 13544 14900 13596 14952
rect 13912 14832 13964 14884
rect 15108 14900 15160 14952
rect 16764 14943 16816 14952
rect 16764 14909 16773 14943
rect 16773 14909 16807 14943
rect 16807 14909 16816 14943
rect 16764 14900 16816 14909
rect 17960 14900 18012 14952
rect 14096 14764 14148 14816
rect 15752 14764 15804 14816
rect 16672 14764 16724 14816
rect 17132 14764 17184 14816
rect 18604 14764 18656 14816
rect 18880 15011 18932 15020
rect 18880 14977 18889 15011
rect 18889 14977 18923 15011
rect 18923 14977 18932 15011
rect 18880 14968 18932 14977
rect 19064 14968 19116 15020
rect 24216 15104 24268 15156
rect 26516 15104 26568 15156
rect 26792 15104 26844 15156
rect 21180 15036 21232 15088
rect 25504 15079 25556 15088
rect 25504 15045 25513 15079
rect 25513 15045 25547 15079
rect 25547 15045 25556 15079
rect 25504 15036 25556 15045
rect 26148 15079 26200 15088
rect 26148 15045 26157 15079
rect 26157 15045 26191 15079
rect 26191 15045 26200 15079
rect 26148 15036 26200 15045
rect 27436 15036 27488 15088
rect 18972 14943 19024 14952
rect 18972 14909 18981 14943
rect 18981 14909 19015 14943
rect 19015 14909 19024 14943
rect 18972 14900 19024 14909
rect 19340 14900 19392 14952
rect 19892 14943 19944 14952
rect 19892 14909 19901 14943
rect 19901 14909 19935 14943
rect 19935 14909 19944 14943
rect 19892 14900 19944 14909
rect 21088 14900 21140 14952
rect 21364 14968 21416 15020
rect 22284 14968 22336 15020
rect 22376 15011 22428 15020
rect 22376 14977 22385 15011
rect 22385 14977 22419 15011
rect 22419 14977 22428 15011
rect 22376 14968 22428 14977
rect 22836 14968 22888 15020
rect 23204 15011 23256 15020
rect 23204 14977 23213 15011
rect 23213 14977 23247 15011
rect 23247 14977 23256 15011
rect 23204 14968 23256 14977
rect 23480 14968 23532 15020
rect 24216 15011 24268 15020
rect 21272 14900 21324 14952
rect 22192 14943 22244 14952
rect 22192 14909 22201 14943
rect 22201 14909 22235 14943
rect 22235 14909 22244 14943
rect 22192 14900 22244 14909
rect 23112 14900 23164 14952
rect 24216 14977 24225 15011
rect 24225 14977 24259 15011
rect 24259 14977 24268 15011
rect 24216 14968 24268 14977
rect 25596 14968 25648 15020
rect 26516 14968 26568 15020
rect 28448 14968 28500 15020
rect 29000 15011 29052 15020
rect 29000 14977 29034 15011
rect 29034 14977 29052 15011
rect 29000 14968 29052 14977
rect 26332 14832 26384 14884
rect 26424 14832 26476 14884
rect 27712 14832 27764 14884
rect 20904 14764 20956 14816
rect 22376 14764 22428 14816
rect 23756 14807 23808 14816
rect 23756 14773 23765 14807
rect 23765 14773 23799 14807
rect 23799 14773 23808 14807
rect 23756 14764 23808 14773
rect 29092 14764 29144 14816
rect 5915 14662 5967 14714
rect 5979 14662 6031 14714
rect 6043 14662 6095 14714
rect 6107 14662 6159 14714
rect 6171 14662 6223 14714
rect 15846 14662 15898 14714
rect 15910 14662 15962 14714
rect 15974 14662 16026 14714
rect 16038 14662 16090 14714
rect 16102 14662 16154 14714
rect 25776 14662 25828 14714
rect 25840 14662 25892 14714
rect 25904 14662 25956 14714
rect 25968 14662 26020 14714
rect 26032 14662 26084 14714
rect 9312 14560 9364 14612
rect 11428 14560 11480 14612
rect 12164 14560 12216 14612
rect 12348 14603 12400 14612
rect 12348 14569 12357 14603
rect 12357 14569 12391 14603
rect 12391 14569 12400 14603
rect 12348 14560 12400 14569
rect 12808 14560 12860 14612
rect 15292 14603 15344 14612
rect 15292 14569 15301 14603
rect 15301 14569 15335 14603
rect 15335 14569 15344 14603
rect 15292 14560 15344 14569
rect 16580 14560 16632 14612
rect 16764 14560 16816 14612
rect 17316 14560 17368 14612
rect 18144 14560 18196 14612
rect 15752 14492 15804 14544
rect 12624 14424 12676 14476
rect 14096 14424 14148 14476
rect 15016 14424 15068 14476
rect 16488 14424 16540 14476
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 11612 14356 11664 14408
rect 13544 14356 13596 14408
rect 13728 14356 13780 14408
rect 15200 14356 15252 14408
rect 15660 14356 15712 14408
rect 18052 14492 18104 14544
rect 17960 14399 18012 14408
rect 10232 14288 10284 14340
rect 11796 14288 11848 14340
rect 15108 14220 15160 14272
rect 17960 14365 17969 14399
rect 17969 14365 18003 14399
rect 18003 14365 18012 14399
rect 17960 14356 18012 14365
rect 18512 14560 18564 14612
rect 20628 14560 20680 14612
rect 18328 14492 18380 14544
rect 18972 14492 19024 14544
rect 21272 14492 21324 14544
rect 18328 14399 18380 14408
rect 18328 14365 18337 14399
rect 18337 14365 18371 14399
rect 18371 14365 18380 14399
rect 18328 14356 18380 14365
rect 18512 14399 18564 14408
rect 18512 14365 18521 14399
rect 18521 14365 18555 14399
rect 18555 14365 18564 14399
rect 18512 14356 18564 14365
rect 19340 14356 19392 14408
rect 19984 14356 20036 14408
rect 20076 14356 20128 14408
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 21272 14399 21324 14408
rect 21272 14365 21281 14399
rect 21281 14365 21315 14399
rect 21315 14365 21324 14399
rect 21272 14356 21324 14365
rect 22008 14560 22060 14612
rect 26976 14560 27028 14612
rect 27620 14560 27672 14612
rect 27436 14424 27488 14476
rect 27712 14424 27764 14476
rect 23480 14356 23532 14408
rect 19708 14220 19760 14272
rect 21824 14263 21876 14272
rect 21824 14229 21833 14263
rect 21833 14229 21867 14263
rect 21867 14229 21876 14263
rect 21824 14220 21876 14229
rect 23572 14288 23624 14340
rect 25136 14288 25188 14340
rect 26792 14356 26844 14408
rect 27252 14399 27304 14408
rect 26976 14288 27028 14340
rect 27252 14365 27261 14399
rect 27261 14365 27295 14399
rect 27295 14365 27304 14399
rect 27252 14356 27304 14365
rect 28540 14356 28592 14408
rect 30104 14356 30156 14408
rect 27988 14288 28040 14340
rect 23388 14220 23440 14272
rect 25688 14220 25740 14272
rect 10880 14118 10932 14170
rect 10944 14118 10996 14170
rect 11008 14118 11060 14170
rect 11072 14118 11124 14170
rect 11136 14118 11188 14170
rect 20811 14118 20863 14170
rect 20875 14118 20927 14170
rect 20939 14118 20991 14170
rect 21003 14118 21055 14170
rect 21067 14118 21119 14170
rect 10232 14059 10284 14068
rect 10232 14025 10241 14059
rect 10241 14025 10275 14059
rect 10275 14025 10284 14059
rect 10232 14016 10284 14025
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 15660 14059 15712 14068
rect 15660 14025 15669 14059
rect 15669 14025 15703 14059
rect 15703 14025 15712 14059
rect 15660 14016 15712 14025
rect 16948 14016 17000 14068
rect 9496 13923 9548 13932
rect 9496 13889 9505 13923
rect 9505 13889 9539 13923
rect 9539 13889 9548 13923
rect 9496 13880 9548 13889
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 15476 13948 15528 14000
rect 18512 14016 18564 14068
rect 21916 14059 21968 14068
rect 21916 14025 21925 14059
rect 21925 14025 21959 14059
rect 21959 14025 21968 14059
rect 21916 14016 21968 14025
rect 24216 14016 24268 14068
rect 28172 14059 28224 14068
rect 28172 14025 28181 14059
rect 28181 14025 28215 14059
rect 28215 14025 28224 14059
rect 28172 14016 28224 14025
rect 11796 13923 11848 13932
rect 11796 13889 11805 13923
rect 11805 13889 11839 13923
rect 11839 13889 11848 13923
rect 11796 13880 11848 13889
rect 12164 13880 12216 13932
rect 14556 13923 14608 13932
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 20352 13948 20404 14000
rect 16580 13880 16632 13932
rect 17500 13923 17552 13932
rect 10140 13812 10192 13864
rect 10784 13855 10836 13864
rect 10784 13821 10793 13855
rect 10793 13821 10827 13855
rect 10827 13821 10836 13855
rect 10784 13812 10836 13821
rect 11612 13812 11664 13864
rect 15200 13812 15252 13864
rect 9956 13744 10008 13796
rect 15660 13744 15712 13796
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 17500 13880 17552 13889
rect 19892 13880 19944 13932
rect 20076 13880 20128 13932
rect 22376 13880 22428 13932
rect 23480 13948 23532 14000
rect 23940 13948 23992 14000
rect 24492 13948 24544 14000
rect 23756 13880 23808 13932
rect 24676 13880 24728 13932
rect 25596 13923 25648 13932
rect 17316 13812 17368 13864
rect 19340 13812 19392 13864
rect 25596 13889 25605 13923
rect 25605 13889 25639 13923
rect 25639 13889 25648 13923
rect 25596 13880 25648 13889
rect 25688 13880 25740 13932
rect 29920 13948 29972 14000
rect 26332 13923 26384 13932
rect 26332 13889 26341 13923
rect 26341 13889 26375 13923
rect 26375 13889 26384 13923
rect 26332 13880 26384 13889
rect 26516 13880 26568 13932
rect 27160 13880 27212 13932
rect 27896 13880 27948 13932
rect 28080 13880 28132 13932
rect 29736 13880 29788 13932
rect 21732 13744 21784 13796
rect 22100 13744 22152 13796
rect 12256 13676 12308 13728
rect 27528 13812 27580 13864
rect 28724 13855 28776 13864
rect 27620 13744 27672 13796
rect 28724 13821 28733 13855
rect 28733 13821 28767 13855
rect 28767 13821 28776 13855
rect 28724 13812 28776 13821
rect 27988 13744 28040 13796
rect 28172 13744 28224 13796
rect 28632 13744 28684 13796
rect 26608 13676 26660 13728
rect 26976 13676 27028 13728
rect 27712 13676 27764 13728
rect 28264 13676 28316 13728
rect 30104 13719 30156 13728
rect 30104 13685 30113 13719
rect 30113 13685 30147 13719
rect 30147 13685 30156 13719
rect 30104 13676 30156 13685
rect 5915 13574 5967 13626
rect 5979 13574 6031 13626
rect 6043 13574 6095 13626
rect 6107 13574 6159 13626
rect 6171 13574 6223 13626
rect 15846 13574 15898 13626
rect 15910 13574 15962 13626
rect 15974 13574 16026 13626
rect 16038 13574 16090 13626
rect 16102 13574 16154 13626
rect 25776 13574 25828 13626
rect 25840 13574 25892 13626
rect 25904 13574 25956 13626
rect 25968 13574 26020 13626
rect 26032 13574 26084 13626
rect 11428 13515 11480 13524
rect 11428 13481 11437 13515
rect 11437 13481 11471 13515
rect 11471 13481 11480 13515
rect 11428 13472 11480 13481
rect 11612 13472 11664 13524
rect 12348 13472 12400 13524
rect 14556 13472 14608 13524
rect 17500 13472 17552 13524
rect 19892 13515 19944 13524
rect 19892 13481 19901 13515
rect 19901 13481 19935 13515
rect 19935 13481 19944 13515
rect 19892 13472 19944 13481
rect 22744 13472 22796 13524
rect 23664 13472 23716 13524
rect 24860 13472 24912 13524
rect 25136 13515 25188 13524
rect 25136 13481 25145 13515
rect 25145 13481 25179 13515
rect 25179 13481 25188 13515
rect 25136 13472 25188 13481
rect 25228 13472 25280 13524
rect 1768 13268 1820 13320
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 11980 13404 12032 13456
rect 15016 13404 15068 13456
rect 18236 13447 18288 13456
rect 10692 13336 10744 13388
rect 12348 13336 12400 13388
rect 15200 13379 15252 13388
rect 15200 13345 15209 13379
rect 15209 13345 15243 13379
rect 15243 13345 15252 13379
rect 15200 13336 15252 13345
rect 18236 13413 18245 13447
rect 18245 13413 18279 13447
rect 18279 13413 18288 13447
rect 18236 13404 18288 13413
rect 20168 13404 20220 13456
rect 21456 13404 21508 13456
rect 19892 13336 19944 13388
rect 20536 13336 20588 13388
rect 21732 13336 21784 13388
rect 23204 13336 23256 13388
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 9956 13175 10008 13184
rect 9956 13141 9965 13175
rect 9965 13141 9999 13175
rect 9999 13141 10008 13175
rect 9956 13132 10008 13141
rect 10784 13268 10836 13320
rect 11796 13268 11848 13320
rect 11980 13268 12032 13320
rect 12256 13311 12308 13320
rect 12256 13277 12265 13311
rect 12265 13277 12299 13311
rect 12299 13277 12308 13311
rect 12256 13268 12308 13277
rect 13912 13268 13964 13320
rect 14648 13268 14700 13320
rect 15660 13268 15712 13320
rect 19248 13268 19300 13320
rect 20352 13268 20404 13320
rect 20444 13311 20496 13320
rect 20444 13277 20453 13311
rect 20453 13277 20487 13311
rect 20487 13277 20496 13311
rect 21364 13311 21416 13320
rect 20444 13268 20496 13277
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 21456 13268 21508 13320
rect 24400 13311 24452 13320
rect 12624 13200 12676 13252
rect 15568 13200 15620 13252
rect 17960 13200 18012 13252
rect 21180 13200 21232 13252
rect 21824 13200 21876 13252
rect 24400 13277 24409 13311
rect 24409 13277 24443 13311
rect 24443 13277 24452 13311
rect 24400 13268 24452 13277
rect 24676 13379 24728 13388
rect 24676 13345 24685 13379
rect 24685 13345 24719 13379
rect 24719 13345 24728 13379
rect 24676 13336 24728 13345
rect 24768 13311 24820 13320
rect 24768 13277 24777 13311
rect 24777 13277 24811 13311
rect 24811 13277 24820 13311
rect 24768 13268 24820 13277
rect 25688 13268 25740 13320
rect 26332 13268 26384 13320
rect 26792 13268 26844 13320
rect 26976 13268 27028 13320
rect 28172 13472 28224 13524
rect 28540 13472 28592 13524
rect 29000 13515 29052 13524
rect 29000 13481 29009 13515
rect 29009 13481 29043 13515
rect 29043 13481 29052 13515
rect 29000 13472 29052 13481
rect 28632 13404 28684 13456
rect 27436 13311 27488 13320
rect 27436 13277 27445 13311
rect 27445 13277 27479 13311
rect 27479 13277 27488 13311
rect 27436 13268 27488 13277
rect 27620 13311 27672 13320
rect 27620 13277 27629 13311
rect 27629 13277 27663 13311
rect 27663 13277 27672 13311
rect 27620 13268 27672 13277
rect 28264 13311 28316 13320
rect 28264 13277 28273 13311
rect 28273 13277 28307 13311
rect 28307 13277 28316 13311
rect 28264 13268 28316 13277
rect 28448 13311 28500 13320
rect 28448 13277 28461 13311
rect 28461 13277 28495 13311
rect 28495 13277 28500 13311
rect 28448 13268 28500 13277
rect 25596 13200 25648 13252
rect 11612 13132 11664 13184
rect 11796 13132 11848 13184
rect 15108 13175 15160 13184
rect 15108 13141 15117 13175
rect 15117 13141 15151 13175
rect 15151 13141 15160 13175
rect 15108 13132 15160 13141
rect 15384 13132 15436 13184
rect 18696 13132 18748 13184
rect 21272 13132 21324 13184
rect 24860 13132 24912 13184
rect 25320 13132 25372 13184
rect 27896 13200 27948 13252
rect 29092 13268 29144 13320
rect 29552 13311 29604 13320
rect 29552 13277 29561 13311
rect 29561 13277 29595 13311
rect 29595 13277 29604 13311
rect 29552 13268 29604 13277
rect 27804 13175 27856 13184
rect 27804 13141 27813 13175
rect 27813 13141 27847 13175
rect 27847 13141 27856 13175
rect 27804 13132 27856 13141
rect 27988 13132 28040 13184
rect 28816 13132 28868 13184
rect 10880 13030 10932 13082
rect 10944 13030 10996 13082
rect 11008 13030 11060 13082
rect 11072 13030 11124 13082
rect 11136 13030 11188 13082
rect 20811 13030 20863 13082
rect 20875 13030 20927 13082
rect 20939 13030 20991 13082
rect 21003 13030 21055 13082
rect 21067 13030 21119 13082
rect 10048 12971 10100 12980
rect 10048 12937 10057 12971
rect 10057 12937 10091 12971
rect 10091 12937 10100 12971
rect 10048 12928 10100 12937
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 13820 12928 13872 12937
rect 15108 12928 15160 12980
rect 15568 12971 15620 12980
rect 15568 12937 15577 12971
rect 15577 12937 15611 12971
rect 15611 12937 15620 12971
rect 15568 12928 15620 12937
rect 10600 12860 10652 12912
rect 11428 12860 11480 12912
rect 10140 12792 10192 12844
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 12716 12835 12768 12844
rect 12716 12801 12725 12835
rect 12725 12801 12759 12835
rect 12759 12801 12768 12835
rect 12716 12792 12768 12801
rect 16580 12928 16632 12980
rect 18328 12928 18380 12980
rect 16212 12860 16264 12912
rect 11520 12724 11572 12776
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 15016 12724 15068 12776
rect 16304 12792 16356 12844
rect 17040 12860 17092 12912
rect 18420 12860 18472 12912
rect 16856 12724 16908 12776
rect 12164 12588 12216 12640
rect 12348 12631 12400 12640
rect 12348 12597 12357 12631
rect 12357 12597 12391 12631
rect 12391 12597 12400 12631
rect 12348 12588 12400 12597
rect 16212 12588 16264 12640
rect 18052 12792 18104 12844
rect 18236 12792 18288 12844
rect 18696 12928 18748 12980
rect 18696 12835 18748 12844
rect 18696 12801 18705 12835
rect 18705 12801 18739 12835
rect 18739 12801 18748 12835
rect 18696 12792 18748 12801
rect 19708 12792 19760 12844
rect 20076 12792 20128 12844
rect 20628 12860 20680 12912
rect 19156 12724 19208 12776
rect 20904 12724 20956 12776
rect 18696 12588 18748 12640
rect 18880 12631 18932 12640
rect 18880 12597 18889 12631
rect 18889 12597 18923 12631
rect 18923 12597 18932 12631
rect 18880 12588 18932 12597
rect 19616 12588 19668 12640
rect 20076 12588 20128 12640
rect 20352 12631 20404 12640
rect 20352 12597 20361 12631
rect 20361 12597 20395 12631
rect 20395 12597 20404 12631
rect 20352 12588 20404 12597
rect 20628 12588 20680 12640
rect 21456 12792 21508 12844
rect 24216 12860 24268 12912
rect 24400 12860 24452 12912
rect 24768 12860 24820 12912
rect 22192 12724 22244 12776
rect 24492 12835 24544 12844
rect 24492 12801 24501 12835
rect 24501 12801 24535 12835
rect 24535 12801 24544 12835
rect 24492 12792 24544 12801
rect 24860 12792 24912 12844
rect 26240 12928 26292 12980
rect 27620 12928 27672 12980
rect 29552 12928 29604 12980
rect 29736 12971 29788 12980
rect 29736 12937 29745 12971
rect 29745 12937 29779 12971
rect 29779 12937 29788 12971
rect 29736 12928 29788 12937
rect 25412 12860 25464 12912
rect 25596 12835 25648 12844
rect 25596 12801 25605 12835
rect 25605 12801 25639 12835
rect 25639 12801 25648 12835
rect 25596 12792 25648 12801
rect 25412 12724 25464 12776
rect 26792 12792 26844 12844
rect 28724 12860 28776 12912
rect 28816 12860 28868 12912
rect 27804 12792 27856 12844
rect 28264 12792 28316 12844
rect 29184 12835 29236 12844
rect 29184 12801 29193 12835
rect 29193 12801 29227 12835
rect 29227 12801 29236 12835
rect 29184 12792 29236 12801
rect 30104 12792 30156 12844
rect 21456 12656 21508 12708
rect 22284 12656 22336 12708
rect 24676 12656 24728 12708
rect 21916 12588 21968 12640
rect 24860 12631 24912 12640
rect 24860 12597 24869 12631
rect 24869 12597 24903 12631
rect 24903 12597 24912 12631
rect 24860 12588 24912 12597
rect 28540 12724 28592 12776
rect 30012 12588 30064 12640
rect 5915 12486 5967 12538
rect 5979 12486 6031 12538
rect 6043 12486 6095 12538
rect 6107 12486 6159 12538
rect 6171 12486 6223 12538
rect 15846 12486 15898 12538
rect 15910 12486 15962 12538
rect 15974 12486 16026 12538
rect 16038 12486 16090 12538
rect 16102 12486 16154 12538
rect 25776 12486 25828 12538
rect 25840 12486 25892 12538
rect 25904 12486 25956 12538
rect 25968 12486 26020 12538
rect 26032 12486 26084 12538
rect 10140 12384 10192 12436
rect 12072 12384 12124 12436
rect 12348 12384 12400 12436
rect 15660 12384 15712 12436
rect 10600 12316 10652 12368
rect 10784 12291 10836 12300
rect 10784 12257 10793 12291
rect 10793 12257 10827 12291
rect 10827 12257 10836 12291
rect 10784 12248 10836 12257
rect 11888 12316 11940 12368
rect 17960 12384 18012 12436
rect 18696 12427 18748 12436
rect 18696 12393 18705 12427
rect 18705 12393 18739 12427
rect 18739 12393 18748 12427
rect 18696 12384 18748 12393
rect 19616 12384 19668 12436
rect 20628 12316 20680 12368
rect 21824 12384 21876 12436
rect 21548 12316 21600 12368
rect 24400 12316 24452 12368
rect 26516 12359 26568 12368
rect 11520 12248 11572 12300
rect 12256 12248 12308 12300
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 11336 12180 11388 12232
rect 12348 12180 12400 12232
rect 15016 12248 15068 12300
rect 16580 12248 16632 12300
rect 17316 12291 17368 12300
rect 17316 12257 17325 12291
rect 17325 12257 17359 12291
rect 17359 12257 17368 12291
rect 17316 12248 17368 12257
rect 20904 12248 20956 12300
rect 21364 12291 21416 12300
rect 15384 12223 15436 12232
rect 15384 12189 15393 12223
rect 15393 12189 15427 12223
rect 15427 12189 15436 12223
rect 15384 12180 15436 12189
rect 13912 12112 13964 12164
rect 14004 12112 14056 12164
rect 14924 12112 14976 12164
rect 16488 12155 16540 12164
rect 16488 12121 16497 12155
rect 16497 12121 16531 12155
rect 16531 12121 16540 12155
rect 16488 12112 16540 12121
rect 17040 12112 17092 12164
rect 11888 12087 11940 12096
rect 11888 12053 11897 12087
rect 11897 12053 11931 12087
rect 11931 12053 11940 12087
rect 11888 12044 11940 12053
rect 12072 12044 12124 12096
rect 13084 12087 13136 12096
rect 13084 12053 13093 12087
rect 13093 12053 13127 12087
rect 13127 12053 13136 12087
rect 13084 12044 13136 12053
rect 13728 12044 13780 12096
rect 15108 12044 15160 12096
rect 15660 12087 15712 12096
rect 15660 12053 15669 12087
rect 15669 12053 15703 12087
rect 15703 12053 15712 12087
rect 15660 12044 15712 12053
rect 16948 12044 17000 12096
rect 18880 12180 18932 12232
rect 19340 12180 19392 12232
rect 21364 12257 21373 12291
rect 21373 12257 21407 12291
rect 21407 12257 21416 12291
rect 21364 12248 21416 12257
rect 19524 12155 19576 12164
rect 19524 12121 19558 12155
rect 19558 12121 19576 12155
rect 22744 12180 22796 12232
rect 24216 12180 24268 12232
rect 26516 12325 26525 12359
rect 26525 12325 26559 12359
rect 26559 12325 26568 12359
rect 26516 12316 26568 12325
rect 24676 12291 24728 12300
rect 24676 12257 24685 12291
rect 24685 12257 24719 12291
rect 24719 12257 24728 12291
rect 24676 12248 24728 12257
rect 26240 12223 26292 12232
rect 19524 12112 19576 12121
rect 19800 12044 19852 12096
rect 22100 12112 22152 12164
rect 22284 12155 22336 12164
rect 22284 12121 22318 12155
rect 22318 12121 22336 12155
rect 22284 12112 22336 12121
rect 23756 12112 23808 12164
rect 24492 12112 24544 12164
rect 26240 12189 26249 12223
rect 26249 12189 26283 12223
rect 26283 12189 26292 12223
rect 26240 12180 26292 12189
rect 27804 12316 27856 12368
rect 26792 12223 26844 12232
rect 25688 12112 25740 12164
rect 26792 12189 26801 12223
rect 26801 12189 26835 12223
rect 26835 12189 26844 12223
rect 26792 12180 26844 12189
rect 21456 12044 21508 12096
rect 22376 12044 22428 12096
rect 25136 12087 25188 12096
rect 25136 12053 25145 12087
rect 25145 12053 25179 12087
rect 25179 12053 25188 12087
rect 25136 12044 25188 12053
rect 26148 12044 26200 12096
rect 27712 12180 27764 12232
rect 28264 12180 28316 12232
rect 29184 12180 29236 12232
rect 30196 12180 30248 12232
rect 27712 12044 27764 12096
rect 28908 12044 28960 12096
rect 10880 11942 10932 11994
rect 10944 11942 10996 11994
rect 11008 11942 11060 11994
rect 11072 11942 11124 11994
rect 11136 11942 11188 11994
rect 20811 11942 20863 11994
rect 20875 11942 20927 11994
rect 20939 11942 20991 11994
rect 21003 11942 21055 11994
rect 21067 11942 21119 11994
rect 12072 11883 12124 11892
rect 12072 11849 12081 11883
rect 12081 11849 12115 11883
rect 12115 11849 12124 11883
rect 12072 11840 12124 11849
rect 12716 11840 12768 11892
rect 13360 11840 13412 11892
rect 13728 11840 13780 11892
rect 14188 11840 14240 11892
rect 14740 11840 14792 11892
rect 15108 11883 15160 11892
rect 9864 11815 9916 11824
rect 9864 11781 9873 11815
rect 9873 11781 9907 11815
rect 9907 11781 9916 11815
rect 9864 11772 9916 11781
rect 14464 11772 14516 11824
rect 14648 11772 14700 11824
rect 11428 11704 11480 11756
rect 12164 11747 12216 11756
rect 12164 11713 12173 11747
rect 12173 11713 12207 11747
rect 12207 11713 12216 11747
rect 12164 11704 12216 11713
rect 13084 11747 13136 11756
rect 13084 11713 13093 11747
rect 13093 11713 13127 11747
rect 13127 11713 13136 11747
rect 13084 11704 13136 11713
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 16488 11840 16540 11892
rect 19524 11883 19576 11892
rect 19524 11849 19533 11883
rect 19533 11849 19567 11883
rect 19567 11849 19576 11883
rect 19524 11840 19576 11849
rect 14004 11679 14056 11688
rect 14004 11645 14013 11679
rect 14013 11645 14047 11679
rect 14047 11645 14056 11679
rect 14004 11636 14056 11645
rect 14188 11679 14240 11688
rect 14188 11645 14197 11679
rect 14197 11645 14231 11679
rect 14231 11645 14240 11679
rect 14188 11636 14240 11645
rect 15016 11636 15068 11688
rect 16212 11704 16264 11756
rect 16672 11747 16724 11756
rect 16672 11713 16681 11747
rect 16681 11713 16715 11747
rect 16715 11713 16724 11747
rect 16672 11704 16724 11713
rect 16304 11636 16356 11688
rect 16948 11747 17000 11756
rect 16948 11713 16982 11747
rect 16982 11713 17000 11747
rect 16948 11704 17000 11713
rect 18236 11772 18288 11824
rect 18052 11704 18104 11756
rect 18788 11747 18840 11756
rect 18788 11713 18797 11747
rect 18797 11713 18831 11747
rect 18831 11713 18840 11747
rect 18788 11704 18840 11713
rect 20352 11772 20404 11824
rect 19156 11679 19208 11688
rect 19156 11645 19165 11679
rect 19165 11645 19199 11679
rect 19199 11645 19208 11679
rect 19156 11636 19208 11645
rect 19800 11704 19852 11756
rect 22284 11840 22336 11892
rect 25320 11883 25372 11892
rect 21824 11772 21876 11824
rect 21916 11772 21968 11824
rect 25320 11849 25329 11883
rect 25329 11849 25363 11883
rect 25363 11849 25372 11883
rect 25320 11840 25372 11849
rect 24860 11772 24912 11824
rect 25504 11772 25556 11824
rect 20996 11704 21048 11756
rect 21456 11704 21508 11756
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22100 11704 22152 11713
rect 22376 11747 22428 11756
rect 22376 11713 22410 11747
rect 22410 11713 22428 11747
rect 23940 11747 23992 11756
rect 22376 11704 22428 11713
rect 23940 11713 23949 11747
rect 23949 11713 23983 11747
rect 23983 11713 23992 11747
rect 23940 11704 23992 11713
rect 27712 11747 27764 11756
rect 20812 11679 20864 11688
rect 20812 11645 20821 11679
rect 20821 11645 20855 11679
rect 20855 11645 20864 11679
rect 20812 11636 20864 11645
rect 27712 11713 27721 11747
rect 27721 11713 27755 11747
rect 27755 11713 27764 11747
rect 27712 11704 27764 11713
rect 28540 11772 28592 11824
rect 28080 11747 28132 11756
rect 28080 11713 28089 11747
rect 28089 11713 28123 11747
rect 28123 11713 28132 11747
rect 28080 11704 28132 11713
rect 29000 11747 29052 11756
rect 29000 11713 29034 11747
rect 29034 11713 29052 11747
rect 29000 11704 29052 11713
rect 27620 11636 27672 11688
rect 28724 11679 28776 11688
rect 21272 11568 21324 11620
rect 9588 11500 9640 11552
rect 15292 11500 15344 11552
rect 15660 11500 15712 11552
rect 26884 11568 26936 11620
rect 28724 11645 28733 11679
rect 28733 11645 28767 11679
rect 28767 11645 28776 11679
rect 28724 11636 28776 11645
rect 28632 11568 28684 11620
rect 25596 11500 25648 11552
rect 29092 11500 29144 11552
rect 30104 11543 30156 11552
rect 30104 11509 30113 11543
rect 30113 11509 30147 11543
rect 30147 11509 30156 11543
rect 30104 11500 30156 11509
rect 5915 11398 5967 11450
rect 5979 11398 6031 11450
rect 6043 11398 6095 11450
rect 6107 11398 6159 11450
rect 6171 11398 6223 11450
rect 15846 11398 15898 11450
rect 15910 11398 15962 11450
rect 15974 11398 16026 11450
rect 16038 11398 16090 11450
rect 16102 11398 16154 11450
rect 25776 11398 25828 11450
rect 25840 11398 25892 11450
rect 25904 11398 25956 11450
rect 25968 11398 26020 11450
rect 26032 11398 26084 11450
rect 10416 11296 10468 11348
rect 11888 11339 11940 11348
rect 11888 11305 11897 11339
rect 11897 11305 11931 11339
rect 11931 11305 11940 11339
rect 11888 11296 11940 11305
rect 9956 11160 10008 11212
rect 12532 11296 12584 11348
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 16212 11296 16264 11348
rect 16856 11339 16908 11348
rect 16856 11305 16865 11339
rect 16865 11305 16899 11339
rect 16899 11305 16908 11339
rect 16856 11296 16908 11305
rect 21364 11296 21416 11348
rect 22376 11296 22428 11348
rect 24032 11296 24084 11348
rect 25688 11296 25740 11348
rect 26792 11296 26844 11348
rect 19432 11228 19484 11280
rect 20628 11228 20680 11280
rect 21456 11228 21508 11280
rect 26700 11271 26752 11280
rect 26700 11237 26709 11271
rect 26709 11237 26743 11271
rect 26743 11237 26752 11271
rect 26700 11228 26752 11237
rect 28724 11296 28776 11348
rect 29000 11271 29052 11280
rect 9588 11135 9640 11144
rect 9588 11101 9597 11135
rect 9597 11101 9631 11135
rect 9631 11101 9640 11135
rect 9588 11092 9640 11101
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 11244 11160 11296 11212
rect 10692 11135 10744 11144
rect 2228 11067 2280 11076
rect 2228 11033 2237 11067
rect 2237 11033 2271 11067
rect 2271 11033 2280 11067
rect 2228 11024 2280 11033
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 12992 11160 13044 11212
rect 14188 11160 14240 11212
rect 10600 11024 10652 11076
rect 11796 11135 11848 11144
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 12072 11135 12124 11144
rect 11796 11092 11848 11101
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 15568 11092 15620 11144
rect 16488 11160 16540 11212
rect 18512 11160 18564 11212
rect 19156 11160 19208 11212
rect 20812 11160 20864 11212
rect 22192 11160 22244 11212
rect 23940 11160 23992 11212
rect 26516 11160 26568 11212
rect 16304 11092 16356 11144
rect 18788 11092 18840 11144
rect 19248 11135 19300 11144
rect 19248 11101 19257 11135
rect 19257 11101 19291 11135
rect 19291 11101 19300 11135
rect 19248 11092 19300 11101
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 14924 11024 14976 11076
rect 18236 11024 18288 11076
rect 18972 11024 19024 11076
rect 19708 11092 19760 11144
rect 20720 11135 20772 11144
rect 20720 11101 20729 11135
rect 20729 11101 20763 11135
rect 20763 11101 20772 11135
rect 20720 11092 20772 11101
rect 21272 11092 21324 11144
rect 21548 11135 21600 11144
rect 21548 11101 21557 11135
rect 21557 11101 21591 11135
rect 21591 11101 21600 11135
rect 21548 11092 21600 11101
rect 21916 11135 21968 11144
rect 21180 11024 21232 11076
rect 21916 11101 21925 11135
rect 21925 11101 21959 11135
rect 21959 11101 21968 11135
rect 21916 11092 21968 11101
rect 22376 11092 22428 11144
rect 22744 11092 22796 11144
rect 25136 11092 25188 11144
rect 25596 11092 25648 11144
rect 26608 11135 26660 11144
rect 26608 11101 26617 11135
rect 26617 11101 26651 11135
rect 26651 11101 26660 11135
rect 26608 11092 26660 11101
rect 27804 11135 27856 11144
rect 21824 11024 21876 11076
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 15568 10956 15620 11008
rect 19524 10956 19576 11008
rect 27804 11101 27813 11135
rect 27813 11101 27847 11135
rect 27847 11101 27856 11135
rect 27804 11092 27856 11101
rect 28264 11135 28316 11144
rect 28264 11101 28273 11135
rect 28273 11101 28307 11135
rect 28307 11101 28316 11135
rect 28264 11092 28316 11101
rect 28540 11203 28592 11212
rect 28540 11169 28549 11203
rect 28549 11169 28583 11203
rect 28583 11169 28592 11203
rect 29000 11237 29009 11271
rect 29009 11237 29043 11271
rect 29043 11237 29052 11271
rect 29000 11228 29052 11237
rect 28540 11160 28592 11169
rect 28632 11135 28684 11144
rect 28632 11101 28641 11135
rect 28641 11101 28675 11135
rect 28675 11101 28684 11135
rect 28632 11092 28684 11101
rect 30104 11160 30156 11212
rect 26884 11024 26936 11076
rect 28080 10956 28132 11008
rect 10880 10854 10932 10906
rect 10944 10854 10996 10906
rect 11008 10854 11060 10906
rect 11072 10854 11124 10906
rect 11136 10854 11188 10906
rect 20811 10854 20863 10906
rect 20875 10854 20927 10906
rect 20939 10854 20991 10906
rect 21003 10854 21055 10906
rect 21067 10854 21119 10906
rect 10140 10752 10192 10804
rect 11520 10752 11572 10804
rect 12072 10752 12124 10804
rect 12716 10795 12768 10804
rect 12716 10761 12725 10795
rect 12725 10761 12759 10795
rect 12759 10761 12768 10795
rect 12716 10752 12768 10761
rect 22008 10752 22060 10804
rect 26516 10752 26568 10804
rect 10508 10684 10560 10736
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 12440 10616 12492 10668
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 15568 10659 15620 10668
rect 15568 10625 15577 10659
rect 15577 10625 15611 10659
rect 15611 10625 15620 10659
rect 15568 10616 15620 10625
rect 19708 10684 19760 10736
rect 19984 10684 20036 10736
rect 12808 10591 12860 10600
rect 12808 10557 12817 10591
rect 12817 10557 12851 10591
rect 12851 10557 12860 10591
rect 12808 10548 12860 10557
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 15476 10548 15528 10600
rect 15844 10616 15896 10668
rect 16948 10616 17000 10668
rect 18512 10659 18564 10668
rect 18512 10625 18521 10659
rect 18521 10625 18555 10659
rect 18555 10625 18564 10659
rect 18512 10616 18564 10625
rect 19248 10616 19300 10668
rect 20628 10616 20680 10668
rect 25596 10659 25648 10668
rect 18604 10548 18656 10600
rect 19064 10548 19116 10600
rect 20444 10548 20496 10600
rect 21916 10548 21968 10600
rect 18972 10480 19024 10532
rect 24216 10548 24268 10600
rect 25596 10625 25605 10659
rect 25605 10625 25639 10659
rect 25639 10625 25648 10659
rect 25596 10616 25648 10625
rect 25688 10616 25740 10668
rect 26056 10548 26108 10600
rect 26516 10616 26568 10668
rect 27160 10659 27212 10668
rect 27160 10625 27169 10659
rect 27169 10625 27203 10659
rect 27203 10625 27212 10659
rect 27160 10616 27212 10625
rect 28080 10752 28132 10804
rect 29092 10684 29144 10736
rect 26792 10548 26844 10600
rect 27068 10591 27120 10600
rect 27068 10557 27077 10591
rect 27077 10557 27111 10591
rect 27111 10557 27120 10591
rect 27068 10548 27120 10557
rect 28540 10548 28592 10600
rect 28724 10591 28776 10600
rect 28724 10557 28733 10591
rect 28733 10557 28767 10591
rect 28767 10557 28776 10591
rect 28724 10548 28776 10557
rect 24584 10480 24636 10532
rect 15660 10412 15712 10464
rect 16212 10412 16264 10464
rect 5915 10310 5967 10362
rect 5979 10310 6031 10362
rect 6043 10310 6095 10362
rect 6107 10310 6159 10362
rect 6171 10310 6223 10362
rect 15846 10310 15898 10362
rect 15910 10310 15962 10362
rect 15974 10310 16026 10362
rect 16038 10310 16090 10362
rect 16102 10310 16154 10362
rect 25776 10310 25828 10362
rect 25840 10310 25892 10362
rect 25904 10310 25956 10362
rect 25968 10310 26020 10362
rect 26032 10310 26084 10362
rect 10692 10208 10744 10260
rect 12440 10251 12492 10260
rect 12440 10217 12449 10251
rect 12449 10217 12483 10251
rect 12483 10217 12492 10251
rect 12440 10208 12492 10217
rect 10692 10072 10744 10124
rect 12992 10208 13044 10260
rect 14280 10208 14332 10260
rect 14832 10208 14884 10260
rect 16580 10251 16632 10260
rect 12992 10115 13044 10124
rect 12992 10081 13001 10115
rect 13001 10081 13035 10115
rect 13035 10081 13044 10115
rect 14740 10115 14792 10124
rect 12992 10072 13044 10081
rect 14740 10081 14749 10115
rect 14749 10081 14783 10115
rect 14783 10081 14792 10115
rect 14740 10072 14792 10081
rect 10508 10004 10560 10056
rect 10876 10004 10928 10056
rect 12716 10004 12768 10056
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 16212 10072 16264 10124
rect 15752 10047 15804 10056
rect 15752 10013 15766 10047
rect 15766 10013 15800 10047
rect 15800 10013 15804 10047
rect 16580 10217 16589 10251
rect 16589 10217 16623 10251
rect 16623 10217 16632 10251
rect 16580 10208 16632 10217
rect 18420 10251 18472 10260
rect 18420 10217 18429 10251
rect 18429 10217 18463 10251
rect 18463 10217 18472 10251
rect 18420 10208 18472 10217
rect 19432 10208 19484 10260
rect 20628 10208 20680 10260
rect 28540 10251 28592 10260
rect 28540 10217 28549 10251
rect 28549 10217 28583 10251
rect 28583 10217 28592 10251
rect 28540 10208 28592 10217
rect 15752 10004 15804 10013
rect 16948 10004 17000 10056
rect 17132 10047 17184 10056
rect 17132 10013 17141 10047
rect 17141 10013 17175 10047
rect 17175 10013 17184 10047
rect 17132 10004 17184 10013
rect 10784 9936 10836 9988
rect 15200 9936 15252 9988
rect 14096 9868 14148 9920
rect 14924 9868 14976 9920
rect 15660 9979 15712 9988
rect 15660 9945 15669 9979
rect 15669 9945 15703 9979
rect 15703 9945 15712 9979
rect 18052 10072 18104 10124
rect 21180 10072 21232 10124
rect 22192 10140 22244 10192
rect 21824 10072 21876 10124
rect 26976 10072 27028 10124
rect 19064 10004 19116 10056
rect 19340 10004 19392 10056
rect 19524 10047 19576 10056
rect 19524 10013 19558 10047
rect 19558 10013 19576 10047
rect 19524 10004 19576 10013
rect 21272 10004 21324 10056
rect 21456 10004 21508 10056
rect 25228 10047 25280 10056
rect 15660 9936 15712 9945
rect 17960 9936 18012 9988
rect 18328 9979 18380 9988
rect 18328 9945 18337 9979
rect 18337 9945 18371 9979
rect 18371 9945 18380 9979
rect 18328 9936 18380 9945
rect 25228 10013 25237 10047
rect 25237 10013 25271 10047
rect 25271 10013 25280 10047
rect 25228 10004 25280 10013
rect 26884 10004 26936 10056
rect 28724 10004 28776 10056
rect 30104 10047 30156 10056
rect 30104 10013 30113 10047
rect 30113 10013 30147 10047
rect 30147 10013 30156 10047
rect 30104 10004 30156 10013
rect 27528 9936 27580 9988
rect 17776 9911 17828 9920
rect 17776 9877 17785 9911
rect 17785 9877 17819 9911
rect 17819 9877 17828 9911
rect 17776 9868 17828 9877
rect 19708 9868 19760 9920
rect 21272 9868 21324 9920
rect 22284 9868 22336 9920
rect 23940 9868 23992 9920
rect 29276 9868 29328 9920
rect 10880 9766 10932 9818
rect 10944 9766 10996 9818
rect 11008 9766 11060 9818
rect 11072 9766 11124 9818
rect 11136 9766 11188 9818
rect 20811 9766 20863 9818
rect 20875 9766 20927 9818
rect 20939 9766 20991 9818
rect 21003 9766 21055 9818
rect 21067 9766 21119 9818
rect 10600 9664 10652 9716
rect 12808 9664 12860 9716
rect 15200 9664 15252 9716
rect 18052 9707 18104 9716
rect 18052 9673 18061 9707
rect 18061 9673 18095 9707
rect 18095 9673 18104 9707
rect 18052 9664 18104 9673
rect 10692 9596 10744 9648
rect 10508 9528 10560 9580
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 14096 9528 14148 9580
rect 14648 9528 14700 9580
rect 15200 9528 15252 9580
rect 12716 9460 12768 9512
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 14740 9460 14792 9512
rect 15384 9571 15436 9580
rect 15384 9537 15393 9571
rect 15393 9537 15427 9571
rect 15427 9537 15436 9571
rect 17776 9596 17828 9648
rect 17960 9596 18012 9648
rect 15384 9528 15436 9537
rect 18236 9528 18288 9580
rect 18604 9571 18656 9580
rect 18604 9537 18614 9571
rect 18614 9537 18648 9571
rect 18648 9537 18656 9571
rect 18788 9571 18840 9580
rect 18604 9528 18656 9537
rect 18788 9537 18797 9571
rect 18797 9537 18831 9571
rect 18831 9537 18840 9571
rect 18788 9528 18840 9537
rect 15752 9460 15804 9512
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 19064 9528 19116 9580
rect 19340 9528 19392 9580
rect 21364 9528 21416 9580
rect 22376 9596 22428 9648
rect 26976 9596 27028 9648
rect 22100 9528 22152 9580
rect 22284 9571 22336 9580
rect 22284 9537 22318 9571
rect 22318 9537 22336 9571
rect 22284 9528 22336 9537
rect 23940 9571 23992 9580
rect 23940 9537 23949 9571
rect 23949 9537 23983 9571
rect 23983 9537 23992 9571
rect 23940 9528 23992 9537
rect 24032 9528 24084 9580
rect 26148 9528 26200 9580
rect 27620 9528 27672 9580
rect 29552 9528 29604 9580
rect 21272 9460 21324 9512
rect 28724 9503 28776 9512
rect 19156 9367 19208 9376
rect 19156 9333 19165 9367
rect 19165 9333 19199 9367
rect 19199 9333 19208 9367
rect 19156 9324 19208 9333
rect 20628 9324 20680 9376
rect 20812 9324 20864 9376
rect 20996 9324 21048 9376
rect 28724 9469 28733 9503
rect 28733 9469 28767 9503
rect 28767 9469 28776 9503
rect 28724 9460 28776 9469
rect 23204 9392 23256 9444
rect 28080 9392 28132 9444
rect 30012 9392 30064 9444
rect 24216 9324 24268 9376
rect 5915 9222 5967 9274
rect 5979 9222 6031 9274
rect 6043 9222 6095 9274
rect 6107 9222 6159 9274
rect 6171 9222 6223 9274
rect 15846 9222 15898 9274
rect 15910 9222 15962 9274
rect 15974 9222 16026 9274
rect 16038 9222 16090 9274
rect 16102 9222 16154 9274
rect 25776 9222 25828 9274
rect 25840 9222 25892 9274
rect 25904 9222 25956 9274
rect 25968 9222 26020 9274
rect 26032 9222 26084 9274
rect 10784 9120 10836 9172
rect 12164 9120 12216 9172
rect 14004 9120 14056 9172
rect 15384 9120 15436 9172
rect 18328 9120 18380 9172
rect 19064 9120 19116 9172
rect 22192 9120 22244 9172
rect 24032 9120 24084 9172
rect 28172 9120 28224 9172
rect 21364 9095 21416 9104
rect 21364 9061 21373 9095
rect 21373 9061 21407 9095
rect 21407 9061 21416 9095
rect 21364 9052 21416 9061
rect 13268 8984 13320 9036
rect 14740 8984 14792 9036
rect 2228 8916 2280 8968
rect 11704 8916 11756 8968
rect 14648 8916 14700 8968
rect 12716 8848 12768 8900
rect 15476 8984 15528 9036
rect 15568 8959 15620 8968
rect 15568 8925 15577 8959
rect 15577 8925 15611 8959
rect 15611 8925 15620 8959
rect 15568 8916 15620 8925
rect 16948 8984 17000 9036
rect 17500 8984 17552 9036
rect 18604 8984 18656 9036
rect 18328 8916 18380 8968
rect 19248 8916 19300 8968
rect 20536 8916 20588 8968
rect 20904 8959 20956 8968
rect 20904 8925 20911 8959
rect 20911 8925 20956 8959
rect 20904 8916 20956 8925
rect 20996 8959 21048 8968
rect 20996 8925 21005 8959
rect 21005 8925 21039 8959
rect 21039 8925 21048 8959
rect 20996 8916 21048 8925
rect 21824 8916 21876 8968
rect 23112 9052 23164 9104
rect 22192 8984 22244 9036
rect 24952 8984 25004 9036
rect 27344 9027 27396 9036
rect 27344 8993 27353 9027
rect 27353 8993 27387 9027
rect 27387 8993 27396 9027
rect 27344 8984 27396 8993
rect 27988 8984 28040 9036
rect 28632 8984 28684 9036
rect 19892 8848 19944 8900
rect 20628 8848 20680 8900
rect 23204 8916 23256 8968
rect 23480 8959 23532 8968
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 10784 8780 10836 8832
rect 11428 8823 11480 8832
rect 11428 8789 11437 8823
rect 11437 8789 11471 8823
rect 11471 8789 11480 8823
rect 14556 8823 14608 8832
rect 11428 8780 11480 8789
rect 14556 8789 14565 8823
rect 14565 8789 14599 8823
rect 14599 8789 14608 8823
rect 14556 8780 14608 8789
rect 15476 8780 15528 8832
rect 15568 8780 15620 8832
rect 20720 8780 20772 8832
rect 22560 8848 22612 8900
rect 22744 8848 22796 8900
rect 23480 8925 23489 8959
rect 23489 8925 23523 8959
rect 23523 8925 23532 8959
rect 23480 8916 23532 8925
rect 25320 8916 25372 8968
rect 26148 8916 26200 8968
rect 26976 8916 27028 8968
rect 28816 8959 28868 8968
rect 28816 8925 28825 8959
rect 28825 8925 28859 8959
rect 28859 8925 28868 8959
rect 28816 8916 28868 8925
rect 30104 8959 30156 8968
rect 30104 8925 30113 8959
rect 30113 8925 30147 8959
rect 30147 8925 30156 8959
rect 30104 8916 30156 8925
rect 24124 8848 24176 8900
rect 25136 8848 25188 8900
rect 22376 8780 22428 8832
rect 24216 8780 24268 8832
rect 28816 8780 28868 8832
rect 10880 8678 10932 8730
rect 10944 8678 10996 8730
rect 11008 8678 11060 8730
rect 11072 8678 11124 8730
rect 11136 8678 11188 8730
rect 20811 8678 20863 8730
rect 20875 8678 20927 8730
rect 20939 8678 20991 8730
rect 21003 8678 21055 8730
rect 21067 8678 21119 8730
rect 10784 8619 10836 8628
rect 10784 8585 10793 8619
rect 10793 8585 10827 8619
rect 10827 8585 10836 8619
rect 10784 8576 10836 8585
rect 14556 8576 14608 8628
rect 16396 8576 16448 8628
rect 18788 8576 18840 8628
rect 20076 8576 20128 8628
rect 24124 8576 24176 8628
rect 29920 8576 29972 8628
rect 11704 8551 11756 8560
rect 11704 8517 11713 8551
rect 11713 8517 11747 8551
rect 11747 8517 11756 8551
rect 11704 8508 11756 8517
rect 11428 8440 11480 8492
rect 11980 8440 12032 8492
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 19156 8508 19208 8560
rect 19248 8508 19300 8560
rect 22100 8551 22152 8560
rect 22100 8517 22109 8551
rect 22109 8517 22143 8551
rect 22143 8517 22152 8551
rect 22100 8508 22152 8517
rect 22468 8508 22520 8560
rect 24216 8508 24268 8560
rect 15752 8483 15804 8492
rect 14648 8440 14700 8449
rect 15752 8449 15761 8483
rect 15761 8449 15795 8483
rect 15795 8449 15804 8483
rect 15752 8440 15804 8449
rect 16764 8440 16816 8492
rect 21916 8483 21968 8492
rect 21916 8449 21925 8483
rect 21925 8449 21959 8483
rect 21959 8449 21968 8483
rect 21916 8440 21968 8449
rect 23020 8483 23072 8492
rect 15476 8372 15528 8424
rect 15568 8372 15620 8424
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 20628 8372 20680 8424
rect 22468 8372 22520 8424
rect 12440 8304 12492 8356
rect 16672 8304 16724 8356
rect 23020 8449 23029 8483
rect 23029 8449 23063 8483
rect 23063 8449 23072 8483
rect 23020 8440 23072 8449
rect 23112 8483 23164 8492
rect 23112 8449 23121 8483
rect 23121 8449 23155 8483
rect 23155 8449 23164 8483
rect 23112 8440 23164 8449
rect 23480 8372 23532 8424
rect 23756 8372 23808 8424
rect 23940 8440 23992 8492
rect 27160 8508 27212 8560
rect 26148 8440 26200 8492
rect 29000 8483 29052 8492
rect 29000 8449 29034 8483
rect 29034 8449 29052 8483
rect 29000 8440 29052 8449
rect 26240 8372 26292 8424
rect 27344 8372 27396 8424
rect 27712 8372 27764 8424
rect 28724 8415 28776 8424
rect 28724 8381 28733 8415
rect 28733 8381 28767 8415
rect 28767 8381 28776 8415
rect 28724 8372 28776 8381
rect 17040 8279 17092 8288
rect 17040 8245 17049 8279
rect 17049 8245 17083 8279
rect 17083 8245 17092 8279
rect 17040 8236 17092 8245
rect 17960 8236 18012 8288
rect 18236 8236 18288 8288
rect 25320 8304 25372 8356
rect 24952 8236 25004 8288
rect 5915 8134 5967 8186
rect 5979 8134 6031 8186
rect 6043 8134 6095 8186
rect 6107 8134 6159 8186
rect 6171 8134 6223 8186
rect 15846 8134 15898 8186
rect 15910 8134 15962 8186
rect 15974 8134 16026 8186
rect 16038 8134 16090 8186
rect 16102 8134 16154 8186
rect 25776 8134 25828 8186
rect 25840 8134 25892 8186
rect 25904 8134 25956 8186
rect 25968 8134 26020 8186
rect 26032 8134 26084 8186
rect 12532 8032 12584 8084
rect 15752 8032 15804 8084
rect 12900 7896 12952 7948
rect 17960 8032 18012 8084
rect 18052 8032 18104 8084
rect 18604 8075 18656 8084
rect 18604 8041 18613 8075
rect 18613 8041 18647 8075
rect 18647 8041 18656 8075
rect 18604 8032 18656 8041
rect 19432 8032 19484 8084
rect 19892 8032 19944 8084
rect 20168 8032 20220 8084
rect 12532 7828 12584 7880
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 17040 7828 17092 7880
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 17316 7828 17368 7837
rect 17500 7871 17552 7880
rect 17500 7837 17507 7871
rect 17507 7837 17552 7871
rect 17500 7828 17552 7837
rect 19524 7964 19576 8016
rect 18420 7828 18472 7880
rect 19892 7896 19944 7948
rect 21272 8032 21324 8084
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 20076 7828 20128 7880
rect 20720 7828 20772 7880
rect 22284 7964 22336 8016
rect 23296 8032 23348 8084
rect 24308 8032 24360 8084
rect 27160 8032 27212 8084
rect 27528 8032 27580 8084
rect 23940 7964 23992 8016
rect 22836 7896 22888 7948
rect 27620 7964 27672 8016
rect 28724 7964 28776 8016
rect 23204 7828 23256 7880
rect 23572 7828 23624 7880
rect 24308 7828 24360 7880
rect 25136 7828 25188 7880
rect 27620 7871 27672 7880
rect 27620 7837 27629 7871
rect 27629 7837 27663 7871
rect 27663 7837 27672 7871
rect 27620 7828 27672 7837
rect 28908 7896 28960 7948
rect 12808 7760 12860 7812
rect 13636 7760 13688 7812
rect 12348 7692 12400 7744
rect 13360 7692 13412 7744
rect 21916 7760 21968 7812
rect 22376 7803 22428 7812
rect 17684 7692 17736 7744
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 18052 7692 18104 7744
rect 19432 7692 19484 7744
rect 22376 7769 22385 7803
rect 22385 7769 22419 7803
rect 22419 7769 22428 7803
rect 22376 7760 22428 7769
rect 22468 7803 22520 7812
rect 22468 7769 22477 7803
rect 22477 7769 22511 7803
rect 22511 7769 22520 7803
rect 22468 7760 22520 7769
rect 23480 7760 23532 7812
rect 27988 7871 28040 7880
rect 27988 7837 27997 7871
rect 27997 7837 28031 7871
rect 28031 7837 28040 7871
rect 27988 7828 28040 7837
rect 28540 7828 28592 7880
rect 30104 7871 30156 7880
rect 30104 7837 30113 7871
rect 30113 7837 30147 7871
rect 30147 7837 30156 7871
rect 30104 7828 30156 7837
rect 28080 7760 28132 7812
rect 22284 7692 22336 7744
rect 27620 7692 27672 7744
rect 10880 7590 10932 7642
rect 10944 7590 10996 7642
rect 11008 7590 11060 7642
rect 11072 7590 11124 7642
rect 11136 7590 11188 7642
rect 20811 7590 20863 7642
rect 20875 7590 20927 7642
rect 20939 7590 20991 7642
rect 21003 7590 21055 7642
rect 21067 7590 21119 7642
rect 13360 7488 13412 7540
rect 14280 7488 14332 7540
rect 19524 7488 19576 7540
rect 23020 7488 23072 7540
rect 24308 7488 24360 7540
rect 27896 7488 27948 7540
rect 29552 7531 29604 7540
rect 29552 7497 29561 7531
rect 29561 7497 29595 7531
rect 29595 7497 29604 7531
rect 29552 7488 29604 7497
rect 14096 7420 14148 7472
rect 17960 7420 18012 7472
rect 20168 7420 20220 7472
rect 21548 7420 21600 7472
rect 1860 7352 1912 7404
rect 12348 7395 12400 7404
rect 12348 7361 12357 7395
rect 12357 7361 12391 7395
rect 12391 7361 12400 7395
rect 12348 7352 12400 7361
rect 12440 7352 12492 7404
rect 13268 7395 13320 7404
rect 13268 7361 13277 7395
rect 13277 7361 13311 7395
rect 13311 7361 13320 7395
rect 14832 7395 14884 7404
rect 13268 7352 13320 7361
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 14832 7352 14884 7361
rect 16672 7352 16724 7404
rect 18604 7352 18656 7404
rect 20444 7352 20496 7404
rect 20720 7352 20772 7404
rect 22928 7420 22980 7472
rect 23480 7420 23532 7472
rect 24400 7420 24452 7472
rect 29092 7420 29144 7472
rect 22100 7352 22152 7404
rect 23388 7352 23440 7404
rect 23756 7352 23808 7404
rect 27252 7395 27304 7404
rect 27252 7361 27286 7395
rect 27286 7361 27304 7395
rect 27252 7352 27304 7361
rect 28356 7352 28408 7404
rect 28724 7352 28776 7404
rect 29276 7352 29328 7404
rect 30012 7352 30064 7404
rect 13360 7327 13412 7336
rect 13360 7293 13394 7327
rect 13394 7293 13412 7327
rect 13360 7284 13412 7293
rect 13544 7327 13596 7336
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 26240 7284 26292 7336
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 15568 7148 15620 7200
rect 16580 7148 16632 7200
rect 17684 7148 17736 7200
rect 20076 7148 20128 7200
rect 20812 7148 20864 7200
rect 28080 7284 28132 7336
rect 28632 7284 28684 7336
rect 27988 7216 28040 7268
rect 28724 7216 28776 7268
rect 27712 7148 27764 7200
rect 5915 7046 5967 7098
rect 5979 7046 6031 7098
rect 6043 7046 6095 7098
rect 6107 7046 6159 7098
rect 6171 7046 6223 7098
rect 15846 7046 15898 7098
rect 15910 7046 15962 7098
rect 15974 7046 16026 7098
rect 16038 7046 16090 7098
rect 16102 7046 16154 7098
rect 25776 7046 25828 7098
rect 25840 7046 25892 7098
rect 25904 7046 25956 7098
rect 25968 7046 26020 7098
rect 26032 7046 26084 7098
rect 12164 6944 12216 6996
rect 15476 6987 15528 6996
rect 15476 6953 15485 6987
rect 15485 6953 15519 6987
rect 15519 6953 15528 6987
rect 15476 6944 15528 6953
rect 10600 6851 10652 6860
rect 10600 6817 10609 6851
rect 10609 6817 10643 6851
rect 10643 6817 10652 6851
rect 10600 6808 10652 6817
rect 12348 6808 12400 6860
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 11704 6740 11756 6792
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 14740 6876 14792 6928
rect 16856 6876 16908 6928
rect 14832 6808 14884 6860
rect 13544 6740 13596 6792
rect 16580 6808 16632 6860
rect 20260 6944 20312 6996
rect 20444 6987 20496 6996
rect 20444 6953 20453 6987
rect 20453 6953 20487 6987
rect 20487 6953 20496 6987
rect 20444 6944 20496 6953
rect 22376 6944 22428 6996
rect 23388 6987 23440 6996
rect 23388 6953 23397 6987
rect 23397 6953 23431 6987
rect 23431 6953 23440 6987
rect 23388 6944 23440 6953
rect 27252 6944 27304 6996
rect 18420 6876 18472 6928
rect 18052 6808 18104 6860
rect 20720 6876 20772 6928
rect 15752 6672 15804 6724
rect 16488 6672 16540 6724
rect 17500 6740 17552 6792
rect 17960 6783 18012 6792
rect 17960 6749 17969 6783
rect 17969 6749 18003 6783
rect 18003 6749 18012 6783
rect 17960 6740 18012 6749
rect 18880 6740 18932 6792
rect 19340 6672 19392 6724
rect 12440 6647 12492 6656
rect 12440 6613 12449 6647
rect 12449 6613 12483 6647
rect 12483 6613 12492 6647
rect 15844 6647 15896 6656
rect 12440 6604 12492 6613
rect 15844 6613 15853 6647
rect 15853 6613 15887 6647
rect 15887 6613 15896 6647
rect 15844 6604 15896 6613
rect 16672 6647 16724 6656
rect 16672 6613 16681 6647
rect 16681 6613 16715 6647
rect 16715 6613 16724 6647
rect 16672 6604 16724 6613
rect 18236 6604 18288 6656
rect 18512 6604 18564 6656
rect 20444 6740 20496 6792
rect 20812 6808 20864 6860
rect 25320 6808 25372 6860
rect 26148 6808 26200 6860
rect 27896 6944 27948 6996
rect 20720 6740 20772 6792
rect 22100 6740 22152 6792
rect 22192 6740 22244 6792
rect 22836 6783 22888 6792
rect 22836 6749 22846 6783
rect 22846 6749 22880 6783
rect 22880 6749 22888 6783
rect 22836 6740 22888 6749
rect 23020 6783 23072 6792
rect 23020 6749 23029 6783
rect 23029 6749 23063 6783
rect 23063 6749 23072 6783
rect 23020 6740 23072 6749
rect 23204 6783 23256 6792
rect 23204 6749 23218 6783
rect 23218 6749 23252 6783
rect 23252 6749 23256 6783
rect 23204 6740 23256 6749
rect 24952 6740 25004 6792
rect 25412 6783 25464 6792
rect 20076 6715 20128 6724
rect 20076 6681 20085 6715
rect 20085 6681 20119 6715
rect 20119 6681 20128 6715
rect 20076 6672 20128 6681
rect 20168 6715 20220 6724
rect 20168 6681 20177 6715
rect 20177 6681 20211 6715
rect 20211 6681 20220 6715
rect 20168 6672 20220 6681
rect 22284 6672 22336 6724
rect 23112 6715 23164 6724
rect 23112 6681 23121 6715
rect 23121 6681 23155 6715
rect 23155 6681 23164 6715
rect 23112 6672 23164 6681
rect 25412 6749 25421 6783
rect 25421 6749 25455 6783
rect 25455 6749 25464 6783
rect 25412 6740 25464 6749
rect 26332 6740 26384 6792
rect 26700 6783 26752 6792
rect 26700 6749 26709 6783
rect 26709 6749 26743 6783
rect 26743 6749 26752 6783
rect 26700 6740 26752 6749
rect 27712 6740 27764 6792
rect 30104 6783 30156 6792
rect 27896 6715 27948 6724
rect 27896 6681 27930 6715
rect 27930 6681 27948 6715
rect 27896 6672 27948 6681
rect 21916 6604 21968 6656
rect 22192 6604 22244 6656
rect 22744 6604 22796 6656
rect 22928 6604 22980 6656
rect 27344 6604 27396 6656
rect 27804 6604 27856 6656
rect 30104 6749 30113 6783
rect 30113 6749 30147 6783
rect 30147 6749 30156 6783
rect 30104 6740 30156 6749
rect 10880 6502 10932 6554
rect 10944 6502 10996 6554
rect 11008 6502 11060 6554
rect 11072 6502 11124 6554
rect 11136 6502 11188 6554
rect 20811 6502 20863 6554
rect 20875 6502 20927 6554
rect 20939 6502 20991 6554
rect 21003 6502 21055 6554
rect 21067 6502 21119 6554
rect 11980 6443 12032 6452
rect 11980 6409 11989 6443
rect 11989 6409 12023 6443
rect 12023 6409 12032 6443
rect 11980 6400 12032 6409
rect 12440 6443 12492 6452
rect 12440 6409 12449 6443
rect 12449 6409 12483 6443
rect 12483 6409 12492 6443
rect 12440 6400 12492 6409
rect 12900 6400 12952 6452
rect 13820 6400 13872 6452
rect 15844 6400 15896 6452
rect 19156 6400 19208 6452
rect 21640 6400 21692 6452
rect 25688 6443 25740 6452
rect 25688 6409 25697 6443
rect 25697 6409 25731 6443
rect 25731 6409 25740 6443
rect 25688 6400 25740 6409
rect 27896 6443 27948 6452
rect 27896 6409 27905 6443
rect 27905 6409 27939 6443
rect 27939 6409 27948 6443
rect 27896 6400 27948 6409
rect 29000 6400 29052 6452
rect 16856 6332 16908 6384
rect 17684 6375 17736 6384
rect 17684 6341 17693 6375
rect 17693 6341 17727 6375
rect 17727 6341 17736 6375
rect 17684 6332 17736 6341
rect 12440 6264 12492 6316
rect 14188 6264 14240 6316
rect 17316 6264 17368 6316
rect 17500 6307 17552 6316
rect 17500 6273 17510 6307
rect 17510 6273 17544 6307
rect 17544 6273 17552 6307
rect 17500 6264 17552 6273
rect 18420 6332 18472 6384
rect 13544 6196 13596 6248
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 14280 6239 14332 6248
rect 14280 6205 14289 6239
rect 14289 6205 14323 6239
rect 14323 6205 14332 6239
rect 14280 6196 14332 6205
rect 15016 6239 15068 6248
rect 15016 6205 15025 6239
rect 15025 6205 15059 6239
rect 15059 6205 15068 6239
rect 15016 6196 15068 6205
rect 15108 6239 15160 6248
rect 15108 6205 15142 6239
rect 15142 6205 15160 6239
rect 15108 6196 15160 6205
rect 15476 6196 15528 6248
rect 11244 6128 11296 6180
rect 11796 6128 11848 6180
rect 12808 6128 12860 6180
rect 14832 6128 14884 6180
rect 18052 6264 18104 6316
rect 18696 6307 18748 6316
rect 18696 6273 18705 6307
rect 18705 6273 18739 6307
rect 18739 6273 18748 6307
rect 18696 6264 18748 6273
rect 19708 6332 19760 6384
rect 25412 6332 25464 6384
rect 18972 6307 19024 6316
rect 18972 6273 18981 6307
rect 18981 6273 19015 6307
rect 19015 6273 19024 6307
rect 18972 6264 19024 6273
rect 19156 6264 19208 6316
rect 20444 6307 20496 6316
rect 20444 6273 20453 6307
rect 20453 6273 20487 6307
rect 20487 6273 20496 6307
rect 20444 6264 20496 6273
rect 21824 6307 21876 6316
rect 21824 6273 21833 6307
rect 21833 6273 21867 6307
rect 21867 6273 21876 6307
rect 21824 6264 21876 6273
rect 22100 6264 22152 6316
rect 22744 6307 22796 6316
rect 22744 6273 22778 6307
rect 22778 6273 22796 6307
rect 22744 6264 22796 6273
rect 23940 6264 23992 6316
rect 25596 6264 25648 6316
rect 27620 6264 27672 6316
rect 27804 6264 27856 6316
rect 28356 6307 28408 6316
rect 28356 6273 28365 6307
rect 28365 6273 28399 6307
rect 28399 6273 28408 6307
rect 28356 6264 28408 6273
rect 28816 6264 28868 6316
rect 29920 6264 29972 6316
rect 30104 6307 30156 6316
rect 30104 6273 30113 6307
rect 30113 6273 30147 6307
rect 30147 6273 30156 6307
rect 30104 6264 30156 6273
rect 19340 6196 19392 6248
rect 19984 6196 20036 6248
rect 21180 6196 21232 6248
rect 26700 6196 26752 6248
rect 27436 6239 27488 6248
rect 27436 6205 27445 6239
rect 27445 6205 27479 6239
rect 27479 6205 27488 6239
rect 27436 6196 27488 6205
rect 28632 6239 28684 6248
rect 21364 6128 21416 6180
rect 22284 6128 22336 6180
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 19432 6103 19484 6112
rect 19432 6069 19441 6103
rect 19441 6069 19475 6103
rect 19475 6069 19484 6103
rect 19432 6060 19484 6069
rect 26148 6128 26200 6180
rect 28632 6205 28641 6239
rect 28641 6205 28675 6239
rect 28675 6205 28684 6239
rect 28632 6196 28684 6205
rect 28724 6239 28776 6248
rect 28724 6205 28733 6239
rect 28733 6205 28767 6239
rect 28767 6205 28776 6239
rect 28724 6196 28776 6205
rect 27620 6128 27672 6180
rect 23572 6060 23624 6112
rect 28356 6060 28408 6112
rect 5915 5958 5967 6010
rect 5979 5958 6031 6010
rect 6043 5958 6095 6010
rect 6107 5958 6159 6010
rect 6171 5958 6223 6010
rect 15846 5958 15898 6010
rect 15910 5958 15962 6010
rect 15974 5958 16026 6010
rect 16038 5958 16090 6010
rect 16102 5958 16154 6010
rect 25776 5958 25828 6010
rect 25840 5958 25892 6010
rect 25904 5958 25956 6010
rect 25968 5958 26020 6010
rect 26032 5958 26084 6010
rect 12440 5899 12492 5908
rect 12440 5865 12449 5899
rect 12449 5865 12483 5899
rect 12483 5865 12492 5899
rect 12440 5856 12492 5865
rect 14556 5856 14608 5908
rect 15108 5856 15160 5908
rect 15752 5856 15804 5908
rect 18236 5856 18288 5908
rect 21180 5856 21232 5908
rect 10600 5788 10652 5840
rect 10784 5763 10836 5772
rect 10784 5729 10793 5763
rect 10793 5729 10827 5763
rect 10827 5729 10836 5763
rect 10784 5720 10836 5729
rect 11244 5763 11296 5772
rect 11244 5729 11253 5763
rect 11253 5729 11287 5763
rect 11287 5729 11296 5763
rect 11244 5720 11296 5729
rect 19524 5788 19576 5840
rect 20076 5788 20128 5840
rect 11520 5763 11572 5772
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 11612 5763 11664 5772
rect 11612 5729 11646 5763
rect 11646 5729 11664 5763
rect 11612 5720 11664 5729
rect 12348 5720 12400 5772
rect 13820 5720 13872 5772
rect 14740 5763 14792 5772
rect 14740 5729 14749 5763
rect 14749 5729 14783 5763
rect 14783 5729 14792 5763
rect 14740 5720 14792 5729
rect 15108 5763 15160 5772
rect 15108 5729 15142 5763
rect 15142 5729 15160 5763
rect 15108 5720 15160 5729
rect 15476 5720 15528 5772
rect 21180 5763 21232 5772
rect 21180 5729 21189 5763
rect 21189 5729 21223 5763
rect 21223 5729 21232 5763
rect 21180 5720 21232 5729
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 13636 5652 13688 5704
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 15016 5695 15068 5704
rect 15016 5661 15025 5695
rect 15025 5661 15059 5695
rect 15059 5661 15068 5695
rect 16396 5695 16448 5704
rect 15016 5652 15068 5661
rect 16396 5661 16405 5695
rect 16405 5661 16439 5695
rect 16439 5661 16448 5695
rect 16396 5652 16448 5661
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 19800 5652 19852 5704
rect 20984 5695 21036 5704
rect 11888 5516 11940 5568
rect 12992 5516 13044 5568
rect 15016 5516 15068 5568
rect 15292 5516 15344 5568
rect 16488 5559 16540 5568
rect 16488 5525 16497 5559
rect 16497 5525 16531 5559
rect 16531 5525 16540 5559
rect 16488 5516 16540 5525
rect 20984 5661 20993 5695
rect 20993 5661 21027 5695
rect 21027 5661 21036 5695
rect 20984 5652 21036 5661
rect 21824 5788 21876 5840
rect 22744 5856 22796 5908
rect 26608 5856 26660 5908
rect 26332 5788 26384 5840
rect 23940 5720 23992 5772
rect 21364 5695 21416 5704
rect 21364 5661 21373 5695
rect 21373 5661 21407 5695
rect 21407 5661 21416 5695
rect 21364 5652 21416 5661
rect 21916 5652 21968 5704
rect 22284 5695 22336 5704
rect 21272 5584 21324 5636
rect 22284 5661 22293 5695
rect 22293 5661 22327 5695
rect 22327 5661 22336 5695
rect 22284 5652 22336 5661
rect 22560 5652 22612 5704
rect 23204 5652 23256 5704
rect 27712 5652 27764 5704
rect 22928 5584 22980 5636
rect 21180 5516 21232 5568
rect 21548 5559 21600 5568
rect 21548 5525 21557 5559
rect 21557 5525 21591 5559
rect 21591 5525 21600 5559
rect 21548 5516 21600 5525
rect 22100 5516 22152 5568
rect 26148 5584 26200 5636
rect 27344 5584 27396 5636
rect 29920 5627 29972 5636
rect 29920 5593 29929 5627
rect 29929 5593 29963 5627
rect 29963 5593 29972 5627
rect 29920 5584 29972 5593
rect 29184 5516 29236 5568
rect 30012 5559 30064 5568
rect 30012 5525 30021 5559
rect 30021 5525 30055 5559
rect 30055 5525 30064 5559
rect 30012 5516 30064 5525
rect 10880 5414 10932 5466
rect 10944 5414 10996 5466
rect 11008 5414 11060 5466
rect 11072 5414 11124 5466
rect 11136 5414 11188 5466
rect 20811 5414 20863 5466
rect 20875 5414 20927 5466
rect 20939 5414 20991 5466
rect 21003 5414 21055 5466
rect 21067 5414 21119 5466
rect 11888 5355 11940 5364
rect 11888 5321 11897 5355
rect 11897 5321 11931 5355
rect 11931 5321 11940 5355
rect 11888 5312 11940 5321
rect 14280 5312 14332 5364
rect 17684 5312 17736 5364
rect 19156 5312 19208 5364
rect 25596 5312 25648 5364
rect 1492 5176 1544 5228
rect 12992 5176 13044 5228
rect 12440 5040 12492 5092
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 14372 5176 14424 5228
rect 13820 5108 13872 5160
rect 15292 5176 15344 5228
rect 18236 5244 18288 5296
rect 18604 5244 18656 5296
rect 19432 5244 19484 5296
rect 19800 5244 19852 5296
rect 15476 5176 15528 5228
rect 17040 5219 17092 5228
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 13268 4972 13320 5024
rect 15384 5040 15436 5092
rect 14372 4972 14424 5024
rect 16396 4972 16448 5024
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 18052 5176 18104 5228
rect 21180 5176 21232 5228
rect 21732 5176 21784 5228
rect 22008 5219 22060 5228
rect 22008 5185 22017 5219
rect 22017 5185 22051 5219
rect 22051 5185 22060 5219
rect 22008 5176 22060 5185
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 23848 5244 23900 5296
rect 22100 5176 22152 5185
rect 23204 5176 23256 5228
rect 24952 5176 25004 5228
rect 30012 5244 30064 5296
rect 25688 5176 25740 5228
rect 29920 5219 29972 5228
rect 29920 5185 29929 5219
rect 29929 5185 29963 5219
rect 29963 5185 29972 5219
rect 29920 5176 29972 5185
rect 22560 5108 22612 5160
rect 25320 5151 25372 5160
rect 25320 5117 25329 5151
rect 25329 5117 25363 5151
rect 25363 5117 25372 5151
rect 25320 5108 25372 5117
rect 25780 5108 25832 5160
rect 26056 5108 26108 5160
rect 29000 5040 29052 5092
rect 18144 4972 18196 5024
rect 22560 5015 22612 5024
rect 22560 4981 22569 5015
rect 22569 4981 22603 5015
rect 22603 4981 22612 5015
rect 22560 4972 22612 4981
rect 30012 5015 30064 5024
rect 30012 4981 30021 5015
rect 30021 4981 30055 5015
rect 30055 4981 30064 5015
rect 30012 4972 30064 4981
rect 5915 4870 5967 4922
rect 5979 4870 6031 4922
rect 6043 4870 6095 4922
rect 6107 4870 6159 4922
rect 6171 4870 6223 4922
rect 15846 4870 15898 4922
rect 15910 4870 15962 4922
rect 15974 4870 16026 4922
rect 16038 4870 16090 4922
rect 16102 4870 16154 4922
rect 25776 4870 25828 4922
rect 25840 4870 25892 4922
rect 25904 4870 25956 4922
rect 25968 4870 26020 4922
rect 26032 4870 26084 4922
rect 12716 4811 12768 4820
rect 12716 4777 12725 4811
rect 12725 4777 12759 4811
rect 12759 4777 12768 4811
rect 12716 4768 12768 4777
rect 11520 4700 11572 4752
rect 14556 4700 14608 4752
rect 13544 4632 13596 4684
rect 14740 4632 14792 4684
rect 17040 4768 17092 4820
rect 21364 4811 21416 4820
rect 21364 4777 21373 4811
rect 21373 4777 21407 4811
rect 21407 4777 21416 4811
rect 21364 4768 21416 4777
rect 22744 4768 22796 4820
rect 23204 4811 23256 4820
rect 23204 4777 23213 4811
rect 23213 4777 23247 4811
rect 23247 4777 23256 4811
rect 23204 4768 23256 4777
rect 26148 4811 26200 4820
rect 26148 4777 26157 4811
rect 26157 4777 26191 4811
rect 26191 4777 26200 4811
rect 26148 4768 26200 4777
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 15476 4564 15528 4616
rect 16672 4564 16724 4616
rect 20720 4564 20772 4616
rect 22560 4564 22612 4616
rect 24952 4564 25004 4616
rect 30012 4700 30064 4752
rect 25780 4675 25832 4684
rect 25780 4641 25789 4675
rect 25789 4641 25823 4675
rect 25823 4641 25832 4675
rect 25780 4632 25832 4641
rect 13084 4471 13136 4480
rect 13084 4437 13093 4471
rect 13093 4437 13127 4471
rect 13127 4437 13136 4471
rect 13084 4428 13136 4437
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 21548 4496 21600 4548
rect 25320 4496 25372 4548
rect 26608 4564 26660 4616
rect 29920 4539 29972 4548
rect 29920 4505 29929 4539
rect 29929 4505 29963 4539
rect 29963 4505 29972 4539
rect 29920 4496 29972 4505
rect 13176 4428 13228 4437
rect 15384 4428 15436 4480
rect 16396 4428 16448 4480
rect 23112 4428 23164 4480
rect 10880 4326 10932 4378
rect 10944 4326 10996 4378
rect 11008 4326 11060 4378
rect 11072 4326 11124 4378
rect 11136 4326 11188 4378
rect 20811 4326 20863 4378
rect 20875 4326 20927 4378
rect 20939 4326 20991 4378
rect 21003 4326 21055 4378
rect 21067 4326 21119 4378
rect 10508 4088 10560 4140
rect 13268 4088 13320 4140
rect 13820 4088 13872 4140
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 15384 4131 15436 4140
rect 12256 3952 12308 4004
rect 14188 4063 14240 4072
rect 14188 4029 14197 4063
rect 14197 4029 14231 4063
rect 14231 4029 14240 4063
rect 14188 4020 14240 4029
rect 14740 4063 14792 4072
rect 14740 4029 14749 4063
rect 14749 4029 14783 4063
rect 14783 4029 14792 4063
rect 15384 4097 15393 4131
rect 15393 4097 15427 4131
rect 15427 4097 15436 4131
rect 15384 4088 15436 4097
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 18512 4131 18564 4140
rect 18512 4097 18546 4131
rect 18546 4097 18564 4131
rect 18512 4088 18564 4097
rect 30012 4088 30064 4140
rect 14740 4020 14792 4029
rect 16580 4020 16632 4072
rect 17132 4063 17184 4072
rect 11152 3884 11204 3936
rect 11612 3884 11664 3936
rect 15016 3952 15068 4004
rect 15384 3952 15436 4004
rect 16764 3952 16816 4004
rect 17132 4029 17141 4063
rect 17141 4029 17175 4063
rect 17175 4029 17184 4063
rect 17132 4020 17184 4029
rect 29184 3952 29236 4004
rect 14280 3884 14332 3936
rect 18880 3884 18932 3936
rect 5915 3782 5967 3834
rect 5979 3782 6031 3834
rect 6043 3782 6095 3834
rect 6107 3782 6159 3834
rect 6171 3782 6223 3834
rect 15846 3782 15898 3834
rect 15910 3782 15962 3834
rect 15974 3782 16026 3834
rect 16038 3782 16090 3834
rect 16102 3782 16154 3834
rect 25776 3782 25828 3834
rect 25840 3782 25892 3834
rect 25904 3782 25956 3834
rect 25968 3782 26020 3834
rect 26032 3782 26084 3834
rect 10508 3723 10560 3732
rect 10508 3689 10517 3723
rect 10517 3689 10551 3723
rect 10551 3689 10560 3723
rect 10508 3680 10560 3689
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 12440 3680 12492 3732
rect 13084 3680 13136 3732
rect 17040 3680 17092 3732
rect 11612 3612 11664 3664
rect 11796 3655 11848 3664
rect 11796 3621 11805 3655
rect 11805 3621 11839 3655
rect 11839 3621 11848 3655
rect 11796 3612 11848 3621
rect 14372 3612 14424 3664
rect 12256 3544 12308 3596
rect 12532 3544 12584 3596
rect 14832 3612 14884 3664
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 14188 3476 14240 3528
rect 15108 3544 15160 3596
rect 18880 3544 18932 3596
rect 15384 3519 15436 3528
rect 15384 3485 15418 3519
rect 15418 3485 15436 3519
rect 15568 3519 15620 3528
rect 15384 3476 15436 3485
rect 15568 3485 15577 3519
rect 15577 3485 15611 3519
rect 15611 3485 15620 3519
rect 15568 3476 15620 3485
rect 29828 3519 29880 3528
rect 29828 3485 29837 3519
rect 29837 3485 29871 3519
rect 29871 3485 29880 3519
rect 29828 3476 29880 3485
rect 12348 3340 12400 3392
rect 12900 3340 12952 3392
rect 21456 3340 21508 3392
rect 10880 3238 10932 3290
rect 10944 3238 10996 3290
rect 11008 3238 11060 3290
rect 11072 3238 11124 3290
rect 11136 3238 11188 3290
rect 20811 3238 20863 3290
rect 20875 3238 20927 3290
rect 20939 3238 20991 3290
rect 21003 3238 21055 3290
rect 21067 3238 21119 3290
rect 1676 3000 1728 3052
rect 11244 3000 11296 3052
rect 12440 3136 12492 3188
rect 13176 3136 13228 3188
rect 12532 3043 12584 3052
rect 12532 3009 12566 3043
rect 12566 3009 12584 3043
rect 12532 3000 12584 3009
rect 11612 2932 11664 2984
rect 12900 2932 12952 2984
rect 15476 3136 15528 3188
rect 17132 3136 17184 3188
rect 29092 3136 29144 3188
rect 14188 3000 14240 3052
rect 14372 3000 14424 3052
rect 15200 3043 15252 3052
rect 15200 3009 15209 3043
rect 15209 3009 15243 3043
rect 15243 3009 15252 3043
rect 15200 3000 15252 3009
rect 15384 3000 15436 3052
rect 29920 3000 29972 3052
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 1584 2907 1636 2916
rect 1584 2873 1593 2907
rect 1593 2873 1627 2907
rect 1627 2873 1636 2907
rect 1584 2864 1636 2873
rect 12164 2907 12216 2916
rect 12164 2873 12173 2907
rect 12173 2873 12207 2907
rect 12207 2873 12216 2907
rect 12164 2864 12216 2873
rect 5915 2694 5967 2746
rect 5979 2694 6031 2746
rect 6043 2694 6095 2746
rect 6107 2694 6159 2746
rect 6171 2694 6223 2746
rect 15846 2694 15898 2746
rect 15910 2694 15962 2746
rect 15974 2694 16026 2746
rect 16038 2694 16090 2746
rect 16102 2694 16154 2746
rect 25776 2694 25828 2746
rect 25840 2694 25892 2746
rect 25904 2694 25956 2746
rect 25968 2694 26020 2746
rect 26032 2694 26084 2746
rect 13268 2635 13320 2644
rect 13268 2601 13277 2635
rect 13277 2601 13311 2635
rect 13311 2601 13320 2635
rect 13268 2592 13320 2601
rect 14740 2592 14792 2644
rect 20168 2592 20220 2644
rect 29000 2592 29052 2644
rect 9496 2388 9548 2440
rect 12440 2388 12492 2440
rect 14188 2388 14240 2440
rect 14372 2388 14424 2440
rect 28724 2431 28776 2440
rect 28724 2397 28733 2431
rect 28733 2397 28767 2431
rect 28767 2397 28776 2431
rect 28724 2388 28776 2397
rect 29736 2363 29788 2372
rect 29736 2329 29745 2363
rect 29745 2329 29779 2363
rect 29779 2329 29788 2363
rect 29736 2320 29788 2329
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 10880 2150 10932 2202
rect 10944 2150 10996 2202
rect 11008 2150 11060 2202
rect 11072 2150 11124 2202
rect 11136 2150 11188 2202
rect 20811 2150 20863 2202
rect 20875 2150 20927 2202
rect 20939 2150 20991 2202
rect 21003 2150 21055 2202
rect 21067 2150 21119 2202
<< metal2 >>
rect 386 47200 442 48000
rect 1122 47200 1178 48000
rect 1858 47200 1914 48000
rect 2594 47200 2650 48000
rect 3422 47200 3478 48000
rect 4158 47200 4214 48000
rect 4894 47200 4950 48000
rect 5722 47200 5778 48000
rect 6458 47200 6514 48000
rect 6564 47246 6868 47274
rect 400 43790 428 47200
rect 1136 45554 1164 47200
rect 1136 45526 1348 45554
rect 388 43784 440 43790
rect 388 43726 440 43732
rect 1320 25702 1348 45526
rect 1584 45484 1636 45490
rect 1584 45426 1636 45432
rect 1400 45280 1452 45286
rect 1400 45222 1452 45228
rect 1412 44946 1440 45222
rect 1596 44985 1624 45426
rect 1582 44976 1638 44985
rect 1400 44940 1452 44946
rect 1582 44911 1638 44920
rect 1400 44882 1452 44888
rect 1872 44878 1900 47200
rect 2608 45490 2636 47200
rect 2778 47016 2834 47025
rect 2778 46951 2834 46960
rect 2596 45484 2648 45490
rect 2596 45426 2648 45432
rect 2688 45416 2740 45422
rect 2688 45358 2740 45364
rect 1860 44872 1912 44878
rect 1860 44814 1912 44820
rect 2412 44804 2464 44810
rect 2412 44746 2464 44752
rect 2424 44402 2452 44746
rect 2044 44396 2096 44402
rect 2044 44338 2096 44344
rect 2412 44396 2464 44402
rect 2412 44338 2464 44344
rect 2056 43994 2084 44338
rect 2044 43988 2096 43994
rect 2044 43930 2096 43936
rect 1584 43308 1636 43314
rect 1584 43250 1636 43256
rect 1596 42945 1624 43250
rect 1582 42936 1638 42945
rect 1582 42871 1638 42880
rect 1584 41132 1636 41138
rect 1584 41074 1636 41080
rect 1596 41041 1624 41074
rect 1582 41032 1638 41041
rect 1582 40967 1638 40976
rect 1584 39432 1636 39438
rect 1584 39374 1636 39380
rect 1596 39001 1624 39374
rect 1582 38992 1638 39001
rect 1582 38927 1638 38936
rect 1584 37256 1636 37262
rect 1584 37198 1636 37204
rect 1596 36961 1624 37198
rect 1582 36952 1638 36961
rect 1582 36887 1638 36896
rect 1584 35080 1636 35086
rect 1582 35048 1584 35057
rect 1636 35048 1638 35057
rect 1582 34983 1638 34992
rect 1400 34196 1452 34202
rect 1400 34138 1452 34144
rect 1412 33658 1440 34138
rect 1400 33652 1452 33658
rect 1400 33594 1452 33600
rect 1584 33516 1636 33522
rect 1584 33458 1636 33464
rect 1596 33017 1624 33458
rect 1582 33008 1638 33017
rect 1582 32943 1638 32952
rect 1400 31272 1452 31278
rect 1400 31214 1452 31220
rect 1412 30977 1440 31214
rect 1398 30968 1454 30977
rect 1398 30903 1454 30912
rect 2320 29164 2372 29170
rect 2320 29106 2372 29112
rect 1584 29028 1636 29034
rect 1584 28970 1636 28976
rect 1596 28937 1624 28970
rect 1582 28928 1638 28937
rect 1582 28863 1638 28872
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1412 26042 1440 27406
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1596 27033 1624 27270
rect 1582 27024 1638 27033
rect 1582 26959 1638 26968
rect 1676 26852 1728 26858
rect 1676 26794 1728 26800
rect 1400 26036 1452 26042
rect 1400 25978 1452 25984
rect 1308 25696 1360 25702
rect 1308 25638 1360 25644
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1412 24954 1440 25230
rect 1584 25152 1636 25158
rect 1584 25094 1636 25100
rect 1596 24993 1624 25094
rect 1582 24984 1638 24993
rect 1400 24948 1452 24954
rect 1582 24919 1638 24928
rect 1400 24890 1452 24896
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1596 24342 1624 24754
rect 1584 24336 1636 24342
rect 1584 24278 1636 24284
rect 1584 22976 1636 22982
rect 1582 22944 1584 22953
rect 1636 22944 1638 22953
rect 1582 22879 1638 22888
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1596 21049 1624 21286
rect 1582 21040 1638 21049
rect 1582 20975 1638 20984
rect 1584 20392 1636 20398
rect 1584 20334 1636 20340
rect 1596 19854 1624 20334
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1400 19712 1452 19718
rect 1400 19654 1452 19660
rect 1412 19378 1440 19654
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1596 19009 1624 19110
rect 1582 19000 1638 19009
rect 1582 18935 1638 18944
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1400 17536 1452 17542
rect 1400 17478 1452 17484
rect 1412 17202 1440 17478
rect 1596 17338 1624 17614
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1400 15360 1452 15366
rect 1400 15302 1452 15308
rect 1412 15026 1440 15302
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1504 5234 1532 17138
rect 1584 16992 1636 16998
rect 1582 16960 1584 16969
rect 1636 16960 1638 16969
rect 1582 16895 1638 16904
rect 1582 14920 1638 14929
rect 1582 14855 1584 14864
rect 1636 14855 1638 14864
rect 1584 14826 1636 14832
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 13025 1624 13126
rect 1582 13016 1638 13025
rect 1582 12951 1638 12960
rect 1584 11008 1636 11014
rect 1582 10976 1584 10985
rect 1636 10976 1638 10985
rect 1582 10911 1638 10920
rect 1582 8936 1638 8945
rect 1582 8871 1638 8880
rect 1596 8838 1624 8871
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 7041 1624 7142
rect 1582 7032 1638 7041
rect 1582 6967 1638 6976
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1584 5024 1636 5030
rect 1582 4992 1584 5001
rect 1636 4992 1638 5001
rect 1582 4927 1638 4936
rect 1688 3058 1716 26794
rect 2228 26240 2280 26246
rect 2228 26182 2280 26188
rect 2240 25906 2268 26182
rect 2332 26042 2360 29106
rect 2320 26036 2372 26042
rect 2320 25978 2372 25984
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 2228 25900 2280 25906
rect 2228 25842 2280 25848
rect 1780 24818 1808 25842
rect 1768 24812 1820 24818
rect 1768 24754 1820 24760
rect 2320 24812 2372 24818
rect 2320 24754 2372 24760
rect 2332 23118 2360 24754
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 2136 22092 2188 22098
rect 2136 22034 2188 22040
rect 2148 21554 2176 22034
rect 2332 21554 2360 23054
rect 2136 21548 2188 21554
rect 2136 21490 2188 21496
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 2332 19854 2360 21490
rect 2424 21078 2452 44338
rect 2700 44334 2728 45358
rect 2792 44470 2820 46951
rect 3436 45490 3464 47200
rect 4172 45490 4200 47200
rect 3424 45484 3476 45490
rect 3424 45426 3476 45432
rect 4160 45484 4212 45490
rect 4160 45426 4212 45432
rect 4908 44878 4936 47200
rect 5736 45490 5764 47200
rect 6472 47138 6500 47200
rect 6564 47138 6592 47246
rect 6472 47110 6592 47138
rect 6840 45506 6868 47246
rect 7194 47200 7250 48000
rect 7930 47200 7986 48000
rect 8758 47200 8814 48000
rect 9494 47200 9550 48000
rect 10230 47200 10286 48000
rect 11058 47200 11114 48000
rect 11794 47200 11850 48000
rect 12530 47200 12586 48000
rect 13266 47200 13322 48000
rect 14094 47200 14150 48000
rect 14830 47200 14886 48000
rect 15566 47200 15622 48000
rect 16394 47200 16450 48000
rect 17130 47200 17186 48000
rect 17866 47200 17922 48000
rect 18602 47200 18658 48000
rect 19430 47200 19486 48000
rect 20166 47200 20222 48000
rect 20902 47200 20958 48000
rect 21008 47246 21220 47274
rect 6840 45490 6960 45506
rect 5724 45484 5776 45490
rect 6840 45484 6972 45490
rect 6840 45478 6920 45484
rect 5724 45426 5776 45432
rect 6920 45426 6972 45432
rect 5356 45416 5408 45422
rect 5356 45358 5408 45364
rect 4896 44872 4948 44878
rect 4896 44814 4948 44820
rect 5172 44736 5224 44742
rect 5172 44678 5224 44684
rect 5184 44538 5212 44678
rect 5172 44532 5224 44538
rect 5172 44474 5224 44480
rect 2780 44464 2832 44470
rect 2780 44406 2832 44412
rect 2596 44328 2648 44334
rect 2596 44270 2648 44276
rect 2688 44328 2740 44334
rect 2688 44270 2740 44276
rect 2608 41546 2636 44270
rect 2596 41540 2648 41546
rect 2596 41482 2648 41488
rect 5368 40662 5396 45358
rect 7012 45280 7064 45286
rect 7012 45222 7064 45228
rect 5915 45180 6223 45200
rect 5915 45178 5921 45180
rect 5977 45178 6001 45180
rect 6057 45178 6081 45180
rect 6137 45178 6161 45180
rect 6217 45178 6223 45180
rect 5977 45126 5979 45178
rect 6159 45126 6161 45178
rect 5915 45124 5921 45126
rect 5977 45124 6001 45126
rect 6057 45124 6081 45126
rect 6137 45124 6161 45126
rect 6217 45124 6223 45126
rect 5915 45104 6223 45124
rect 5915 44092 6223 44112
rect 5915 44090 5921 44092
rect 5977 44090 6001 44092
rect 6057 44090 6081 44092
rect 6137 44090 6161 44092
rect 6217 44090 6223 44092
rect 5977 44038 5979 44090
rect 6159 44038 6161 44090
rect 5915 44036 5921 44038
rect 5977 44036 6001 44038
rect 6057 44036 6081 44038
rect 6137 44036 6161 44038
rect 6217 44036 6223 44038
rect 5915 44016 6223 44036
rect 5915 43004 6223 43024
rect 5915 43002 5921 43004
rect 5977 43002 6001 43004
rect 6057 43002 6081 43004
rect 6137 43002 6161 43004
rect 6217 43002 6223 43004
rect 5977 42950 5979 43002
rect 6159 42950 6161 43002
rect 5915 42948 5921 42950
rect 5977 42948 6001 42950
rect 6057 42948 6081 42950
rect 6137 42948 6161 42950
rect 6217 42948 6223 42950
rect 5915 42928 6223 42948
rect 5915 41916 6223 41936
rect 5915 41914 5921 41916
rect 5977 41914 6001 41916
rect 6057 41914 6081 41916
rect 6137 41914 6161 41916
rect 6217 41914 6223 41916
rect 5977 41862 5979 41914
rect 6159 41862 6161 41914
rect 5915 41860 5921 41862
rect 5977 41860 6001 41862
rect 6057 41860 6081 41862
rect 6137 41860 6161 41862
rect 6217 41860 6223 41862
rect 5915 41840 6223 41860
rect 5915 40828 6223 40848
rect 5915 40826 5921 40828
rect 5977 40826 6001 40828
rect 6057 40826 6081 40828
rect 6137 40826 6161 40828
rect 6217 40826 6223 40828
rect 5977 40774 5979 40826
rect 6159 40774 6161 40826
rect 5915 40772 5921 40774
rect 5977 40772 6001 40774
rect 6057 40772 6081 40774
rect 6137 40772 6161 40774
rect 6217 40772 6223 40774
rect 5915 40752 6223 40772
rect 5356 40656 5408 40662
rect 5356 40598 5408 40604
rect 5915 39740 6223 39760
rect 5915 39738 5921 39740
rect 5977 39738 6001 39740
rect 6057 39738 6081 39740
rect 6137 39738 6161 39740
rect 6217 39738 6223 39740
rect 5977 39686 5979 39738
rect 6159 39686 6161 39738
rect 5915 39684 5921 39686
rect 5977 39684 6001 39686
rect 6057 39684 6081 39686
rect 6137 39684 6161 39686
rect 6217 39684 6223 39686
rect 5915 39664 6223 39684
rect 5915 38652 6223 38672
rect 5915 38650 5921 38652
rect 5977 38650 6001 38652
rect 6057 38650 6081 38652
rect 6137 38650 6161 38652
rect 6217 38650 6223 38652
rect 5977 38598 5979 38650
rect 6159 38598 6161 38650
rect 5915 38596 5921 38598
rect 5977 38596 6001 38598
rect 6057 38596 6081 38598
rect 6137 38596 6161 38598
rect 6217 38596 6223 38598
rect 5915 38576 6223 38596
rect 7024 37942 7052 45222
rect 7208 44878 7236 47200
rect 7944 45490 7972 47200
rect 8772 45490 8800 47200
rect 9508 45490 9536 47200
rect 7932 45484 7984 45490
rect 7932 45426 7984 45432
rect 8760 45484 8812 45490
rect 8760 45426 8812 45432
rect 9496 45484 9548 45490
rect 9496 45426 9548 45432
rect 8852 45416 8904 45422
rect 8852 45358 8904 45364
rect 7196 44872 7248 44878
rect 7196 44814 7248 44820
rect 7012 37936 7064 37942
rect 7012 37878 7064 37884
rect 5915 37564 6223 37584
rect 5915 37562 5921 37564
rect 5977 37562 6001 37564
rect 6057 37562 6081 37564
rect 6137 37562 6161 37564
rect 6217 37562 6223 37564
rect 5977 37510 5979 37562
rect 6159 37510 6161 37562
rect 5915 37508 5921 37510
rect 5977 37508 6001 37510
rect 6057 37508 6081 37510
rect 6137 37508 6161 37510
rect 6217 37508 6223 37510
rect 5915 37488 6223 37508
rect 8864 36786 8892 45358
rect 8944 45348 8996 45354
rect 8944 45290 8996 45296
rect 8956 45082 8984 45290
rect 9864 45280 9916 45286
rect 9864 45222 9916 45228
rect 8944 45076 8996 45082
rect 8944 45018 8996 45024
rect 9772 45008 9824 45014
rect 9772 44950 9824 44956
rect 8852 36780 8904 36786
rect 8852 36722 8904 36728
rect 9680 36780 9732 36786
rect 9680 36722 9732 36728
rect 9312 36576 9364 36582
rect 9312 36518 9364 36524
rect 5915 36476 6223 36496
rect 5915 36474 5921 36476
rect 5977 36474 6001 36476
rect 6057 36474 6081 36476
rect 6137 36474 6161 36476
rect 6217 36474 6223 36476
rect 5977 36422 5979 36474
rect 6159 36422 6161 36474
rect 5915 36420 5921 36422
rect 5977 36420 6001 36422
rect 6057 36420 6081 36422
rect 6137 36420 6161 36422
rect 6217 36420 6223 36422
rect 5915 36400 6223 36420
rect 9324 35698 9352 36518
rect 9692 36038 9720 36722
rect 9680 36032 9732 36038
rect 9680 35974 9732 35980
rect 9312 35692 9364 35698
rect 9312 35634 9364 35640
rect 9692 35494 9720 35974
rect 9680 35488 9732 35494
rect 9680 35430 9732 35436
rect 5915 35388 6223 35408
rect 5915 35386 5921 35388
rect 5977 35386 6001 35388
rect 6057 35386 6081 35388
rect 6137 35386 6161 35388
rect 6217 35386 6223 35388
rect 5977 35334 5979 35386
rect 6159 35334 6161 35386
rect 5915 35332 5921 35334
rect 5977 35332 6001 35334
rect 6057 35332 6081 35334
rect 6137 35332 6161 35334
rect 6217 35332 6223 35334
rect 5915 35312 6223 35332
rect 5915 34300 6223 34320
rect 5915 34298 5921 34300
rect 5977 34298 6001 34300
rect 6057 34298 6081 34300
rect 6137 34298 6161 34300
rect 6217 34298 6223 34300
rect 5977 34246 5979 34298
rect 6159 34246 6161 34298
rect 5915 34244 5921 34246
rect 5977 34244 6001 34246
rect 6057 34244 6081 34246
rect 6137 34244 6161 34246
rect 6217 34244 6223 34246
rect 5915 34224 6223 34244
rect 9680 33312 9732 33318
rect 9680 33254 9732 33260
rect 5915 33212 6223 33232
rect 5915 33210 5921 33212
rect 5977 33210 6001 33212
rect 6057 33210 6081 33212
rect 6137 33210 6161 33212
rect 6217 33210 6223 33212
rect 5977 33158 5979 33210
rect 6159 33158 6161 33210
rect 5915 33156 5921 33158
rect 5977 33156 6001 33158
rect 6057 33156 6081 33158
rect 6137 33156 6161 33158
rect 6217 33156 6223 33158
rect 5915 33136 6223 33156
rect 9588 32224 9640 32230
rect 9588 32166 9640 32172
rect 5915 32124 6223 32144
rect 5915 32122 5921 32124
rect 5977 32122 6001 32124
rect 6057 32122 6081 32124
rect 6137 32122 6161 32124
rect 6217 32122 6223 32124
rect 5977 32070 5979 32122
rect 6159 32070 6161 32122
rect 5915 32068 5921 32070
rect 5977 32068 6001 32070
rect 6057 32068 6081 32070
rect 6137 32068 6161 32070
rect 6217 32068 6223 32070
rect 5915 32048 6223 32068
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 8852 31340 8904 31346
rect 8852 31282 8904 31288
rect 5915 31036 6223 31056
rect 5915 31034 5921 31036
rect 5977 31034 6001 31036
rect 6057 31034 6081 31036
rect 6137 31034 6161 31036
rect 6217 31034 6223 31036
rect 5977 30982 5979 31034
rect 6159 30982 6161 31034
rect 5915 30980 5921 30982
rect 5977 30980 6001 30982
rect 6057 30980 6081 30982
rect 6137 30980 6161 30982
rect 6217 30980 6223 30982
rect 5915 30960 6223 30980
rect 5915 29948 6223 29968
rect 5915 29946 5921 29948
rect 5977 29946 6001 29948
rect 6057 29946 6081 29948
rect 6137 29946 6161 29948
rect 6217 29946 6223 29948
rect 5977 29894 5979 29946
rect 6159 29894 6161 29946
rect 5915 29892 5921 29894
rect 5977 29892 6001 29894
rect 6057 29892 6081 29894
rect 6137 29892 6161 29894
rect 6217 29892 6223 29894
rect 5915 29872 6223 29892
rect 7840 29232 7892 29238
rect 7840 29174 7892 29180
rect 5915 28860 6223 28880
rect 5915 28858 5921 28860
rect 5977 28858 6001 28860
rect 6057 28858 6081 28860
rect 6137 28858 6161 28860
rect 6217 28858 6223 28860
rect 5977 28806 5979 28858
rect 6159 28806 6161 28858
rect 5915 28804 5921 28806
rect 5977 28804 6001 28806
rect 6057 28804 6081 28806
rect 6137 28804 6161 28806
rect 6217 28804 6223 28806
rect 5915 28784 6223 28804
rect 7852 28082 7880 29174
rect 7932 28960 7984 28966
rect 7932 28902 7984 28908
rect 7944 28558 7972 28902
rect 8220 28626 8248 31282
rect 8864 30394 8892 31282
rect 9496 30592 9548 30598
rect 9496 30534 9548 30540
rect 8852 30388 8904 30394
rect 8852 30330 8904 30336
rect 8852 30252 8904 30258
rect 8852 30194 8904 30200
rect 9312 30252 9364 30258
rect 9312 30194 9364 30200
rect 8864 29850 8892 30194
rect 8852 29844 8904 29850
rect 8852 29786 8904 29792
rect 9324 29646 9352 30194
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 8392 29504 8444 29510
rect 8392 29446 8444 29452
rect 8404 29170 8432 29446
rect 8392 29164 8444 29170
rect 8392 29106 8444 29112
rect 9324 29102 9352 29582
rect 8300 29096 8352 29102
rect 8300 29038 8352 29044
rect 9312 29096 9364 29102
rect 9312 29038 9364 29044
rect 9508 29050 9536 30534
rect 9600 29646 9628 32166
rect 9588 29640 9640 29646
rect 9588 29582 9640 29588
rect 9692 29170 9720 33254
rect 9784 30598 9812 44950
rect 9772 30592 9824 30598
rect 9772 30534 9824 30540
rect 9772 30320 9824 30326
rect 9772 30262 9824 30268
rect 9784 29510 9812 30262
rect 9876 30002 9904 45222
rect 10244 44878 10272 47200
rect 11072 46458 11100 47200
rect 11072 46430 11284 46458
rect 10880 45724 11188 45744
rect 10880 45722 10886 45724
rect 10942 45722 10966 45724
rect 11022 45722 11046 45724
rect 11102 45722 11126 45724
rect 11182 45722 11188 45724
rect 10942 45670 10944 45722
rect 11124 45670 11126 45722
rect 10880 45668 10886 45670
rect 10942 45668 10966 45670
rect 11022 45668 11046 45670
rect 11102 45668 11126 45670
rect 11182 45668 11188 45670
rect 10880 45648 11188 45668
rect 11256 45490 11284 46430
rect 11244 45484 11296 45490
rect 11244 45426 11296 45432
rect 11704 45280 11756 45286
rect 11704 45222 11756 45228
rect 11244 44940 11296 44946
rect 11244 44882 11296 44888
rect 10232 44872 10284 44878
rect 10232 44814 10284 44820
rect 10048 44736 10100 44742
rect 10048 44678 10100 44684
rect 9956 37868 10008 37874
rect 9956 37810 10008 37816
rect 9968 37194 9996 37810
rect 9956 37188 10008 37194
rect 9956 37130 10008 37136
rect 9968 36854 9996 37130
rect 9956 36848 10008 36854
rect 9956 36790 10008 36796
rect 10060 36786 10088 44678
rect 10880 44636 11188 44656
rect 10880 44634 10886 44636
rect 10942 44634 10966 44636
rect 11022 44634 11046 44636
rect 11102 44634 11126 44636
rect 11182 44634 11188 44636
rect 10942 44582 10944 44634
rect 11124 44582 11126 44634
rect 10880 44580 10886 44582
rect 10942 44580 10966 44582
rect 11022 44580 11046 44582
rect 11102 44580 11126 44582
rect 11182 44580 11188 44582
rect 10880 44560 11188 44580
rect 10876 44260 10928 44266
rect 10876 44202 10928 44208
rect 10888 43858 10916 44202
rect 11256 43858 11284 44882
rect 10876 43852 10928 43858
rect 10876 43794 10928 43800
rect 11244 43852 11296 43858
rect 11244 43794 11296 43800
rect 11336 43784 11388 43790
rect 11336 43726 11388 43732
rect 11244 43648 11296 43654
rect 11244 43590 11296 43596
rect 10880 43548 11188 43568
rect 10880 43546 10886 43548
rect 10942 43546 10966 43548
rect 11022 43546 11046 43548
rect 11102 43546 11126 43548
rect 11182 43546 11188 43548
rect 10942 43494 10944 43546
rect 11124 43494 11126 43546
rect 10880 43492 10886 43494
rect 10942 43492 10966 43494
rect 11022 43492 11046 43494
rect 11102 43492 11126 43494
rect 11182 43492 11188 43494
rect 10880 43472 11188 43492
rect 11256 43178 11284 43590
rect 11244 43172 11296 43178
rect 11244 43114 11296 43120
rect 10876 43104 10928 43110
rect 10876 43046 10928 43052
rect 10888 42770 10916 43046
rect 10876 42764 10928 42770
rect 10876 42706 10928 42712
rect 11348 42702 11376 43726
rect 11336 42696 11388 42702
rect 11336 42638 11388 42644
rect 11244 42560 11296 42566
rect 11244 42502 11296 42508
rect 10880 42460 11188 42480
rect 10880 42458 10886 42460
rect 10942 42458 10966 42460
rect 11022 42458 11046 42460
rect 11102 42458 11126 42460
rect 11182 42458 11188 42460
rect 10942 42406 10944 42458
rect 11124 42406 11126 42458
rect 10880 42404 10886 42406
rect 10942 42404 10966 42406
rect 11022 42404 11046 42406
rect 11102 42404 11126 42406
rect 11182 42404 11188 42406
rect 10880 42384 11188 42404
rect 11256 42294 11284 42502
rect 11244 42288 11296 42294
rect 11244 42230 11296 42236
rect 10880 41372 11188 41392
rect 10880 41370 10886 41372
rect 10942 41370 10966 41372
rect 11022 41370 11046 41372
rect 11102 41370 11126 41372
rect 11182 41370 11188 41372
rect 10942 41318 10944 41370
rect 11124 41318 11126 41370
rect 10880 41316 10886 41318
rect 10942 41316 10966 41318
rect 11022 41316 11046 41318
rect 11102 41316 11126 41318
rect 11182 41316 11188 41318
rect 10880 41296 11188 41316
rect 10880 40284 11188 40304
rect 10880 40282 10886 40284
rect 10942 40282 10966 40284
rect 11022 40282 11046 40284
rect 11102 40282 11126 40284
rect 11182 40282 11188 40284
rect 10942 40230 10944 40282
rect 11124 40230 11126 40282
rect 10880 40228 10886 40230
rect 10942 40228 10966 40230
rect 11022 40228 11046 40230
rect 11102 40228 11126 40230
rect 11182 40228 11188 40230
rect 10880 40208 11188 40228
rect 10880 39196 11188 39216
rect 10880 39194 10886 39196
rect 10942 39194 10966 39196
rect 11022 39194 11046 39196
rect 11102 39194 11126 39196
rect 11182 39194 11188 39196
rect 10942 39142 10944 39194
rect 11124 39142 11126 39194
rect 10880 39140 10886 39142
rect 10942 39140 10966 39142
rect 11022 39140 11046 39142
rect 11102 39140 11126 39142
rect 11182 39140 11188 39142
rect 10880 39120 11188 39140
rect 10140 38344 10192 38350
rect 10140 38286 10192 38292
rect 10152 37262 10180 38286
rect 10600 38276 10652 38282
rect 10600 38218 10652 38224
rect 10324 37800 10376 37806
rect 10324 37742 10376 37748
rect 10508 37800 10560 37806
rect 10508 37742 10560 37748
rect 10140 37256 10192 37262
rect 10140 37198 10192 37204
rect 10336 36786 10364 37742
rect 10416 37256 10468 37262
rect 10416 37198 10468 37204
rect 10048 36780 10100 36786
rect 10048 36722 10100 36728
rect 10324 36780 10376 36786
rect 10324 36722 10376 36728
rect 10428 36650 10456 37198
rect 10416 36644 10468 36650
rect 10416 36586 10468 36592
rect 10428 35766 10456 36586
rect 10520 36582 10548 37742
rect 10612 36922 10640 38218
rect 11244 38208 11296 38214
rect 11244 38150 11296 38156
rect 10880 38108 11188 38128
rect 10880 38106 10886 38108
rect 10942 38106 10966 38108
rect 11022 38106 11046 38108
rect 11102 38106 11126 38108
rect 11182 38106 11188 38108
rect 10942 38054 10944 38106
rect 11124 38054 11126 38106
rect 10880 38052 10886 38054
rect 10942 38052 10966 38054
rect 11022 38052 11046 38054
rect 11102 38052 11126 38054
rect 11182 38052 11188 38054
rect 10880 38032 11188 38052
rect 10784 37868 10836 37874
rect 10784 37810 10836 37816
rect 10692 37664 10744 37670
rect 10692 37606 10744 37612
rect 10704 37262 10732 37606
rect 10692 37256 10744 37262
rect 10692 37198 10744 37204
rect 10796 37126 10824 37810
rect 10692 37120 10744 37126
rect 10692 37062 10744 37068
rect 10784 37120 10836 37126
rect 10784 37062 10836 37068
rect 10704 36922 10732 37062
rect 10600 36916 10652 36922
rect 10600 36858 10652 36864
rect 10692 36916 10744 36922
rect 10692 36858 10744 36864
rect 10508 36576 10560 36582
rect 10508 36518 10560 36524
rect 10416 35760 10468 35766
rect 10416 35702 10468 35708
rect 10140 35080 10192 35086
rect 10140 35022 10192 35028
rect 10048 34604 10100 34610
rect 10048 34546 10100 34552
rect 10060 33930 10088 34546
rect 10048 33924 10100 33930
rect 10048 33866 10100 33872
rect 9956 33448 10008 33454
rect 9956 33390 10008 33396
rect 9968 33114 9996 33390
rect 9956 33108 10008 33114
rect 9956 33050 10008 33056
rect 9956 32904 10008 32910
rect 9956 32846 10008 32852
rect 9968 31210 9996 32846
rect 9956 31204 10008 31210
rect 9956 31146 10008 31152
rect 10060 30784 10088 33866
rect 9968 30756 10088 30784
rect 9968 30161 9996 30756
rect 10048 30660 10100 30666
rect 10048 30602 10100 30608
rect 9954 30152 10010 30161
rect 9954 30087 10010 30096
rect 9876 29974 9996 30002
rect 9864 29572 9916 29578
rect 9864 29514 9916 29520
rect 9772 29504 9824 29510
rect 9772 29446 9824 29452
rect 9784 29306 9812 29446
rect 9772 29300 9824 29306
rect 9772 29242 9824 29248
rect 9680 29164 9732 29170
rect 9680 29106 9732 29112
rect 8312 28762 8340 29038
rect 9508 29022 9720 29050
rect 9876 29034 9904 29514
rect 8300 28756 8352 28762
rect 8300 28698 8352 28704
rect 8208 28620 8260 28626
rect 8208 28562 8260 28568
rect 7932 28552 7984 28558
rect 7932 28494 7984 28500
rect 7840 28076 7892 28082
rect 7840 28018 7892 28024
rect 8024 27872 8076 27878
rect 8024 27814 8076 27820
rect 5915 27772 6223 27792
rect 5915 27770 5921 27772
rect 5977 27770 6001 27772
rect 6057 27770 6081 27772
rect 6137 27770 6161 27772
rect 6217 27770 6223 27772
rect 5977 27718 5979 27770
rect 6159 27718 6161 27770
rect 5915 27716 5921 27718
rect 5977 27716 6001 27718
rect 6057 27716 6081 27718
rect 6137 27716 6161 27718
rect 6217 27716 6223 27718
rect 5915 27696 6223 27716
rect 8036 27470 8064 27814
rect 8024 27464 8076 27470
rect 8024 27406 8076 27412
rect 9588 27396 9640 27402
rect 9588 27338 9640 27344
rect 7748 27328 7800 27334
rect 7748 27270 7800 27276
rect 5915 26684 6223 26704
rect 5915 26682 5921 26684
rect 5977 26682 6001 26684
rect 6057 26682 6081 26684
rect 6137 26682 6161 26684
rect 6217 26682 6223 26684
rect 5977 26630 5979 26682
rect 6159 26630 6161 26682
rect 5915 26628 5921 26630
rect 5977 26628 6001 26630
rect 6057 26628 6081 26630
rect 6137 26628 6161 26630
rect 6217 26628 6223 26630
rect 5915 26608 6223 26628
rect 5264 25968 5316 25974
rect 5264 25910 5316 25916
rect 5276 25430 5304 25910
rect 5915 25596 6223 25616
rect 5915 25594 5921 25596
rect 5977 25594 6001 25596
rect 6057 25594 6081 25596
rect 6137 25594 6161 25596
rect 6217 25594 6223 25596
rect 5977 25542 5979 25594
rect 6159 25542 6161 25594
rect 5915 25540 5921 25542
rect 5977 25540 6001 25542
rect 6057 25540 6081 25542
rect 6137 25540 6161 25542
rect 6217 25540 6223 25542
rect 5915 25520 6223 25540
rect 5264 25424 5316 25430
rect 5264 25366 5316 25372
rect 5915 24508 6223 24528
rect 5915 24506 5921 24508
rect 5977 24506 6001 24508
rect 6057 24506 6081 24508
rect 6137 24506 6161 24508
rect 6217 24506 6223 24508
rect 5977 24454 5979 24506
rect 6159 24454 6161 24506
rect 5915 24452 5921 24454
rect 5977 24452 6001 24454
rect 6057 24452 6081 24454
rect 6137 24452 6161 24454
rect 6217 24452 6223 24454
rect 5915 24432 6223 24452
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7576 23730 7604 24006
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7288 23656 7340 23662
rect 7288 23598 7340 23604
rect 5915 23420 6223 23440
rect 5915 23418 5921 23420
rect 5977 23418 6001 23420
rect 6057 23418 6081 23420
rect 6137 23418 6161 23420
rect 6217 23418 6223 23420
rect 5977 23366 5979 23418
rect 6159 23366 6161 23418
rect 5915 23364 5921 23366
rect 5977 23364 6001 23366
rect 6057 23364 6081 23366
rect 6137 23364 6161 23366
rect 6217 23364 6223 23366
rect 5915 23344 6223 23364
rect 5915 22332 6223 22352
rect 5915 22330 5921 22332
rect 5977 22330 6001 22332
rect 6057 22330 6081 22332
rect 6137 22330 6161 22332
rect 6217 22330 6223 22332
rect 5977 22278 5979 22330
rect 6159 22278 6161 22330
rect 5915 22276 5921 22278
rect 5977 22276 6001 22278
rect 6057 22276 6081 22278
rect 6137 22276 6161 22278
rect 6217 22276 6223 22278
rect 5915 22256 6223 22276
rect 7300 21554 7328 23598
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 5915 21244 6223 21264
rect 5915 21242 5921 21244
rect 5977 21242 6001 21244
rect 6057 21242 6081 21244
rect 6137 21242 6161 21244
rect 6217 21242 6223 21244
rect 5977 21190 5979 21242
rect 6159 21190 6161 21242
rect 5915 21188 5921 21190
rect 5977 21188 6001 21190
rect 6057 21188 6081 21190
rect 6137 21188 6161 21190
rect 6217 21188 6223 21190
rect 5915 21168 6223 21188
rect 2412 21072 2464 21078
rect 2412 21014 2464 21020
rect 5915 20156 6223 20176
rect 5915 20154 5921 20156
rect 5977 20154 6001 20156
rect 6057 20154 6081 20156
rect 6137 20154 6161 20156
rect 6217 20154 6223 20156
rect 5977 20102 5979 20154
rect 6159 20102 6161 20154
rect 5915 20100 5921 20102
rect 5977 20100 6001 20102
rect 6057 20100 6081 20102
rect 6137 20100 6161 20102
rect 6217 20100 6223 20102
rect 5915 20080 6223 20100
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 2320 19848 2372 19854
rect 2320 19790 2372 19796
rect 1780 17678 1808 19790
rect 5915 19068 6223 19088
rect 5915 19066 5921 19068
rect 5977 19066 6001 19068
rect 6057 19066 6081 19068
rect 6137 19066 6161 19068
rect 6217 19066 6223 19068
rect 5977 19014 5979 19066
rect 6159 19014 6161 19066
rect 5915 19012 5921 19014
rect 5977 19012 6001 19014
rect 6057 19012 6081 19014
rect 6137 19012 6161 19014
rect 6217 19012 6223 19014
rect 5915 18992 6223 19012
rect 2688 18352 2740 18358
rect 2688 18294 2740 18300
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1780 15502 1808 17614
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 13326 1808 15438
rect 1768 13320 1820 13326
rect 1768 13262 1820 13268
rect 1872 7410 1900 16934
rect 2700 15570 2728 18294
rect 7760 18290 7788 27270
rect 9312 26988 9364 26994
rect 9312 26930 9364 26936
rect 8852 26920 8904 26926
rect 8852 26862 8904 26868
rect 8864 25226 8892 26862
rect 8944 26784 8996 26790
rect 8944 26726 8996 26732
rect 8956 26450 8984 26726
rect 8944 26444 8996 26450
rect 8944 26386 8996 26392
rect 9036 26376 9088 26382
rect 9036 26318 9088 26324
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 9048 25498 9076 26318
rect 9140 25906 9168 26318
rect 9128 25900 9180 25906
rect 9128 25842 9180 25848
rect 9220 25900 9272 25906
rect 9220 25842 9272 25848
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 8852 25220 8904 25226
rect 8852 25162 8904 25168
rect 8864 24886 8892 25162
rect 9232 24954 9260 25842
rect 9324 25226 9352 26930
rect 9600 26586 9628 27338
rect 9588 26580 9640 26586
rect 9588 26522 9640 26528
rect 9692 26518 9720 29022
rect 9864 29028 9916 29034
rect 9864 28970 9916 28976
rect 9864 28552 9916 28558
rect 9864 28494 9916 28500
rect 9772 27872 9824 27878
rect 9772 27814 9824 27820
rect 9784 27282 9812 27814
rect 9876 27402 9904 28494
rect 9968 28218 9996 29974
rect 10060 29646 10088 30602
rect 10048 29640 10100 29646
rect 10048 29582 10100 29588
rect 10060 28422 10088 29582
rect 10152 29238 10180 35022
rect 10232 33992 10284 33998
rect 10230 33960 10232 33969
rect 10284 33960 10286 33969
rect 10230 33895 10286 33904
rect 10414 33960 10470 33969
rect 10414 33895 10470 33904
rect 10232 33856 10284 33862
rect 10232 33798 10284 33804
rect 10244 32910 10272 33798
rect 10324 33448 10376 33454
rect 10324 33390 10376 33396
rect 10336 33046 10364 33390
rect 10324 33040 10376 33046
rect 10324 32982 10376 32988
rect 10232 32904 10284 32910
rect 10232 32846 10284 32852
rect 10244 31958 10272 32846
rect 10336 32450 10364 32982
rect 10428 32910 10456 33895
rect 10416 32904 10468 32910
rect 10416 32846 10468 32852
rect 10336 32422 10456 32450
rect 10324 32360 10376 32366
rect 10324 32302 10376 32308
rect 10336 32026 10364 32302
rect 10324 32020 10376 32026
rect 10324 31962 10376 31968
rect 10232 31952 10284 31958
rect 10232 31894 10284 31900
rect 10428 31822 10456 32422
rect 10416 31816 10468 31822
rect 10416 31758 10468 31764
rect 10520 31686 10548 36518
rect 10796 36106 10824 37062
rect 10880 37020 11188 37040
rect 10880 37018 10886 37020
rect 10942 37018 10966 37020
rect 11022 37018 11046 37020
rect 11102 37018 11126 37020
rect 11182 37018 11188 37020
rect 10942 36966 10944 37018
rect 11124 36966 11126 37018
rect 10880 36964 10886 36966
rect 10942 36964 10966 36966
rect 11022 36964 11046 36966
rect 11102 36964 11126 36966
rect 11182 36964 11188 36966
rect 10880 36944 11188 36964
rect 11256 36786 11284 38150
rect 11244 36780 11296 36786
rect 11244 36722 11296 36728
rect 11256 36174 11284 36722
rect 11244 36168 11296 36174
rect 11244 36110 11296 36116
rect 10784 36100 10836 36106
rect 10784 36042 10836 36048
rect 10880 35932 11188 35952
rect 10880 35930 10886 35932
rect 10942 35930 10966 35932
rect 11022 35930 11046 35932
rect 11102 35930 11126 35932
rect 11182 35930 11188 35932
rect 10942 35878 10944 35930
rect 11124 35878 11126 35930
rect 10880 35876 10886 35878
rect 10942 35876 10966 35878
rect 11022 35876 11046 35878
rect 11102 35876 11126 35878
rect 11182 35876 11188 35878
rect 10880 35856 11188 35876
rect 11244 34944 11296 34950
rect 11244 34886 11296 34892
rect 10880 34844 11188 34864
rect 10880 34842 10886 34844
rect 10942 34842 10966 34844
rect 11022 34842 11046 34844
rect 11102 34842 11126 34844
rect 11182 34842 11188 34844
rect 10942 34790 10944 34842
rect 11124 34790 11126 34842
rect 10880 34788 10886 34790
rect 10942 34788 10966 34790
rect 11022 34788 11046 34790
rect 11102 34788 11126 34790
rect 11182 34788 11188 34790
rect 10880 34768 11188 34788
rect 10692 34740 10744 34746
rect 10692 34682 10744 34688
rect 10600 33992 10652 33998
rect 10600 33934 10652 33940
rect 10612 32774 10640 33934
rect 10704 33386 10732 34682
rect 11256 33998 11284 34886
rect 11348 34746 11376 42638
rect 11716 40594 11744 45222
rect 11808 44878 11836 47200
rect 12544 44878 12572 47200
rect 11796 44872 11848 44878
rect 11796 44814 11848 44820
rect 12532 44872 12584 44878
rect 12532 44814 12584 44820
rect 12624 44532 12676 44538
rect 12624 44474 12676 44480
rect 12072 40928 12124 40934
rect 12072 40870 12124 40876
rect 11704 40588 11756 40594
rect 11704 40530 11756 40536
rect 12084 40050 12112 40870
rect 12636 40730 12664 44474
rect 13280 43790 13308 47200
rect 13452 45484 13504 45490
rect 13452 45426 13504 45432
rect 13820 45484 13872 45490
rect 13820 45426 13872 45432
rect 13464 44742 13492 45426
rect 13544 44872 13596 44878
rect 13544 44814 13596 44820
rect 13452 44736 13504 44742
rect 13452 44678 13504 44684
rect 13556 44305 13584 44814
rect 13542 44296 13598 44305
rect 13542 44231 13598 44240
rect 13832 43994 13860 45426
rect 13912 45076 13964 45082
rect 13912 45018 13964 45024
rect 13820 43988 13872 43994
rect 13820 43930 13872 43936
rect 13268 43784 13320 43790
rect 13268 43726 13320 43732
rect 13544 43784 13596 43790
rect 13544 43726 13596 43732
rect 13556 43450 13584 43726
rect 13544 43444 13596 43450
rect 13544 43386 13596 43392
rect 13924 41274 13952 45018
rect 14004 44396 14056 44402
rect 14004 44338 14056 44344
rect 14016 43897 14044 44338
rect 14002 43888 14058 43897
rect 14002 43823 14058 43832
rect 14108 43314 14136 47200
rect 14188 45824 14240 45830
rect 14188 45766 14240 45772
rect 14200 44402 14228 45766
rect 14280 45280 14332 45286
rect 14280 45222 14332 45228
rect 14464 45280 14516 45286
rect 14464 45222 14516 45228
rect 14292 44985 14320 45222
rect 14476 45014 14504 45222
rect 14740 45076 14792 45082
rect 14740 45018 14792 45024
rect 14372 45008 14424 45014
rect 14278 44976 14334 44985
rect 14372 44950 14424 44956
rect 14464 45008 14516 45014
rect 14464 44950 14516 44956
rect 14278 44911 14334 44920
rect 14188 44396 14240 44402
rect 14188 44338 14240 44344
rect 14188 44192 14240 44198
rect 14186 44160 14188 44169
rect 14240 44160 14242 44169
rect 14186 44095 14242 44104
rect 14188 43716 14240 43722
rect 14188 43658 14240 43664
rect 14200 43450 14228 43658
rect 14188 43444 14240 43450
rect 14188 43386 14240 43392
rect 14096 43308 14148 43314
rect 14096 43250 14148 43256
rect 14384 42226 14412 44950
rect 14752 44878 14780 45018
rect 14740 44872 14792 44878
rect 14646 44840 14702 44849
rect 14740 44814 14792 44820
rect 14646 44775 14648 44784
rect 14700 44775 14702 44784
rect 14648 44746 14700 44752
rect 14464 44736 14516 44742
rect 14464 44678 14516 44684
rect 14476 43858 14504 44678
rect 14740 44192 14792 44198
rect 14740 44134 14792 44140
rect 14464 43852 14516 43858
rect 14464 43794 14516 43800
rect 14464 43648 14516 43654
rect 14464 43590 14516 43596
rect 14556 43648 14608 43654
rect 14556 43590 14608 43596
rect 14476 42702 14504 43590
rect 14464 42696 14516 42702
rect 14464 42638 14516 42644
rect 14372 42220 14424 42226
rect 14372 42162 14424 42168
rect 14476 41682 14504 42638
rect 14464 41676 14516 41682
rect 14464 41618 14516 41624
rect 14280 41472 14332 41478
rect 14280 41414 14332 41420
rect 13912 41268 13964 41274
rect 13912 41210 13964 41216
rect 14188 40928 14240 40934
rect 14188 40870 14240 40876
rect 12624 40724 12676 40730
rect 12624 40666 12676 40672
rect 12072 40044 12124 40050
rect 12072 39986 12124 39992
rect 12256 40044 12308 40050
rect 12256 39986 12308 39992
rect 12072 39296 12124 39302
rect 12072 39238 12124 39244
rect 12084 38962 12112 39238
rect 12268 38962 12296 39986
rect 12072 38956 12124 38962
rect 12072 38898 12124 38904
rect 12256 38956 12308 38962
rect 12256 38898 12308 38904
rect 12164 37120 12216 37126
rect 12164 37062 12216 37068
rect 12072 36916 12124 36922
rect 12072 36858 12124 36864
rect 11796 36576 11848 36582
rect 11796 36518 11848 36524
rect 11612 36168 11664 36174
rect 11612 36110 11664 36116
rect 11336 34740 11388 34746
rect 11336 34682 11388 34688
rect 11520 34536 11572 34542
rect 11520 34478 11572 34484
rect 11532 34202 11560 34478
rect 11520 34196 11572 34202
rect 11520 34138 11572 34144
rect 11244 33992 11296 33998
rect 11244 33934 11296 33940
rect 11520 33856 11572 33862
rect 11520 33798 11572 33804
rect 10880 33756 11188 33776
rect 10880 33754 10886 33756
rect 10942 33754 10966 33756
rect 11022 33754 11046 33756
rect 11102 33754 11126 33756
rect 11182 33754 11188 33756
rect 10942 33702 10944 33754
rect 11124 33702 11126 33754
rect 10880 33700 10886 33702
rect 10942 33700 10966 33702
rect 11022 33700 11046 33702
rect 11102 33700 11126 33702
rect 11182 33700 11188 33702
rect 10880 33680 11188 33700
rect 11428 33652 11480 33658
rect 11428 33594 11480 33600
rect 10692 33380 10744 33386
rect 10692 33322 10744 33328
rect 10600 32768 10652 32774
rect 10600 32710 10652 32716
rect 10508 31680 10560 31686
rect 10508 31622 10560 31628
rect 10416 31476 10468 31482
rect 10416 31418 10468 31424
rect 10428 31346 10456 31418
rect 10416 31340 10468 31346
rect 10416 31282 10468 31288
rect 10428 30598 10456 31282
rect 10508 31204 10560 31210
rect 10508 31146 10560 31152
rect 10232 30592 10284 30598
rect 10232 30534 10284 30540
rect 10416 30592 10468 30598
rect 10416 30534 10468 30540
rect 10244 30258 10272 30534
rect 10324 30388 10376 30394
rect 10324 30330 10376 30336
rect 10336 30258 10364 30330
rect 10232 30252 10284 30258
rect 10232 30194 10284 30200
rect 10324 30252 10376 30258
rect 10324 30194 10376 30200
rect 10244 29714 10272 30194
rect 10232 29708 10284 29714
rect 10232 29650 10284 29656
rect 10230 29608 10286 29617
rect 10230 29543 10286 29552
rect 10140 29232 10192 29238
rect 10140 29174 10192 29180
rect 10048 28416 10100 28422
rect 10048 28358 10100 28364
rect 9956 28212 10008 28218
rect 9956 28154 10008 28160
rect 10244 28098 10272 29543
rect 10336 28762 10364 30194
rect 10324 28756 10376 28762
rect 10324 28698 10376 28704
rect 10060 28070 10272 28098
rect 9956 27600 10008 27606
rect 9956 27542 10008 27548
rect 9864 27396 9916 27402
rect 9864 27338 9916 27344
rect 9784 27254 9904 27282
rect 9680 26512 9732 26518
rect 9680 26454 9732 26460
rect 9496 25696 9548 25702
rect 9496 25638 9548 25644
rect 9312 25220 9364 25226
rect 9312 25162 9364 25168
rect 9220 24948 9272 24954
rect 9220 24890 9272 24896
rect 9324 24886 9352 25162
rect 8852 24880 8904 24886
rect 8852 24822 8904 24828
rect 9036 24880 9088 24886
rect 9036 24822 9088 24828
rect 9312 24880 9364 24886
rect 9312 24822 9364 24828
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8312 23322 8340 24346
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 8312 22778 8340 23122
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8312 22234 8340 22714
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 8404 20466 8432 22578
rect 8576 22500 8628 22506
rect 8576 22442 8628 22448
rect 8484 22432 8536 22438
rect 8484 22374 8536 22380
rect 8496 21622 8524 22374
rect 8588 22030 8616 22442
rect 8680 22030 8708 24754
rect 9048 24206 9076 24822
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 9140 24410 9168 24754
rect 9128 24404 9180 24410
rect 9128 24346 9180 24352
rect 9324 24290 9352 24822
rect 9324 24262 9444 24290
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 8852 24132 8904 24138
rect 8852 24074 8904 24080
rect 8864 23798 8892 24074
rect 8852 23792 8904 23798
rect 8852 23734 8904 23740
rect 8956 23118 8984 24142
rect 9048 23866 9076 24142
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 8944 22636 8996 22642
rect 9048 22624 9076 23802
rect 9232 23186 9260 24142
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 9416 23118 9444 24262
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 9508 22710 9536 25638
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 9588 24404 9640 24410
rect 9588 24346 9640 24352
rect 9496 22704 9548 22710
rect 9496 22646 9548 22652
rect 9128 22636 9180 22642
rect 9048 22596 9128 22624
rect 8944 22578 8996 22584
rect 9128 22578 9180 22584
rect 8956 22234 8984 22578
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 9600 22098 9628 24346
rect 9784 24206 9812 24754
rect 9876 24426 9904 27254
rect 9968 26994 9996 27542
rect 10060 27538 10088 28070
rect 10140 28008 10192 28014
rect 10140 27950 10192 27956
rect 10428 27962 10456 30534
rect 10520 30258 10548 31146
rect 10612 31142 10640 32710
rect 10704 32366 10732 33322
rect 11244 32904 11296 32910
rect 11244 32846 11296 32852
rect 10880 32668 11188 32688
rect 10880 32666 10886 32668
rect 10942 32666 10966 32668
rect 11022 32666 11046 32668
rect 11102 32666 11126 32668
rect 11182 32666 11188 32668
rect 10942 32614 10944 32666
rect 11124 32614 11126 32666
rect 10880 32612 10886 32614
rect 10942 32612 10966 32614
rect 11022 32612 11046 32614
rect 11102 32612 11126 32614
rect 11182 32612 11188 32614
rect 10880 32592 11188 32612
rect 10692 32360 10744 32366
rect 10692 32302 10744 32308
rect 10692 31884 10744 31890
rect 10692 31826 10744 31832
rect 10704 31482 10732 31826
rect 11256 31822 11284 32846
rect 11336 32836 11388 32842
rect 11336 32778 11388 32784
rect 10784 31816 10836 31822
rect 10784 31758 10836 31764
rect 11244 31816 11296 31822
rect 11244 31758 11296 31764
rect 10692 31476 10744 31482
rect 10692 31418 10744 31424
rect 10796 31278 10824 31758
rect 10880 31580 11188 31600
rect 10880 31578 10886 31580
rect 10942 31578 10966 31580
rect 11022 31578 11046 31580
rect 11102 31578 11126 31580
rect 11182 31578 11188 31580
rect 10942 31526 10944 31578
rect 11124 31526 11126 31578
rect 10880 31524 10886 31526
rect 10942 31524 10966 31526
rect 11022 31524 11046 31526
rect 11102 31524 11126 31526
rect 11182 31524 11188 31526
rect 10880 31504 11188 31524
rect 10784 31272 10836 31278
rect 10784 31214 10836 31220
rect 10600 31136 10652 31142
rect 10600 31078 10652 31084
rect 10612 30938 10640 31078
rect 10600 30932 10652 30938
rect 10600 30874 10652 30880
rect 10508 30252 10560 30258
rect 10508 30194 10560 30200
rect 10520 28082 10548 30194
rect 10612 30122 10640 30874
rect 10880 30492 11188 30512
rect 10880 30490 10886 30492
rect 10942 30490 10966 30492
rect 11022 30490 11046 30492
rect 11102 30490 11126 30492
rect 11182 30490 11188 30492
rect 10942 30438 10944 30490
rect 11124 30438 11126 30490
rect 10880 30436 10886 30438
rect 10942 30436 10966 30438
rect 11022 30436 11046 30438
rect 11102 30436 11126 30438
rect 11182 30436 11188 30438
rect 10880 30416 11188 30436
rect 11256 30394 11284 31758
rect 11348 31482 11376 32778
rect 11440 32774 11468 33594
rect 11532 33590 11560 33798
rect 11520 33584 11572 33590
rect 11520 33526 11572 33532
rect 11428 32768 11480 32774
rect 11428 32710 11480 32716
rect 11336 31476 11388 31482
rect 11336 31418 11388 31424
rect 11440 31362 11468 32710
rect 11520 32360 11572 32366
rect 11520 32302 11572 32308
rect 11348 31334 11468 31362
rect 11532 31346 11560 32302
rect 11520 31340 11572 31346
rect 11244 30388 11296 30394
rect 11244 30330 11296 30336
rect 10600 30116 10652 30122
rect 10600 30058 10652 30064
rect 10612 29646 10640 30058
rect 11348 29730 11376 31334
rect 11520 31282 11572 31288
rect 11428 31204 11480 31210
rect 11428 31146 11480 31152
rect 11440 30734 11468 31146
rect 11428 30728 11480 30734
rect 11428 30670 11480 30676
rect 11440 29782 11468 30670
rect 11520 29844 11572 29850
rect 11520 29786 11572 29792
rect 10692 29708 10744 29714
rect 10692 29650 10744 29656
rect 11256 29702 11376 29730
rect 11428 29776 11480 29782
rect 11428 29718 11480 29724
rect 10600 29640 10652 29646
rect 10600 29582 10652 29588
rect 10612 28966 10640 29582
rect 10704 29170 10732 29650
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10796 29170 10824 29446
rect 10880 29404 11188 29424
rect 10880 29402 10886 29404
rect 10942 29402 10966 29404
rect 11022 29402 11046 29404
rect 11102 29402 11126 29404
rect 11182 29402 11188 29404
rect 10942 29350 10944 29402
rect 11124 29350 11126 29402
rect 10880 29348 10886 29350
rect 10942 29348 10966 29350
rect 11022 29348 11046 29350
rect 11102 29348 11126 29350
rect 11182 29348 11188 29350
rect 10880 29328 11188 29348
rect 11256 29306 11284 29702
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 11244 29300 11296 29306
rect 11244 29242 11296 29248
rect 11150 29200 11206 29209
rect 10692 29164 10744 29170
rect 10692 29106 10744 29112
rect 10784 29164 10836 29170
rect 11150 29135 11206 29144
rect 10784 29106 10836 29112
rect 10600 28960 10652 28966
rect 10600 28902 10652 28908
rect 10612 28490 10640 28902
rect 10600 28484 10652 28490
rect 10600 28426 10652 28432
rect 10692 28416 10744 28422
rect 10612 28364 10692 28370
rect 10612 28358 10744 28364
rect 10612 28342 10732 28358
rect 10508 28076 10560 28082
rect 10508 28018 10560 28024
rect 10612 28014 10640 28342
rect 10600 28008 10652 28014
rect 10048 27532 10100 27538
rect 10048 27474 10100 27480
rect 10060 26994 10088 27474
rect 10152 27470 10180 27950
rect 10428 27934 10548 27962
rect 10600 27950 10652 27956
rect 10140 27464 10192 27470
rect 10140 27406 10192 27412
rect 10232 27396 10284 27402
rect 10284 27356 10364 27384
rect 10232 27338 10284 27344
rect 9956 26988 10008 26994
rect 9956 26930 10008 26936
rect 10048 26988 10100 26994
rect 10100 26948 10180 26976
rect 10048 26930 10100 26936
rect 9968 25158 9996 26930
rect 10048 25220 10100 25226
rect 10048 25162 10100 25168
rect 9956 25152 10008 25158
rect 9956 25094 10008 25100
rect 9968 24562 9996 25094
rect 10060 24886 10088 25162
rect 10048 24880 10100 24886
rect 10048 24822 10100 24828
rect 10060 24682 10088 24822
rect 10152 24721 10180 26948
rect 10232 26784 10284 26790
rect 10232 26726 10284 26732
rect 10138 24712 10194 24721
rect 10048 24676 10100 24682
rect 10138 24647 10194 24656
rect 10048 24618 10100 24624
rect 10140 24608 10192 24614
rect 9968 24534 10088 24562
rect 10140 24550 10192 24556
rect 9876 24398 9996 24426
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 9692 23322 9720 23666
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9678 23216 9734 23225
rect 9678 23151 9734 23160
rect 9692 22574 9720 23151
rect 9784 22778 9812 24142
rect 9864 24132 9916 24138
rect 9864 24074 9916 24080
rect 9876 23118 9904 24074
rect 9864 23112 9916 23118
rect 9968 23100 9996 24398
rect 10060 23225 10088 24534
rect 10046 23216 10102 23225
rect 10152 23186 10180 24550
rect 10046 23151 10102 23160
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 9968 23072 10088 23100
rect 9864 23054 9916 23060
rect 9876 22794 9904 23054
rect 9772 22772 9824 22778
rect 9876 22766 9996 22794
rect 9772 22714 9824 22720
rect 9784 22642 9812 22714
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 9968 22506 9996 22766
rect 9956 22500 10008 22506
rect 9956 22442 10008 22448
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 8576 22024 8628 22030
rect 8576 21966 8628 21972
rect 8668 22024 8720 22030
rect 8668 21966 8720 21972
rect 8680 21690 8708 21966
rect 8668 21684 8720 21690
rect 8668 21626 8720 21632
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 9128 20800 9180 20806
rect 9128 20742 9180 20748
rect 9140 20466 9168 20742
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9140 20330 9168 20402
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 9312 19780 9364 19786
rect 9312 19722 9364 19728
rect 9232 19514 9260 19722
rect 9220 19508 9272 19514
rect 9220 19450 9272 19456
rect 9324 18766 9352 19722
rect 9692 19378 9720 20538
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 5915 17980 6223 18000
rect 5915 17978 5921 17980
rect 5977 17978 6001 17980
rect 6057 17978 6081 17980
rect 6137 17978 6161 17980
rect 6217 17978 6223 17980
rect 5977 17926 5979 17978
rect 6159 17926 6161 17978
rect 5915 17924 5921 17926
rect 5977 17924 6001 17926
rect 6057 17924 6081 17926
rect 6137 17924 6161 17926
rect 6217 17924 6223 17926
rect 5915 17904 6223 17924
rect 8036 17882 8064 18226
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 8404 17202 8432 18022
rect 9324 17202 9352 18702
rect 9784 18154 9812 22170
rect 9876 22166 9904 22374
rect 9864 22160 9916 22166
rect 9864 22102 9916 22108
rect 9968 21418 9996 22442
rect 10060 22030 10088 23072
rect 10048 22024 10100 22030
rect 10100 21984 10180 22012
rect 10048 21966 10100 21972
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10060 21457 10088 21830
rect 10046 21448 10102 21457
rect 9956 21412 10008 21418
rect 10046 21383 10102 21392
rect 9956 21354 10008 21360
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9968 20534 9996 20878
rect 10152 20806 10180 21984
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 10140 20800 10192 20806
rect 10140 20742 10192 20748
rect 10060 20534 10088 20742
rect 9956 20528 10008 20534
rect 9876 20488 9956 20516
rect 9876 19378 9904 20488
rect 9956 20470 10008 20476
rect 10048 20528 10100 20534
rect 10100 20488 10180 20516
rect 10048 20470 10100 20476
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9968 18873 9996 20198
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10060 19378 10088 19654
rect 10152 19378 10180 20488
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10048 19236 10100 19242
rect 10048 19178 10100 19184
rect 9954 18864 10010 18873
rect 9954 18799 10010 18808
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9784 17626 9812 18090
rect 9692 17610 9812 17626
rect 9680 17604 9812 17610
rect 9732 17598 9812 17604
rect 9680 17546 9732 17552
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 5915 16892 6223 16912
rect 5915 16890 5921 16892
rect 5977 16890 6001 16892
rect 6057 16890 6081 16892
rect 6137 16890 6161 16892
rect 6217 16890 6223 16892
rect 5977 16838 5979 16890
rect 6159 16838 6161 16890
rect 5915 16836 5921 16838
rect 5977 16836 6001 16838
rect 6057 16836 6081 16838
rect 6137 16836 6161 16838
rect 6217 16836 6223 16838
rect 5915 16816 6223 16836
rect 5915 15804 6223 15824
rect 5915 15802 5921 15804
rect 5977 15802 6001 15804
rect 6057 15802 6081 15804
rect 6137 15802 6161 15804
rect 6217 15802 6223 15804
rect 5977 15750 5979 15802
rect 6159 15750 6161 15802
rect 5915 15748 5921 15750
rect 5977 15748 6001 15750
rect 6057 15748 6081 15750
rect 6137 15748 6161 15750
rect 6217 15748 6223 15750
rect 5915 15728 6223 15748
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 9324 14958 9352 17138
rect 9784 16998 9812 17478
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9876 16794 9904 16934
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9876 16590 9904 16730
rect 9968 16658 9996 18799
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9692 15178 9720 16526
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9508 15150 9720 15178
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 5915 14716 6223 14736
rect 5915 14714 5921 14716
rect 5977 14714 6001 14716
rect 6057 14714 6081 14716
rect 6137 14714 6161 14716
rect 6217 14714 6223 14716
rect 5977 14662 5979 14714
rect 6159 14662 6161 14714
rect 5915 14660 5921 14662
rect 5977 14660 6001 14662
rect 6057 14660 6081 14662
rect 6137 14660 6161 14662
rect 6217 14660 6223 14662
rect 5915 14640 6223 14660
rect 9324 14618 9352 14894
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9508 13938 9536 15150
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 5915 13628 6223 13648
rect 5915 13626 5921 13628
rect 5977 13626 6001 13628
rect 6057 13626 6081 13628
rect 6137 13626 6161 13628
rect 6217 13626 6223 13628
rect 5977 13574 5979 13626
rect 6159 13574 6161 13626
rect 5915 13572 5921 13574
rect 5977 13572 6001 13574
rect 6057 13572 6081 13574
rect 6137 13572 6161 13574
rect 6217 13572 6223 13574
rect 5915 13552 6223 13572
rect 5915 12540 6223 12560
rect 5915 12538 5921 12540
rect 5977 12538 6001 12540
rect 6057 12538 6081 12540
rect 6137 12538 6161 12540
rect 6217 12538 6223 12540
rect 5977 12486 5979 12538
rect 6159 12486 6161 12538
rect 5915 12484 5921 12486
rect 5977 12484 6001 12486
rect 6057 12484 6081 12486
rect 6137 12484 6161 12486
rect 6217 12484 6223 12486
rect 5915 12464 6223 12484
rect 5915 11452 6223 11472
rect 5915 11450 5921 11452
rect 5977 11450 6001 11452
rect 6057 11450 6081 11452
rect 6137 11450 6161 11452
rect 6217 11450 6223 11452
rect 5977 11398 5979 11450
rect 6159 11398 6161 11450
rect 5915 11396 5921 11398
rect 5977 11396 6001 11398
rect 6057 11396 6081 11398
rect 6137 11396 6161 11398
rect 6217 11396 6223 11398
rect 5915 11376 6223 11396
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2240 8974 2268 11018
rect 5915 10364 6223 10384
rect 5915 10362 5921 10364
rect 5977 10362 6001 10364
rect 6057 10362 6081 10364
rect 6137 10362 6161 10364
rect 6217 10362 6223 10364
rect 5977 10310 5979 10362
rect 6159 10310 6161 10362
rect 5915 10308 5921 10310
rect 5977 10308 6001 10310
rect 6057 10308 6081 10310
rect 6137 10308 6161 10310
rect 6217 10308 6223 10310
rect 5915 10288 6223 10308
rect 5915 9276 6223 9296
rect 5915 9274 5921 9276
rect 5977 9274 6001 9276
rect 6057 9274 6081 9276
rect 6137 9274 6161 9276
rect 6217 9274 6223 9276
rect 5977 9222 5979 9274
rect 6159 9222 6161 9274
rect 5915 9220 5921 9222
rect 5977 9220 6001 9222
rect 6057 9220 6081 9222
rect 6137 9220 6161 9222
rect 6217 9220 6223 9222
rect 5915 9200 6223 9220
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 5915 8188 6223 8208
rect 5915 8186 5921 8188
rect 5977 8186 6001 8188
rect 6057 8186 6081 8188
rect 6137 8186 6161 8188
rect 6217 8186 6223 8188
rect 5977 8134 5979 8186
rect 6159 8134 6161 8186
rect 5915 8132 5921 8134
rect 5977 8132 6001 8134
rect 6057 8132 6081 8134
rect 6137 8132 6161 8134
rect 6217 8132 6223 8134
rect 5915 8112 6223 8132
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 5915 7100 6223 7120
rect 5915 7098 5921 7100
rect 5977 7098 6001 7100
rect 6057 7098 6081 7100
rect 6137 7098 6161 7100
rect 6217 7098 6223 7100
rect 5977 7046 5979 7098
rect 6159 7046 6161 7098
rect 5915 7044 5921 7046
rect 5977 7044 6001 7046
rect 6057 7044 6081 7046
rect 6137 7044 6161 7046
rect 6217 7044 6223 7046
rect 5915 7024 6223 7044
rect 5915 6012 6223 6032
rect 5915 6010 5921 6012
rect 5977 6010 6001 6012
rect 6057 6010 6081 6012
rect 6137 6010 6161 6012
rect 6217 6010 6223 6012
rect 5977 5958 5979 6010
rect 6159 5958 6161 6010
rect 5915 5956 5921 5958
rect 5977 5956 6001 5958
rect 6057 5956 6081 5958
rect 6137 5956 6161 5958
rect 6217 5956 6223 5958
rect 5915 5936 6223 5956
rect 5915 4924 6223 4944
rect 5915 4922 5921 4924
rect 5977 4922 6001 4924
rect 6057 4922 6081 4924
rect 6137 4922 6161 4924
rect 6217 4922 6223 4924
rect 5977 4870 5979 4922
rect 6159 4870 6161 4922
rect 5915 4868 5921 4870
rect 5977 4868 6001 4870
rect 6057 4868 6081 4870
rect 6137 4868 6161 4870
rect 6217 4868 6223 4870
rect 5915 4848 6223 4868
rect 5915 3836 6223 3856
rect 5915 3834 5921 3836
rect 5977 3834 6001 3836
rect 6057 3834 6081 3836
rect 6137 3834 6161 3836
rect 6217 3834 6223 3836
rect 5977 3782 5979 3834
rect 6159 3782 6161 3834
rect 5915 3780 5921 3782
rect 5977 3780 6001 3782
rect 6057 3780 6081 3782
rect 6137 3780 6161 3782
rect 6217 3780 6223 3782
rect 5915 3760 6223 3780
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1582 2952 1638 2961
rect 1582 2887 1584 2896
rect 1636 2887 1638 2896
rect 1584 2858 1636 2864
rect 5915 2748 6223 2768
rect 5915 2746 5921 2748
rect 5977 2746 6001 2748
rect 6057 2746 6081 2748
rect 6137 2746 6161 2748
rect 6217 2746 6223 2748
rect 5977 2694 5979 2746
rect 6159 2694 6161 2746
rect 5915 2692 5921 2694
rect 5977 2692 6001 2694
rect 6057 2692 6081 2694
rect 6137 2692 6161 2694
rect 6217 2692 6223 2694
rect 5915 2672 6223 2692
rect 9508 2446 9536 13874
rect 9876 11830 9904 15438
rect 9968 15366 9996 16594
rect 10060 15502 10088 19178
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10152 16590 10180 18906
rect 10244 17678 10272 26726
rect 10336 25158 10364 27356
rect 10520 27334 10548 27934
rect 10508 27328 10560 27334
rect 10508 27270 10560 27276
rect 10520 27130 10548 27270
rect 10508 27124 10560 27130
rect 10508 27066 10560 27072
rect 10508 26920 10560 26926
rect 10612 26874 10640 27950
rect 10692 27328 10744 27334
rect 10796 27282 10824 29106
rect 11164 29102 11192 29135
rect 11152 29096 11204 29102
rect 11152 29038 11204 29044
rect 10880 28316 11188 28336
rect 10880 28314 10886 28316
rect 10942 28314 10966 28316
rect 11022 28314 11046 28316
rect 11102 28314 11126 28316
rect 11182 28314 11188 28316
rect 10942 28262 10944 28314
rect 11124 28262 11126 28314
rect 10880 28260 10886 28262
rect 10942 28260 10966 28262
rect 11022 28260 11046 28262
rect 11102 28260 11126 28262
rect 11182 28260 11188 28262
rect 10880 28240 11188 28260
rect 11256 28098 11284 29242
rect 11348 29102 11376 29582
rect 11428 29504 11480 29510
rect 11428 29446 11480 29452
rect 11336 29096 11388 29102
rect 11336 29038 11388 29044
rect 11348 28642 11376 29038
rect 11440 28762 11468 29446
rect 11532 29170 11560 29786
rect 11520 29164 11572 29170
rect 11520 29106 11572 29112
rect 11428 28756 11480 28762
rect 11428 28698 11480 28704
rect 11532 28694 11560 29106
rect 11520 28688 11572 28694
rect 11348 28614 11468 28642
rect 11520 28630 11572 28636
rect 11256 28070 11376 28098
rect 11244 27532 11296 27538
rect 11244 27474 11296 27480
rect 10744 27276 10824 27282
rect 10692 27270 10824 27276
rect 10704 27254 10824 27270
rect 10704 26994 10732 27254
rect 10880 27228 11188 27248
rect 10880 27226 10886 27228
rect 10942 27226 10966 27228
rect 11022 27226 11046 27228
rect 11102 27226 11126 27228
rect 11182 27226 11188 27228
rect 10942 27174 10944 27226
rect 11124 27174 11126 27226
rect 10880 27172 10886 27174
rect 10942 27172 10966 27174
rect 11022 27172 11046 27174
rect 11102 27172 11126 27174
rect 11182 27172 11188 27174
rect 10880 27152 11188 27172
rect 10692 26988 10744 26994
rect 10692 26930 10744 26936
rect 10784 26988 10836 26994
rect 10784 26930 10836 26936
rect 10796 26874 10824 26930
rect 10560 26868 10824 26874
rect 10508 26862 10824 26868
rect 10520 26846 10824 26862
rect 11256 26382 11284 27474
rect 11348 26586 11376 28070
rect 11440 27606 11468 28614
rect 11520 28416 11572 28422
rect 11520 28358 11572 28364
rect 11428 27600 11480 27606
rect 11428 27542 11480 27548
rect 11440 27402 11468 27542
rect 11428 27396 11480 27402
rect 11428 27338 11480 27344
rect 11336 26580 11388 26586
rect 11336 26522 11388 26528
rect 11244 26376 11296 26382
rect 11244 26318 11296 26324
rect 10508 26240 10560 26246
rect 10508 26182 10560 26188
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10336 23168 10364 25094
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 10428 23526 10456 24754
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10416 23180 10468 23186
rect 10336 23140 10416 23168
rect 10416 23122 10468 23128
rect 10324 23044 10376 23050
rect 10324 22986 10376 22992
rect 10336 21010 10364 22986
rect 10520 22094 10548 26182
rect 10880 26140 11188 26160
rect 10880 26138 10886 26140
rect 10942 26138 10966 26140
rect 11022 26138 11046 26140
rect 11102 26138 11126 26140
rect 11182 26138 11188 26140
rect 10942 26086 10944 26138
rect 11124 26086 11126 26138
rect 10880 26084 10886 26086
rect 10942 26084 10966 26086
rect 11022 26084 11046 26086
rect 11102 26084 11126 26086
rect 11182 26084 11188 26086
rect 10880 26064 11188 26084
rect 11152 25832 11204 25838
rect 11152 25774 11204 25780
rect 10600 25764 10652 25770
rect 10600 25706 10652 25712
rect 10612 25226 10640 25706
rect 10692 25356 10744 25362
rect 10692 25298 10744 25304
rect 10600 25220 10652 25226
rect 10600 25162 10652 25168
rect 10612 24818 10640 25162
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10598 24712 10654 24721
rect 10598 24647 10654 24656
rect 10612 23730 10640 24647
rect 10704 24206 10732 25298
rect 11164 25294 11192 25774
rect 11152 25288 11204 25294
rect 11204 25236 11284 25242
rect 11152 25230 11284 25236
rect 11164 25214 11284 25230
rect 10880 25052 11188 25072
rect 10880 25050 10886 25052
rect 10942 25050 10966 25052
rect 11022 25050 11046 25052
rect 11102 25050 11126 25052
rect 11182 25050 11188 25052
rect 10942 24998 10944 25050
rect 11124 24998 11126 25050
rect 10880 24996 10886 24998
rect 10942 24996 10966 24998
rect 11022 24996 11046 24998
rect 11102 24996 11126 24998
rect 11182 24996 11188 24998
rect 10880 24976 11188 24996
rect 11256 24886 11284 25214
rect 11244 24880 11296 24886
rect 11244 24822 11296 24828
rect 10784 24608 10836 24614
rect 10784 24550 10836 24556
rect 10692 24200 10744 24206
rect 10692 24142 10744 24148
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10428 22066 10548 22094
rect 10428 21554 10456 22066
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10428 20942 10456 21490
rect 10508 21140 10560 21146
rect 10508 21082 10560 21088
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 10324 20868 10376 20874
rect 10324 20810 10376 20816
rect 10336 20262 10364 20810
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10324 20256 10376 20262
rect 10324 20198 10376 20204
rect 10428 19334 10456 20742
rect 10520 20534 10548 21082
rect 10612 20942 10640 23122
rect 10704 22030 10732 24142
rect 10796 22234 10824 24550
rect 11334 24304 11390 24313
rect 11334 24239 11336 24248
rect 11388 24239 11390 24248
rect 11336 24210 11388 24216
rect 11244 24200 11296 24206
rect 11532 24154 11560 28358
rect 11244 24142 11296 24148
rect 10880 23964 11188 23984
rect 10880 23962 10886 23964
rect 10942 23962 10966 23964
rect 11022 23962 11046 23964
rect 11102 23962 11126 23964
rect 11182 23962 11188 23964
rect 10942 23910 10944 23962
rect 11124 23910 11126 23962
rect 10880 23908 10886 23910
rect 10942 23908 10966 23910
rect 11022 23908 11046 23910
rect 11102 23908 11126 23910
rect 11182 23908 11188 23910
rect 10880 23888 11188 23908
rect 11256 23769 11284 24142
rect 11440 24126 11560 24154
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11242 23760 11298 23769
rect 10968 23724 11020 23730
rect 11242 23695 11298 23704
rect 10968 23666 11020 23672
rect 10876 23588 10928 23594
rect 10876 23530 10928 23536
rect 10888 23118 10916 23530
rect 10980 23186 11008 23666
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 10880 22876 11188 22896
rect 10880 22874 10886 22876
rect 10942 22874 10966 22876
rect 11022 22874 11046 22876
rect 11102 22874 11126 22876
rect 11182 22874 11188 22876
rect 10942 22822 10944 22874
rect 11124 22822 11126 22874
rect 10880 22820 10886 22822
rect 10942 22820 10966 22822
rect 11022 22820 11046 22822
rect 11102 22820 11126 22822
rect 11182 22820 11188 22822
rect 10880 22800 11188 22820
rect 11256 22642 11284 23695
rect 11348 23118 11376 24006
rect 11440 23798 11468 24126
rect 11428 23792 11480 23798
rect 11428 23734 11480 23740
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 11348 22574 11376 23054
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 11334 22400 11390 22409
rect 11334 22335 11390 22344
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 11152 22024 11204 22030
rect 11204 21984 11284 22012
rect 11152 21966 11204 21972
rect 10704 21690 10732 21966
rect 10880 21788 11188 21808
rect 10880 21786 10886 21788
rect 10942 21786 10966 21788
rect 11022 21786 11046 21788
rect 11102 21786 11126 21788
rect 11182 21786 11188 21788
rect 10942 21734 10944 21786
rect 11124 21734 11126 21786
rect 10880 21732 10886 21734
rect 10942 21732 10966 21734
rect 11022 21732 11046 21734
rect 11102 21732 11126 21734
rect 11182 21732 11188 21734
rect 10880 21712 11188 21732
rect 11256 21690 11284 21984
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 10704 20942 10732 21626
rect 11058 21584 11114 21593
rect 11058 21519 11114 21528
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10980 20874 11008 21354
rect 11072 21078 11100 21519
rect 11060 21072 11112 21078
rect 11060 21014 11112 21020
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10508 20528 10560 20534
rect 10508 20470 10560 20476
rect 10336 19306 10456 19334
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9968 13802 9996 15302
rect 10152 14822 10180 16526
rect 10336 16046 10364 19306
rect 10520 18970 10548 20470
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10704 18426 10732 20742
rect 10880 20700 11188 20720
rect 10880 20698 10886 20700
rect 10942 20698 10966 20700
rect 11022 20698 11046 20700
rect 11102 20698 11126 20700
rect 11182 20698 11188 20700
rect 10942 20646 10944 20698
rect 11124 20646 11126 20698
rect 10880 20644 10886 20646
rect 10942 20644 10966 20646
rect 11022 20644 11046 20646
rect 11102 20644 11126 20646
rect 11182 20644 11188 20646
rect 10880 20624 11188 20644
rect 11256 20330 11284 21626
rect 11244 20324 11296 20330
rect 11244 20266 11296 20272
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10704 17626 10732 18362
rect 10796 18222 10824 19858
rect 10880 19612 11188 19632
rect 10880 19610 10886 19612
rect 10942 19610 10966 19612
rect 11022 19610 11046 19612
rect 11102 19610 11126 19612
rect 11182 19610 11188 19612
rect 10942 19558 10944 19610
rect 11124 19558 11126 19610
rect 10880 19556 10886 19558
rect 10942 19556 10966 19558
rect 11022 19556 11046 19558
rect 11102 19556 11126 19558
rect 11182 19556 11188 19558
rect 10880 19536 11188 19556
rect 10880 18524 11188 18544
rect 10880 18522 10886 18524
rect 10942 18522 10966 18524
rect 11022 18522 11046 18524
rect 11102 18522 11126 18524
rect 11182 18522 11188 18524
rect 10942 18470 10944 18522
rect 11124 18470 11126 18522
rect 10880 18468 10886 18470
rect 10942 18468 10966 18470
rect 11022 18468 11046 18470
rect 11102 18468 11126 18470
rect 11182 18468 11188 18470
rect 10880 18448 11188 18468
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10612 17610 10732 17626
rect 10600 17604 10732 17610
rect 10652 17598 10732 17604
rect 10600 17546 10652 17552
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10428 16794 10456 17070
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10520 16522 10548 16934
rect 10508 16516 10560 16522
rect 10508 16458 10560 16464
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11150 9628 11494
rect 9968 11218 9996 13126
rect 10060 12986 10088 13874
rect 10152 13870 10180 14758
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 10244 14074 10272 14282
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10152 12850 10180 13262
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10152 12442 10180 12786
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10428 11354 10456 12786
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10152 10810 10180 11086
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10520 10742 10548 15846
rect 10612 15638 10640 17546
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10600 15632 10652 15638
rect 10600 15574 10652 15580
rect 10704 15484 10732 16730
rect 10796 16658 10824 18158
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11348 17626 11376 22335
rect 11440 21554 11468 23734
rect 11624 22080 11652 36110
rect 11808 35766 11836 36518
rect 11980 36032 12032 36038
rect 11980 35974 12032 35980
rect 11796 35760 11848 35766
rect 11796 35702 11848 35708
rect 11888 33652 11940 33658
rect 11888 33594 11940 33600
rect 11704 32904 11756 32910
rect 11704 32846 11756 32852
rect 11716 32570 11744 32846
rect 11900 32774 11928 33594
rect 11888 32768 11940 32774
rect 11888 32710 11940 32716
rect 11704 32564 11756 32570
rect 11704 32506 11756 32512
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 11808 32026 11836 32370
rect 11796 32020 11848 32026
rect 11796 31962 11848 31968
rect 11900 31890 11928 32710
rect 11888 31884 11940 31890
rect 11888 31826 11940 31832
rect 11796 31816 11848 31822
rect 11796 31758 11848 31764
rect 11808 31346 11836 31758
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11796 31340 11848 31346
rect 11796 31282 11848 31288
rect 11716 28422 11744 31282
rect 11900 31278 11928 31826
rect 11888 31272 11940 31278
rect 11888 31214 11940 31220
rect 11888 31136 11940 31142
rect 11888 31078 11940 31084
rect 11796 30592 11848 30598
rect 11796 30534 11848 30540
rect 11808 29170 11836 30534
rect 11900 30258 11928 31078
rect 11992 30870 12020 35974
rect 12084 35698 12112 36858
rect 12176 36718 12204 37062
rect 12164 36712 12216 36718
rect 12164 36654 12216 36660
rect 12176 36038 12204 36654
rect 12164 36032 12216 36038
rect 12164 35974 12216 35980
rect 12268 35698 12296 38898
rect 12636 37398 12664 40666
rect 14096 38888 14148 38894
rect 14096 38830 14148 38836
rect 14108 38350 14136 38830
rect 14096 38344 14148 38350
rect 14096 38286 14148 38292
rect 14108 37942 14136 38286
rect 14096 37936 14148 37942
rect 14096 37878 14148 37884
rect 13084 37868 13136 37874
rect 13084 37810 13136 37816
rect 13096 37466 13124 37810
rect 13636 37664 13688 37670
rect 13636 37606 13688 37612
rect 13084 37460 13136 37466
rect 13084 37402 13136 37408
rect 12624 37392 12676 37398
rect 12624 37334 12676 37340
rect 13268 37324 13320 37330
rect 13268 37266 13320 37272
rect 12900 37256 12952 37262
rect 12900 37198 12952 37204
rect 12532 37188 12584 37194
rect 12584 37148 12664 37176
rect 12532 37130 12584 37136
rect 12636 36718 12664 37148
rect 12624 36712 12676 36718
rect 12624 36654 12676 36660
rect 12636 36174 12664 36654
rect 12624 36168 12676 36174
rect 12624 36110 12676 36116
rect 12912 36106 12940 37198
rect 13176 36780 13228 36786
rect 13176 36722 13228 36728
rect 12900 36100 12952 36106
rect 12900 36042 12952 36048
rect 12072 35692 12124 35698
rect 12072 35634 12124 35640
rect 12256 35692 12308 35698
rect 12256 35634 12308 35640
rect 12268 35086 12296 35634
rect 12256 35080 12308 35086
rect 12256 35022 12308 35028
rect 12164 34604 12216 34610
rect 12164 34546 12216 34552
rect 12072 33516 12124 33522
rect 12072 33458 12124 33464
rect 12084 32910 12112 33458
rect 12072 32904 12124 32910
rect 12072 32846 12124 32852
rect 11980 30864 12032 30870
rect 11980 30806 12032 30812
rect 11980 30728 12032 30734
rect 11980 30670 12032 30676
rect 11888 30252 11940 30258
rect 11888 30194 11940 30200
rect 11992 30138 12020 30670
rect 12072 30660 12124 30666
rect 12072 30602 12124 30608
rect 12084 30258 12112 30602
rect 12176 30326 12204 34546
rect 12268 34134 12296 35022
rect 13188 35018 13216 36722
rect 13280 36378 13308 37266
rect 13648 37262 13676 37606
rect 13636 37256 13688 37262
rect 13636 37198 13688 37204
rect 13268 36372 13320 36378
rect 13268 36314 13320 36320
rect 13280 36174 13308 36314
rect 13820 36304 13872 36310
rect 13820 36246 13872 36252
rect 13268 36168 13320 36174
rect 13268 36110 13320 36116
rect 13544 36168 13596 36174
rect 13544 36110 13596 36116
rect 13268 36032 13320 36038
rect 13268 35974 13320 35980
rect 13280 35630 13308 35974
rect 13556 35698 13584 36110
rect 13544 35692 13596 35698
rect 13544 35634 13596 35640
rect 13268 35624 13320 35630
rect 13268 35566 13320 35572
rect 13176 35012 13228 35018
rect 13176 34954 13228 34960
rect 12900 34400 12952 34406
rect 12900 34342 12952 34348
rect 12256 34128 12308 34134
rect 12256 34070 12308 34076
rect 12268 33998 12296 34070
rect 12256 33992 12308 33998
rect 12256 33934 12308 33940
rect 12716 33924 12768 33930
rect 12716 33866 12768 33872
rect 12728 33658 12756 33866
rect 12716 33652 12768 33658
rect 12716 33594 12768 33600
rect 12728 33318 12756 33594
rect 12256 33312 12308 33318
rect 12256 33254 12308 33260
rect 12716 33312 12768 33318
rect 12716 33254 12768 33260
rect 12268 30734 12296 33254
rect 12808 32768 12860 32774
rect 12808 32710 12860 32716
rect 12820 32434 12848 32710
rect 12348 32428 12400 32434
rect 12348 32370 12400 32376
rect 12440 32428 12492 32434
rect 12440 32370 12492 32376
rect 12808 32428 12860 32434
rect 12808 32370 12860 32376
rect 12360 32026 12388 32370
rect 12348 32020 12400 32026
rect 12348 31962 12400 31968
rect 12452 31414 12480 32370
rect 12624 32292 12676 32298
rect 12624 32234 12676 32240
rect 12636 31890 12664 32234
rect 12624 31884 12676 31890
rect 12624 31826 12676 31832
rect 12532 31748 12584 31754
rect 12532 31690 12584 31696
rect 12440 31408 12492 31414
rect 12440 31350 12492 31356
rect 12348 30864 12400 30870
rect 12348 30806 12400 30812
rect 12256 30728 12308 30734
rect 12256 30670 12308 30676
rect 12164 30320 12216 30326
rect 12164 30262 12216 30268
rect 12072 30252 12124 30258
rect 12072 30194 12124 30200
rect 11900 30110 12020 30138
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11900 29102 11928 30110
rect 11980 30048 12032 30054
rect 11980 29990 12032 29996
rect 11992 29578 12020 29990
rect 12072 29640 12124 29646
rect 12072 29582 12124 29588
rect 11980 29572 12032 29578
rect 11980 29514 12032 29520
rect 11888 29096 11940 29102
rect 11888 29038 11940 29044
rect 11796 29028 11848 29034
rect 11796 28970 11848 28976
rect 11808 28558 11836 28970
rect 11796 28552 11848 28558
rect 11796 28494 11848 28500
rect 11900 28506 11928 29038
rect 11992 29034 12020 29514
rect 12084 29170 12112 29582
rect 12256 29300 12308 29306
rect 12256 29242 12308 29248
rect 12072 29164 12124 29170
rect 12072 29106 12124 29112
rect 11980 29028 12032 29034
rect 11980 28970 12032 28976
rect 12268 28762 12296 29242
rect 12256 28756 12308 28762
rect 12256 28698 12308 28704
rect 12164 28552 12216 28558
rect 11900 28500 12164 28506
rect 11900 28494 12216 28500
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 11808 27878 11836 28494
rect 11900 28478 12204 28494
rect 11900 28150 11928 28478
rect 12256 28416 12308 28422
rect 12256 28358 12308 28364
rect 11888 28144 11940 28150
rect 11888 28086 11940 28092
rect 11796 27872 11848 27878
rect 11796 27814 11848 27820
rect 11900 27606 11928 28086
rect 12072 27668 12124 27674
rect 12072 27610 12124 27616
rect 11888 27600 11940 27606
rect 11888 27542 11940 27548
rect 12084 27334 12112 27610
rect 12268 27538 12296 28358
rect 12256 27532 12308 27538
rect 12256 27474 12308 27480
rect 12072 27328 12124 27334
rect 12072 27270 12124 27276
rect 11980 25832 12032 25838
rect 11980 25774 12032 25780
rect 11992 25226 12020 25774
rect 11980 25220 12032 25226
rect 11980 25162 12032 25168
rect 11992 24954 12020 25162
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 11888 24880 11940 24886
rect 11888 24822 11940 24828
rect 11796 24608 11848 24614
rect 11796 24550 11848 24556
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11716 23798 11744 24006
rect 11704 23792 11756 23798
rect 11704 23734 11756 23740
rect 11808 22624 11836 24550
rect 11900 24274 11928 24822
rect 11888 24268 11940 24274
rect 11888 24210 11940 24216
rect 11900 23322 11928 24210
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 11992 23526 12020 24142
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 11888 23316 11940 23322
rect 11888 23258 11940 23264
rect 11992 22778 12020 23462
rect 12084 23050 12112 27270
rect 12164 26376 12216 26382
rect 12164 26318 12216 26324
rect 12176 25242 12204 26318
rect 12176 25214 12296 25242
rect 12164 24608 12216 24614
rect 12164 24550 12216 24556
rect 12176 24410 12204 24550
rect 12164 24404 12216 24410
rect 12164 24346 12216 24352
rect 12072 23044 12124 23050
rect 12072 22986 12124 22992
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11888 22636 11940 22642
rect 11808 22596 11888 22624
rect 11888 22578 11940 22584
rect 11624 22052 11836 22080
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11428 21548 11480 21554
rect 11428 21490 11480 21496
rect 11428 21344 11480 21350
rect 11426 21312 11428 21321
rect 11480 21312 11482 21321
rect 11426 21247 11482 21256
rect 11440 17746 11468 21247
rect 11532 21185 11560 21830
rect 11716 21418 11744 21830
rect 11704 21412 11756 21418
rect 11704 21354 11756 21360
rect 11518 21176 11574 21185
rect 11518 21111 11574 21120
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11624 20534 11652 20878
rect 11808 20534 11836 22052
rect 11612 20528 11664 20534
rect 11612 20470 11664 20476
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 11624 18766 11652 19110
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11532 17678 11560 18022
rect 11520 17672 11572 17678
rect 10880 17436 11188 17456
rect 10880 17434 10886 17436
rect 10942 17434 10966 17436
rect 11022 17434 11046 17436
rect 11102 17434 11126 17436
rect 11182 17434 11188 17436
rect 10942 17382 10944 17434
rect 11124 17382 11126 17434
rect 10880 17380 10886 17382
rect 10942 17380 10966 17382
rect 11022 17380 11046 17382
rect 11102 17380 11126 17382
rect 11182 17380 11188 17382
rect 10880 17360 11188 17380
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 11256 16590 11284 17614
rect 11348 17598 11468 17626
rect 11520 17614 11572 17620
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11348 16658 11376 17478
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11440 16436 11468 17598
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11256 16408 11468 16436
rect 10880 16348 11188 16368
rect 10880 16346 10886 16348
rect 10942 16346 10966 16348
rect 11022 16346 11046 16348
rect 11102 16346 11126 16348
rect 11182 16346 11188 16348
rect 10942 16294 10944 16346
rect 11124 16294 11126 16346
rect 10880 16292 10886 16294
rect 10942 16292 10966 16294
rect 11022 16292 11046 16294
rect 11102 16292 11126 16294
rect 11182 16292 11188 16294
rect 10880 16272 11188 16292
rect 10612 15456 10732 15484
rect 10612 12918 10640 15456
rect 10880 15260 11188 15280
rect 10880 15258 10886 15260
rect 10942 15258 10966 15260
rect 11022 15258 11046 15260
rect 11102 15258 11126 15260
rect 11182 15258 11188 15260
rect 10942 15206 10944 15258
rect 11124 15206 11126 15258
rect 10880 15204 10886 15206
rect 10942 15204 10966 15206
rect 11022 15204 11046 15206
rect 11102 15204 11126 15206
rect 11182 15204 11188 15206
rect 10880 15184 11188 15204
rect 10880 14172 11188 14192
rect 10880 14170 10886 14172
rect 10942 14170 10966 14172
rect 11022 14170 11046 14172
rect 11102 14170 11126 14172
rect 11182 14170 11188 14172
rect 10942 14118 10944 14170
rect 11124 14118 11126 14170
rect 10880 14116 10886 14118
rect 10942 14116 10966 14118
rect 11022 14116 11046 14118
rect 11102 14116 11126 14118
rect 11182 14116 11188 14118
rect 10880 14096 11188 14116
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10612 11082 10640 12310
rect 10704 12238 10732 13330
rect 10796 13326 10824 13806
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10796 12306 10824 13262
rect 10880 13084 11188 13104
rect 10880 13082 10886 13084
rect 10942 13082 10966 13084
rect 11022 13082 11046 13084
rect 11102 13082 11126 13084
rect 11182 13082 11188 13084
rect 10942 13030 10944 13082
rect 11124 13030 11126 13082
rect 10880 13028 10886 13030
rect 10942 13028 10966 13030
rect 11022 13028 11046 13030
rect 11102 13028 11126 13030
rect 11182 13028 11188 13030
rect 10880 13008 11188 13028
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11234 10732 12174
rect 10880 11996 11188 12016
rect 10880 11994 10886 11996
rect 10942 11994 10966 11996
rect 11022 11994 11046 11996
rect 11102 11994 11126 11996
rect 11182 11994 11188 11996
rect 10942 11942 10944 11994
rect 11124 11942 11126 11994
rect 10880 11940 10886 11942
rect 10942 11940 10966 11942
rect 11022 11940 11046 11942
rect 11102 11940 11126 11942
rect 11182 11940 11188 11942
rect 10880 11920 11188 11940
rect 10704 11206 10824 11234
rect 11256 11218 11284 16408
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11348 12238 11376 16186
rect 11532 15706 11560 17478
rect 11624 16998 11652 18702
rect 11716 18578 11744 20266
rect 11808 18970 11836 20470
rect 11900 19310 11928 22578
rect 12176 22506 12204 24346
rect 12164 22500 12216 22506
rect 12164 22442 12216 22448
rect 12268 22094 12296 25214
rect 12360 22409 12388 30806
rect 12440 30660 12492 30666
rect 12440 30602 12492 30608
rect 12452 29238 12480 30602
rect 12440 29232 12492 29238
rect 12440 29174 12492 29180
rect 12452 28490 12480 29174
rect 12440 28484 12492 28490
rect 12440 28426 12492 28432
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12452 25770 12480 26930
rect 12440 25764 12492 25770
rect 12440 25706 12492 25712
rect 12440 24200 12492 24206
rect 12544 24188 12572 31690
rect 12636 30326 12664 31826
rect 12820 31482 12848 32370
rect 12808 31476 12860 31482
rect 12808 31418 12860 31424
rect 12912 31346 12940 34342
rect 13188 34202 13216 34954
rect 13556 34610 13584 35634
rect 13544 34604 13596 34610
rect 13544 34546 13596 34552
rect 13176 34196 13228 34202
rect 13176 34138 13228 34144
rect 13360 33380 13412 33386
rect 13360 33322 13412 33328
rect 13268 33312 13320 33318
rect 13268 33254 13320 33260
rect 13280 32910 13308 33254
rect 13268 32904 13320 32910
rect 13268 32846 13320 32852
rect 12992 32836 13044 32842
rect 12992 32778 13044 32784
rect 13004 32570 13032 32778
rect 12992 32564 13044 32570
rect 12992 32506 13044 32512
rect 13372 32434 13400 33322
rect 13452 32496 13504 32502
rect 13452 32438 13504 32444
rect 13360 32428 13412 32434
rect 13360 32370 13412 32376
rect 13464 32230 13492 32438
rect 13452 32224 13504 32230
rect 13452 32166 13504 32172
rect 13464 31414 13492 32166
rect 13452 31408 13504 31414
rect 13452 31350 13504 31356
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 13084 31272 13136 31278
rect 13084 31214 13136 31220
rect 12716 30796 12768 30802
rect 12716 30738 12768 30744
rect 12728 30394 12756 30738
rect 13096 30734 13124 31214
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 12992 30592 13044 30598
rect 12992 30534 13044 30540
rect 12716 30388 12768 30394
rect 12716 30330 12768 30336
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12624 30320 12676 30326
rect 12624 30262 12676 30268
rect 12716 30116 12768 30122
rect 12716 30058 12768 30064
rect 12624 29164 12676 29170
rect 12624 29106 12676 29112
rect 12636 27402 12664 29106
rect 12624 27396 12676 27402
rect 12624 27338 12676 27344
rect 12636 26858 12664 27338
rect 12624 26852 12676 26858
rect 12624 26794 12676 26800
rect 12728 25838 12756 30058
rect 12820 29782 12848 30330
rect 12808 29776 12860 29782
rect 12808 29718 12860 29724
rect 13004 29646 13032 30534
rect 13268 30184 13320 30190
rect 13268 30126 13320 30132
rect 12992 29640 13044 29646
rect 12992 29582 13044 29588
rect 13176 29640 13228 29646
rect 13176 29582 13228 29588
rect 12806 29336 12862 29345
rect 13188 29306 13216 29582
rect 13280 29481 13308 30126
rect 13266 29472 13322 29481
rect 13266 29407 13322 29416
rect 12806 29271 12862 29280
rect 13176 29300 13228 29306
rect 12820 29034 12848 29271
rect 13176 29242 13228 29248
rect 12898 29200 12954 29209
rect 12898 29135 12954 29144
rect 12808 29028 12860 29034
rect 12808 28970 12860 28976
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12820 26586 12848 26930
rect 12808 26580 12860 26586
rect 12808 26522 12860 26528
rect 12912 26466 12940 29135
rect 13280 29102 13308 29407
rect 13268 29096 13320 29102
rect 13268 29038 13320 29044
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 12992 27464 13044 27470
rect 12992 27406 13044 27412
rect 13004 27130 13032 27406
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 12992 27124 13044 27130
rect 12992 27066 13044 27072
rect 13096 26926 13124 27270
rect 13280 27130 13308 28018
rect 13268 27124 13320 27130
rect 13268 27066 13320 27072
rect 13268 26988 13320 26994
rect 13268 26930 13320 26936
rect 13084 26920 13136 26926
rect 13084 26862 13136 26868
rect 13280 26466 13308 26930
rect 12820 26438 13308 26466
rect 12716 25832 12768 25838
rect 12716 25774 12768 25780
rect 12492 24160 12572 24188
rect 12716 24200 12768 24206
rect 12440 24142 12492 24148
rect 12716 24142 12768 24148
rect 12452 23662 12480 24142
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12452 23118 12480 23598
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12532 22432 12584 22438
rect 12346 22400 12402 22409
rect 12532 22374 12584 22380
rect 12346 22335 12402 22344
rect 12544 22234 12572 22374
rect 12532 22228 12584 22234
rect 12532 22170 12584 22176
rect 12176 22066 12296 22094
rect 12438 22128 12494 22137
rect 12176 21690 12204 22066
rect 12438 22063 12494 22072
rect 12452 22030 12480 22063
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12072 21480 12124 21486
rect 12256 21480 12308 21486
rect 12254 21448 12256 21457
rect 12308 21448 12310 21457
rect 12124 21428 12204 21434
rect 12072 21422 12204 21428
rect 12084 21406 12204 21422
rect 12176 21146 12204 21406
rect 12254 21383 12310 21392
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12452 20924 12480 21966
rect 12544 21842 12572 22170
rect 12636 22030 12664 23258
rect 12728 23186 12756 24142
rect 12716 23180 12768 23186
rect 12716 23122 12768 23128
rect 12728 22642 12756 23122
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12544 21814 12664 21842
rect 12530 21176 12586 21185
rect 12530 21111 12586 21120
rect 12544 21078 12572 21111
rect 12532 21072 12584 21078
rect 12532 21014 12584 21020
rect 11992 20896 12480 20924
rect 11888 19304 11940 19310
rect 11888 19246 11940 19252
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 18970 11928 19110
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11808 18748 11836 18906
rect 11888 18760 11940 18766
rect 11808 18720 11888 18748
rect 11888 18702 11940 18708
rect 11716 18550 11836 18578
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11716 17338 11744 18226
rect 11808 18086 11836 18550
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11428 15496 11480 15502
rect 11624 15484 11652 16662
rect 11716 16114 11744 17274
rect 11808 17270 11836 17682
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11808 16794 11836 17206
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11900 16658 11928 17682
rect 11888 16652 11940 16658
rect 11808 16612 11888 16640
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11716 15502 11744 15914
rect 11480 15456 11652 15484
rect 11704 15496 11756 15502
rect 11428 15438 11480 15444
rect 11704 15438 11756 15444
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11440 14890 11468 15302
rect 11808 15042 11836 16612
rect 11888 16594 11940 16600
rect 11992 16250 12020 20896
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12176 20058 12204 20402
rect 12348 20324 12400 20330
rect 12348 20266 12400 20272
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11532 15014 11836 15042
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11440 14414 11468 14554
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11440 13530 11468 14350
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11428 12912 11480 12918
rect 11428 12854 11480 12860
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11440 11762 11468 12854
rect 11532 12782 11560 15014
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11624 14414 11652 14894
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11624 13870 11652 14350
rect 11796 14340 11848 14346
rect 11796 14282 11848 14288
rect 11808 13938 11836 14282
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11612 13864 11664 13870
rect 11664 13824 11744 13852
rect 11612 13806 11664 13812
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11624 13190 11652 13466
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11716 12850 11744 13824
rect 11808 13326 11836 13874
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11532 12306 11560 12718
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10508 10736 10560 10742
rect 10508 10678 10560 10684
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10520 9586 10548 9998
rect 10612 9722 10640 10610
rect 10704 10266 10732 11086
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10796 10146 10824 11206
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11808 11150 11836 13126
rect 11900 12374 11928 15982
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11992 15502 12020 15642
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 12084 15178 12112 19654
rect 11992 15150 12112 15178
rect 11992 13462 12020 15150
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11992 13326 12020 13398
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 12084 12442 12112 14962
rect 12176 14618 12204 19994
rect 12360 19854 12388 20266
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12254 18864 12310 18873
rect 12254 18799 12310 18808
rect 12268 18766 12296 18799
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12268 18426 12296 18566
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12176 13938 12204 14554
rect 12268 14498 12296 18022
rect 12360 14618 12388 19790
rect 12452 19786 12480 20470
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12636 19718 12664 21814
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12728 20942 12756 21286
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12820 20618 12848 26438
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 13004 25974 13032 26318
rect 12992 25968 13044 25974
rect 12992 25910 13044 25916
rect 13084 25900 13136 25906
rect 13084 25842 13136 25848
rect 12900 25764 12952 25770
rect 12900 25706 12952 25712
rect 12912 23202 12940 25706
rect 13096 25498 13124 25842
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 13096 25294 13124 25434
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 13084 25152 13136 25158
rect 13084 25094 13136 25100
rect 13096 24818 13124 25094
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13096 24206 13124 24754
rect 13188 24682 13216 26318
rect 13360 26308 13412 26314
rect 13360 26250 13412 26256
rect 13372 25906 13400 26250
rect 13360 25900 13412 25906
rect 13360 25842 13412 25848
rect 13358 25800 13414 25809
rect 13268 25764 13320 25770
rect 13358 25735 13414 25744
rect 13268 25706 13320 25712
rect 13280 24954 13308 25706
rect 13372 25129 13400 25735
rect 13358 25120 13414 25129
rect 13358 25055 13414 25064
rect 13268 24948 13320 24954
rect 13268 24890 13320 24896
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 13188 24410 13216 24618
rect 13176 24404 13228 24410
rect 13176 24346 13228 24352
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 12992 23656 13044 23662
rect 12992 23598 13044 23604
rect 13004 23322 13032 23598
rect 13084 23520 13136 23526
rect 13084 23462 13136 23468
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 12912 23174 13032 23202
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 12912 20874 12940 23054
rect 13004 22166 13032 23174
rect 13096 22438 13124 23462
rect 13188 23118 13216 24346
rect 13280 23202 13308 24890
rect 13372 23730 13400 25055
rect 13464 24614 13492 31350
rect 13636 30184 13688 30190
rect 13636 30126 13688 30132
rect 13544 30048 13596 30054
rect 13544 29990 13596 29996
rect 13556 29578 13584 29990
rect 13544 29572 13596 29578
rect 13544 29514 13596 29520
rect 13556 25242 13584 29514
rect 13648 29102 13676 30126
rect 13636 29096 13688 29102
rect 13636 29038 13688 29044
rect 13648 25344 13676 29038
rect 13832 26874 13860 36246
rect 13912 36100 13964 36106
rect 13912 36042 13964 36048
rect 13924 35494 13952 36042
rect 13912 35488 13964 35494
rect 13912 35430 13964 35436
rect 13924 28558 13952 35430
rect 14004 33652 14056 33658
rect 14004 33594 14056 33600
rect 14016 32502 14044 33594
rect 14200 32994 14228 40870
rect 14292 34610 14320 41414
rect 14372 41268 14424 41274
rect 14372 41210 14424 41216
rect 14384 40050 14412 41210
rect 14476 41002 14504 41618
rect 14464 40996 14516 41002
rect 14464 40938 14516 40944
rect 14568 40882 14596 43590
rect 14648 42560 14700 42566
rect 14648 42502 14700 42508
rect 14660 41614 14688 42502
rect 14648 41608 14700 41614
rect 14648 41550 14700 41556
rect 14648 41132 14700 41138
rect 14648 41074 14700 41080
rect 14476 40854 14596 40882
rect 14372 40044 14424 40050
rect 14372 39986 14424 39992
rect 14476 35630 14504 40854
rect 14556 40588 14608 40594
rect 14556 40530 14608 40536
rect 14568 40118 14596 40530
rect 14660 40186 14688 41074
rect 14648 40180 14700 40186
rect 14648 40122 14700 40128
rect 14556 40112 14608 40118
rect 14556 40054 14608 40060
rect 14752 37194 14780 44134
rect 14844 43382 14872 47200
rect 15580 45830 15608 47200
rect 15568 45824 15620 45830
rect 15568 45766 15620 45772
rect 16408 45558 16436 47200
rect 16672 45620 16724 45626
rect 16724 45580 16896 45608
rect 16672 45562 16724 45568
rect 16396 45552 16448 45558
rect 16396 45494 16448 45500
rect 15292 45484 15344 45490
rect 15292 45426 15344 45432
rect 15198 45384 15254 45393
rect 14936 45342 15198 45370
rect 14936 44878 14964 45342
rect 15198 45319 15254 45328
rect 15212 45286 15240 45319
rect 15108 45280 15160 45286
rect 15108 45222 15160 45228
rect 15200 45280 15252 45286
rect 15200 45222 15252 45228
rect 15016 45076 15068 45082
rect 15016 45018 15068 45024
rect 14924 44872 14976 44878
rect 14924 44814 14976 44820
rect 14924 44736 14976 44742
rect 14924 44678 14976 44684
rect 14936 44470 14964 44678
rect 14924 44464 14976 44470
rect 14924 44406 14976 44412
rect 15028 44334 15056 45018
rect 15016 44328 15068 44334
rect 15016 44270 15068 44276
rect 15028 44010 15056 44270
rect 14936 43982 15056 44010
rect 14936 43722 14964 43982
rect 15016 43852 15068 43858
rect 15016 43794 15068 43800
rect 14924 43716 14976 43722
rect 14924 43658 14976 43664
rect 14832 43376 14884 43382
rect 14832 43318 14884 43324
rect 15028 43110 15056 43794
rect 15120 43450 15148 45222
rect 15304 44810 15332 45426
rect 16672 45416 16724 45422
rect 16672 45358 16724 45364
rect 16580 45348 16632 45354
rect 16580 45290 16632 45296
rect 15660 45280 15712 45286
rect 15660 45222 15712 45228
rect 15292 44804 15344 44810
rect 15292 44746 15344 44752
rect 15200 44328 15252 44334
rect 15200 44270 15252 44276
rect 15212 43858 15240 44270
rect 15304 44169 15332 44746
rect 15672 44538 15700 45222
rect 15846 45180 16154 45200
rect 15846 45178 15852 45180
rect 15908 45178 15932 45180
rect 15988 45178 16012 45180
rect 16068 45178 16092 45180
rect 16148 45178 16154 45180
rect 15908 45126 15910 45178
rect 16090 45126 16092 45178
rect 15846 45124 15852 45126
rect 15908 45124 15932 45126
rect 15988 45124 16012 45126
rect 16068 45124 16092 45126
rect 16148 45124 16154 45126
rect 15846 45104 16154 45124
rect 16592 45082 16620 45290
rect 16580 45076 16632 45082
rect 16580 45018 16632 45024
rect 16212 44940 16264 44946
rect 16212 44882 16264 44888
rect 15752 44872 15804 44878
rect 15752 44814 15804 44820
rect 15660 44532 15712 44538
rect 15660 44474 15712 44480
rect 15290 44160 15346 44169
rect 15290 44095 15346 44104
rect 15200 43852 15252 43858
rect 15200 43794 15252 43800
rect 15108 43444 15160 43450
rect 15108 43386 15160 43392
rect 15212 43246 15240 43794
rect 15304 43450 15332 44095
rect 15764 43790 15792 44814
rect 15846 44092 16154 44112
rect 15846 44090 15852 44092
rect 15908 44090 15932 44092
rect 15988 44090 16012 44092
rect 16068 44090 16092 44092
rect 16148 44090 16154 44092
rect 15908 44038 15910 44090
rect 16090 44038 16092 44090
rect 15846 44036 15852 44038
rect 15908 44036 15932 44038
rect 15988 44036 16012 44038
rect 16068 44036 16092 44038
rect 16148 44036 16154 44038
rect 15846 44016 16154 44036
rect 16224 43858 16252 44882
rect 16684 44742 16712 45358
rect 16868 44878 16896 45580
rect 16948 45484 17000 45490
rect 16948 45426 17000 45432
rect 16960 45082 16988 45426
rect 17038 45384 17094 45393
rect 17038 45319 17094 45328
rect 17052 45286 17080 45319
rect 17040 45280 17092 45286
rect 17040 45222 17092 45228
rect 16948 45076 17000 45082
rect 16948 45018 17000 45024
rect 16856 44872 16908 44878
rect 16856 44814 16908 44820
rect 16672 44736 16724 44742
rect 16672 44678 16724 44684
rect 16396 44396 16448 44402
rect 16396 44338 16448 44344
rect 16488 44396 16540 44402
rect 16488 44338 16540 44344
rect 16304 44192 16356 44198
rect 16304 44134 16356 44140
rect 16212 43852 16264 43858
rect 16212 43794 16264 43800
rect 15752 43784 15804 43790
rect 15752 43726 15804 43732
rect 15476 43716 15528 43722
rect 15476 43658 15528 43664
rect 15384 43648 15436 43654
rect 15384 43590 15436 43596
rect 15292 43444 15344 43450
rect 15292 43386 15344 43392
rect 15200 43240 15252 43246
rect 15252 43188 15332 43194
rect 15200 43182 15332 43188
rect 15212 43166 15332 43182
rect 14924 43104 14976 43110
rect 14924 43046 14976 43052
rect 15016 43104 15068 43110
rect 15016 43046 15068 43052
rect 14832 42016 14884 42022
rect 14832 41958 14884 41964
rect 14844 40526 14872 41958
rect 14832 40520 14884 40526
rect 14832 40462 14884 40468
rect 14936 37874 14964 43046
rect 15108 42696 15160 42702
rect 15108 42638 15160 42644
rect 15016 42220 15068 42226
rect 15016 42162 15068 42168
rect 15028 41138 15056 42162
rect 15120 42158 15148 42638
rect 15200 42628 15252 42634
rect 15200 42570 15252 42576
rect 15212 42226 15240 42570
rect 15200 42220 15252 42226
rect 15200 42162 15252 42168
rect 15108 42152 15160 42158
rect 15108 42094 15160 42100
rect 15016 41132 15068 41138
rect 15016 41074 15068 41080
rect 15028 40662 15056 41074
rect 15016 40656 15068 40662
rect 15016 40598 15068 40604
rect 15120 40050 15148 42094
rect 15108 40044 15160 40050
rect 15108 39986 15160 39992
rect 15212 39982 15240 42162
rect 15304 41682 15332 43166
rect 15292 41676 15344 41682
rect 15292 41618 15344 41624
rect 15304 41070 15332 41618
rect 15292 41064 15344 41070
rect 15292 41006 15344 41012
rect 15304 40594 15332 41006
rect 15292 40588 15344 40594
rect 15292 40530 15344 40536
rect 15292 40384 15344 40390
rect 15292 40326 15344 40332
rect 15200 39976 15252 39982
rect 15200 39918 15252 39924
rect 15200 38412 15252 38418
rect 15200 38354 15252 38360
rect 15108 37936 15160 37942
rect 15212 37890 15240 38354
rect 15160 37884 15240 37890
rect 15108 37878 15240 37884
rect 14924 37868 14976 37874
rect 15120 37862 15240 37878
rect 14924 37810 14976 37816
rect 15108 37460 15160 37466
rect 15108 37402 15160 37408
rect 15016 37256 15068 37262
rect 15016 37198 15068 37204
rect 14740 37188 14792 37194
rect 14740 37130 14792 37136
rect 14464 35624 14516 35630
rect 14464 35566 14516 35572
rect 14464 35488 14516 35494
rect 14464 35430 14516 35436
rect 14476 35290 14504 35430
rect 14464 35284 14516 35290
rect 14464 35226 14516 35232
rect 14924 34944 14976 34950
rect 14924 34886 14976 34892
rect 14280 34604 14332 34610
rect 14280 34546 14332 34552
rect 14556 33652 14608 33658
rect 14556 33594 14608 33600
rect 14464 33380 14516 33386
rect 14464 33322 14516 33328
rect 14200 32966 14320 32994
rect 14188 32904 14240 32910
rect 14188 32846 14240 32852
rect 14004 32496 14056 32502
rect 14004 32438 14056 32444
rect 14016 30802 14044 32438
rect 14004 30796 14056 30802
rect 14004 30738 14056 30744
rect 14200 30258 14228 32846
rect 14292 32366 14320 32966
rect 14476 32434 14504 33322
rect 14464 32428 14516 32434
rect 14464 32370 14516 32376
rect 14280 32360 14332 32366
rect 14280 32302 14332 32308
rect 14568 32298 14596 33594
rect 14556 32292 14608 32298
rect 14556 32234 14608 32240
rect 14372 30728 14424 30734
rect 14372 30670 14424 30676
rect 14188 30252 14240 30258
rect 14188 30194 14240 30200
rect 14096 29504 14148 29510
rect 14096 29446 14148 29452
rect 14108 28694 14136 29446
rect 14200 29238 14228 30194
rect 14384 29850 14412 30670
rect 14372 29844 14424 29850
rect 14372 29786 14424 29792
rect 14188 29232 14240 29238
rect 14188 29174 14240 29180
rect 14096 28688 14148 28694
rect 14096 28630 14148 28636
rect 13912 28552 13964 28558
rect 13912 28494 13964 28500
rect 13832 26846 14044 26874
rect 13728 26784 13780 26790
rect 13728 26726 13780 26732
rect 13912 26784 13964 26790
rect 13912 26726 13964 26732
rect 13740 26314 13768 26726
rect 13924 26518 13952 26726
rect 13912 26512 13964 26518
rect 13912 26454 13964 26460
rect 13820 26444 13872 26450
rect 13820 26386 13872 26392
rect 13728 26308 13780 26314
rect 13728 26250 13780 26256
rect 13832 26042 13860 26386
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13728 25900 13780 25906
rect 13728 25842 13780 25848
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13740 25498 13768 25842
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13832 25362 13860 25842
rect 13924 25770 13952 26454
rect 14016 25809 14044 26846
rect 14002 25800 14058 25809
rect 13912 25764 13964 25770
rect 14002 25735 14058 25744
rect 13912 25706 13964 25712
rect 13924 25430 13952 25706
rect 14004 25696 14056 25702
rect 14004 25638 14056 25644
rect 13912 25424 13964 25430
rect 13912 25366 13964 25372
rect 13820 25356 13872 25362
rect 13648 25316 13768 25344
rect 13556 25214 13676 25242
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13360 23724 13412 23730
rect 13412 23684 13492 23712
rect 13360 23666 13412 23672
rect 13280 23174 13400 23202
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13268 23044 13320 23050
rect 13268 22986 13320 22992
rect 13280 22778 13308 22986
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 12992 22160 13044 22166
rect 12992 22102 13044 22108
rect 13004 21622 13032 22102
rect 12992 21616 13044 21622
rect 12992 21558 13044 21564
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 13004 21321 13032 21354
rect 12990 21312 13046 21321
rect 12990 21247 13046 21256
rect 13096 21162 13124 22374
rect 13372 22094 13400 23174
rect 13004 21134 13124 21162
rect 13280 22066 13400 22094
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12728 20602 12848 20618
rect 12716 20596 12848 20602
rect 12768 20590 12848 20596
rect 12716 20538 12768 20544
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12544 19174 12572 19450
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12452 17338 12480 18022
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12544 17218 12572 19110
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12728 17882 12756 18702
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12452 17190 12572 17218
rect 12452 16658 12480 17190
rect 12624 17128 12676 17134
rect 12544 17088 12624 17116
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12544 16538 12572 17088
rect 12624 17070 12676 17076
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12728 16726 12756 17002
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12452 16510 12572 16538
rect 12452 16454 12480 16510
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 15638 12480 16390
rect 12532 15972 12584 15978
rect 12532 15914 12584 15920
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12268 14470 12388 14498
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12268 13326 12296 13670
rect 12360 13530 12388 14470
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11900 11354 11928 12038
rect 12084 11898 12112 12038
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12176 11762 12204 12582
rect 12268 12306 12296 13262
rect 12360 12646 12388 13330
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12360 12238 12388 12378
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12544 11354 12572 15914
rect 12636 14482 12664 16594
rect 13004 15910 13032 21134
rect 13084 19780 13136 19786
rect 13084 19722 13136 19728
rect 13096 19378 13124 19722
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 13096 18834 13124 19314
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 13084 18352 13136 18358
rect 13082 18320 13084 18329
rect 13136 18320 13138 18329
rect 13188 18290 13216 19110
rect 13082 18255 13138 18264
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 13280 15722 13308 22066
rect 13464 21690 13492 23684
rect 13544 23520 13596 23526
rect 13544 23462 13596 23468
rect 13556 23050 13584 23462
rect 13544 23044 13596 23050
rect 13544 22986 13596 22992
rect 13556 22642 13584 22986
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13464 21146 13492 21626
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13452 20868 13504 20874
rect 13452 20810 13504 20816
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13372 18902 13400 19790
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13372 18766 13400 18838
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13358 17776 13414 17785
rect 13358 17711 13360 17720
rect 13412 17711 13414 17720
rect 13360 17682 13412 17688
rect 13464 17678 13492 20810
rect 13556 20058 13584 22578
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13556 19514 13584 19994
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13464 16794 13492 17138
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13188 15694 13308 15722
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 12820 14618 12848 15438
rect 13004 15162 13032 15438
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 13188 15094 13216 15694
rect 13372 15638 13400 15982
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 13280 15026 13308 15574
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12636 13258 12664 14418
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12728 11898 12756 12786
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 10880 10908 11188 10928
rect 10880 10906 10886 10908
rect 10942 10906 10966 10908
rect 11022 10906 11046 10908
rect 11102 10906 11126 10908
rect 11182 10906 11188 10908
rect 10942 10854 10944 10906
rect 11124 10854 11126 10906
rect 10880 10852 10886 10854
rect 10942 10852 10966 10854
rect 11022 10852 11046 10854
rect 11102 10852 11126 10854
rect 11182 10852 11188 10854
rect 10880 10832 11188 10852
rect 11532 10810 11560 11086
rect 12084 10810 12112 11086
rect 12728 10810 12756 11834
rect 13096 11762 13124 12038
rect 13372 11898 13400 15438
rect 13556 14958 13584 18090
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13556 14414 13584 14894
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12452 10266 12480 10610
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 10692 10124 10744 10130
rect 10796 10118 10916 10146
rect 10692 10066 10744 10072
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10704 9654 10732 10066
rect 10888 10062 10916 10118
rect 12728 10062 12756 10746
rect 13004 10606 13032 11154
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10796 9178 10824 9930
rect 10880 9820 11188 9840
rect 10880 9818 10886 9820
rect 10942 9818 10966 9820
rect 11022 9818 11046 9820
rect 11102 9818 11126 9820
rect 11182 9818 11188 9820
rect 10942 9766 10944 9818
rect 11124 9766 11126 9818
rect 10880 9764 10886 9766
rect 10942 9764 10966 9766
rect 11022 9764 11046 9766
rect 11102 9764 11126 9766
rect 11182 9764 11188 9766
rect 10880 9744 11188 9764
rect 12820 9722 12848 10542
rect 13004 10266 13032 10542
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13004 10130 13032 10202
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12176 9178 12204 9522
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 10796 8634 10824 8774
rect 10880 8732 11188 8752
rect 10880 8730 10886 8732
rect 10942 8730 10966 8732
rect 11022 8730 11046 8732
rect 11102 8730 11126 8732
rect 11182 8730 11188 8732
rect 10942 8678 10944 8730
rect 11124 8678 11126 8730
rect 10880 8676 10886 8678
rect 10942 8676 10966 8678
rect 11022 8676 11046 8678
rect 11102 8676 11126 8678
rect 11182 8676 11188 8678
rect 10880 8656 11188 8676
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 11440 8498 11468 8774
rect 11716 8566 11744 8910
rect 12728 8906 12756 9454
rect 13280 9042 13308 9454
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 10880 7644 11188 7664
rect 10880 7642 10886 7644
rect 10942 7642 10966 7644
rect 11022 7642 11046 7644
rect 11102 7642 11126 7644
rect 11182 7642 11188 7644
rect 10942 7590 10944 7642
rect 11124 7590 11126 7642
rect 10880 7588 10886 7590
rect 10942 7588 10966 7590
rect 11022 7588 11046 7590
rect 11102 7588 11126 7590
rect 11182 7588 11188 7590
rect 10880 7568 11188 7588
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10612 5846 10640 6802
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10612 5710 10640 5782
rect 10796 5778 10824 6734
rect 10880 6556 11188 6576
rect 10880 6554 10886 6556
rect 10942 6554 10966 6556
rect 11022 6554 11046 6556
rect 11102 6554 11126 6556
rect 11182 6554 11188 6556
rect 10942 6502 10944 6554
rect 11124 6502 11126 6554
rect 10880 6500 10886 6502
rect 10942 6500 10966 6502
rect 11022 6500 11046 6502
rect 11102 6500 11126 6502
rect 11182 6500 11188 6502
rect 10880 6480 11188 6500
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 11256 5778 11284 6122
rect 11716 5930 11744 6734
rect 11992 6458 12020 8434
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12452 7868 12480 8298
rect 12544 8090 12572 8434
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12532 7880 12584 7886
rect 12452 7840 12532 7868
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12360 7410 12388 7686
rect 12452 7410 12480 7840
rect 12532 7822 12584 7828
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11624 5902 11744 5930
rect 11624 5778 11652 5902
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10880 5468 11188 5488
rect 10880 5466 10886 5468
rect 10942 5466 10966 5468
rect 11022 5466 11046 5468
rect 11102 5466 11126 5468
rect 11182 5466 11188 5468
rect 10942 5414 10944 5466
rect 11124 5414 11126 5466
rect 10880 5412 10886 5414
rect 10942 5412 10966 5414
rect 11022 5412 11046 5414
rect 11102 5412 11126 5414
rect 11182 5412 11188 5414
rect 10880 5392 11188 5412
rect 11532 4758 11560 5714
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 10880 4380 11188 4400
rect 10880 4378 10886 4380
rect 10942 4378 10966 4380
rect 11022 4378 11046 4380
rect 11102 4378 11126 4380
rect 11182 4378 11188 4380
rect 10942 4326 10944 4378
rect 11124 4326 11126 4378
rect 10880 4324 10886 4326
rect 10942 4324 10966 4326
rect 11022 4324 11046 4326
rect 11102 4324 11126 4326
rect 11182 4324 11188 4326
rect 10880 4304 11188 4324
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10520 3738 10548 4082
rect 11624 3942 11652 5714
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 11164 3602 11192 3878
rect 11624 3670 11652 3878
rect 11808 3670 11836 6122
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11900 5370 11928 5510
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11164 3482 11192 3538
rect 11164 3454 11284 3482
rect 10880 3292 11188 3312
rect 10880 3290 10886 3292
rect 10942 3290 10966 3292
rect 11022 3290 11046 3292
rect 11102 3290 11126 3292
rect 11182 3290 11188 3292
rect 10942 3238 10944 3290
rect 11124 3238 11126 3290
rect 10880 3236 10886 3238
rect 10942 3236 10966 3238
rect 11022 3236 11046 3238
rect 11102 3236 11126 3238
rect 11182 3236 11188 3238
rect 10880 3216 11188 3236
rect 11256 3058 11284 3454
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11624 2990 11652 3606
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 12176 2922 12204 6938
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12360 5778 12388 6802
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12452 6458 12480 6598
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12452 5914 12480 6258
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12256 4004 12308 4010
rect 12256 3946 12308 3952
rect 12268 3602 12296 3946
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12360 3534 12388 5714
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12452 3738 12480 5034
rect 12728 4826 12756 8842
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12820 6186 12848 7754
rect 12912 6798 12940 7890
rect 13648 7818 13676 25214
rect 13740 24886 13768 25316
rect 13820 25298 13872 25304
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13728 24880 13780 24886
rect 13728 24822 13780 24828
rect 13924 24274 13952 25230
rect 14016 25226 14044 25638
rect 14004 25220 14056 25226
rect 14004 25162 14056 25168
rect 14108 25106 14136 28630
rect 14200 28082 14228 29174
rect 14188 28076 14240 28082
rect 14188 28018 14240 28024
rect 14200 25294 14228 28018
rect 14280 27872 14332 27878
rect 14280 27814 14332 27820
rect 14292 27606 14320 27814
rect 14280 27600 14332 27606
rect 14280 27542 14332 27548
rect 14292 26994 14320 27542
rect 14372 27532 14424 27538
rect 14372 27474 14424 27480
rect 14280 26988 14332 26994
rect 14280 26930 14332 26936
rect 14280 26444 14332 26450
rect 14280 26386 14332 26392
rect 14188 25288 14240 25294
rect 14188 25230 14240 25236
rect 14016 25078 14136 25106
rect 13912 24268 13964 24274
rect 13912 24210 13964 24216
rect 13820 21956 13872 21962
rect 13820 21898 13872 21904
rect 13832 21554 13860 21898
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13740 19258 13768 21014
rect 13832 20602 13860 21490
rect 13912 20868 13964 20874
rect 13912 20810 13964 20816
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13820 20460 13872 20466
rect 13924 20448 13952 20810
rect 13872 20420 13952 20448
rect 13820 20402 13872 20408
rect 13832 19922 13860 20402
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13832 19360 13860 19858
rect 13912 19372 13964 19378
rect 13832 19332 13912 19360
rect 13912 19314 13964 19320
rect 13740 19230 13952 19258
rect 13820 19168 13872 19174
rect 13818 19136 13820 19145
rect 13872 19136 13874 19145
rect 13818 19071 13874 19080
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13740 17338 13768 17478
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13728 16176 13780 16182
rect 13728 16118 13780 16124
rect 13740 16046 13768 16118
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13740 15162 13768 15982
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13740 14414 13768 14962
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 12102 13768 14350
rect 13832 12986 13860 16050
rect 13924 15570 13952 19230
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13924 14890 13952 15506
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13924 12170 13952 13262
rect 14016 12170 14044 25078
rect 14292 24154 14320 26386
rect 14200 24126 14320 24154
rect 14096 23248 14148 23254
rect 14094 23216 14096 23225
rect 14148 23216 14150 23225
rect 14094 23151 14150 23160
rect 14200 21962 14228 24126
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 14188 21956 14240 21962
rect 14188 21898 14240 21904
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14108 20058 14136 20538
rect 14200 20466 14228 21082
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 14108 18766 14136 19858
rect 14200 19786 14228 20402
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14200 19378 14228 19450
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14188 18896 14240 18902
rect 14188 18838 14240 18844
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14108 16658 14136 18702
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14108 15502 14136 16390
rect 14200 16266 14228 18838
rect 14292 18714 14320 23802
rect 14384 23186 14412 27474
rect 14464 27396 14516 27402
rect 14464 27338 14516 27344
rect 14476 27062 14504 27338
rect 14464 27056 14516 27062
rect 14464 26998 14516 27004
rect 14568 26234 14596 32234
rect 14740 30252 14792 30258
rect 14740 30194 14792 30200
rect 14752 29850 14780 30194
rect 14740 29844 14792 29850
rect 14740 29786 14792 29792
rect 14936 29578 14964 34886
rect 15028 34610 15056 37198
rect 15016 34604 15068 34610
rect 15016 34546 15068 34552
rect 15028 33522 15056 34546
rect 15120 33998 15148 37402
rect 15212 37330 15240 37862
rect 15200 37324 15252 37330
rect 15200 37266 15252 37272
rect 15212 36786 15240 37266
rect 15200 36780 15252 36786
rect 15200 36722 15252 36728
rect 15200 36032 15252 36038
rect 15200 35974 15252 35980
rect 15212 35086 15240 35974
rect 15200 35080 15252 35086
rect 15200 35022 15252 35028
rect 15108 33992 15160 33998
rect 15108 33934 15160 33940
rect 15304 33590 15332 40326
rect 15396 39438 15424 43590
rect 15488 42770 15516 43658
rect 15476 42764 15528 42770
rect 15476 42706 15528 42712
rect 15764 42702 15792 43726
rect 16212 43648 16264 43654
rect 16212 43590 16264 43596
rect 15846 43004 16154 43024
rect 15846 43002 15852 43004
rect 15908 43002 15932 43004
rect 15988 43002 16012 43004
rect 16068 43002 16092 43004
rect 16148 43002 16154 43004
rect 15908 42950 15910 43002
rect 16090 42950 16092 43002
rect 15846 42948 15852 42950
rect 15908 42948 15932 42950
rect 15988 42948 16012 42950
rect 16068 42948 16092 42950
rect 16148 42948 16154 42950
rect 15846 42928 16154 42948
rect 16224 42906 16252 43590
rect 16212 42900 16264 42906
rect 16212 42842 16264 42848
rect 15752 42696 15804 42702
rect 15752 42638 15804 42644
rect 15846 41916 16154 41936
rect 15846 41914 15852 41916
rect 15908 41914 15932 41916
rect 15988 41914 16012 41916
rect 16068 41914 16092 41916
rect 16148 41914 16154 41916
rect 15908 41862 15910 41914
rect 16090 41862 16092 41914
rect 15846 41860 15852 41862
rect 15908 41860 15932 41862
rect 15988 41860 16012 41862
rect 16068 41860 16092 41862
rect 16148 41860 16154 41862
rect 15846 41840 16154 41860
rect 15568 41472 15620 41478
rect 15568 41414 15620 41420
rect 15384 39432 15436 39438
rect 15384 39374 15436 39380
rect 15476 39432 15528 39438
rect 15476 39374 15528 39380
rect 15488 38418 15516 39374
rect 15476 38412 15528 38418
rect 15476 38354 15528 38360
rect 15384 38276 15436 38282
rect 15384 38218 15436 38224
rect 15396 37806 15424 38218
rect 15384 37800 15436 37806
rect 15384 37742 15436 37748
rect 15384 37256 15436 37262
rect 15384 37198 15436 37204
rect 15396 36938 15424 37198
rect 15396 36910 15516 36938
rect 15384 36780 15436 36786
rect 15384 36722 15436 36728
rect 15396 35698 15424 36722
rect 15384 35692 15436 35698
rect 15384 35634 15436 35640
rect 15488 35630 15516 36910
rect 15476 35624 15528 35630
rect 15476 35566 15528 35572
rect 15384 35080 15436 35086
rect 15384 35022 15436 35028
rect 15396 34066 15424 35022
rect 15488 34474 15516 35566
rect 15476 34468 15528 34474
rect 15476 34410 15528 34416
rect 15384 34060 15436 34066
rect 15384 34002 15436 34008
rect 15108 33584 15160 33590
rect 15108 33526 15160 33532
rect 15292 33584 15344 33590
rect 15292 33526 15344 33532
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 15016 32768 15068 32774
rect 15016 32710 15068 32716
rect 15028 32434 15056 32710
rect 15120 32570 15148 33526
rect 15488 33522 15516 34410
rect 15580 33538 15608 41414
rect 15846 40828 16154 40848
rect 15846 40826 15852 40828
rect 15908 40826 15932 40828
rect 15988 40826 16012 40828
rect 16068 40826 16092 40828
rect 16148 40826 16154 40828
rect 15908 40774 15910 40826
rect 16090 40774 16092 40826
rect 15846 40772 15852 40774
rect 15908 40772 15932 40774
rect 15988 40772 16012 40774
rect 16068 40772 16092 40774
rect 16148 40772 16154 40774
rect 15846 40752 16154 40772
rect 15846 39740 16154 39760
rect 15846 39738 15852 39740
rect 15908 39738 15932 39740
rect 15988 39738 16012 39740
rect 16068 39738 16092 39740
rect 16148 39738 16154 39740
rect 15908 39686 15910 39738
rect 16090 39686 16092 39738
rect 15846 39684 15852 39686
rect 15908 39684 15932 39686
rect 15988 39684 16012 39686
rect 16068 39684 16092 39686
rect 16148 39684 16154 39686
rect 15846 39664 16154 39684
rect 15660 39432 15712 39438
rect 15660 39374 15712 39380
rect 16028 39432 16080 39438
rect 16028 39374 16080 39380
rect 15672 38486 15700 39374
rect 15936 39296 15988 39302
rect 15936 39238 15988 39244
rect 15752 39092 15804 39098
rect 15752 39034 15804 39040
rect 15660 38480 15712 38486
rect 15660 38422 15712 38428
rect 15672 38010 15700 38422
rect 15660 38004 15712 38010
rect 15660 37946 15712 37952
rect 15764 37874 15792 39034
rect 15948 38962 15976 39238
rect 16040 39098 16068 39374
rect 16028 39092 16080 39098
rect 16028 39034 16080 39040
rect 15936 38956 15988 38962
rect 15936 38898 15988 38904
rect 15846 38652 16154 38672
rect 15846 38650 15852 38652
rect 15908 38650 15932 38652
rect 15988 38650 16012 38652
rect 16068 38650 16092 38652
rect 16148 38650 16154 38652
rect 15908 38598 15910 38650
rect 16090 38598 16092 38650
rect 15846 38596 15852 38598
rect 15908 38596 15932 38598
rect 15988 38596 16012 38598
rect 16068 38596 16092 38598
rect 16148 38596 16154 38598
rect 15846 38576 16154 38596
rect 16316 38350 16344 44134
rect 16408 43654 16436 44338
rect 16500 43874 16528 44338
rect 16764 44328 16816 44334
rect 16764 44270 16816 44276
rect 16500 43858 16620 43874
rect 16500 43852 16632 43858
rect 16500 43846 16580 43852
rect 16580 43794 16632 43800
rect 16488 43784 16540 43790
rect 16488 43726 16540 43732
rect 16396 43648 16448 43654
rect 16396 43590 16448 43596
rect 16500 42702 16528 43726
rect 16776 43450 16804 44270
rect 16764 43444 16816 43450
rect 16764 43386 16816 43392
rect 16488 42696 16540 42702
rect 16488 42638 16540 42644
rect 16488 41676 16540 41682
rect 16488 41618 16540 41624
rect 16396 40928 16448 40934
rect 16396 40870 16448 40876
rect 16304 38344 16356 38350
rect 16304 38286 16356 38292
rect 16028 38208 16080 38214
rect 16028 38150 16080 38156
rect 16040 37874 16068 38150
rect 15752 37868 15804 37874
rect 15752 37810 15804 37816
rect 16028 37868 16080 37874
rect 16028 37810 16080 37816
rect 15846 37564 16154 37584
rect 15846 37562 15852 37564
rect 15908 37562 15932 37564
rect 15988 37562 16012 37564
rect 16068 37562 16092 37564
rect 16148 37562 16154 37564
rect 15908 37510 15910 37562
rect 16090 37510 16092 37562
rect 15846 37508 15852 37510
rect 15908 37508 15932 37510
rect 15988 37508 16012 37510
rect 16068 37508 16092 37510
rect 16148 37508 16154 37510
rect 15846 37488 16154 37508
rect 15660 37324 15712 37330
rect 15660 37266 15712 37272
rect 15672 35018 15700 37266
rect 15846 36476 16154 36496
rect 15846 36474 15852 36476
rect 15908 36474 15932 36476
rect 15988 36474 16012 36476
rect 16068 36474 16092 36476
rect 16148 36474 16154 36476
rect 15908 36422 15910 36474
rect 16090 36422 16092 36474
rect 15846 36420 15852 36422
rect 15908 36420 15932 36422
rect 15988 36420 16012 36422
rect 16068 36420 16092 36422
rect 16148 36420 16154 36422
rect 15846 36400 16154 36420
rect 15844 36100 15896 36106
rect 15844 36042 15896 36048
rect 15752 36032 15804 36038
rect 15752 35974 15804 35980
rect 15764 35766 15792 35974
rect 15752 35760 15804 35766
rect 15752 35702 15804 35708
rect 15856 35630 15884 36042
rect 15844 35624 15896 35630
rect 15844 35566 15896 35572
rect 15846 35388 16154 35408
rect 15846 35386 15852 35388
rect 15908 35386 15932 35388
rect 15988 35386 16012 35388
rect 16068 35386 16092 35388
rect 16148 35386 16154 35388
rect 15908 35334 15910 35386
rect 16090 35334 16092 35386
rect 15846 35332 15852 35334
rect 15908 35332 15932 35334
rect 15988 35332 16012 35334
rect 16068 35332 16092 35334
rect 16148 35332 16154 35334
rect 15846 35312 16154 35332
rect 15660 35012 15712 35018
rect 15660 34954 15712 34960
rect 16212 34536 16264 34542
rect 16212 34478 16264 34484
rect 15846 34300 16154 34320
rect 15846 34298 15852 34300
rect 15908 34298 15932 34300
rect 15988 34298 16012 34300
rect 16068 34298 16092 34300
rect 16148 34298 16154 34300
rect 15908 34246 15910 34298
rect 16090 34246 16092 34298
rect 15846 34244 15852 34246
rect 15908 34244 15932 34246
rect 15988 34244 16012 34246
rect 16068 34244 16092 34246
rect 16148 34244 16154 34246
rect 15846 34224 16154 34244
rect 15844 33924 15896 33930
rect 15844 33866 15896 33872
rect 15476 33516 15528 33522
rect 15580 33510 15792 33538
rect 15856 33522 15884 33866
rect 15476 33458 15528 33464
rect 15292 33448 15344 33454
rect 15292 33390 15344 33396
rect 15304 33318 15332 33390
rect 15292 33312 15344 33318
rect 15292 33254 15344 33260
rect 15200 32836 15252 32842
rect 15200 32778 15252 32784
rect 15108 32564 15160 32570
rect 15108 32506 15160 32512
rect 15212 32434 15240 32778
rect 15016 32428 15068 32434
rect 15016 32370 15068 32376
rect 15200 32428 15252 32434
rect 15200 32370 15252 32376
rect 15028 31822 15056 32370
rect 15304 32298 15332 33254
rect 15488 32366 15516 33458
rect 15476 32360 15528 32366
rect 15476 32302 15528 32308
rect 15292 32292 15344 32298
rect 15292 32234 15344 32240
rect 15660 32292 15712 32298
rect 15660 32234 15712 32240
rect 15672 32026 15700 32234
rect 15660 32020 15712 32026
rect 15660 31962 15712 31968
rect 15016 31816 15068 31822
rect 15016 31758 15068 31764
rect 15658 31784 15714 31793
rect 15658 31719 15714 31728
rect 15384 31680 15436 31686
rect 15384 31622 15436 31628
rect 15396 31521 15424 31622
rect 15382 31512 15438 31521
rect 15382 31447 15438 31456
rect 15292 31340 15344 31346
rect 15292 31282 15344 31288
rect 15200 30592 15252 30598
rect 15200 30534 15252 30540
rect 15212 30054 15240 30534
rect 15200 30048 15252 30054
rect 15200 29990 15252 29996
rect 15304 29730 15332 31282
rect 15396 29850 15424 31447
rect 15476 30048 15528 30054
rect 15476 29990 15528 29996
rect 15384 29844 15436 29850
rect 15384 29786 15436 29792
rect 15304 29702 15424 29730
rect 15488 29714 15516 29990
rect 14924 29572 14976 29578
rect 14924 29514 14976 29520
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 14924 29164 14976 29170
rect 14844 29124 14924 29152
rect 14740 28552 14792 28558
rect 14740 28494 14792 28500
rect 14752 27674 14780 28494
rect 14844 28422 14872 29124
rect 14924 29106 14976 29112
rect 15108 28484 15160 28490
rect 15108 28426 15160 28432
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14740 27668 14792 27674
rect 14740 27610 14792 27616
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14648 26784 14700 26790
rect 14648 26726 14700 26732
rect 14660 26382 14688 26726
rect 14648 26376 14700 26382
rect 14648 26318 14700 26324
rect 14476 26206 14596 26234
rect 14476 24818 14504 26206
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14476 23866 14504 24754
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14462 23760 14518 23769
rect 14462 23695 14518 23704
rect 14476 23662 14504 23695
rect 14464 23656 14516 23662
rect 14464 23598 14516 23604
rect 14366 23180 14418 23186
rect 14366 23122 14418 23128
rect 14372 23044 14424 23050
rect 14372 22986 14424 22992
rect 14384 22438 14412 22986
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14384 19718 14412 20878
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14372 19346 14424 19352
rect 14372 19288 14424 19294
rect 14384 18873 14412 19288
rect 14476 18902 14504 23598
rect 14568 22094 14596 25842
rect 14752 25294 14780 27406
rect 14740 25288 14792 25294
rect 14740 25230 14792 25236
rect 14752 23798 14780 25230
rect 14844 24682 14872 28358
rect 15016 27124 15068 27130
rect 15016 27066 15068 27072
rect 15028 26450 15056 27066
rect 15016 26444 15068 26450
rect 15016 26386 15068 26392
rect 14924 25900 14976 25906
rect 14924 25842 14976 25848
rect 14936 24886 14964 25842
rect 15120 25770 15148 28426
rect 15212 28150 15240 29446
rect 15396 28966 15424 29702
rect 15476 29708 15528 29714
rect 15476 29650 15528 29656
rect 15488 29170 15516 29650
rect 15672 29646 15700 31719
rect 15568 29640 15620 29646
rect 15568 29582 15620 29588
rect 15660 29640 15712 29646
rect 15660 29582 15712 29588
rect 15476 29164 15528 29170
rect 15476 29106 15528 29112
rect 15580 29050 15608 29582
rect 15488 29022 15608 29050
rect 15384 28960 15436 28966
rect 15384 28902 15436 28908
rect 15200 28144 15252 28150
rect 15200 28086 15252 28092
rect 15292 27872 15344 27878
rect 15292 27814 15344 27820
rect 15200 27600 15252 27606
rect 15200 27542 15252 27548
rect 15212 26858 15240 27542
rect 15304 27538 15332 27814
rect 15292 27532 15344 27538
rect 15292 27474 15344 27480
rect 15200 26852 15252 26858
rect 15200 26794 15252 26800
rect 15212 26586 15240 26794
rect 15304 26790 15332 27474
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15200 26580 15252 26586
rect 15200 26522 15252 26528
rect 15200 26308 15252 26314
rect 15200 26250 15252 26256
rect 15108 25764 15160 25770
rect 15108 25706 15160 25712
rect 14924 24880 14976 24886
rect 14924 24822 14976 24828
rect 14832 24676 14884 24682
rect 14832 24618 14884 24624
rect 14740 23792 14792 23798
rect 14740 23734 14792 23740
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 14660 23254 14688 23462
rect 14648 23248 14700 23254
rect 14648 23190 14700 23196
rect 14752 22574 14780 23734
rect 14844 23594 14872 24618
rect 14924 24268 14976 24274
rect 14924 24210 14976 24216
rect 14936 23866 14964 24210
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 15016 23724 15068 23730
rect 15016 23666 15068 23672
rect 14832 23588 14884 23594
rect 14832 23530 14884 23536
rect 15028 23050 15056 23666
rect 15120 23662 15148 25706
rect 15108 23656 15160 23662
rect 15108 23598 15160 23604
rect 15212 23118 15240 26250
rect 15292 24064 15344 24070
rect 15292 24006 15344 24012
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 14924 23044 14976 23050
rect 14924 22986 14976 22992
rect 15016 23044 15068 23050
rect 15068 23004 15148 23032
rect 15016 22986 15068 22992
rect 14740 22568 14792 22574
rect 14740 22510 14792 22516
rect 14568 22066 14688 22094
rect 14660 21350 14688 22066
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14844 21622 14872 21830
rect 14832 21616 14884 21622
rect 14832 21558 14884 21564
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14832 21344 14884 21350
rect 14832 21286 14884 21292
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14464 18896 14516 18902
rect 14370 18864 14426 18873
rect 14464 18838 14516 18844
rect 14568 18834 14596 20402
rect 14370 18799 14426 18808
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14292 18686 14504 18714
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14292 17678 14320 18566
rect 14280 17672 14332 17678
rect 14332 17632 14412 17660
rect 14280 17614 14332 17620
rect 14384 17202 14412 17632
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14200 16238 14320 16266
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14200 15706 14228 16050
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14292 15586 14320 16238
rect 14200 15558 14320 15586
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 14482 14136 14758
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13740 11898 13768 12038
rect 14200 11898 14228 15558
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14016 9178 14044 11630
rect 14200 11218 14228 11630
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14292 10266 14320 12718
rect 14476 11830 14504 18686
rect 14660 17746 14688 21286
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14752 19378 14780 19654
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14738 18864 14794 18873
rect 14738 18799 14794 18808
rect 14752 18766 14780 18799
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14568 15978 14596 17614
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14568 13530 14596 13874
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14660 13326 14688 17682
rect 14752 16794 14780 18226
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14752 14074 14780 14962
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14648 11824 14700 11830
rect 14648 11766 14700 11772
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9586 14136 9862
rect 14660 9586 14688 11766
rect 14752 10130 14780 11834
rect 14844 10266 14872 21286
rect 14936 20788 14964 22986
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 15028 21010 15056 21830
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 15120 20942 15148 23004
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 15212 22642 15240 22918
rect 15304 22642 15332 24006
rect 15200 22636 15252 22642
rect 15200 22578 15252 22584
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15396 22522 15424 28902
rect 15488 26790 15516 29022
rect 15568 28552 15620 28558
rect 15568 28494 15620 28500
rect 15580 27674 15608 28494
rect 15568 27668 15620 27674
rect 15568 27610 15620 27616
rect 15672 27606 15700 29582
rect 15764 28150 15792 33510
rect 15844 33516 15896 33522
rect 15844 33458 15896 33464
rect 16224 33318 16252 34478
rect 16212 33312 16264 33318
rect 16212 33254 16264 33260
rect 15846 33212 16154 33232
rect 15846 33210 15852 33212
rect 15908 33210 15932 33212
rect 15988 33210 16012 33212
rect 16068 33210 16092 33212
rect 16148 33210 16154 33212
rect 15908 33158 15910 33210
rect 16090 33158 16092 33210
rect 15846 33156 15852 33158
rect 15908 33156 15932 33158
rect 15988 33156 16012 33158
rect 16068 33156 16092 33158
rect 16148 33156 16154 33158
rect 15846 33136 16154 33156
rect 16304 33108 16356 33114
rect 16304 33050 16356 33056
rect 16212 32428 16264 32434
rect 16212 32370 16264 32376
rect 15846 32124 16154 32144
rect 15846 32122 15852 32124
rect 15908 32122 15932 32124
rect 15988 32122 16012 32124
rect 16068 32122 16092 32124
rect 16148 32122 16154 32124
rect 15908 32070 15910 32122
rect 16090 32070 16092 32122
rect 15846 32068 15852 32070
rect 15908 32068 15932 32070
rect 15988 32068 16012 32070
rect 16068 32068 16092 32070
rect 16148 32068 16154 32070
rect 15846 32048 16154 32068
rect 15936 31816 15988 31822
rect 15936 31758 15988 31764
rect 15948 31482 15976 31758
rect 16224 31754 16252 32370
rect 16316 32026 16344 33050
rect 16304 32020 16356 32026
rect 16304 31962 16356 31968
rect 16224 31726 16344 31754
rect 15936 31476 15988 31482
rect 15936 31418 15988 31424
rect 15846 31036 16154 31056
rect 15846 31034 15852 31036
rect 15908 31034 15932 31036
rect 15988 31034 16012 31036
rect 16068 31034 16092 31036
rect 16148 31034 16154 31036
rect 15908 30982 15910 31034
rect 16090 30982 16092 31034
rect 15846 30980 15852 30982
rect 15908 30980 15932 30982
rect 15988 30980 16012 30982
rect 16068 30980 16092 30982
rect 16148 30980 16154 30982
rect 15846 30960 16154 30980
rect 16212 30660 16264 30666
rect 16212 30602 16264 30608
rect 15846 29948 16154 29968
rect 15846 29946 15852 29948
rect 15908 29946 15932 29948
rect 15988 29946 16012 29948
rect 16068 29946 16092 29948
rect 16148 29946 16154 29948
rect 15908 29894 15910 29946
rect 16090 29894 16092 29946
rect 15846 29892 15852 29894
rect 15908 29892 15932 29894
rect 15988 29892 16012 29894
rect 16068 29892 16092 29894
rect 16148 29892 16154 29894
rect 15846 29872 16154 29892
rect 16028 29640 16080 29646
rect 16028 29582 16080 29588
rect 16120 29640 16172 29646
rect 16120 29582 16172 29588
rect 16040 29209 16068 29582
rect 16132 29306 16160 29582
rect 16120 29300 16172 29306
rect 16120 29242 16172 29248
rect 16026 29200 16082 29209
rect 16026 29135 16082 29144
rect 15846 28860 16154 28880
rect 15846 28858 15852 28860
rect 15908 28858 15932 28860
rect 15988 28858 16012 28860
rect 16068 28858 16092 28860
rect 16148 28858 16154 28860
rect 15908 28806 15910 28858
rect 16090 28806 16092 28858
rect 15846 28804 15852 28806
rect 15908 28804 15932 28806
rect 15988 28804 16012 28806
rect 16068 28804 16092 28806
rect 16148 28804 16154 28806
rect 15846 28784 16154 28804
rect 15752 28144 15804 28150
rect 15752 28086 15804 28092
rect 15846 27772 16154 27792
rect 15846 27770 15852 27772
rect 15908 27770 15932 27772
rect 15988 27770 16012 27772
rect 16068 27770 16092 27772
rect 16148 27770 16154 27772
rect 15908 27718 15910 27770
rect 16090 27718 16092 27770
rect 15846 27716 15852 27718
rect 15908 27716 15932 27718
rect 15988 27716 16012 27718
rect 16068 27716 16092 27718
rect 16148 27716 16154 27718
rect 15846 27696 16154 27716
rect 15660 27600 15712 27606
rect 15660 27542 15712 27548
rect 16120 27464 16172 27470
rect 16120 27406 16172 27412
rect 15568 27328 15620 27334
rect 15568 27270 15620 27276
rect 15752 27328 15804 27334
rect 15752 27270 15804 27276
rect 15476 26784 15528 26790
rect 15476 26726 15528 26732
rect 15476 26376 15528 26382
rect 15476 26318 15528 26324
rect 15488 25770 15516 26318
rect 15580 25974 15608 27270
rect 15568 25968 15620 25974
rect 15568 25910 15620 25916
rect 15660 25832 15712 25838
rect 15660 25774 15712 25780
rect 15476 25764 15528 25770
rect 15476 25706 15528 25712
rect 15476 25152 15528 25158
rect 15476 25094 15528 25100
rect 15488 24206 15516 25094
rect 15568 24676 15620 24682
rect 15568 24618 15620 24624
rect 15476 24200 15528 24206
rect 15580 24188 15608 24618
rect 15672 24410 15700 25774
rect 15764 25242 15792 27270
rect 16132 27130 16160 27406
rect 16224 27334 16252 30602
rect 16212 27328 16264 27334
rect 16212 27270 16264 27276
rect 16120 27124 16172 27130
rect 16120 27066 16172 27072
rect 16316 26874 16344 31726
rect 16224 26846 16344 26874
rect 15846 26684 16154 26704
rect 15846 26682 15852 26684
rect 15908 26682 15932 26684
rect 15988 26682 16012 26684
rect 16068 26682 16092 26684
rect 16148 26682 16154 26684
rect 15908 26630 15910 26682
rect 16090 26630 16092 26682
rect 15846 26628 15852 26630
rect 15908 26628 15932 26630
rect 15988 26628 16012 26630
rect 16068 26628 16092 26630
rect 16148 26628 16154 26630
rect 15846 26608 16154 26628
rect 16028 26512 16080 26518
rect 16028 26454 16080 26460
rect 15936 26240 15988 26246
rect 15936 26182 15988 26188
rect 15948 26042 15976 26182
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 16040 25684 16068 26454
rect 16224 25945 16252 26846
rect 16304 26784 16356 26790
rect 16304 26726 16356 26732
rect 16210 25936 16266 25945
rect 16210 25871 16266 25880
rect 16040 25656 16252 25684
rect 15846 25596 16154 25616
rect 15846 25594 15852 25596
rect 15908 25594 15932 25596
rect 15988 25594 16012 25596
rect 16068 25594 16092 25596
rect 16148 25594 16154 25596
rect 15908 25542 15910 25594
rect 16090 25542 16092 25594
rect 15846 25540 15852 25542
rect 15908 25540 15932 25542
rect 15988 25540 16012 25542
rect 16068 25540 16092 25542
rect 16148 25540 16154 25542
rect 15846 25520 16154 25540
rect 15764 25214 15976 25242
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15580 24160 15700 24188
rect 15476 24142 15528 24148
rect 15476 23792 15528 23798
rect 15476 23734 15528 23740
rect 15488 22642 15516 23734
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15200 22500 15252 22506
rect 15200 22442 15252 22448
rect 15304 22494 15424 22522
rect 15108 20936 15160 20942
rect 15108 20878 15160 20884
rect 14936 20760 15148 20788
rect 15014 20632 15070 20641
rect 15014 20567 15070 20576
rect 15028 20534 15056 20567
rect 15016 20528 15068 20534
rect 15016 20470 15068 20476
rect 14924 19984 14976 19990
rect 14924 19926 14976 19932
rect 14936 19378 14964 19926
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 15028 19446 15056 19654
rect 15016 19440 15068 19446
rect 15016 19382 15068 19388
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 15028 19145 15056 19246
rect 15014 19136 15070 19145
rect 15014 19071 15070 19080
rect 15120 18358 15148 20760
rect 15212 18714 15240 22442
rect 15304 21146 15332 22494
rect 15384 22432 15436 22438
rect 15384 22374 15436 22380
rect 15396 22030 15424 22374
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15384 22024 15436 22030
rect 15384 21966 15436 21972
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15488 21026 15516 21966
rect 15304 20998 15516 21026
rect 15304 18850 15332 20998
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15396 20448 15424 20810
rect 15476 20460 15528 20466
rect 15396 20420 15476 20448
rect 15476 20402 15528 20408
rect 15488 20058 15516 20402
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15580 19922 15608 22034
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15396 18970 15424 19654
rect 15580 19446 15608 19722
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15304 18834 15424 18850
rect 15304 18828 15436 18834
rect 15304 18822 15384 18828
rect 15384 18770 15436 18776
rect 15476 18760 15528 18766
rect 15212 18686 15424 18714
rect 15476 18702 15528 18708
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15108 18352 15160 18358
rect 14936 18312 15108 18340
rect 14936 15910 14964 18312
rect 15108 18294 15160 18300
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15120 18086 15148 18158
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 15212 17678 15240 18566
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15304 17882 15332 18226
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15396 17490 15424 18686
rect 15304 17462 15424 17490
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15028 16454 15056 16934
rect 15304 16590 15332 17462
rect 15488 17338 15516 18702
rect 15580 18426 15608 18702
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15672 18170 15700 24160
rect 15764 22642 15792 25094
rect 15948 24682 15976 25214
rect 15936 24676 15988 24682
rect 15936 24618 15988 24624
rect 15846 24508 16154 24528
rect 15846 24506 15852 24508
rect 15908 24506 15932 24508
rect 15988 24506 16012 24508
rect 16068 24506 16092 24508
rect 16148 24506 16154 24508
rect 15908 24454 15910 24506
rect 16090 24454 16092 24506
rect 15846 24452 15852 24454
rect 15908 24452 15932 24454
rect 15988 24452 16012 24454
rect 16068 24452 16092 24454
rect 16148 24452 16154 24454
rect 15846 24432 16154 24452
rect 16224 24206 16252 25656
rect 16316 25242 16344 26726
rect 16408 25838 16436 40870
rect 16500 40594 16528 41618
rect 16672 41540 16724 41546
rect 16672 41482 16724 41488
rect 16684 41274 16712 41482
rect 16868 41478 16896 44814
rect 16960 44334 16988 45018
rect 16948 44328 17000 44334
rect 16948 44270 17000 44276
rect 16948 43784 17000 43790
rect 16948 43726 17000 43732
rect 16960 42158 16988 43726
rect 17052 43246 17080 45222
rect 17144 43314 17172 47200
rect 17500 45620 17552 45626
rect 17500 45562 17552 45568
rect 17408 45416 17460 45422
rect 17408 45358 17460 45364
rect 17314 44976 17370 44985
rect 17224 44940 17276 44946
rect 17314 44911 17370 44920
rect 17224 44882 17276 44888
rect 17236 44849 17264 44882
rect 17222 44840 17278 44849
rect 17328 44810 17356 44911
rect 17222 44775 17278 44784
rect 17316 44804 17368 44810
rect 17316 44746 17368 44752
rect 17222 44296 17278 44305
rect 17222 44231 17278 44240
rect 17236 43382 17264 44231
rect 17328 44198 17356 44746
rect 17316 44192 17368 44198
rect 17316 44134 17368 44140
rect 17420 43858 17448 45358
rect 17512 44538 17540 45562
rect 17592 45280 17644 45286
rect 17592 45222 17644 45228
rect 17500 44532 17552 44538
rect 17500 44474 17552 44480
rect 17408 43852 17460 43858
rect 17408 43794 17460 43800
rect 17224 43376 17276 43382
rect 17420 43330 17448 43794
rect 17604 43790 17632 45222
rect 17880 44962 17908 47200
rect 18420 45484 18472 45490
rect 18420 45426 18472 45432
rect 18512 45484 18564 45490
rect 18512 45426 18564 45432
rect 17696 44934 17908 44962
rect 18432 44946 18460 45426
rect 18420 44940 18472 44946
rect 17592 43784 17644 43790
rect 17592 43726 17644 43732
rect 17592 43648 17644 43654
rect 17592 43590 17644 43596
rect 17604 43450 17632 43590
rect 17592 43444 17644 43450
rect 17592 43386 17644 43392
rect 17224 43318 17276 43324
rect 17132 43308 17184 43314
rect 17132 43250 17184 43256
rect 17328 43302 17448 43330
rect 17040 43240 17092 43246
rect 17040 43182 17092 43188
rect 17052 42906 17080 43182
rect 17040 42900 17092 42906
rect 17040 42842 17092 42848
rect 17052 42634 17080 42842
rect 17328 42770 17356 43302
rect 17408 43240 17460 43246
rect 17408 43182 17460 43188
rect 17420 42906 17448 43182
rect 17408 42900 17460 42906
rect 17408 42842 17460 42848
rect 17316 42764 17368 42770
rect 17316 42706 17368 42712
rect 17040 42628 17092 42634
rect 17040 42570 17092 42576
rect 17224 42560 17276 42566
rect 17224 42502 17276 42508
rect 16948 42152 17000 42158
rect 16948 42094 17000 42100
rect 17132 42152 17184 42158
rect 17132 42094 17184 42100
rect 16960 41750 16988 42094
rect 16948 41744 17000 41750
rect 16948 41686 17000 41692
rect 16856 41472 16908 41478
rect 16856 41414 16908 41420
rect 16672 41268 16724 41274
rect 16672 41210 16724 41216
rect 16868 41138 16896 41414
rect 16856 41132 16908 41138
rect 16856 41074 16908 41080
rect 17144 41070 17172 42094
rect 17132 41064 17184 41070
rect 17132 41006 17184 41012
rect 17040 40928 17092 40934
rect 17040 40870 17092 40876
rect 16856 40656 16908 40662
rect 16856 40598 16908 40604
rect 16488 40588 16540 40594
rect 16488 40530 16540 40536
rect 16580 40384 16632 40390
rect 16580 40326 16632 40332
rect 16592 40186 16620 40326
rect 16580 40180 16632 40186
rect 16580 40122 16632 40128
rect 16580 39500 16632 39506
rect 16580 39442 16632 39448
rect 16592 38282 16620 39442
rect 16672 38956 16724 38962
rect 16672 38898 16724 38904
rect 16580 38276 16632 38282
rect 16580 38218 16632 38224
rect 16592 37738 16620 38218
rect 16580 37732 16632 37738
rect 16580 37674 16632 37680
rect 16488 37664 16540 37670
rect 16488 37606 16540 37612
rect 16500 29850 16528 37606
rect 16580 37256 16632 37262
rect 16580 37198 16632 37204
rect 16592 35630 16620 37198
rect 16684 36242 16712 38898
rect 16764 37188 16816 37194
rect 16764 37130 16816 37136
rect 16672 36236 16724 36242
rect 16672 36178 16724 36184
rect 16580 35624 16632 35630
rect 16580 35566 16632 35572
rect 16592 30977 16620 35566
rect 16684 35290 16712 36178
rect 16776 35290 16804 37130
rect 16672 35284 16724 35290
rect 16672 35226 16724 35232
rect 16764 35284 16816 35290
rect 16764 35226 16816 35232
rect 16776 35086 16804 35226
rect 16764 35080 16816 35086
rect 16764 35022 16816 35028
rect 16672 34128 16724 34134
rect 16672 34070 16724 34076
rect 16684 33930 16712 34070
rect 16672 33924 16724 33930
rect 16672 33866 16724 33872
rect 16764 33856 16816 33862
rect 16764 33798 16816 33804
rect 16776 33590 16804 33798
rect 16764 33584 16816 33590
rect 16764 33526 16816 33532
rect 16672 33108 16724 33114
rect 16672 33050 16724 33056
rect 16684 31958 16712 33050
rect 16776 32774 16804 33526
rect 16868 33522 16896 40598
rect 16948 40384 17000 40390
rect 16948 40326 17000 40332
rect 16960 40050 16988 40326
rect 16948 40044 17000 40050
rect 16948 39986 17000 39992
rect 16960 39846 16988 39986
rect 17052 39982 17080 40870
rect 17144 40186 17172 41006
rect 17132 40180 17184 40186
rect 17132 40122 17184 40128
rect 17040 39976 17092 39982
rect 17040 39918 17092 39924
rect 16948 39840 17000 39846
rect 16948 39782 17000 39788
rect 16948 38956 17000 38962
rect 16948 38898 17000 38904
rect 16960 38554 16988 38898
rect 16948 38548 17000 38554
rect 16948 38490 17000 38496
rect 17132 37732 17184 37738
rect 17132 37674 17184 37680
rect 16948 37664 17000 37670
rect 16948 37606 17000 37612
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 16764 32768 16816 32774
rect 16764 32710 16816 32716
rect 16856 32224 16908 32230
rect 16856 32166 16908 32172
rect 16672 31952 16724 31958
rect 16672 31894 16724 31900
rect 16764 31748 16816 31754
rect 16764 31690 16816 31696
rect 16776 31142 16804 31690
rect 16764 31136 16816 31142
rect 16764 31078 16816 31084
rect 16578 30968 16634 30977
rect 16578 30903 16634 30912
rect 16578 30832 16634 30841
rect 16578 30767 16634 30776
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16488 29028 16540 29034
rect 16488 28970 16540 28976
rect 16500 26314 16528 28970
rect 16488 26308 16540 26314
rect 16488 26250 16540 26256
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 16396 25696 16448 25702
rect 16396 25638 16448 25644
rect 16408 25362 16436 25638
rect 16396 25356 16448 25362
rect 16396 25298 16448 25304
rect 16316 25214 16436 25242
rect 16304 25152 16356 25158
rect 16302 25120 16304 25129
rect 16356 25120 16358 25129
rect 16302 25055 16358 25064
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16316 24313 16344 24346
rect 16302 24304 16358 24313
rect 16302 24239 16358 24248
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16304 23520 16356 23526
rect 16304 23462 16356 23468
rect 15846 23420 16154 23440
rect 15846 23418 15852 23420
rect 15908 23418 15932 23420
rect 15988 23418 16012 23420
rect 16068 23418 16092 23420
rect 16148 23418 16154 23420
rect 15908 23366 15910 23418
rect 16090 23366 16092 23418
rect 15846 23364 15852 23366
rect 15908 23364 15932 23366
rect 15988 23364 16012 23366
rect 16068 23364 16092 23366
rect 16148 23364 16154 23366
rect 15846 23344 16154 23364
rect 15936 23248 15988 23254
rect 15934 23216 15936 23225
rect 15988 23216 15990 23225
rect 15934 23151 15990 23160
rect 16212 23180 16264 23186
rect 16212 23122 16264 23128
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15752 22500 15804 22506
rect 15752 22442 15804 22448
rect 15764 22094 15792 22442
rect 15846 22332 16154 22352
rect 15846 22330 15852 22332
rect 15908 22330 15932 22332
rect 15988 22330 16012 22332
rect 16068 22330 16092 22332
rect 16148 22330 16154 22332
rect 15908 22278 15910 22330
rect 16090 22278 16092 22330
rect 15846 22276 15852 22278
rect 15908 22276 15932 22278
rect 15988 22276 16012 22278
rect 16068 22276 16092 22278
rect 16148 22276 16154 22278
rect 15846 22256 16154 22276
rect 15844 22094 15896 22098
rect 15764 22092 15896 22094
rect 15764 22066 15844 22092
rect 15844 22034 15896 22040
rect 15752 22024 15804 22030
rect 15752 21966 15804 21972
rect 15764 18272 15792 21966
rect 15846 21244 16154 21264
rect 15846 21242 15852 21244
rect 15908 21242 15932 21244
rect 15988 21242 16012 21244
rect 16068 21242 16092 21244
rect 16148 21242 16154 21244
rect 15908 21190 15910 21242
rect 16090 21190 16092 21242
rect 15846 21188 15852 21190
rect 15908 21188 15932 21190
rect 15988 21188 16012 21190
rect 16068 21188 16092 21190
rect 16148 21188 16154 21190
rect 15846 21168 16154 21188
rect 15846 20156 16154 20176
rect 15846 20154 15852 20156
rect 15908 20154 15932 20156
rect 15988 20154 16012 20156
rect 16068 20154 16092 20156
rect 16148 20154 16154 20156
rect 15908 20102 15910 20154
rect 16090 20102 16092 20154
rect 15846 20100 15852 20102
rect 15908 20100 15932 20102
rect 15988 20100 16012 20102
rect 16068 20100 16092 20102
rect 16148 20100 16154 20102
rect 15846 20080 16154 20100
rect 16224 19854 16252 23122
rect 16316 23118 16344 23462
rect 16304 23112 16356 23118
rect 16304 23054 16356 23060
rect 16316 21554 16344 23054
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 16224 19378 16252 19654
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 15846 19068 16154 19088
rect 15846 19066 15852 19068
rect 15908 19066 15932 19068
rect 15988 19066 16012 19068
rect 16068 19066 16092 19068
rect 16148 19066 16154 19068
rect 15908 19014 15910 19066
rect 16090 19014 16092 19066
rect 15846 19012 15852 19014
rect 15908 19012 15932 19014
rect 15988 19012 16012 19014
rect 16068 19012 16092 19014
rect 16148 19012 16154 19014
rect 15846 18992 16154 19012
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 15764 18244 15884 18272
rect 15580 18142 15700 18170
rect 15856 18154 15884 18244
rect 16040 18222 16068 18770
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16132 18290 16160 18702
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15752 18148 15804 18154
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15396 16726 15424 17274
rect 15384 16720 15436 16726
rect 15384 16662 15436 16668
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 15028 15434 15056 16390
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15028 14770 15056 15370
rect 15120 14958 15148 16186
rect 15304 15450 15332 16526
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15396 16250 15424 16458
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15304 15422 15516 15450
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 15028 14742 15148 14770
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 15028 13462 15056 14418
rect 15120 14278 15148 14742
rect 15212 14414 15240 15302
rect 15396 15094 15424 15302
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15304 14618 15332 14962
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15016 13456 15068 13462
rect 15016 13398 15068 13404
rect 15028 12782 15056 13398
rect 15120 13190 15148 14214
rect 15488 14006 15516 15422
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15580 13920 15608 18142
rect 15752 18090 15804 18096
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15672 16998 15700 18022
rect 15764 17882 15792 18090
rect 15846 17980 16154 18000
rect 15846 17978 15852 17980
rect 15908 17978 15932 17980
rect 15988 17978 16012 17980
rect 16068 17978 16092 17980
rect 16148 17978 16154 17980
rect 15908 17926 15910 17978
rect 16090 17926 16092 17978
rect 15846 17924 15852 17926
rect 15908 17924 15932 17926
rect 15988 17924 16012 17926
rect 16068 17924 16092 17926
rect 16148 17924 16154 17926
rect 15846 17904 16154 17924
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 16224 17678 16252 19314
rect 16316 17785 16344 19858
rect 16408 18902 16436 25214
rect 16500 24682 16528 26250
rect 16592 25158 16620 30767
rect 16776 30190 16804 31078
rect 16868 30666 16896 32166
rect 16960 31822 16988 37606
rect 17040 37120 17092 37126
rect 17040 37062 17092 37068
rect 17052 35034 17080 37062
rect 17144 36666 17172 37674
rect 17236 36786 17264 42502
rect 17420 42294 17448 42842
rect 17696 42838 17724 44934
rect 18420 44882 18472 44888
rect 17776 44872 17828 44878
rect 17776 44814 17828 44820
rect 18052 44872 18104 44878
rect 18052 44814 18104 44820
rect 17684 42832 17736 42838
rect 17684 42774 17736 42780
rect 17788 42770 17816 44814
rect 17868 44736 17920 44742
rect 17868 44678 17920 44684
rect 17880 44470 17908 44678
rect 17868 44464 17920 44470
rect 17868 44406 17920 44412
rect 17960 44192 18012 44198
rect 17960 44134 18012 44140
rect 17972 43314 18000 44134
rect 17960 43308 18012 43314
rect 17960 43250 18012 43256
rect 17776 42764 17828 42770
rect 17776 42706 17828 42712
rect 17788 42566 17816 42706
rect 17684 42560 17736 42566
rect 17684 42502 17736 42508
rect 17776 42560 17828 42566
rect 17776 42502 17828 42508
rect 17696 42362 17724 42502
rect 17684 42356 17736 42362
rect 17684 42298 17736 42304
rect 17408 42288 17460 42294
rect 17408 42230 17460 42236
rect 17788 42226 17816 42502
rect 17776 42220 17828 42226
rect 17776 42162 17828 42168
rect 17500 41608 17552 41614
rect 17500 41550 17552 41556
rect 17512 40934 17540 41550
rect 18064 41002 18092 44814
rect 18524 44470 18552 45426
rect 18512 44464 18564 44470
rect 18512 44406 18564 44412
rect 18616 43994 18644 47200
rect 19340 45416 19392 45422
rect 19340 45358 19392 45364
rect 19444 45370 19472 47200
rect 19248 45008 19300 45014
rect 19248 44950 19300 44956
rect 18696 44464 18748 44470
rect 18696 44406 18748 44412
rect 18708 44266 18736 44406
rect 18696 44260 18748 44266
rect 18696 44202 18748 44208
rect 18972 44192 19024 44198
rect 18972 44134 19024 44140
rect 18604 43988 18656 43994
rect 18604 43930 18656 43936
rect 18788 43648 18840 43654
rect 18788 43590 18840 43596
rect 18144 43308 18196 43314
rect 18144 43250 18196 43256
rect 18156 41274 18184 43250
rect 18604 43240 18656 43246
rect 18604 43182 18656 43188
rect 18512 43104 18564 43110
rect 18510 43072 18512 43081
rect 18564 43072 18566 43081
rect 18510 43007 18566 43016
rect 18420 42764 18472 42770
rect 18420 42706 18472 42712
rect 18144 41268 18196 41274
rect 18144 41210 18196 41216
rect 18432 41070 18460 42706
rect 18512 42356 18564 42362
rect 18512 42298 18564 42304
rect 18524 42022 18552 42298
rect 18616 42158 18644 43182
rect 18696 43104 18748 43110
rect 18696 43046 18748 43052
rect 18604 42152 18656 42158
rect 18604 42094 18656 42100
rect 18512 42016 18564 42022
rect 18512 41958 18564 41964
rect 18524 41546 18552 41958
rect 18512 41540 18564 41546
rect 18512 41482 18564 41488
rect 18420 41064 18472 41070
rect 18420 41006 18472 41012
rect 18052 40996 18104 41002
rect 18052 40938 18104 40944
rect 17500 40928 17552 40934
rect 17500 40870 17552 40876
rect 17868 40928 17920 40934
rect 17868 40870 17920 40876
rect 17684 40044 17736 40050
rect 17684 39986 17736 39992
rect 17592 39840 17644 39846
rect 17592 39782 17644 39788
rect 17500 38208 17552 38214
rect 17500 38150 17552 38156
rect 17224 36780 17276 36786
rect 17224 36722 17276 36728
rect 17144 36650 17264 36666
rect 17144 36644 17276 36650
rect 17144 36638 17224 36644
rect 17224 36586 17276 36592
rect 17132 36576 17184 36582
rect 17132 36518 17184 36524
rect 17144 36174 17172 36518
rect 17132 36168 17184 36174
rect 17132 36110 17184 36116
rect 17132 35692 17184 35698
rect 17236 35680 17264 36586
rect 17184 35652 17264 35680
rect 17132 35634 17184 35640
rect 17052 35006 17172 35034
rect 17040 34944 17092 34950
rect 17040 34886 17092 34892
rect 16948 31816 17000 31822
rect 16948 31758 17000 31764
rect 16948 31680 17000 31686
rect 16948 31622 17000 31628
rect 16856 30660 16908 30666
rect 16856 30602 16908 30608
rect 16854 30424 16910 30433
rect 16854 30359 16910 30368
rect 16868 30326 16896 30359
rect 16960 30326 16988 31622
rect 16856 30320 16908 30326
rect 16856 30262 16908 30268
rect 16948 30320 17000 30326
rect 16948 30262 17000 30268
rect 16764 30184 16816 30190
rect 16764 30126 16816 30132
rect 16776 29646 16804 30126
rect 16948 30048 17000 30054
rect 16948 29990 17000 29996
rect 16764 29640 16816 29646
rect 16764 29582 16816 29588
rect 16776 29306 16804 29582
rect 16856 29504 16908 29510
rect 16856 29446 16908 29452
rect 16764 29300 16816 29306
rect 16764 29242 16816 29248
rect 16868 29170 16896 29446
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16764 29096 16816 29102
rect 16764 29038 16816 29044
rect 16672 28960 16724 28966
rect 16672 28902 16724 28908
rect 16684 28558 16712 28902
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 16672 28212 16724 28218
rect 16672 28154 16724 28160
rect 16684 27674 16712 28154
rect 16672 27668 16724 27674
rect 16672 27610 16724 27616
rect 16672 26308 16724 26314
rect 16672 26250 16724 26256
rect 16684 25362 16712 26250
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16488 24676 16540 24682
rect 16488 24618 16540 24624
rect 16684 23882 16712 25298
rect 16592 23854 16712 23882
rect 16592 22642 16620 23854
rect 16672 23792 16724 23798
rect 16672 23734 16724 23740
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16592 22234 16620 22578
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16592 21690 16620 21830
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16592 20398 16620 21286
rect 16684 20874 16712 23734
rect 16776 22545 16804 29038
rect 16856 28552 16908 28558
rect 16856 28494 16908 28500
rect 16868 26994 16896 28494
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 16868 26586 16896 26930
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 16868 25430 16896 25774
rect 16856 25424 16908 25430
rect 16856 25366 16908 25372
rect 16856 24948 16908 24954
rect 16856 24890 16908 24896
rect 16868 24070 16896 24890
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16960 23610 16988 29990
rect 16868 23582 16988 23610
rect 17052 23594 17080 34886
rect 17144 33114 17172 35006
rect 17408 34944 17460 34950
rect 17328 34904 17408 34932
rect 17328 34746 17356 34904
rect 17408 34886 17460 34892
rect 17224 34740 17276 34746
rect 17224 34682 17276 34688
rect 17316 34740 17368 34746
rect 17316 34682 17368 34688
rect 17236 34649 17264 34682
rect 17222 34640 17278 34649
rect 17222 34575 17278 34584
rect 17132 33108 17184 33114
rect 17132 33050 17184 33056
rect 17132 32428 17184 32434
rect 17132 32370 17184 32376
rect 17040 23588 17092 23594
rect 16762 22536 16818 22545
rect 16762 22471 16818 22480
rect 16868 22420 16896 23582
rect 17040 23530 17092 23536
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16960 23322 16988 23462
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 17040 23316 17092 23322
rect 17040 23258 17092 23264
rect 17052 23202 17080 23258
rect 16960 23174 17080 23202
rect 16960 22982 16988 23174
rect 16948 22976 17000 22982
rect 16948 22918 17000 22924
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 16960 22642 16988 22918
rect 17052 22778 17080 22918
rect 17144 22778 17172 32370
rect 17328 30716 17356 34682
rect 17408 33312 17460 33318
rect 17408 33254 17460 33260
rect 17420 32842 17448 33254
rect 17408 32836 17460 32842
rect 17408 32778 17460 32784
rect 17408 31680 17460 31686
rect 17408 31622 17460 31628
rect 17236 30688 17356 30716
rect 17236 29510 17264 30688
rect 17316 30592 17368 30598
rect 17316 30534 17368 30540
rect 17328 30258 17356 30534
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 17224 29504 17276 29510
rect 17222 29472 17224 29481
rect 17276 29472 17278 29481
rect 17222 29407 17278 29416
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17236 24342 17264 29106
rect 17328 28422 17356 30194
rect 17316 28416 17368 28422
rect 17316 28358 17368 28364
rect 17314 28248 17370 28257
rect 17314 28183 17316 28192
rect 17368 28183 17370 28192
rect 17316 28154 17368 28160
rect 17316 27940 17368 27946
rect 17316 27882 17368 27888
rect 17328 27470 17356 27882
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 17316 26580 17368 26586
rect 17316 26522 17368 26528
rect 17224 24336 17276 24342
rect 17224 24278 17276 24284
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17236 23526 17264 24142
rect 17224 23520 17276 23526
rect 17224 23462 17276 23468
rect 17328 23186 17356 26522
rect 17420 25294 17448 31622
rect 17512 30666 17540 38150
rect 17604 33969 17632 39782
rect 17696 39438 17724 39986
rect 17776 39500 17828 39506
rect 17776 39442 17828 39448
rect 17684 39432 17736 39438
rect 17684 39374 17736 39380
rect 17696 38350 17724 39374
rect 17684 38344 17736 38350
rect 17684 38286 17736 38292
rect 17788 38282 17816 39442
rect 17880 39438 17908 40870
rect 17960 40588 18012 40594
rect 17960 40530 18012 40536
rect 17868 39432 17920 39438
rect 17868 39374 17920 39380
rect 17776 38276 17828 38282
rect 17776 38218 17828 38224
rect 17684 36780 17736 36786
rect 17684 36722 17736 36728
rect 17696 36038 17724 36722
rect 17684 36032 17736 36038
rect 17684 35974 17736 35980
rect 17696 33998 17724 35974
rect 17972 35698 18000 40530
rect 18064 40526 18092 40938
rect 18144 40928 18196 40934
rect 18144 40870 18196 40876
rect 18052 40520 18104 40526
rect 18052 40462 18104 40468
rect 18052 38752 18104 38758
rect 18052 38694 18104 38700
rect 18064 38418 18092 38694
rect 18052 38412 18104 38418
rect 18052 38354 18104 38360
rect 18156 38350 18184 40870
rect 18432 40610 18460 41006
rect 18248 40582 18460 40610
rect 18524 40594 18552 41482
rect 18248 40458 18276 40582
rect 18236 40452 18288 40458
rect 18236 40394 18288 40400
rect 18328 40452 18380 40458
rect 18328 40394 18380 40400
rect 18236 39432 18288 39438
rect 18236 39374 18288 39380
rect 18248 38758 18276 39374
rect 18236 38752 18288 38758
rect 18236 38694 18288 38700
rect 18144 38344 18196 38350
rect 18144 38286 18196 38292
rect 18052 38276 18104 38282
rect 18052 38218 18104 38224
rect 18064 36718 18092 38218
rect 18144 37868 18196 37874
rect 18248 37856 18276 38694
rect 18196 37828 18276 37856
rect 18144 37810 18196 37816
rect 18052 36712 18104 36718
rect 18052 36654 18104 36660
rect 18340 35698 18368 40394
rect 18432 40338 18460 40582
rect 18512 40588 18564 40594
rect 18512 40530 18564 40536
rect 18616 40458 18644 42094
rect 18708 41206 18736 43046
rect 18800 42158 18828 43590
rect 18788 42152 18840 42158
rect 18788 42094 18840 42100
rect 18696 41200 18748 41206
rect 18696 41142 18748 41148
rect 18604 40452 18656 40458
rect 18604 40394 18656 40400
rect 18432 40310 18644 40338
rect 18512 39500 18564 39506
rect 18512 39442 18564 39448
rect 18420 39296 18472 39302
rect 18420 39238 18472 39244
rect 18432 39030 18460 39238
rect 18420 39024 18472 39030
rect 18420 38966 18472 38972
rect 18524 38962 18552 39442
rect 18512 38956 18564 38962
rect 18512 38898 18564 38904
rect 18524 38010 18552 38898
rect 18512 38004 18564 38010
rect 18512 37946 18564 37952
rect 18420 37664 18472 37670
rect 18420 37606 18472 37612
rect 17960 35692 18012 35698
rect 17960 35634 18012 35640
rect 18328 35692 18380 35698
rect 18328 35634 18380 35640
rect 18052 35488 18104 35494
rect 18052 35430 18104 35436
rect 17960 35284 18012 35290
rect 17960 35226 18012 35232
rect 17776 35080 17828 35086
rect 17776 35022 17828 35028
rect 17788 34202 17816 35022
rect 17868 34468 17920 34474
rect 17868 34410 17920 34416
rect 17776 34196 17828 34202
rect 17776 34138 17828 34144
rect 17776 34060 17828 34066
rect 17776 34002 17828 34008
rect 17684 33992 17736 33998
rect 17590 33960 17646 33969
rect 17684 33934 17736 33940
rect 17590 33895 17646 33904
rect 17592 33856 17644 33862
rect 17592 33798 17644 33804
rect 17500 30660 17552 30666
rect 17500 30602 17552 30608
rect 17604 30258 17632 33798
rect 17788 33658 17816 34002
rect 17880 33998 17908 34410
rect 17868 33992 17920 33998
rect 17868 33934 17920 33940
rect 17776 33652 17828 33658
rect 17776 33594 17828 33600
rect 17972 33522 18000 35226
rect 17776 33516 17828 33522
rect 17776 33458 17828 33464
rect 17960 33516 18012 33522
rect 17960 33458 18012 33464
rect 17684 33448 17736 33454
rect 17684 33390 17736 33396
rect 17696 31929 17724 33390
rect 17788 33114 17816 33458
rect 17868 33380 17920 33386
rect 17868 33322 17920 33328
rect 17776 33108 17828 33114
rect 17776 33050 17828 33056
rect 17788 32434 17816 33050
rect 17776 32428 17828 32434
rect 17776 32370 17828 32376
rect 17682 31920 17738 31929
rect 17682 31855 17738 31864
rect 17880 31770 17908 33322
rect 17972 32978 18000 33458
rect 17960 32972 18012 32978
rect 17960 32914 18012 32920
rect 17960 32768 18012 32774
rect 17960 32710 18012 32716
rect 17788 31742 17908 31770
rect 17684 31408 17736 31414
rect 17684 31350 17736 31356
rect 17696 30802 17724 31350
rect 17684 30796 17736 30802
rect 17684 30738 17736 30744
rect 17788 30682 17816 31742
rect 17868 31680 17920 31686
rect 17868 31622 17920 31628
rect 17696 30654 17816 30682
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 17590 30152 17646 30161
rect 17590 30087 17646 30096
rect 17498 29744 17554 29753
rect 17498 29679 17554 29688
rect 17512 25906 17540 29679
rect 17604 28082 17632 30087
rect 17592 28076 17644 28082
rect 17592 28018 17644 28024
rect 17500 25900 17552 25906
rect 17604 25888 17632 28018
rect 17696 27606 17724 30654
rect 17776 30592 17828 30598
rect 17776 30534 17828 30540
rect 17684 27600 17736 27606
rect 17684 27542 17736 27548
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 17696 27130 17724 27406
rect 17684 27124 17736 27130
rect 17684 27066 17736 27072
rect 17604 25860 17724 25888
rect 17500 25842 17552 25848
rect 17696 25770 17724 25860
rect 17592 25764 17644 25770
rect 17592 25706 17644 25712
rect 17684 25764 17736 25770
rect 17684 25706 17736 25712
rect 17500 25696 17552 25702
rect 17500 25638 17552 25644
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 17512 24886 17540 25638
rect 17604 25226 17632 25706
rect 17788 25514 17816 30534
rect 17880 30054 17908 31622
rect 17972 31346 18000 32710
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17960 31136 18012 31142
rect 17960 31078 18012 31084
rect 17972 30870 18000 31078
rect 17960 30864 18012 30870
rect 17960 30806 18012 30812
rect 17960 30660 18012 30666
rect 17960 30602 18012 30608
rect 17868 30048 17920 30054
rect 17868 29990 17920 29996
rect 17880 29714 17908 29990
rect 17868 29708 17920 29714
rect 17868 29650 17920 29656
rect 17868 28484 17920 28490
rect 17868 28426 17920 28432
rect 17880 28218 17908 28426
rect 17868 28212 17920 28218
rect 17868 28154 17920 28160
rect 17868 28008 17920 28014
rect 17866 27976 17868 27985
rect 17920 27976 17922 27985
rect 17866 27911 17922 27920
rect 17880 27538 17908 27911
rect 17868 27532 17920 27538
rect 17868 27474 17920 27480
rect 17972 26382 18000 30602
rect 18064 29170 18092 35430
rect 18144 35216 18196 35222
rect 18144 35158 18196 35164
rect 18156 34406 18184 35158
rect 18144 34400 18196 34406
rect 18144 34342 18196 34348
rect 18156 31278 18184 34342
rect 18236 34060 18288 34066
rect 18236 34002 18288 34008
rect 18248 31958 18276 34002
rect 18340 33998 18368 35634
rect 18328 33992 18380 33998
rect 18328 33934 18380 33940
rect 18326 33824 18382 33833
rect 18326 33759 18382 33768
rect 18236 31952 18288 31958
rect 18236 31894 18288 31900
rect 18248 31521 18276 31894
rect 18340 31822 18368 33759
rect 18328 31816 18380 31822
rect 18328 31758 18380 31764
rect 18234 31512 18290 31521
rect 18234 31447 18290 31456
rect 18236 31408 18288 31414
rect 18236 31350 18288 31356
rect 18144 31272 18196 31278
rect 18144 31214 18196 31220
rect 18144 30796 18196 30802
rect 18144 30738 18196 30744
rect 18156 30433 18184 30738
rect 18248 30666 18276 31350
rect 18236 30660 18288 30666
rect 18236 30602 18288 30608
rect 18142 30424 18198 30433
rect 18142 30359 18198 30368
rect 18144 30320 18196 30326
rect 18144 30262 18196 30268
rect 18156 29753 18184 30262
rect 18236 30252 18288 30258
rect 18236 30194 18288 30200
rect 18142 29744 18198 29753
rect 18142 29679 18198 29688
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 17696 25486 17816 25514
rect 17592 25220 17644 25226
rect 17592 25162 17644 25168
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 17604 24750 17632 25162
rect 17592 24744 17644 24750
rect 17592 24686 17644 24692
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17408 24336 17460 24342
rect 17408 24278 17460 24284
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 17420 23050 17448 24278
rect 17512 23730 17540 24550
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17420 22642 17448 22986
rect 16948 22636 17000 22642
rect 16948 22578 17000 22584
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17512 22574 17540 23666
rect 17604 23526 17632 24686
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17500 22568 17552 22574
rect 17328 22516 17500 22522
rect 17328 22510 17552 22516
rect 17328 22494 17540 22510
rect 16776 22392 16896 22420
rect 16948 22432 17000 22438
rect 16672 20868 16724 20874
rect 16672 20810 16724 20816
rect 16580 20392 16632 20398
rect 16580 20334 16632 20340
rect 16488 20256 16540 20262
rect 16672 20256 16724 20262
rect 16540 20204 16620 20210
rect 16488 20198 16620 20204
rect 16672 20198 16724 20204
rect 16500 20182 16620 20198
rect 16592 20058 16620 20182
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16684 19990 16712 20198
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16396 18896 16448 18902
rect 16396 18838 16448 18844
rect 16500 18748 16528 19790
rect 16776 19786 16804 22392
rect 16948 22374 17000 22380
rect 17130 22400 17186 22409
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16868 21418 16896 22034
rect 16856 21412 16908 21418
rect 16856 21354 16908 21360
rect 16868 20398 16896 21354
rect 16856 20392 16908 20398
rect 16856 20334 16908 20340
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16408 18720 16528 18748
rect 16302 17776 16358 17785
rect 16408 17746 16436 18720
rect 16672 18352 16724 18358
rect 16670 18320 16672 18329
rect 16724 18320 16726 18329
rect 16670 18255 16726 18264
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16302 17711 16358 17720
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15764 17105 15792 17138
rect 15750 17096 15806 17105
rect 15750 17031 15806 17040
rect 15934 17096 15990 17105
rect 15934 17031 15936 17040
rect 15988 17031 15990 17040
rect 15936 17002 15988 17008
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15672 15502 15700 16934
rect 15846 16892 16154 16912
rect 15846 16890 15852 16892
rect 15908 16890 15932 16892
rect 15988 16890 16012 16892
rect 16068 16890 16092 16892
rect 16148 16890 16154 16892
rect 15908 16838 15910 16890
rect 16090 16838 16092 16890
rect 15846 16836 15852 16838
rect 15908 16836 15932 16838
rect 15988 16836 16012 16838
rect 16068 16836 16092 16838
rect 16148 16836 16154 16838
rect 15846 16816 16154 16836
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15948 16046 15976 16526
rect 16408 16130 16436 17682
rect 16500 16590 16528 18158
rect 16776 17270 16804 18158
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16316 16102 16436 16130
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15846 15804 16154 15824
rect 15846 15802 15852 15804
rect 15908 15802 15932 15804
rect 15988 15802 16012 15804
rect 16068 15802 16092 15804
rect 16148 15802 16154 15804
rect 15908 15750 15910 15802
rect 16090 15750 16092 15802
rect 15846 15748 15852 15750
rect 15908 15748 15932 15750
rect 15988 15748 16012 15750
rect 16068 15748 16092 15750
rect 16148 15748 16154 15750
rect 15846 15728 16154 15748
rect 16316 15638 16344 16102
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15764 14550 15792 14758
rect 15846 14716 16154 14736
rect 15846 14714 15852 14716
rect 15908 14714 15932 14716
rect 15988 14714 16012 14716
rect 16068 14714 16092 14716
rect 16148 14714 16154 14716
rect 15908 14662 15910 14714
rect 16090 14662 16092 14714
rect 15846 14660 15852 14662
rect 15908 14660 15932 14662
rect 15988 14660 16012 14662
rect 16068 14660 16092 14662
rect 16148 14660 16154 14662
rect 15846 14640 16154 14660
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15672 14074 15700 14350
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15580 13892 15700 13920
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15212 13394 15240 13806
rect 15672 13802 15700 13892
rect 15660 13796 15712 13802
rect 15660 13738 15712 13744
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15672 13326 15700 13738
rect 15846 13628 16154 13648
rect 15846 13626 15852 13628
rect 15908 13626 15932 13628
rect 15988 13626 16012 13628
rect 16068 13626 16092 13628
rect 16148 13626 16154 13628
rect 15908 13574 15910 13626
rect 16090 13574 16092 13626
rect 15846 13572 15852 13574
rect 15908 13572 15932 13574
rect 15988 13572 16012 13574
rect 16068 13572 16092 13574
rect 16148 13572 16154 13574
rect 15846 13552 16154 13572
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15120 12986 15148 13126
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 15028 12306 15056 12718
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 14924 12164 14976 12170
rect 14924 12106 14976 12112
rect 14936 11082 14964 12106
rect 15028 11694 15056 12242
rect 15396 12238 15424 13126
rect 15580 12986 15608 13194
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15672 12594 15700 13262
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16224 12646 16252 12854
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 15488 12566 15700 12594
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 15120 11898 15148 12038
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15304 11354 15332 11494
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15488 11234 15516 12566
rect 15846 12540 16154 12560
rect 15846 12538 15852 12540
rect 15908 12538 15932 12540
rect 15988 12538 16012 12540
rect 16068 12538 16092 12540
rect 16148 12538 16154 12540
rect 15908 12486 15910 12538
rect 16090 12486 16092 12538
rect 15846 12484 15852 12486
rect 15908 12484 15932 12486
rect 15988 12484 16012 12486
rect 16068 12484 16092 12486
rect 16148 12484 16154 12486
rect 15846 12464 16154 12484
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15672 12102 15700 12378
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15672 11558 15700 12038
rect 16224 11762 16252 12582
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15846 11452 16154 11472
rect 15846 11450 15852 11452
rect 15908 11450 15932 11452
rect 15988 11450 16012 11452
rect 16068 11450 16092 11452
rect 16148 11450 16154 11452
rect 15908 11398 15910 11450
rect 16090 11398 16092 11450
rect 15846 11396 15852 11398
rect 15908 11396 15932 11398
rect 15988 11396 16012 11398
rect 16068 11396 16092 11398
rect 16148 11396 16154 11398
rect 15846 11376 16154 11396
rect 16224 11354 16252 11698
rect 16316 11694 16344 12786
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 15304 11206 15516 11234
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13360 7744 13412 7750
rect 13280 7704 13360 7732
rect 13280 7410 13308 7704
rect 13360 7686 13412 7692
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13372 7342 13400 7482
rect 14108 7478 14136 9522
rect 14660 8974 14688 9522
rect 14752 9518 14780 10066
rect 14936 9926 14964 10610
rect 15304 10062 15332 11206
rect 16316 11150 16344 11630
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 15580 11014 15608 11086
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15580 10674 15608 10950
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 15212 9722 15240 9930
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15200 9580 15252 9586
rect 15304 9568 15332 9998
rect 15252 9540 15332 9568
rect 15384 9580 15436 9586
rect 15200 9522 15252 9528
rect 15384 9522 15436 9528
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 9042 14780 9454
rect 15396 9178 15424 9522
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15488 9042 15516 10542
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15580 8974 15608 10610
rect 15856 10554 15884 10610
rect 15764 10526 15884 10554
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15672 9994 15700 10406
rect 15764 10062 15792 10526
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 15846 10364 16154 10384
rect 15846 10362 15852 10364
rect 15908 10362 15932 10364
rect 15988 10362 16012 10364
rect 16068 10362 16092 10364
rect 16148 10362 16154 10364
rect 15908 10310 15910 10362
rect 16090 10310 16092 10362
rect 15846 10308 15852 10310
rect 15908 10308 15932 10310
rect 15988 10308 16012 10310
rect 16068 10308 16092 10310
rect 16148 10308 16154 10310
rect 15846 10288 16154 10308
rect 16224 10130 16252 10406
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15764 9518 15792 9998
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15846 9276 16154 9296
rect 15846 9274 15852 9276
rect 15908 9274 15932 9276
rect 15988 9274 16012 9276
rect 16068 9274 16092 9276
rect 16148 9274 16154 9276
rect 15908 9222 15910 9274
rect 16090 9222 16092 9274
rect 15846 9220 15852 9222
rect 15908 9220 15932 9222
rect 15988 9220 16012 9222
rect 16068 9220 16092 9222
rect 16148 9220 16154 9222
rect 15846 9200 16154 9220
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14568 8634 14596 8774
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14660 8498 14688 8910
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 15488 8430 15516 8774
rect 15580 8430 15608 8774
rect 16408 8634 16436 15982
rect 16592 15910 16620 16594
rect 16684 15978 16712 17138
rect 16868 17134 16896 19654
rect 16960 18290 16988 22374
rect 17130 22335 17186 22344
rect 17040 22160 17092 22166
rect 17040 22102 17092 22108
rect 17052 21146 17080 22102
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17052 19446 17080 20402
rect 17144 20262 17172 22335
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17236 22098 17264 22170
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17328 22030 17356 22494
rect 17406 22264 17462 22273
rect 17406 22199 17462 22208
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17224 20868 17276 20874
rect 17224 20810 17276 20816
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 17144 18698 17172 19790
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17144 18426 17172 18634
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 17144 17660 17172 18362
rect 17236 18290 17264 20810
rect 17420 20330 17448 22199
rect 17500 22092 17552 22098
rect 17500 22034 17552 22040
rect 17408 20324 17460 20330
rect 17408 20266 17460 20272
rect 17420 20058 17448 20266
rect 17316 20052 17368 20058
rect 17316 19994 17368 20000
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17328 19378 17356 19994
rect 17512 19922 17540 22034
rect 17604 21554 17632 23462
rect 17696 22438 17724 25486
rect 17776 25356 17828 25362
rect 17776 25298 17828 25304
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 17328 18766 17356 19314
rect 17512 18834 17540 19858
rect 17604 19854 17632 21490
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17788 19718 17816 25298
rect 17880 25294 17908 25842
rect 17868 25288 17920 25294
rect 17868 25230 17920 25236
rect 17880 24206 17908 25230
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17880 22094 17908 24142
rect 17972 23730 18000 26318
rect 18064 26042 18092 29106
rect 18052 26036 18104 26042
rect 18052 25978 18104 25984
rect 18050 25936 18106 25945
rect 18050 25871 18052 25880
rect 18104 25871 18106 25880
rect 18052 25842 18104 25848
rect 18064 24954 18092 25842
rect 18052 24948 18104 24954
rect 18052 24890 18104 24896
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 17880 22066 18000 22094
rect 17866 21720 17922 21729
rect 17866 21655 17922 21664
rect 17880 21554 17908 21655
rect 17972 21554 18000 22066
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 17972 20942 18000 21490
rect 18064 21010 18092 24686
rect 18156 22094 18184 29582
rect 18248 29238 18276 30194
rect 18236 29232 18288 29238
rect 18236 29174 18288 29180
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18248 27656 18276 28494
rect 18340 27962 18368 31758
rect 18432 31346 18460 37606
rect 18524 35290 18552 37946
rect 18616 36281 18644 40310
rect 18800 39522 18828 42094
rect 18800 39494 18920 39522
rect 18788 39364 18840 39370
rect 18788 39306 18840 39312
rect 18696 38208 18748 38214
rect 18696 38150 18748 38156
rect 18708 37942 18736 38150
rect 18696 37936 18748 37942
rect 18696 37878 18748 37884
rect 18800 37398 18828 39306
rect 18788 37392 18840 37398
rect 18788 37334 18840 37340
rect 18696 37188 18748 37194
rect 18696 37130 18748 37136
rect 18602 36272 18658 36281
rect 18602 36207 18658 36216
rect 18604 36168 18656 36174
rect 18604 36110 18656 36116
rect 18512 35284 18564 35290
rect 18512 35226 18564 35232
rect 18510 35184 18566 35193
rect 18510 35119 18566 35128
rect 18524 34610 18552 35119
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 18524 33522 18552 33798
rect 18512 33516 18564 33522
rect 18512 33458 18564 33464
rect 18512 31884 18564 31890
rect 18512 31826 18564 31832
rect 18524 31498 18552 31826
rect 18616 31754 18644 36110
rect 18708 36038 18736 37130
rect 18800 36650 18828 37334
rect 18788 36644 18840 36650
rect 18788 36586 18840 36592
rect 18696 36032 18748 36038
rect 18696 35974 18748 35980
rect 18892 35714 18920 39494
rect 18708 35686 18920 35714
rect 18708 34490 18736 35686
rect 18880 35624 18932 35630
rect 18880 35566 18932 35572
rect 18892 35222 18920 35566
rect 18880 35216 18932 35222
rect 18800 35176 18880 35204
rect 18800 34678 18828 35176
rect 18984 35193 19012 44134
rect 19064 43104 19116 43110
rect 19064 43046 19116 43052
rect 19076 42362 19104 43046
rect 19064 42356 19116 42362
rect 19064 42298 19116 42304
rect 19064 41608 19116 41614
rect 19064 41550 19116 41556
rect 19076 36174 19104 41550
rect 19260 41478 19288 44950
rect 19352 44742 19380 45358
rect 19444 45342 19564 45370
rect 19432 45280 19484 45286
rect 19432 45222 19484 45228
rect 19340 44736 19392 44742
rect 19340 44678 19392 44684
rect 19352 44402 19380 44678
rect 19340 44396 19392 44402
rect 19340 44338 19392 44344
rect 19352 43858 19380 44338
rect 19444 44334 19472 45222
rect 19432 44328 19484 44334
rect 19432 44270 19484 44276
rect 19444 43994 19472 44270
rect 19432 43988 19484 43994
rect 19432 43930 19484 43936
rect 19340 43852 19392 43858
rect 19340 43794 19392 43800
rect 19536 43382 19564 45342
rect 19616 45280 19668 45286
rect 19616 45222 19668 45228
rect 19524 43376 19576 43382
rect 19524 43318 19576 43324
rect 19628 43314 19656 45222
rect 19984 44940 20036 44946
rect 19984 44882 20036 44888
rect 19892 44872 19944 44878
rect 19892 44814 19944 44820
rect 19904 44470 19932 44814
rect 19892 44464 19944 44470
rect 19720 44412 19892 44418
rect 19720 44406 19944 44412
rect 19720 44402 19932 44406
rect 19708 44396 19932 44402
rect 19760 44390 19932 44396
rect 19708 44338 19760 44344
rect 19996 43654 20024 44882
rect 20076 44736 20128 44742
rect 20076 44678 20128 44684
rect 20088 43790 20116 44678
rect 20076 43784 20128 43790
rect 20076 43726 20128 43732
rect 19984 43648 20036 43654
rect 19984 43590 20036 43596
rect 19616 43308 19668 43314
rect 19616 43250 19668 43256
rect 19338 42392 19394 42401
rect 19338 42327 19394 42336
rect 19352 42158 19380 42327
rect 19432 42288 19484 42294
rect 19430 42256 19432 42265
rect 19484 42256 19486 42265
rect 19430 42191 19486 42200
rect 19524 42220 19576 42226
rect 19524 42162 19576 42168
rect 19340 42152 19392 42158
rect 19340 42094 19392 42100
rect 19248 41472 19300 41478
rect 19248 41414 19300 41420
rect 19536 41256 19564 42162
rect 19628 41546 19656 43250
rect 19708 43104 19760 43110
rect 19708 43046 19760 43052
rect 19720 42906 19748 43046
rect 19708 42900 19760 42906
rect 19708 42842 19760 42848
rect 20076 42696 20128 42702
rect 20076 42638 20128 42644
rect 19800 42560 19852 42566
rect 19800 42502 19852 42508
rect 19812 42294 19840 42502
rect 19890 42392 19946 42401
rect 19890 42327 19946 42336
rect 19708 42288 19760 42294
rect 19708 42230 19760 42236
rect 19800 42288 19852 42294
rect 19800 42230 19852 42236
rect 19720 42072 19748 42230
rect 19904 42226 19932 42327
rect 19892 42220 19944 42226
rect 19892 42162 19944 42168
rect 19984 42220 20036 42226
rect 19984 42162 20036 42168
rect 19892 42084 19944 42090
rect 19720 42044 19892 42072
rect 19892 42026 19944 42032
rect 19996 41750 20024 42162
rect 19984 41744 20036 41750
rect 19984 41686 20036 41692
rect 20088 41682 20116 42638
rect 20076 41676 20128 41682
rect 20076 41618 20128 41624
rect 19616 41540 19668 41546
rect 19616 41482 19668 41488
rect 19536 41228 19932 41256
rect 19798 41168 19854 41177
rect 19248 41132 19300 41138
rect 19798 41103 19854 41112
rect 19248 41074 19300 41080
rect 19260 40730 19288 41074
rect 19524 40996 19576 41002
rect 19524 40938 19576 40944
rect 19248 40724 19300 40730
rect 19248 40666 19300 40672
rect 19536 40662 19564 40938
rect 19708 40724 19760 40730
rect 19708 40666 19760 40672
rect 19524 40656 19576 40662
rect 19524 40598 19576 40604
rect 19614 40488 19670 40497
rect 19614 40423 19670 40432
rect 19628 40390 19656 40423
rect 19616 40384 19668 40390
rect 19616 40326 19668 40332
rect 19720 40118 19748 40666
rect 19812 40526 19840 41103
rect 19800 40520 19852 40526
rect 19800 40462 19852 40468
rect 19708 40112 19760 40118
rect 19708 40054 19760 40060
rect 19524 40044 19576 40050
rect 19524 39986 19576 39992
rect 19156 39296 19208 39302
rect 19156 39238 19208 39244
rect 19168 38962 19196 39238
rect 19536 38962 19564 39986
rect 19708 39976 19760 39982
rect 19708 39918 19760 39924
rect 19614 39672 19670 39681
rect 19614 39607 19616 39616
rect 19668 39607 19670 39616
rect 19616 39578 19668 39584
rect 19720 39574 19748 39918
rect 19708 39568 19760 39574
rect 19708 39510 19760 39516
rect 19156 38956 19208 38962
rect 19156 38898 19208 38904
rect 19524 38956 19576 38962
rect 19524 38898 19576 38904
rect 19720 38894 19748 39510
rect 19708 38888 19760 38894
rect 19708 38830 19760 38836
rect 19616 38480 19668 38486
rect 19616 38422 19668 38428
rect 19628 37670 19656 38422
rect 19616 37664 19668 37670
rect 19616 37606 19668 37612
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 19260 36854 19288 37198
rect 19432 36916 19484 36922
rect 19432 36858 19484 36864
rect 19248 36848 19300 36854
rect 19248 36790 19300 36796
rect 19444 36718 19472 36858
rect 19432 36712 19484 36718
rect 19432 36654 19484 36660
rect 19156 36372 19208 36378
rect 19156 36314 19208 36320
rect 19064 36168 19116 36174
rect 19064 36110 19116 36116
rect 19064 36032 19116 36038
rect 19064 35974 19116 35980
rect 18880 35158 18932 35164
rect 18970 35184 19026 35193
rect 18970 35119 19026 35128
rect 19076 35086 19104 35974
rect 19064 35080 19116 35086
rect 19062 35048 19064 35057
rect 19116 35048 19118 35057
rect 19062 34983 19118 34992
rect 18788 34672 18840 34678
rect 18788 34614 18840 34620
rect 18880 34604 18932 34610
rect 18880 34546 18932 34552
rect 18708 34462 18828 34490
rect 18800 31929 18828 34462
rect 18892 32774 18920 34546
rect 19168 34542 19196 36314
rect 19444 35698 19472 36654
rect 19524 36644 19576 36650
rect 19524 36586 19576 36592
rect 19432 35692 19484 35698
rect 19432 35634 19484 35640
rect 19248 34672 19300 34678
rect 19248 34614 19300 34620
rect 19156 34536 19208 34542
rect 18970 34504 19026 34513
rect 19156 34478 19208 34484
rect 18970 34439 19026 34448
rect 18880 32768 18932 32774
rect 18880 32710 18932 32716
rect 18786 31920 18842 31929
rect 18786 31855 18842 31864
rect 18604 31748 18656 31754
rect 18604 31690 18656 31696
rect 18524 31470 18736 31498
rect 18420 31340 18472 31346
rect 18420 31282 18472 31288
rect 18512 31272 18564 31278
rect 18512 31214 18564 31220
rect 18420 30660 18472 30666
rect 18420 30602 18472 30608
rect 18432 28694 18460 30602
rect 18524 30161 18552 31214
rect 18604 31136 18656 31142
rect 18604 31078 18656 31084
rect 18510 30152 18566 30161
rect 18510 30087 18566 30096
rect 18512 30048 18564 30054
rect 18512 29990 18564 29996
rect 18420 28688 18472 28694
rect 18420 28630 18472 28636
rect 18432 28082 18460 28630
rect 18524 28121 18552 29990
rect 18510 28112 18566 28121
rect 18420 28076 18472 28082
rect 18510 28047 18566 28056
rect 18420 28018 18472 28024
rect 18340 27934 18552 27962
rect 18420 27668 18472 27674
rect 18248 27628 18368 27656
rect 18236 27532 18288 27538
rect 18236 27474 18288 27480
rect 18248 27062 18276 27474
rect 18340 27470 18368 27628
rect 18420 27610 18472 27616
rect 18328 27464 18380 27470
rect 18328 27406 18380 27412
rect 18236 27056 18288 27062
rect 18236 26998 18288 27004
rect 18236 26920 18288 26926
rect 18236 26862 18288 26868
rect 18248 26234 18276 26862
rect 18340 26858 18368 27406
rect 18328 26852 18380 26858
rect 18328 26794 18380 26800
rect 18432 26382 18460 27610
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18248 26206 18460 26234
rect 18328 25832 18380 25838
rect 18328 25774 18380 25780
rect 18340 25430 18368 25774
rect 18328 25424 18380 25430
rect 18328 25366 18380 25372
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18248 24138 18276 24754
rect 18236 24132 18288 24138
rect 18236 24074 18288 24080
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 18340 23322 18368 23734
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18156 22066 18276 22094
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 18156 21418 18184 21966
rect 18144 21412 18196 21418
rect 18144 21354 18196 21360
rect 18248 21078 18276 22066
rect 18236 21072 18288 21078
rect 18236 21014 18288 21020
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17972 19854 18000 20878
rect 18248 20806 18276 21014
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 18340 20466 18368 23054
rect 18432 22506 18460 26206
rect 18420 22500 18472 22506
rect 18420 22442 18472 22448
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 17684 19236 17736 19242
rect 17684 19178 17736 19184
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17328 18170 17356 18702
rect 17052 17632 17172 17660
rect 17236 18142 17356 18170
rect 17052 17270 17080 17632
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17144 17338 17172 17478
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 17040 17264 17092 17270
rect 17040 17206 17092 17212
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 17052 16250 17080 17206
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16672 15972 16724 15978
rect 16672 15914 16724 15920
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 16592 15570 16620 15846
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16592 15450 16620 15506
rect 16500 15422 16620 15450
rect 16500 14482 16528 15422
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16592 14618 16620 15302
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16592 12986 16620 13874
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11898 16528 12106
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16500 11218 16528 11834
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16592 10266 16620 12242
rect 16684 11762 16712 14758
rect 16776 14618 16804 14894
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16960 14074 16988 16050
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 17144 14822 17172 15438
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16868 11354 16896 12718
rect 17052 12170 17080 12854
rect 17236 12434 17264 18142
rect 17512 17134 17540 18770
rect 17696 18630 17724 19178
rect 17788 18766 17816 19314
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17696 18426 17724 18566
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17512 16046 17540 17070
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17328 13870 17356 14554
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17144 12406 17264 12434
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16960 11762 16988 12038
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16960 10062 16988 10610
rect 17144 10062 17172 12406
rect 17328 12306 17356 13806
rect 17512 13530 17540 13874
rect 17788 13784 17816 18702
rect 17868 18692 17920 18698
rect 17868 18634 17920 18640
rect 17880 17542 17908 18634
rect 17972 18290 18000 19110
rect 18064 18766 18092 19314
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 18248 17610 18276 18566
rect 18340 18358 18368 20402
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 18340 17678 18368 18294
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17880 17202 17908 17478
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 18052 16176 18104 16182
rect 18052 16118 18104 16124
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17972 14414 18000 14894
rect 18064 14550 18092 16118
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18156 14618 18184 15098
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 17960 14408 18012 14414
rect 18012 14368 18092 14396
rect 17960 14350 18012 14356
rect 17788 13756 18000 13784
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17972 13258 18000 13756
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 17972 12442 18000 13194
rect 18064 12850 18092 14368
rect 18248 13462 18276 15506
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18340 14414 18368 14486
rect 18328 14408 18380 14414
rect 18328 14350 18380 14356
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 18248 12850 18276 13398
rect 18340 12986 18368 14350
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18432 12918 18460 21966
rect 18524 16454 18552 27934
rect 18616 26568 18644 31078
rect 18708 30258 18736 31470
rect 18892 30666 18920 32710
rect 18880 30660 18932 30666
rect 18880 30602 18932 30608
rect 18878 30560 18934 30569
rect 18878 30495 18934 30504
rect 18696 30252 18748 30258
rect 18696 30194 18748 30200
rect 18788 30252 18840 30258
rect 18788 30194 18840 30200
rect 18694 30152 18750 30161
rect 18694 30087 18750 30096
rect 18708 26926 18736 30087
rect 18800 29850 18828 30194
rect 18788 29844 18840 29850
rect 18788 29786 18840 29792
rect 18892 28626 18920 30495
rect 18880 28620 18932 28626
rect 18880 28562 18932 28568
rect 18788 28416 18840 28422
rect 18788 28358 18840 28364
rect 18696 26920 18748 26926
rect 18696 26862 18748 26868
rect 18616 26540 18736 26568
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18616 21962 18644 22986
rect 18604 21956 18656 21962
rect 18604 21898 18656 21904
rect 18708 21729 18736 26540
rect 18800 22545 18828 28358
rect 18892 26994 18920 28562
rect 18984 28393 19012 34439
rect 19168 34134 19196 34478
rect 19260 34474 19288 34614
rect 19340 34604 19392 34610
rect 19340 34546 19392 34552
rect 19248 34468 19300 34474
rect 19248 34410 19300 34416
rect 19156 34128 19208 34134
rect 19156 34070 19208 34076
rect 19260 33998 19288 34410
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19352 33862 19380 34546
rect 19248 33856 19300 33862
rect 19248 33798 19300 33804
rect 19340 33856 19392 33862
rect 19444 33844 19472 35634
rect 19536 34950 19564 36586
rect 19800 36372 19852 36378
rect 19800 36314 19852 36320
rect 19616 36236 19668 36242
rect 19616 36178 19668 36184
rect 19628 35698 19656 36178
rect 19616 35692 19668 35698
rect 19616 35634 19668 35640
rect 19628 35290 19656 35634
rect 19708 35624 19760 35630
rect 19708 35566 19760 35572
rect 19616 35284 19668 35290
rect 19616 35226 19668 35232
rect 19720 35154 19748 35566
rect 19812 35562 19840 36314
rect 19904 35578 19932 41228
rect 19984 38956 20036 38962
rect 19984 38898 20036 38904
rect 19996 37874 20024 38898
rect 20088 38554 20116 41618
rect 20180 40526 20208 47200
rect 20916 47138 20944 47200
rect 21008 47138 21036 47246
rect 20916 47110 21036 47138
rect 20811 45724 21119 45744
rect 20811 45722 20817 45724
rect 20873 45722 20897 45724
rect 20953 45722 20977 45724
rect 21033 45722 21057 45724
rect 21113 45722 21119 45724
rect 20873 45670 20875 45722
rect 21055 45670 21057 45722
rect 20811 45668 20817 45670
rect 20873 45668 20897 45670
rect 20953 45668 20977 45670
rect 21033 45668 21057 45670
rect 21113 45668 21119 45670
rect 20811 45648 21119 45668
rect 20996 45552 21048 45558
rect 20996 45494 21048 45500
rect 20536 45484 20588 45490
rect 20536 45426 20588 45432
rect 20444 45416 20496 45422
rect 20444 45358 20496 45364
rect 20260 44396 20312 44402
rect 20260 44338 20312 44344
rect 20272 43722 20300 44338
rect 20352 44328 20404 44334
rect 20352 44270 20404 44276
rect 20364 43790 20392 44270
rect 20456 44198 20484 45358
rect 20444 44192 20496 44198
rect 20444 44134 20496 44140
rect 20456 43994 20484 44134
rect 20444 43988 20496 43994
rect 20444 43930 20496 43936
rect 20352 43784 20404 43790
rect 20352 43726 20404 43732
rect 20260 43716 20312 43722
rect 20260 43658 20312 43664
rect 20272 40730 20300 43658
rect 20260 40724 20312 40730
rect 20260 40666 20312 40672
rect 20364 40662 20392 43726
rect 20352 40656 20404 40662
rect 20352 40598 20404 40604
rect 20168 40520 20220 40526
rect 20168 40462 20220 40468
rect 20168 39840 20220 39846
rect 20168 39782 20220 39788
rect 20076 38548 20128 38554
rect 20076 38490 20128 38496
rect 19984 37868 20036 37874
rect 19984 37810 20036 37816
rect 19996 37330 20024 37810
rect 20088 37330 20116 38490
rect 20180 38282 20208 39782
rect 20352 39296 20404 39302
rect 20352 39238 20404 39244
rect 20364 39001 20392 39238
rect 20350 38992 20406 39001
rect 20350 38927 20406 38936
rect 20168 38276 20220 38282
rect 20168 38218 20220 38224
rect 20456 37942 20484 43930
rect 20548 43092 20576 45426
rect 21008 45393 21036 45494
rect 21088 45484 21140 45490
rect 21088 45426 21140 45432
rect 20994 45384 21050 45393
rect 20994 45319 21050 45328
rect 20628 45280 20680 45286
rect 20628 45222 20680 45228
rect 20996 45280 21048 45286
rect 20996 45222 21048 45228
rect 20640 43722 20668 45222
rect 20720 45076 20772 45082
rect 20720 45018 20772 45024
rect 20732 44305 20760 45018
rect 21008 44878 21036 45222
rect 21100 45082 21128 45426
rect 21088 45076 21140 45082
rect 21088 45018 21140 45024
rect 20996 44872 21048 44878
rect 20994 44840 20996 44849
rect 21048 44840 21050 44849
rect 21192 44826 21220 47246
rect 21730 47200 21786 48000
rect 22466 47200 22522 48000
rect 23202 47200 23258 48000
rect 23938 47200 23994 48000
rect 24766 47200 24822 48000
rect 24964 47246 25452 47274
rect 21456 45552 21508 45558
rect 21454 45520 21456 45529
rect 21508 45520 21510 45529
rect 21744 45490 21772 47200
rect 21454 45455 21510 45464
rect 21732 45484 21784 45490
rect 21732 45426 21784 45432
rect 22376 45076 22428 45082
rect 22376 45018 22428 45024
rect 22192 45008 22244 45014
rect 21454 44976 21510 44985
rect 21454 44911 21456 44920
rect 21508 44911 21510 44920
rect 22006 44976 22062 44985
rect 22006 44911 22062 44920
rect 22190 44976 22192 44985
rect 22244 44976 22246 44985
rect 22388 44946 22416 45018
rect 22480 44946 22508 47200
rect 23216 45422 23244 47200
rect 23296 45824 23348 45830
rect 23296 45766 23348 45772
rect 23204 45416 23256 45422
rect 23204 45358 23256 45364
rect 22190 44911 22246 44920
rect 22376 44940 22428 44946
rect 21456 44882 21508 44888
rect 21916 44872 21968 44878
rect 21192 44798 21404 44826
rect 21916 44814 21968 44820
rect 20994 44775 21050 44784
rect 21272 44736 21324 44742
rect 21272 44678 21324 44684
rect 20811 44636 21119 44656
rect 20811 44634 20817 44636
rect 20873 44634 20897 44636
rect 20953 44634 20977 44636
rect 21033 44634 21057 44636
rect 21113 44634 21119 44636
rect 20873 44582 20875 44634
rect 21055 44582 21057 44634
rect 20811 44580 20817 44582
rect 20873 44580 20897 44582
rect 20953 44580 20977 44582
rect 21033 44580 21057 44582
rect 21113 44580 21119 44582
rect 20811 44560 21119 44580
rect 21180 44396 21232 44402
rect 21180 44338 21232 44344
rect 20812 44328 20864 44334
rect 20718 44296 20774 44305
rect 20812 44270 20864 44276
rect 20718 44231 20774 44240
rect 20720 44192 20772 44198
rect 20720 44134 20772 44140
rect 20628 43716 20680 43722
rect 20628 43658 20680 43664
rect 20732 43178 20760 44134
rect 20824 43790 20852 44270
rect 20812 43784 20864 43790
rect 20812 43726 20864 43732
rect 21088 43784 21140 43790
rect 21192 43772 21220 44338
rect 21284 43790 21312 44678
rect 21140 43744 21220 43772
rect 21088 43726 21140 43732
rect 20811 43548 21119 43568
rect 20811 43546 20817 43548
rect 20873 43546 20897 43548
rect 20953 43546 20977 43548
rect 21033 43546 21057 43548
rect 21113 43546 21119 43548
rect 20873 43494 20875 43546
rect 21055 43494 21057 43546
rect 20811 43492 20817 43494
rect 20873 43492 20897 43494
rect 20953 43492 20977 43494
rect 21033 43492 21057 43494
rect 21113 43492 21119 43494
rect 20811 43472 21119 43492
rect 21192 43450 21220 43744
rect 21272 43784 21324 43790
rect 21272 43726 21324 43732
rect 21180 43444 21232 43450
rect 21180 43386 21232 43392
rect 21180 43308 21232 43314
rect 21284 43296 21312 43726
rect 21232 43268 21312 43296
rect 21180 43250 21232 43256
rect 20720 43172 20772 43178
rect 20720 43114 20772 43120
rect 20628 43104 20680 43110
rect 20548 43064 20628 43092
rect 20628 43046 20680 43052
rect 20628 42696 20680 42702
rect 20628 42638 20680 42644
rect 20640 42362 20668 42638
rect 21180 42628 21232 42634
rect 21180 42570 21232 42576
rect 20811 42460 21119 42480
rect 20811 42458 20817 42460
rect 20873 42458 20897 42460
rect 20953 42458 20977 42460
rect 21033 42458 21057 42460
rect 21113 42458 21119 42460
rect 20873 42406 20875 42458
rect 21055 42406 21057 42458
rect 20811 42404 20817 42406
rect 20873 42404 20897 42406
rect 20953 42404 20977 42406
rect 21033 42404 21057 42406
rect 21113 42404 21119 42406
rect 20811 42384 21119 42404
rect 21192 42362 21220 42570
rect 20628 42356 20680 42362
rect 20628 42298 20680 42304
rect 21180 42356 21232 42362
rect 21180 42298 21232 42304
rect 20626 42256 20682 42265
rect 20626 42191 20628 42200
rect 20680 42191 20682 42200
rect 21178 42256 21234 42265
rect 21178 42191 21234 42200
rect 21272 42220 21324 42226
rect 20628 42162 20680 42168
rect 20626 42120 20682 42129
rect 20626 42055 20682 42064
rect 20536 40044 20588 40050
rect 20536 39986 20588 39992
rect 20548 38826 20576 39986
rect 20536 38820 20588 38826
rect 20536 38762 20588 38768
rect 20548 38350 20576 38762
rect 20640 38654 20668 42055
rect 21088 42016 21140 42022
rect 21088 41958 21140 41964
rect 21100 41750 21128 41958
rect 21088 41744 21140 41750
rect 21088 41686 21140 41692
rect 20720 41472 20772 41478
rect 20720 41414 20772 41420
rect 20732 41070 20760 41414
rect 20811 41372 21119 41392
rect 20811 41370 20817 41372
rect 20873 41370 20897 41372
rect 20953 41370 20977 41372
rect 21033 41370 21057 41372
rect 21113 41370 21119 41372
rect 20873 41318 20875 41370
rect 21055 41318 21057 41370
rect 20811 41316 20817 41318
rect 20873 41316 20897 41318
rect 20953 41316 20977 41318
rect 21033 41316 21057 41318
rect 21113 41316 21119 41318
rect 20811 41296 21119 41316
rect 21192 41070 21220 42191
rect 21272 42162 21324 42168
rect 21284 41818 21312 42162
rect 21272 41812 21324 41818
rect 21272 41754 21324 41760
rect 21284 41614 21312 41754
rect 21272 41608 21324 41614
rect 21272 41550 21324 41556
rect 20720 41064 20772 41070
rect 20720 41006 20772 41012
rect 21180 41064 21232 41070
rect 21180 41006 21232 41012
rect 20720 40928 20772 40934
rect 20720 40870 20772 40876
rect 20732 40730 20760 40870
rect 20720 40724 20772 40730
rect 20720 40666 20772 40672
rect 21180 40656 21232 40662
rect 21180 40598 21232 40604
rect 20811 40284 21119 40304
rect 20811 40282 20817 40284
rect 20873 40282 20897 40284
rect 20953 40282 20977 40284
rect 21033 40282 21057 40284
rect 21113 40282 21119 40284
rect 20873 40230 20875 40282
rect 21055 40230 21057 40282
rect 20811 40228 20817 40230
rect 20873 40228 20897 40230
rect 20953 40228 20977 40230
rect 21033 40228 21057 40230
rect 21113 40228 21119 40230
rect 20811 40208 21119 40228
rect 20904 40112 20956 40118
rect 20904 40054 20956 40060
rect 20916 39846 20944 40054
rect 20904 39840 20956 39846
rect 20904 39782 20956 39788
rect 20720 39364 20772 39370
rect 20720 39306 20772 39312
rect 20732 39098 20760 39306
rect 20811 39196 21119 39216
rect 20811 39194 20817 39196
rect 20873 39194 20897 39196
rect 20953 39194 20977 39196
rect 21033 39194 21057 39196
rect 21113 39194 21119 39196
rect 20873 39142 20875 39194
rect 21055 39142 21057 39194
rect 20811 39140 20817 39142
rect 20873 39140 20897 39142
rect 20953 39140 20977 39142
rect 21033 39140 21057 39142
rect 21113 39140 21119 39142
rect 20811 39120 21119 39140
rect 20720 39092 20772 39098
rect 20720 39034 20772 39040
rect 21192 39030 21220 40598
rect 21376 40526 21404 44798
rect 21456 44804 21508 44810
rect 21456 44746 21508 44752
rect 21640 44804 21692 44810
rect 21640 44746 21692 44752
rect 21468 44441 21496 44746
rect 21454 44432 21510 44441
rect 21652 44402 21680 44746
rect 21454 44367 21510 44376
rect 21640 44396 21692 44402
rect 21468 42129 21496 44367
rect 21640 44338 21692 44344
rect 21732 44328 21784 44334
rect 21732 44270 21784 44276
rect 21744 44198 21772 44270
rect 21732 44192 21784 44198
rect 21546 44160 21602 44169
rect 21732 44134 21784 44140
rect 21546 44095 21602 44104
rect 21560 42265 21588 44095
rect 21546 42256 21602 42265
rect 21546 42191 21602 42200
rect 21548 42152 21600 42158
rect 21454 42120 21510 42129
rect 21548 42094 21600 42100
rect 21454 42055 21510 42064
rect 21456 41472 21508 41478
rect 21456 41414 21508 41420
rect 21468 41002 21496 41414
rect 21456 40996 21508 41002
rect 21456 40938 21508 40944
rect 21364 40520 21416 40526
rect 21364 40462 21416 40468
rect 21272 40452 21324 40458
rect 21272 40394 21324 40400
rect 21284 40050 21312 40394
rect 21364 40384 21416 40390
rect 21364 40326 21416 40332
rect 21272 40044 21324 40050
rect 21272 39986 21324 39992
rect 21272 39840 21324 39846
rect 21272 39782 21324 39788
rect 21180 39024 21232 39030
rect 21180 38966 21232 38972
rect 20640 38626 20760 38654
rect 20536 38344 20588 38350
rect 20536 38286 20588 38292
rect 20444 37936 20496 37942
rect 20444 37878 20496 37884
rect 20352 37800 20404 37806
rect 20352 37742 20404 37748
rect 20444 37800 20496 37806
rect 20548 37754 20576 38286
rect 20628 37868 20680 37874
rect 20628 37810 20680 37816
rect 20496 37748 20576 37754
rect 20444 37742 20576 37748
rect 19984 37324 20036 37330
rect 19984 37266 20036 37272
rect 20076 37324 20128 37330
rect 20076 37266 20128 37272
rect 20088 36242 20116 37266
rect 20076 36236 20128 36242
rect 20076 36178 20128 36184
rect 19984 35760 20036 35766
rect 19982 35728 19984 35737
rect 20036 35728 20038 35737
rect 19982 35663 20038 35672
rect 19800 35556 19852 35562
rect 19904 35550 20024 35578
rect 19800 35498 19852 35504
rect 19708 35148 19760 35154
rect 19708 35090 19760 35096
rect 19800 35148 19852 35154
rect 19800 35090 19852 35096
rect 19614 35048 19670 35057
rect 19614 34983 19670 34992
rect 19524 34944 19576 34950
rect 19524 34886 19576 34892
rect 19536 34610 19564 34886
rect 19628 34678 19656 34983
rect 19616 34672 19668 34678
rect 19616 34614 19668 34620
rect 19524 34604 19576 34610
rect 19524 34546 19576 34552
rect 19524 34400 19576 34406
rect 19524 34342 19576 34348
rect 19536 33998 19564 34342
rect 19524 33992 19576 33998
rect 19524 33934 19576 33940
rect 19616 33856 19668 33862
rect 19444 33816 19564 33844
rect 19340 33798 19392 33804
rect 19260 33674 19288 33798
rect 19260 33646 19472 33674
rect 19248 32972 19300 32978
rect 19248 32914 19300 32920
rect 19260 32434 19288 32914
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 19248 31748 19300 31754
rect 19248 31690 19300 31696
rect 19064 31340 19116 31346
rect 19064 31282 19116 31288
rect 19076 28558 19104 31282
rect 19260 30190 19288 31690
rect 19340 31340 19392 31346
rect 19340 31282 19392 31288
rect 19352 30734 19380 31282
rect 19340 30728 19392 30734
rect 19338 30696 19340 30705
rect 19392 30696 19394 30705
rect 19338 30631 19394 30640
rect 19248 30184 19300 30190
rect 19248 30126 19300 30132
rect 19444 30122 19472 33646
rect 19536 30258 19564 33816
rect 19616 33798 19668 33804
rect 19628 32910 19656 33798
rect 19720 33658 19748 35090
rect 19812 34610 19840 35090
rect 19800 34604 19852 34610
rect 19800 34546 19852 34552
rect 19812 33998 19840 34546
rect 19800 33992 19852 33998
rect 19800 33934 19852 33940
rect 19708 33652 19760 33658
rect 19708 33594 19760 33600
rect 19708 33516 19760 33522
rect 19708 33458 19760 33464
rect 19616 32904 19668 32910
rect 19616 32846 19668 32852
rect 19720 32756 19748 33458
rect 19628 32728 19748 32756
rect 19628 32230 19656 32728
rect 19616 32224 19668 32230
rect 19616 32166 19668 32172
rect 19524 30252 19576 30258
rect 19524 30194 19576 30200
rect 19432 30116 19484 30122
rect 19432 30058 19484 30064
rect 19156 29776 19208 29782
rect 19156 29718 19208 29724
rect 19168 29345 19196 29718
rect 19432 29640 19484 29646
rect 19432 29582 19484 29588
rect 19444 29458 19472 29582
rect 19524 29504 19576 29510
rect 19444 29452 19524 29458
rect 19444 29446 19576 29452
rect 19444 29430 19564 29446
rect 19154 29336 19210 29345
rect 19154 29271 19210 29280
rect 19444 29170 19472 29430
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 19168 28665 19196 28970
rect 19154 28656 19210 28665
rect 19154 28591 19210 28600
rect 19338 28656 19394 28665
rect 19338 28591 19394 28600
rect 19352 28558 19380 28591
rect 19064 28552 19116 28558
rect 19064 28494 19116 28500
rect 19156 28552 19208 28558
rect 19156 28494 19208 28500
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 18970 28384 19026 28393
rect 19168 28370 19196 28494
rect 19340 28416 19392 28422
rect 19338 28384 19340 28393
rect 19392 28384 19394 28393
rect 19168 28342 19288 28370
rect 18970 28319 19026 28328
rect 19062 28248 19118 28257
rect 19118 28206 19196 28234
rect 19260 28218 19288 28342
rect 19338 28319 19394 28328
rect 19062 28183 19118 28192
rect 18972 28144 19024 28150
rect 18972 28086 19024 28092
rect 19062 28112 19118 28121
rect 18984 27962 19012 28086
rect 19168 28098 19196 28206
rect 19248 28212 19300 28218
rect 19248 28154 19300 28160
rect 19338 28112 19394 28121
rect 19168 28070 19338 28098
rect 19062 28047 19064 28056
rect 19116 28047 19118 28056
rect 19338 28047 19394 28056
rect 19064 28018 19116 28024
rect 18984 27934 19196 27962
rect 19168 27928 19196 27934
rect 19340 27940 19392 27946
rect 19168 27900 19340 27928
rect 19340 27882 19392 27888
rect 19064 27872 19116 27878
rect 18970 27840 19026 27849
rect 19064 27814 19116 27820
rect 18970 27775 19026 27784
rect 18880 26988 18932 26994
rect 18880 26930 18932 26936
rect 18880 26852 18932 26858
rect 18880 26794 18932 26800
rect 18892 26450 18920 26794
rect 18880 26444 18932 26450
rect 18880 26386 18932 26392
rect 18892 25702 18920 26386
rect 18984 25974 19012 27775
rect 19076 27334 19104 27814
rect 19246 27704 19302 27713
rect 19246 27639 19302 27648
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 19154 27160 19210 27169
rect 19154 27095 19156 27104
rect 19208 27095 19210 27104
rect 19156 27066 19208 27072
rect 19156 26376 19208 26382
rect 19156 26318 19208 26324
rect 18972 25968 19024 25974
rect 18972 25910 19024 25916
rect 18880 25696 18932 25702
rect 18880 25638 18932 25644
rect 18892 25362 18920 25638
rect 18880 25356 18932 25362
rect 18880 25298 18932 25304
rect 18984 25294 19012 25910
rect 19168 25906 19196 26318
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19064 25492 19116 25498
rect 19064 25434 19116 25440
rect 18972 25288 19024 25294
rect 18972 25230 19024 25236
rect 18880 24948 18932 24954
rect 18880 24890 18932 24896
rect 18892 23322 18920 24890
rect 18984 24818 19012 25230
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 19076 24614 19104 25434
rect 19168 25430 19196 25842
rect 19156 25424 19208 25430
rect 19156 25366 19208 25372
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 19168 24682 19196 24754
rect 19156 24676 19208 24682
rect 19156 24618 19208 24624
rect 19064 24608 19116 24614
rect 19064 24550 19116 24556
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18786 22536 18842 22545
rect 18786 22471 18842 22480
rect 18892 22216 18920 22918
rect 18800 22188 18920 22216
rect 18800 22030 18828 22188
rect 19076 22137 19104 23666
rect 19260 22982 19288 27639
rect 19444 27470 19472 29106
rect 19515 28484 19567 28490
rect 19515 28426 19567 28432
rect 19536 28218 19564 28426
rect 19524 28212 19576 28218
rect 19524 28154 19576 28160
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19524 26308 19576 26314
rect 19524 26250 19576 26256
rect 19536 25294 19564 26250
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19352 23730 19380 25094
rect 19444 24954 19472 25162
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 19628 24750 19656 32166
rect 19708 31340 19760 31346
rect 19708 31282 19760 31288
rect 19720 29850 19748 31282
rect 19892 30592 19944 30598
rect 19892 30534 19944 30540
rect 19800 30252 19852 30258
rect 19800 30194 19852 30200
rect 19708 29844 19760 29850
rect 19708 29786 19760 29792
rect 19812 29730 19840 30194
rect 19720 29702 19840 29730
rect 19720 27402 19748 29702
rect 19904 28422 19932 30534
rect 19996 28966 20024 35550
rect 20260 35488 20312 35494
rect 20260 35430 20312 35436
rect 20168 35012 20220 35018
rect 20168 34954 20220 34960
rect 20180 34746 20208 34954
rect 20168 34740 20220 34746
rect 20168 34682 20220 34688
rect 20168 34536 20220 34542
rect 20272 34524 20300 35430
rect 20364 35154 20392 37742
rect 20456 37726 20576 37742
rect 20456 35193 20484 37726
rect 20536 37664 20588 37670
rect 20536 37606 20588 37612
rect 20442 35184 20498 35193
rect 20352 35148 20404 35154
rect 20442 35119 20498 35128
rect 20352 35090 20404 35096
rect 20456 35086 20484 35119
rect 20444 35080 20496 35086
rect 20444 35022 20496 35028
rect 20548 34678 20576 37606
rect 20640 37233 20668 37810
rect 20626 37224 20682 37233
rect 20626 37159 20628 37168
rect 20680 37159 20682 37168
rect 20628 37130 20680 37136
rect 20640 37099 20668 37130
rect 20628 35828 20680 35834
rect 20628 35770 20680 35776
rect 20444 34672 20496 34678
rect 20444 34614 20496 34620
rect 20536 34672 20588 34678
rect 20536 34614 20588 34620
rect 20220 34496 20300 34524
rect 20168 34478 20220 34484
rect 20456 34490 20484 34614
rect 20640 34490 20668 35770
rect 20732 35057 20760 38626
rect 21284 38214 21312 39782
rect 21376 38214 21404 40326
rect 21454 40216 21510 40225
rect 21454 40151 21456 40160
rect 21508 40151 21510 40160
rect 21456 40122 21508 40128
rect 21456 39500 21508 39506
rect 21456 39442 21508 39448
rect 21272 38208 21324 38214
rect 21272 38150 21324 38156
rect 21364 38208 21416 38214
rect 21364 38150 21416 38156
rect 20811 38108 21119 38128
rect 20811 38106 20817 38108
rect 20873 38106 20897 38108
rect 20953 38106 20977 38108
rect 21033 38106 21057 38108
rect 21113 38106 21119 38108
rect 20873 38054 20875 38106
rect 21055 38054 21057 38106
rect 20811 38052 20817 38054
rect 20873 38052 20897 38054
rect 20953 38052 20977 38054
rect 21033 38052 21057 38054
rect 21113 38052 21119 38054
rect 20811 38032 21119 38052
rect 21180 37664 21232 37670
rect 21180 37606 21232 37612
rect 21192 37274 21220 37606
rect 21284 37466 21312 38150
rect 21272 37460 21324 37466
rect 21272 37402 21324 37408
rect 20916 37246 21220 37274
rect 20916 37194 20944 37246
rect 21362 37224 21418 37233
rect 20904 37188 20956 37194
rect 21362 37159 21418 37168
rect 20904 37130 20956 37136
rect 21376 37126 21404 37159
rect 21364 37120 21416 37126
rect 21364 37062 21416 37068
rect 20811 37020 21119 37040
rect 20811 37018 20817 37020
rect 20873 37018 20897 37020
rect 20953 37018 20977 37020
rect 21033 37018 21057 37020
rect 21113 37018 21119 37020
rect 20873 36966 20875 37018
rect 21055 36966 21057 37018
rect 20811 36964 20817 36966
rect 20873 36964 20897 36966
rect 20953 36964 20977 36966
rect 21033 36964 21057 36966
rect 21113 36964 21119 36966
rect 20811 36944 21119 36964
rect 21272 36100 21324 36106
rect 21272 36042 21324 36048
rect 20811 35932 21119 35952
rect 20811 35930 20817 35932
rect 20873 35930 20897 35932
rect 20953 35930 20977 35932
rect 21033 35930 21057 35932
rect 21113 35930 21119 35932
rect 20873 35878 20875 35930
rect 21055 35878 21057 35930
rect 20811 35876 20817 35878
rect 20873 35876 20897 35878
rect 20953 35876 20977 35878
rect 21033 35876 21057 35878
rect 21113 35876 21119 35878
rect 20811 35856 21119 35876
rect 20812 35760 20864 35766
rect 20810 35728 20812 35737
rect 20864 35728 20866 35737
rect 20810 35663 20866 35672
rect 21284 35222 21312 36042
rect 21364 36032 21416 36038
rect 21364 35974 21416 35980
rect 21272 35216 21324 35222
rect 20902 35184 20958 35193
rect 21272 35158 21324 35164
rect 20902 35119 20958 35128
rect 20916 35086 20944 35119
rect 21376 35086 21404 35974
rect 20904 35080 20956 35086
rect 20718 35048 20774 35057
rect 20904 35022 20956 35028
rect 21364 35080 21416 35086
rect 21364 35022 21416 35028
rect 20718 34983 20774 34992
rect 20811 34844 21119 34864
rect 20811 34842 20817 34844
rect 20873 34842 20897 34844
rect 20953 34842 20977 34844
rect 21033 34842 21057 34844
rect 21113 34842 21119 34844
rect 20873 34790 20875 34842
rect 21055 34790 21057 34842
rect 20811 34788 20817 34790
rect 20873 34788 20897 34790
rect 20953 34788 20977 34790
rect 21033 34788 21057 34790
rect 21113 34788 21119 34790
rect 20811 34768 21119 34788
rect 21180 34604 21232 34610
rect 21180 34546 21232 34552
rect 20076 33856 20128 33862
rect 20076 33798 20128 33804
rect 20088 32434 20116 33798
rect 20076 32428 20128 32434
rect 20076 32370 20128 32376
rect 20180 31414 20208 34478
rect 20456 34462 20668 34490
rect 20444 33992 20496 33998
rect 20444 33934 20496 33940
rect 20260 33652 20312 33658
rect 20260 33594 20312 33600
rect 20168 31408 20220 31414
rect 20168 31350 20220 31356
rect 20272 30274 20300 33594
rect 20456 32298 20484 33934
rect 20811 33756 21119 33776
rect 20811 33754 20817 33756
rect 20873 33754 20897 33756
rect 20953 33754 20977 33756
rect 21033 33754 21057 33756
rect 21113 33754 21119 33756
rect 20873 33702 20875 33754
rect 21055 33702 21057 33754
rect 20811 33700 20817 33702
rect 20873 33700 20897 33702
rect 20953 33700 20977 33702
rect 21033 33700 21057 33702
rect 21113 33700 21119 33702
rect 20811 33680 21119 33700
rect 20810 33552 20866 33561
rect 20720 33516 20772 33522
rect 20810 33487 20812 33496
rect 20720 33458 20772 33464
rect 20864 33487 20866 33496
rect 20812 33458 20864 33464
rect 20732 32842 20760 33458
rect 20720 32836 20772 32842
rect 20720 32778 20772 32784
rect 20811 32668 21119 32688
rect 20811 32666 20817 32668
rect 20873 32666 20897 32668
rect 20953 32666 20977 32668
rect 21033 32666 21057 32668
rect 21113 32666 21119 32668
rect 20873 32614 20875 32666
rect 21055 32614 21057 32666
rect 20811 32612 20817 32614
rect 20873 32612 20897 32614
rect 20953 32612 20977 32614
rect 21033 32612 21057 32614
rect 21113 32612 21119 32614
rect 20811 32592 21119 32612
rect 20720 32564 20772 32570
rect 20720 32506 20772 32512
rect 20444 32292 20496 32298
rect 20444 32234 20496 32240
rect 20352 31136 20404 31142
rect 20352 31078 20404 31084
rect 20364 30802 20392 31078
rect 20352 30796 20404 30802
rect 20352 30738 20404 30744
rect 20456 30666 20484 32234
rect 20732 31414 20760 32506
rect 20811 31580 21119 31600
rect 20811 31578 20817 31580
rect 20873 31578 20897 31580
rect 20953 31578 20977 31580
rect 21033 31578 21057 31580
rect 21113 31578 21119 31580
rect 20873 31526 20875 31578
rect 21055 31526 21057 31578
rect 20811 31524 20817 31526
rect 20873 31524 20897 31526
rect 20953 31524 20977 31526
rect 21033 31524 21057 31526
rect 21113 31524 21119 31526
rect 20811 31504 21119 31524
rect 20720 31408 20772 31414
rect 20720 31350 20772 31356
rect 21192 31142 21220 34546
rect 21272 33992 21324 33998
rect 21272 33934 21324 33940
rect 21284 32570 21312 33934
rect 21376 33538 21404 35022
rect 21468 34406 21496 39442
rect 21456 34400 21508 34406
rect 21456 34342 21508 34348
rect 21456 33924 21508 33930
rect 21456 33866 21508 33872
rect 21468 33658 21496 33866
rect 21456 33652 21508 33658
rect 21456 33594 21508 33600
rect 21376 33510 21496 33538
rect 21364 32836 21416 32842
rect 21364 32778 21416 32784
rect 21272 32564 21324 32570
rect 21272 32506 21324 32512
rect 21376 32366 21404 32778
rect 21364 32360 21416 32366
rect 21364 32302 21416 32308
rect 21376 31890 21404 32302
rect 21468 31958 21496 33510
rect 21456 31952 21508 31958
rect 21456 31894 21508 31900
rect 21364 31884 21416 31890
rect 21364 31826 21416 31832
rect 21272 31816 21324 31822
rect 21272 31758 21324 31764
rect 21180 31136 21232 31142
rect 21180 31078 21232 31084
rect 20444 30660 20496 30666
rect 20444 30602 20496 30608
rect 20811 30492 21119 30512
rect 20811 30490 20817 30492
rect 20873 30490 20897 30492
rect 20953 30490 20977 30492
rect 21033 30490 21057 30492
rect 21113 30490 21119 30492
rect 20873 30438 20875 30490
rect 21055 30438 21057 30490
rect 20811 30436 20817 30438
rect 20873 30436 20897 30438
rect 20953 30436 20977 30438
rect 21033 30436 21057 30438
rect 21113 30436 21119 30438
rect 20811 30416 21119 30436
rect 20272 30246 20392 30274
rect 20168 30184 20220 30190
rect 20168 30126 20220 30132
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 20088 29170 20116 29990
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 19984 28960 20036 28966
rect 19984 28902 20036 28908
rect 19892 28416 19944 28422
rect 20180 28393 20208 30126
rect 20272 29306 20300 30126
rect 20364 29646 20392 30246
rect 20720 30252 20772 30258
rect 20720 30194 20772 30200
rect 20444 30116 20496 30122
rect 20444 30058 20496 30064
rect 20352 29640 20404 29646
rect 20352 29582 20404 29588
rect 20260 29300 20312 29306
rect 20260 29242 20312 29248
rect 19892 28358 19944 28364
rect 20166 28384 20222 28393
rect 19904 28082 19932 28358
rect 20166 28319 20222 28328
rect 19982 28112 20038 28121
rect 19892 28076 19944 28082
rect 19982 28047 20038 28056
rect 19892 28018 19944 28024
rect 19800 27872 19852 27878
rect 19800 27814 19852 27820
rect 19708 27396 19760 27402
rect 19708 27338 19760 27344
rect 19708 25152 19760 25158
rect 19708 25094 19760 25100
rect 19720 24818 19748 25094
rect 19708 24812 19760 24818
rect 19708 24754 19760 24760
rect 19616 24744 19668 24750
rect 19616 24686 19668 24692
rect 19432 24676 19484 24682
rect 19432 24618 19484 24624
rect 19444 24070 19472 24618
rect 19812 24342 19840 27814
rect 19892 27464 19944 27470
rect 19892 27406 19944 27412
rect 19904 27062 19932 27406
rect 19892 27056 19944 27062
rect 19892 26998 19944 27004
rect 19800 24336 19852 24342
rect 19800 24278 19852 24284
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 19062 22128 19118 22137
rect 19062 22063 19118 22072
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 18694 21720 18750 21729
rect 18694 21655 18750 21664
rect 18970 21584 19026 21593
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18788 21548 18840 21554
rect 18970 21519 19026 21528
rect 18788 21490 18840 21496
rect 18616 20874 18644 21490
rect 18800 21078 18828 21490
rect 18984 21486 19012 21519
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 18604 20868 18656 20874
rect 18604 20810 18656 20816
rect 18788 20868 18840 20874
rect 18788 20810 18840 20816
rect 18800 19854 18828 20810
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18524 15706 18552 16050
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18524 14618 18552 14962
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18616 14498 18644 14758
rect 18524 14470 18644 14498
rect 18524 14414 18552 14470
rect 18512 14408 18564 14414
rect 18708 14396 18736 18702
rect 18800 16114 18828 19790
rect 18880 19780 18932 19786
rect 18880 19722 18932 19728
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18800 15502 18828 16050
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18512 14350 18564 14356
rect 18616 14368 18736 14396
rect 18524 14074 18552 14350
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 18064 11762 18092 12786
rect 18248 11830 18276 12786
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 7546 14320 7822
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14096 7472 14148 7478
rect 14096 7414 14148 7420
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13556 6798 13584 7278
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 12912 6458 12940 6734
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 13556 6254 13584 6734
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 13004 5234 13032 5510
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13280 5030 13308 5646
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 13556 4690 13584 6190
rect 13832 5778 13860 6394
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13648 5234 13676 5646
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13832 5166 13860 5714
rect 14108 5710 14136 6190
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13096 3738 13124 4422
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12360 3398 12388 3470
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12452 3194 12480 3674
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 12452 2446 12480 3130
rect 12544 3058 12572 3538
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12912 2990 12940 3334
rect 13188 3194 13216 4422
rect 13832 4146 13860 5102
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 13280 2650 13308 4082
rect 14200 4078 14228 6258
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14292 5710 14320 6190
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14292 5370 14320 5646
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14384 5030 14412 5170
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14200 3534 14228 4014
rect 14292 3942 14320 4558
rect 14384 4146 14412 4966
rect 14568 4758 14596 5850
rect 14752 5778 14780 6870
rect 14844 6866 14872 7346
rect 15488 7002 15516 8366
rect 15580 7206 15608 8366
rect 15764 8090 15792 8434
rect 16684 8362 16712 9454
rect 16960 9042 16988 9998
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17788 9654 17816 9862
rect 17972 9654 18000 9930
rect 18064 9722 18092 10066
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 15846 8188 16154 8208
rect 15846 8186 15852 8188
rect 15908 8186 15932 8188
rect 15988 8186 16012 8188
rect 16068 8186 16092 8188
rect 16148 8186 16154 8188
rect 15908 8134 15910 8186
rect 16090 8134 16092 8186
rect 15846 8132 15852 8134
rect 15908 8132 15932 8134
rect 15988 8132 16012 8134
rect 16068 8132 16092 8134
rect 16148 8132 16154 8134
rect 15846 8112 16154 8132
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 16684 7410 16712 8298
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15476 6248 15528 6254
rect 15580 6236 15608 7142
rect 15846 7100 16154 7120
rect 15846 7098 15852 7100
rect 15908 7098 15932 7100
rect 15988 7098 16012 7100
rect 16068 7098 16092 7100
rect 16148 7098 16154 7100
rect 15908 7046 15910 7098
rect 16090 7046 16092 7098
rect 15846 7044 15852 7046
rect 15908 7044 15932 7046
rect 15988 7044 16012 7046
rect 16068 7044 16092 7046
rect 16148 7044 16154 7046
rect 15846 7024 16154 7044
rect 16592 6866 16620 7142
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 15752 6724 15804 6730
rect 15752 6666 15804 6672
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 15528 6208 15608 6236
rect 15476 6190 15528 6196
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14384 3670 14412 4082
rect 14752 4078 14780 4626
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14200 3058 14228 3470
rect 14384 3058 14412 3606
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 14200 2446 14228 2994
rect 14384 2446 14412 2994
rect 14752 2650 14780 4014
rect 14844 3670 14872 6122
rect 15028 5710 15056 6190
rect 15120 5914 15148 6190
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15120 5778 15148 5850
rect 15488 5778 15516 6190
rect 15764 5914 15792 6666
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15856 6458 15884 6598
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15846 6012 16154 6032
rect 15846 6010 15852 6012
rect 15908 6010 15932 6012
rect 15988 6010 16012 6012
rect 16068 6010 16092 6012
rect 16148 6010 16154 6012
rect 15908 5958 15910 6010
rect 16090 5958 16092 6010
rect 15846 5956 15852 5958
rect 15908 5956 15932 5958
rect 15988 5956 16012 5958
rect 16068 5956 16092 5958
rect 16148 5956 16154 5958
rect 15846 5936 16154 5956
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15476 5772 15528 5778
rect 15528 5732 15608 5760
rect 15476 5714 15528 5720
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 15028 5574 15056 5646
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15028 4010 15056 5510
rect 15304 5234 15332 5510
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15384 5092 15436 5098
rect 15384 5034 15436 5040
rect 15396 4486 15424 5034
rect 15488 4622 15516 5170
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15396 4146 15424 4422
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15120 3040 15148 3538
rect 15396 3534 15424 3946
rect 15580 3534 15608 5732
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16408 5030 16436 5646
rect 16500 5574 16528 6666
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 15846 4924 16154 4944
rect 15846 4922 15852 4924
rect 15908 4922 15932 4924
rect 15988 4922 16012 4924
rect 16068 4922 16092 4924
rect 16148 4922 16154 4924
rect 15908 4870 15910 4922
rect 16090 4870 16092 4922
rect 15846 4868 15852 4870
rect 15908 4868 15932 4870
rect 15988 4868 16012 4870
rect 16068 4868 16092 4870
rect 16148 4868 16154 4870
rect 15846 4848 16154 4868
rect 16408 4486 16436 4966
rect 16396 4480 16448 4486
rect 16396 4422 16448 4428
rect 16592 4078 16620 6802
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16684 4622 16712 6598
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16776 4010 16804 8434
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 17052 7886 17080 8230
rect 17512 7886 17540 8978
rect 18064 8514 18092 9658
rect 18248 9586 18276 11018
rect 18432 10266 18460 12854
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 18524 10674 18552 11154
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18616 10606 18644 14368
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18708 12986 18736 13126
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18708 12646 18736 12786
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18708 12442 18736 12582
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18800 11880 18828 15438
rect 18892 15162 18920 19722
rect 19076 16114 19104 21830
rect 19168 21554 19196 22510
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19168 19242 19196 19858
rect 19352 19854 19380 23054
rect 19432 21616 19484 21622
rect 19432 21558 19484 21564
rect 19444 20942 19472 21558
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19536 20602 19564 24142
rect 19904 24138 19932 26998
rect 19996 24313 20024 28047
rect 20076 27532 20128 27538
rect 20076 27474 20128 27480
rect 20088 26586 20116 27474
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20088 25226 20116 25842
rect 20076 25220 20128 25226
rect 20076 25162 20128 25168
rect 19982 24304 20038 24313
rect 19982 24239 20038 24248
rect 19892 24132 19944 24138
rect 19892 24074 19944 24080
rect 20076 24132 20128 24138
rect 20076 24074 20128 24080
rect 19892 23588 19944 23594
rect 19892 23530 19944 23536
rect 19616 23520 19668 23526
rect 19616 23462 19668 23468
rect 19628 23322 19656 23462
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19628 21049 19656 21286
rect 19614 21040 19670 21049
rect 19614 20975 19670 20984
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 19444 20058 19472 20266
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19430 19816 19486 19825
rect 19430 19751 19486 19760
rect 19444 19718 19472 19751
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19156 19236 19208 19242
rect 19156 19178 19208 19184
rect 19536 19174 19564 20198
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19352 18358 19380 18566
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19522 18184 19578 18193
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 19064 16108 19116 16114
rect 19116 16068 19196 16096
rect 19064 16050 19116 16056
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18892 15026 18920 15098
rect 19076 15026 19104 15642
rect 19168 15570 19196 16068
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19156 15428 19208 15434
rect 19156 15370 19208 15376
rect 19168 15162 19196 15370
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 18892 14396 18920 14962
rect 18972 14952 19024 14958
rect 18972 14894 19024 14900
rect 18984 14550 19012 14894
rect 18972 14544 19024 14550
rect 18972 14486 19024 14492
rect 18892 14368 19012 14396
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18892 12238 18920 12582
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18708 11852 18828 11880
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18064 8486 18184 8514
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17972 8090 18000 8230
rect 18064 8090 18092 8366
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16868 6390 16896 6870
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 17328 6322 17356 7822
rect 17512 6798 17540 7822
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17696 7206 17724 7686
rect 17972 7478 18000 7686
rect 17960 7472 18012 7478
rect 17960 7414 18012 7420
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 18064 6866 18092 7686
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17512 6322 17540 6734
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17696 5370 17724 6326
rect 17972 6304 18000 6734
rect 18052 6316 18104 6322
rect 17972 6276 18052 6304
rect 18052 6258 18104 6264
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 18064 5234 18092 6054
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 17052 4826 17080 5170
rect 18156 5030 18184 8486
rect 18248 8294 18276 9522
rect 18340 9178 18368 9930
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18340 8974 18368 9114
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18432 7886 18460 10202
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18616 9042 18644 9522
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18432 6934 18460 7822
rect 18616 7410 18644 8026
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18420 6928 18472 6934
rect 18420 6870 18472 6876
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18248 5914 18276 6598
rect 18432 6390 18460 6870
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18236 5296 18288 5302
rect 18236 5238 18288 5244
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 18248 4146 18276 5238
rect 18524 4146 18552 6598
rect 18616 5302 18644 7346
rect 18708 6322 18736 11852
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18800 11150 18828 11698
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18984 11082 19012 14368
rect 19260 13326 19288 17682
rect 19352 16590 19380 18158
rect 19432 18148 19484 18154
rect 19522 18119 19578 18128
rect 19432 18090 19484 18096
rect 19444 18057 19472 18090
rect 19430 18048 19486 18057
rect 19430 17983 19486 17992
rect 19536 17814 19564 18119
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19444 15502 19472 17138
rect 19524 16516 19576 16522
rect 19524 16458 19576 16464
rect 19536 16250 19564 16458
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19628 16046 19656 19790
rect 19720 16182 19748 22714
rect 19800 21888 19852 21894
rect 19800 21830 19852 21836
rect 19812 21418 19840 21830
rect 19800 21412 19852 21418
rect 19800 21354 19852 21360
rect 19800 20596 19852 20602
rect 19800 20538 19852 20544
rect 19812 19854 19840 20538
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19812 17377 19840 18702
rect 19798 17368 19854 17377
rect 19798 17303 19854 17312
rect 19904 17218 19932 23530
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19996 21622 20024 21830
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19996 21010 20024 21558
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 20088 20806 20116 24074
rect 20180 21554 20208 28319
rect 20352 28008 20404 28014
rect 20352 27950 20404 27956
rect 20364 27674 20392 27950
rect 20352 27668 20404 27674
rect 20352 27610 20404 27616
rect 20456 26330 20484 30058
rect 20732 29510 20760 30194
rect 20720 29504 20772 29510
rect 20720 29446 20772 29452
rect 20732 28082 20760 29446
rect 20811 29404 21119 29424
rect 20811 29402 20817 29404
rect 20873 29402 20897 29404
rect 20953 29402 20977 29404
rect 21033 29402 21057 29404
rect 21113 29402 21119 29404
rect 20873 29350 20875 29402
rect 21055 29350 21057 29402
rect 20811 29348 20817 29350
rect 20873 29348 20897 29350
rect 20953 29348 20977 29350
rect 21033 29348 21057 29350
rect 21113 29348 21119 29350
rect 20811 29328 21119 29348
rect 21192 29170 21220 31078
rect 21284 29646 21312 31758
rect 21364 31136 21416 31142
rect 21364 31078 21416 31084
rect 21376 30734 21404 31078
rect 21364 30728 21416 30734
rect 21364 30670 21416 30676
rect 21456 30728 21508 30734
rect 21456 30670 21508 30676
rect 21364 30320 21416 30326
rect 21364 30262 21416 30268
rect 21272 29640 21324 29646
rect 21272 29582 21324 29588
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 21180 29028 21232 29034
rect 21180 28970 21232 28976
rect 20811 28316 21119 28336
rect 20811 28314 20817 28316
rect 20873 28314 20897 28316
rect 20953 28314 20977 28316
rect 21033 28314 21057 28316
rect 21113 28314 21119 28316
rect 20873 28262 20875 28314
rect 21055 28262 21057 28314
rect 20811 28260 20817 28262
rect 20873 28260 20897 28262
rect 20953 28260 20977 28262
rect 21033 28260 21057 28262
rect 21113 28260 21119 28262
rect 20811 28240 21119 28260
rect 20812 28144 20864 28150
rect 20812 28086 20864 28092
rect 20720 28076 20772 28082
rect 20720 28018 20772 28024
rect 20536 27532 20588 27538
rect 20536 27474 20588 27480
rect 20548 26994 20576 27474
rect 20628 27396 20680 27402
rect 20824 27384 20852 28086
rect 20628 27338 20680 27344
rect 20732 27356 20852 27384
rect 20640 26994 20668 27338
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20628 26988 20680 26994
rect 20628 26930 20680 26936
rect 20536 26852 20588 26858
rect 20536 26794 20588 26800
rect 20548 26450 20576 26794
rect 20536 26444 20588 26450
rect 20536 26386 20588 26392
rect 20260 26308 20312 26314
rect 20456 26302 20576 26330
rect 20260 26250 20312 26256
rect 20272 25974 20300 26250
rect 20260 25968 20312 25974
rect 20260 25910 20312 25916
rect 20352 25696 20404 25702
rect 20352 25638 20404 25644
rect 20364 25158 20392 25638
rect 20352 25152 20404 25158
rect 20352 25094 20404 25100
rect 20364 23118 20392 25094
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20456 24206 20484 24754
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20444 23656 20496 23662
rect 20444 23598 20496 23604
rect 20352 23112 20404 23118
rect 20272 23060 20352 23066
rect 20272 23054 20404 23060
rect 20272 23038 20392 23054
rect 20272 21622 20300 23038
rect 20456 22964 20484 23598
rect 20364 22936 20484 22964
rect 20364 21622 20392 22936
rect 20548 22094 20576 26302
rect 20732 26042 20760 27356
rect 20811 27228 21119 27248
rect 20811 27226 20817 27228
rect 20873 27226 20897 27228
rect 20953 27226 20977 27228
rect 21033 27226 21057 27228
rect 21113 27226 21119 27228
rect 20873 27174 20875 27226
rect 21055 27174 21057 27226
rect 20811 27172 20817 27174
rect 20873 27172 20897 27174
rect 20953 27172 20977 27174
rect 21033 27172 21057 27174
rect 21113 27172 21119 27174
rect 20811 27152 21119 27172
rect 20904 27056 20956 27062
rect 20904 26998 20956 27004
rect 20916 26926 20944 26998
rect 21192 26994 21220 28970
rect 21284 28626 21312 29582
rect 21376 29578 21404 30262
rect 21364 29572 21416 29578
rect 21364 29514 21416 29520
rect 21272 28620 21324 28626
rect 21272 28562 21324 28568
rect 21284 28150 21312 28562
rect 21468 28558 21496 30670
rect 21456 28552 21508 28558
rect 21456 28494 21508 28500
rect 21272 28144 21324 28150
rect 21272 28086 21324 28092
rect 21284 27402 21312 28086
rect 21468 28082 21496 28494
rect 21456 28076 21508 28082
rect 21456 28018 21508 28024
rect 21468 27674 21496 28018
rect 21456 27668 21508 27674
rect 21456 27610 21508 27616
rect 21272 27396 21324 27402
rect 21272 27338 21324 27344
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 21192 26382 21220 26930
rect 21272 26784 21324 26790
rect 21272 26726 21324 26732
rect 21180 26376 21232 26382
rect 21180 26318 21232 26324
rect 21284 26314 21312 26726
rect 21272 26308 21324 26314
rect 21272 26250 21324 26256
rect 20811 26140 21119 26160
rect 20811 26138 20817 26140
rect 20873 26138 20897 26140
rect 20953 26138 20977 26140
rect 21033 26138 21057 26140
rect 21113 26138 21119 26140
rect 20873 26086 20875 26138
rect 21055 26086 21057 26138
rect 20811 26084 20817 26086
rect 20873 26084 20897 26086
rect 20953 26084 20977 26086
rect 21033 26084 21057 26086
rect 21113 26084 21119 26086
rect 20811 26064 21119 26084
rect 20628 26036 20680 26042
rect 20628 25978 20680 25984
rect 20720 26036 20772 26042
rect 20720 25978 20772 25984
rect 20640 25770 20668 25978
rect 20628 25764 20680 25770
rect 20628 25706 20680 25712
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 20720 25492 20772 25498
rect 20720 25434 20772 25440
rect 20732 24750 20760 25434
rect 21468 25430 21496 25638
rect 21456 25424 21508 25430
rect 21456 25366 21508 25372
rect 21560 25362 21588 42094
rect 21744 41256 21772 44134
rect 21928 43330 21956 44814
rect 22020 44402 22048 44911
rect 22376 44882 22428 44888
rect 22468 44940 22520 44946
rect 22468 44882 22520 44888
rect 22836 44872 22888 44878
rect 22836 44814 22888 44820
rect 22192 44804 22244 44810
rect 22192 44746 22244 44752
rect 22100 44736 22152 44742
rect 22100 44678 22152 44684
rect 22008 44396 22060 44402
rect 22008 44338 22060 44344
rect 21836 43302 21956 43330
rect 21836 41478 21864 43302
rect 21916 43240 21968 43246
rect 21914 43208 21916 43217
rect 21968 43208 21970 43217
rect 21914 43143 21970 43152
rect 21824 41472 21876 41478
rect 21824 41414 21876 41420
rect 21744 41228 21956 41256
rect 21824 41132 21876 41138
rect 21824 41074 21876 41080
rect 21640 41064 21692 41070
rect 21640 41006 21692 41012
rect 21652 39506 21680 41006
rect 21732 40928 21784 40934
rect 21732 40870 21784 40876
rect 21640 39500 21692 39506
rect 21640 39442 21692 39448
rect 21640 39296 21692 39302
rect 21640 39238 21692 39244
rect 21652 38962 21680 39238
rect 21640 38956 21692 38962
rect 21640 38898 21692 38904
rect 21652 38350 21680 38898
rect 21640 38344 21692 38350
rect 21640 38286 21692 38292
rect 21640 38208 21692 38214
rect 21640 38150 21692 38156
rect 21652 28665 21680 38150
rect 21744 31754 21772 40870
rect 21836 40730 21864 41074
rect 21824 40724 21876 40730
rect 21824 40666 21876 40672
rect 21822 40624 21878 40633
rect 21822 40559 21878 40568
rect 21836 35329 21864 40559
rect 21928 40066 21956 41228
rect 22020 40186 22048 44338
rect 22112 44334 22140 44678
rect 22100 44328 22152 44334
rect 22204 44305 22232 44746
rect 22100 44270 22152 44276
rect 22190 44296 22246 44305
rect 22190 44231 22246 44240
rect 22848 44198 22876 44814
rect 22928 44396 22980 44402
rect 22928 44338 22980 44344
rect 22836 44192 22888 44198
rect 22836 44134 22888 44140
rect 22836 43920 22888 43926
rect 22836 43862 22888 43868
rect 22652 43852 22704 43858
rect 22652 43794 22704 43800
rect 22468 43784 22520 43790
rect 22468 43726 22520 43732
rect 22560 43784 22612 43790
rect 22560 43726 22612 43732
rect 22376 43648 22428 43654
rect 22376 43590 22428 43596
rect 22192 43308 22244 43314
rect 22192 43250 22244 43256
rect 22100 43104 22152 43110
rect 22100 43046 22152 43052
rect 22112 42809 22140 43046
rect 22098 42800 22154 42809
rect 22098 42735 22154 42744
rect 22204 41002 22232 43250
rect 22282 43208 22338 43217
rect 22282 43143 22338 43152
rect 22296 43110 22324 43143
rect 22284 43104 22336 43110
rect 22284 43046 22336 43052
rect 22388 41414 22416 43590
rect 22480 43450 22508 43726
rect 22468 43444 22520 43450
rect 22468 43386 22520 43392
rect 22572 41414 22600 43726
rect 22664 42294 22692 43794
rect 22744 43308 22796 43314
rect 22744 43250 22796 43256
rect 22756 42702 22784 43250
rect 22744 42696 22796 42702
rect 22744 42638 22796 42644
rect 22652 42288 22704 42294
rect 22652 42230 22704 42236
rect 22296 41386 22416 41414
rect 22480 41386 22600 41414
rect 22192 40996 22244 41002
rect 22192 40938 22244 40944
rect 22100 40384 22152 40390
rect 22100 40326 22152 40332
rect 22008 40180 22060 40186
rect 22008 40122 22060 40128
rect 21928 40038 22048 40066
rect 22112 40050 22140 40326
rect 21916 38208 21968 38214
rect 21916 38150 21968 38156
rect 21822 35320 21878 35329
rect 21822 35255 21878 35264
rect 21824 35012 21876 35018
rect 21824 34954 21876 34960
rect 21836 34746 21864 34954
rect 21824 34740 21876 34746
rect 21824 34682 21876 34688
rect 21744 31726 21864 31754
rect 21732 31408 21784 31414
rect 21732 31350 21784 31356
rect 21744 30326 21772 31350
rect 21732 30320 21784 30326
rect 21732 30262 21784 30268
rect 21732 29504 21784 29510
rect 21732 29446 21784 29452
rect 21638 28656 21694 28665
rect 21744 28626 21772 29446
rect 21638 28591 21694 28600
rect 21732 28620 21784 28626
rect 21732 28562 21784 28568
rect 21640 28552 21692 28558
rect 21640 28494 21692 28500
rect 21652 28218 21680 28494
rect 21640 28212 21692 28218
rect 21640 28154 21692 28160
rect 21744 28014 21772 28562
rect 21732 28008 21784 28014
rect 21732 27950 21784 27956
rect 21548 25356 21600 25362
rect 21548 25298 21600 25304
rect 21640 25220 21692 25226
rect 21640 25162 21692 25168
rect 20811 25052 21119 25072
rect 20811 25050 20817 25052
rect 20873 25050 20897 25052
rect 20953 25050 20977 25052
rect 21033 25050 21057 25052
rect 21113 25050 21119 25052
rect 20873 24998 20875 25050
rect 21055 24998 21057 25050
rect 20811 24996 20817 24998
rect 20873 24996 20897 24998
rect 20953 24996 20977 24998
rect 21033 24996 21057 24998
rect 21113 24996 21119 24998
rect 20811 24976 21119 24996
rect 20720 24744 20772 24750
rect 20720 24686 20772 24692
rect 20732 23186 20760 24686
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 20811 23964 21119 23984
rect 20811 23962 20817 23964
rect 20873 23962 20897 23964
rect 20953 23962 20977 23964
rect 21033 23962 21057 23964
rect 21113 23962 21119 23964
rect 20873 23910 20875 23962
rect 21055 23910 21057 23962
rect 20811 23908 20817 23910
rect 20873 23908 20897 23910
rect 20953 23908 20977 23910
rect 21033 23908 21057 23910
rect 21113 23908 21119 23910
rect 20811 23888 21119 23908
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20628 22568 20680 22574
rect 20628 22510 20680 22516
rect 20456 22066 20576 22094
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 20168 21548 20220 21554
rect 20168 21490 20220 21496
rect 20166 21312 20222 21321
rect 20166 21247 20222 21256
rect 20180 20874 20208 21247
rect 20456 20890 20484 22066
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20364 20862 20484 20890
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 20076 20528 20128 20534
rect 20074 20496 20076 20505
rect 20128 20496 20130 20505
rect 19984 20460 20036 20466
rect 20074 20431 20130 20440
rect 19984 20402 20036 20408
rect 19996 20058 20024 20402
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19996 18329 20024 19790
rect 19982 18320 20038 18329
rect 19982 18255 20038 18264
rect 20088 17610 20116 20334
rect 20180 20330 20208 20538
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20180 17882 20208 19858
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 19812 17190 19932 17218
rect 19708 16176 19760 16182
rect 19708 16118 19760 16124
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19524 15972 19576 15978
rect 19524 15914 19576 15920
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19536 15162 19564 15914
rect 19628 15502 19656 15982
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19352 14414 19380 14894
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19352 13870 19380 14350
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19168 11694 19196 12718
rect 19628 12646 19656 15438
rect 19720 14278 19748 15438
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19616 12436 19668 12442
rect 19720 12434 19748 12786
rect 19668 12406 19748 12434
rect 19616 12378 19668 12384
rect 19812 12288 19840 17190
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19904 15910 19932 16526
rect 19996 15978 20024 17070
rect 19984 15972 20036 15978
rect 19984 15914 20036 15920
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19904 14958 19932 15846
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19996 14414 20024 15302
rect 20088 14414 20116 17546
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19904 13530 19932 13874
rect 19892 13524 19944 13530
rect 19944 13484 20024 13512
rect 19892 13466 19944 13472
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 19628 12260 19840 12288
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19168 11218 19196 11630
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 18972 11076 19024 11082
rect 18972 11018 19024 11024
rect 18984 10538 19012 11018
rect 19260 10674 19288 11086
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 18972 10532 19024 10538
rect 18972 10474 19024 10480
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18800 8634 18828 9522
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18604 5296 18656 5302
rect 18604 5238 18656 5244
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 15846 3836 16154 3856
rect 15846 3834 15852 3836
rect 15908 3834 15932 3836
rect 15988 3834 16012 3836
rect 16068 3834 16092 3836
rect 16148 3834 16154 3836
rect 15908 3782 15910 3834
rect 16090 3782 16092 3834
rect 15846 3780 15852 3782
rect 15908 3780 15932 3782
rect 15988 3780 16012 3782
rect 16068 3780 16092 3782
rect 16148 3780 16154 3782
rect 15846 3760 16154 3780
rect 17052 3738 17080 4082
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 15384 3528 15436 3534
rect 15568 3528 15620 3534
rect 15384 3470 15436 3476
rect 15488 3488 15568 3516
rect 15396 3058 15424 3470
rect 15488 3194 15516 3488
rect 15568 3470 15620 3476
rect 17144 3194 17172 4014
rect 18892 3942 18920 6734
rect 18984 6322 19012 10474
rect 19076 10062 19104 10542
rect 19352 10062 19380 12174
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 19536 11898 19564 12106
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19432 11280 19484 11286
rect 19432 11222 19484 11228
rect 19444 11150 19472 11222
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19076 9586 19104 9998
rect 19352 9586 19380 9998
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19076 9178 19104 9522
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 19168 8566 19196 9318
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19260 8566 19288 8910
rect 19156 8560 19208 8566
rect 19156 8502 19208 8508
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19444 8090 19472 10202
rect 19536 10062 19564 10950
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19628 9674 19656 12260
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11762 19840 12038
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19720 10742 19748 11086
rect 19708 10736 19760 10742
rect 19708 10678 19760 10684
rect 19720 9926 19748 10678
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19628 9646 19840 9674
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19444 7750 19472 8026
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19168 6322 19196 6394
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19168 5370 19196 6258
rect 19352 6254 19380 6666
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19444 6202 19472 7686
rect 19536 7546 19564 7958
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19720 6390 19748 7822
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19444 6174 19564 6202
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19444 5302 19472 6054
rect 19536 5846 19564 6174
rect 19524 5840 19576 5846
rect 19524 5782 19576 5788
rect 19616 5704 19668 5710
rect 19720 5692 19748 6326
rect 19812 5710 19840 9646
rect 19904 8906 19932 13330
rect 19996 10742 20024 13484
rect 20088 12850 20116 13874
rect 20168 13456 20220 13462
rect 20168 13398 20220 13404
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 19984 10736 20036 10742
rect 19984 10678 20036 10684
rect 19892 8900 19944 8906
rect 19892 8842 19944 8848
rect 20088 8634 20116 12582
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19904 7954 19932 8026
rect 20088 7970 20116 8570
rect 20180 8090 20208 13398
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19996 7942 20116 7970
rect 19996 6254 20024 7942
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 20088 7206 20116 7822
rect 20168 7472 20220 7478
rect 20168 7414 20220 7420
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 20088 6730 20116 7142
rect 20180 6730 20208 7414
rect 20272 7002 20300 20742
rect 20364 19854 20392 20862
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20456 20534 20484 20742
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 20456 20398 20484 20470
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 20548 19854 20576 21626
rect 20640 20913 20668 22510
rect 20732 22234 20760 23122
rect 20811 22876 21119 22896
rect 20811 22874 20817 22876
rect 20873 22874 20897 22876
rect 20953 22874 20977 22876
rect 21033 22874 21057 22876
rect 21113 22874 21119 22876
rect 20873 22822 20875 22874
rect 21055 22822 21057 22874
rect 20811 22820 20817 22822
rect 20873 22820 20897 22822
rect 20953 22820 20977 22822
rect 21033 22820 21057 22822
rect 21113 22820 21119 22822
rect 20811 22800 21119 22820
rect 21284 22642 21312 24142
rect 21652 23186 21680 25162
rect 21836 24206 21864 31726
rect 21928 31414 21956 38150
rect 22020 34950 22048 40038
rect 22100 40044 22152 40050
rect 22100 39986 22152 39992
rect 22296 39438 22324 41386
rect 22284 39432 22336 39438
rect 22284 39374 22336 39380
rect 22100 39296 22152 39302
rect 22100 39238 22152 39244
rect 22112 39098 22140 39238
rect 22100 39092 22152 39098
rect 22100 39034 22152 39040
rect 22100 38344 22152 38350
rect 22100 38286 22152 38292
rect 22112 38010 22140 38286
rect 22100 38004 22152 38010
rect 22100 37946 22152 37952
rect 22100 37868 22152 37874
rect 22100 37810 22152 37816
rect 22112 37194 22140 37810
rect 22192 37256 22244 37262
rect 22192 37198 22244 37204
rect 22100 37188 22152 37194
rect 22100 37130 22152 37136
rect 22112 36786 22140 37130
rect 22100 36780 22152 36786
rect 22100 36722 22152 36728
rect 22204 36666 22232 37198
rect 22112 36638 22232 36666
rect 22376 36712 22428 36718
rect 22376 36654 22428 36660
rect 22112 36174 22140 36638
rect 22388 36378 22416 36654
rect 22376 36372 22428 36378
rect 22376 36314 22428 36320
rect 22388 36258 22416 36314
rect 22296 36230 22416 36258
rect 22100 36168 22152 36174
rect 22100 36110 22152 36116
rect 22112 35630 22140 36110
rect 22100 35624 22152 35630
rect 22100 35566 22152 35572
rect 22008 34944 22060 34950
rect 22008 34886 22060 34892
rect 22296 34490 22324 36230
rect 22376 34944 22428 34950
rect 22376 34886 22428 34892
rect 22388 34610 22416 34886
rect 22376 34604 22428 34610
rect 22376 34546 22428 34552
rect 22296 34462 22416 34490
rect 22284 33992 22336 33998
rect 22284 33934 22336 33940
rect 22296 33658 22324 33934
rect 22284 33652 22336 33658
rect 22284 33594 22336 33600
rect 22192 33584 22244 33590
rect 22192 33526 22244 33532
rect 22100 33516 22152 33522
rect 22100 33458 22152 33464
rect 22112 32570 22140 33458
rect 22100 32564 22152 32570
rect 22100 32506 22152 32512
rect 22100 32428 22152 32434
rect 22100 32370 22152 32376
rect 22008 31884 22060 31890
rect 22008 31826 22060 31832
rect 21916 31408 21968 31414
rect 21916 31350 21968 31356
rect 22020 31346 22048 31826
rect 22112 31822 22140 32370
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 21916 31272 21968 31278
rect 21916 31214 21968 31220
rect 21928 30734 21956 31214
rect 22020 30802 22048 31282
rect 22008 30796 22060 30802
rect 22008 30738 22060 30744
rect 21916 30728 21968 30734
rect 21916 30670 21968 30676
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 22112 28422 22140 29106
rect 22204 28558 22232 33526
rect 22388 31754 22416 34462
rect 22296 31726 22416 31754
rect 22296 28966 22324 31726
rect 22376 30592 22428 30598
rect 22376 30534 22428 30540
rect 22388 30326 22416 30534
rect 22376 30320 22428 30326
rect 22376 30262 22428 30268
rect 22284 28960 22336 28966
rect 22284 28902 22336 28908
rect 22192 28552 22244 28558
rect 22192 28494 22244 28500
rect 22100 28416 22152 28422
rect 22100 28358 22152 28364
rect 22296 28082 22324 28902
rect 22374 28520 22430 28529
rect 22374 28455 22430 28464
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 21916 28008 21968 28014
rect 21916 27950 21968 27956
rect 21928 27130 21956 27950
rect 22284 27940 22336 27946
rect 22284 27882 22336 27888
rect 22296 27402 22324 27882
rect 22284 27396 22336 27402
rect 22284 27338 22336 27344
rect 22388 27130 22416 28455
rect 22480 28200 22508 41386
rect 22560 40588 22612 40594
rect 22560 40530 22612 40536
rect 22572 40186 22600 40530
rect 22560 40180 22612 40186
rect 22560 40122 22612 40128
rect 22756 39642 22784 42638
rect 22848 41041 22876 43862
rect 22940 42566 22968 44338
rect 23112 44192 23164 44198
rect 23112 44134 23164 44140
rect 23124 43314 23152 44134
rect 23204 43784 23256 43790
rect 23204 43726 23256 43732
rect 23216 43450 23244 43726
rect 23204 43444 23256 43450
rect 23204 43386 23256 43392
rect 23112 43308 23164 43314
rect 23112 43250 23164 43256
rect 23308 43081 23336 45766
rect 23846 45656 23902 45665
rect 23846 45591 23848 45600
rect 23900 45591 23902 45600
rect 23848 45562 23900 45568
rect 23848 45484 23900 45490
rect 23848 45426 23900 45432
rect 23388 44328 23440 44334
rect 23386 44296 23388 44305
rect 23572 44328 23624 44334
rect 23440 44296 23442 44305
rect 23572 44270 23624 44276
rect 23386 44231 23442 44240
rect 23386 44160 23442 44169
rect 23386 44095 23442 44104
rect 23400 43654 23428 44095
rect 23584 43994 23612 44270
rect 23572 43988 23624 43994
rect 23572 43930 23624 43936
rect 23664 43988 23716 43994
rect 23664 43930 23716 43936
rect 23676 43874 23704 43930
rect 23492 43846 23704 43874
rect 23388 43648 23440 43654
rect 23388 43590 23440 43596
rect 23492 43314 23520 43846
rect 23572 43784 23624 43790
rect 23570 43752 23572 43761
rect 23624 43752 23626 43761
rect 23860 43738 23888 45426
rect 23952 44946 23980 47200
rect 23940 44940 23992 44946
rect 23940 44882 23992 44888
rect 24780 44384 24808 47200
rect 24860 44396 24912 44402
rect 24780 44356 24860 44384
rect 24860 44338 24912 44344
rect 24964 44282 24992 47246
rect 25424 47138 25452 47246
rect 25502 47200 25558 48000
rect 26238 47200 26294 48000
rect 27066 47200 27122 48000
rect 27802 47200 27858 48000
rect 28538 47200 28594 48000
rect 29274 47200 29330 48000
rect 30010 47560 30066 47569
rect 30010 47495 30066 47504
rect 25516 47138 25544 47200
rect 25424 47110 25544 47138
rect 26146 45656 26202 45665
rect 26146 45591 26202 45600
rect 26160 45490 26188 45591
rect 26148 45484 26200 45490
rect 26148 45426 26200 45432
rect 25776 45180 26084 45200
rect 25776 45178 25782 45180
rect 25838 45178 25862 45180
rect 25918 45178 25942 45180
rect 25998 45178 26022 45180
rect 26078 45178 26084 45180
rect 25838 45126 25840 45178
rect 26020 45126 26022 45178
rect 25776 45124 25782 45126
rect 25838 45124 25862 45126
rect 25918 45124 25942 45126
rect 25998 45124 26022 45126
rect 26078 45124 26084 45126
rect 25776 45104 26084 45124
rect 25044 44872 25096 44878
rect 25044 44814 25096 44820
rect 24872 44254 24992 44282
rect 24492 43852 24544 43858
rect 24492 43794 24544 43800
rect 24400 43784 24452 43790
rect 23860 43710 23980 43738
rect 24136 43722 24348 43738
rect 24400 43726 24452 43732
rect 23570 43687 23626 43696
rect 23952 43654 23980 43710
rect 24124 43716 24360 43722
rect 24176 43710 24308 43716
rect 24124 43658 24176 43664
rect 24308 43658 24360 43664
rect 23848 43648 23900 43654
rect 23848 43590 23900 43596
rect 23940 43648 23992 43654
rect 23940 43590 23992 43596
rect 23860 43382 23888 43590
rect 24412 43450 24440 43726
rect 24504 43450 24532 43794
rect 24584 43784 24636 43790
rect 24676 43784 24728 43790
rect 24584 43726 24636 43732
rect 24674 43752 24676 43761
rect 24728 43752 24730 43761
rect 24400 43444 24452 43450
rect 24400 43386 24452 43392
rect 24492 43444 24544 43450
rect 24492 43386 24544 43392
rect 23848 43376 23900 43382
rect 23848 43318 23900 43324
rect 23480 43308 23532 43314
rect 23480 43250 23532 43256
rect 23386 43208 23442 43217
rect 23386 43143 23388 43152
rect 23440 43143 23442 43152
rect 23388 43114 23440 43120
rect 24596 43110 24624 43726
rect 24730 43710 24808 43738
rect 24674 43687 24730 43696
rect 24584 43104 24636 43110
rect 23294 43072 23350 43081
rect 24584 43046 24636 43052
rect 23294 43007 23350 43016
rect 22928 42560 22980 42566
rect 22928 42502 22980 42508
rect 23388 42560 23440 42566
rect 23388 42502 23440 42508
rect 23400 42294 23428 42502
rect 23848 42356 23900 42362
rect 23848 42298 23900 42304
rect 23388 42288 23440 42294
rect 23860 42265 23888 42298
rect 23388 42230 23440 42236
rect 23846 42256 23902 42265
rect 23020 42220 23072 42226
rect 23846 42191 23902 42200
rect 24032 42220 24084 42226
rect 23020 42162 23072 42168
rect 24032 42162 24084 42168
rect 24124 42220 24176 42226
rect 24124 42162 24176 42168
rect 23032 41313 23060 42162
rect 24044 41750 24072 42162
rect 24032 41744 24084 41750
rect 23846 41712 23902 41721
rect 24032 41686 24084 41692
rect 23846 41647 23848 41656
rect 23900 41647 23902 41656
rect 23848 41618 23900 41624
rect 24136 41614 24164 42162
rect 24216 42152 24268 42158
rect 24216 42094 24268 42100
rect 23388 41608 23440 41614
rect 23388 41550 23440 41556
rect 24124 41608 24176 41614
rect 24124 41550 24176 41556
rect 23018 41304 23074 41313
rect 23018 41239 23074 41248
rect 22834 41032 22890 41041
rect 22834 40967 22890 40976
rect 23112 40996 23164 41002
rect 23112 40938 23164 40944
rect 22928 40520 22980 40526
rect 22928 40462 22980 40468
rect 22940 40186 22968 40462
rect 22928 40180 22980 40186
rect 22928 40122 22980 40128
rect 22836 40044 22888 40050
rect 22836 39986 22888 39992
rect 22744 39636 22796 39642
rect 22744 39578 22796 39584
rect 22560 38208 22612 38214
rect 22560 38150 22612 38156
rect 22572 37874 22600 38150
rect 22756 38010 22784 39578
rect 22848 39438 22876 39986
rect 22836 39432 22888 39438
rect 22836 39374 22888 39380
rect 22744 38004 22796 38010
rect 22744 37946 22796 37952
rect 22560 37868 22612 37874
rect 22560 37810 22612 37816
rect 22652 36780 22704 36786
rect 22652 36722 22704 36728
rect 22664 36310 22692 36722
rect 22744 36576 22796 36582
rect 22744 36518 22796 36524
rect 22652 36304 22704 36310
rect 22652 36246 22704 36252
rect 22756 36174 22784 36518
rect 22744 36168 22796 36174
rect 22744 36110 22796 36116
rect 22652 35760 22704 35766
rect 22652 35702 22704 35708
rect 22664 34746 22692 35702
rect 22848 35494 22876 39374
rect 23018 39128 23074 39137
rect 23018 39063 23020 39072
rect 23072 39063 23074 39072
rect 23020 39034 23072 39040
rect 22928 37664 22980 37670
rect 22928 37606 22980 37612
rect 22940 37262 22968 37606
rect 22928 37256 22980 37262
rect 22928 37198 22980 37204
rect 23020 37256 23072 37262
rect 23020 37198 23072 37204
rect 22928 37120 22980 37126
rect 22928 37062 22980 37068
rect 22940 36786 22968 37062
rect 22928 36780 22980 36786
rect 22928 36722 22980 36728
rect 22940 36242 22968 36722
rect 23032 36310 23060 37198
rect 23020 36304 23072 36310
rect 23020 36246 23072 36252
rect 22928 36236 22980 36242
rect 22928 36178 22980 36184
rect 23124 36106 23152 40938
rect 23204 40452 23256 40458
rect 23204 40394 23256 40400
rect 23296 40452 23348 40458
rect 23296 40394 23348 40400
rect 23216 40361 23244 40394
rect 23202 40352 23258 40361
rect 23202 40287 23258 40296
rect 23308 40118 23336 40394
rect 23400 40118 23428 41550
rect 23572 41472 23624 41478
rect 23572 41414 23624 41420
rect 23480 41064 23532 41070
rect 23480 41006 23532 41012
rect 23492 40730 23520 41006
rect 23480 40724 23532 40730
rect 23480 40666 23532 40672
rect 23584 40526 23612 41414
rect 23848 41200 23900 41206
rect 23848 41142 23900 41148
rect 23572 40520 23624 40526
rect 23572 40462 23624 40468
rect 23296 40112 23348 40118
rect 23296 40054 23348 40060
rect 23388 40112 23440 40118
rect 23388 40054 23440 40060
rect 23296 39976 23348 39982
rect 23296 39918 23348 39924
rect 23204 39908 23256 39914
rect 23204 39850 23256 39856
rect 23216 39642 23244 39850
rect 23204 39636 23256 39642
rect 23204 39578 23256 39584
rect 23308 38196 23336 39918
rect 23400 39914 23428 40054
rect 23860 40050 23888 41142
rect 23848 40044 23900 40050
rect 23848 39986 23900 39992
rect 23388 39908 23440 39914
rect 23388 39850 23440 39856
rect 23664 39840 23716 39846
rect 23664 39782 23716 39788
rect 23478 39536 23534 39545
rect 23478 39471 23480 39480
rect 23532 39471 23534 39480
rect 23480 39442 23532 39448
rect 23572 39364 23624 39370
rect 23572 39306 23624 39312
rect 23584 38654 23612 39306
rect 23676 39098 23704 39782
rect 23860 39438 23888 39986
rect 24124 39976 24176 39982
rect 24228 39964 24256 42094
rect 24308 41608 24360 41614
rect 24308 41550 24360 41556
rect 24320 39982 24348 41550
rect 24596 41478 24624 43046
rect 24780 42566 24808 43710
rect 24676 42560 24728 42566
rect 24674 42528 24676 42537
rect 24768 42560 24820 42566
rect 24728 42528 24730 42537
rect 24768 42502 24820 42508
rect 24674 42463 24730 42472
rect 24780 42158 24808 42502
rect 24768 42152 24820 42158
rect 24768 42094 24820 42100
rect 24584 41472 24636 41478
rect 24584 41414 24636 41420
rect 24768 41472 24820 41478
rect 24768 41414 24820 41420
rect 24584 41132 24636 41138
rect 24584 41074 24636 41080
rect 24400 40928 24452 40934
rect 24400 40870 24452 40876
rect 24412 40050 24440 40870
rect 24596 40050 24624 41074
rect 24400 40044 24452 40050
rect 24400 39986 24452 39992
rect 24584 40044 24636 40050
rect 24584 39986 24636 39992
rect 24176 39936 24256 39964
rect 24124 39918 24176 39924
rect 23848 39432 23900 39438
rect 23848 39374 23900 39380
rect 24228 39370 24256 39936
rect 24308 39976 24360 39982
rect 24308 39918 24360 39924
rect 24492 39976 24544 39982
rect 24492 39918 24544 39924
rect 24320 39522 24348 39918
rect 24504 39681 24532 39918
rect 24780 39846 24808 41414
rect 24872 40390 24900 44254
rect 24952 44192 25004 44198
rect 24952 44134 25004 44140
rect 24964 43790 24992 44134
rect 24952 43784 25004 43790
rect 24952 43726 25004 43732
rect 24964 43382 24992 43726
rect 24952 43376 25004 43382
rect 24952 43318 25004 43324
rect 25056 42770 25084 44814
rect 25320 44736 25372 44742
rect 25320 44678 25372 44684
rect 25136 44328 25188 44334
rect 25136 44270 25188 44276
rect 25226 44296 25282 44305
rect 25148 43926 25176 44270
rect 25226 44231 25282 44240
rect 25240 44198 25268 44231
rect 25228 44192 25280 44198
rect 25228 44134 25280 44140
rect 25136 43920 25188 43926
rect 25136 43862 25188 43868
rect 25332 43450 25360 44678
rect 25686 44432 25742 44441
rect 25686 44367 25688 44376
rect 25740 44367 25742 44376
rect 25688 44338 25740 44344
rect 26252 44305 26280 47200
rect 27080 45830 27108 47200
rect 27068 45824 27120 45830
rect 27068 45766 27120 45772
rect 27436 45484 27488 45490
rect 27436 45426 27488 45432
rect 27620 45484 27672 45490
rect 27620 45426 27672 45432
rect 27160 45280 27212 45286
rect 27160 45222 27212 45228
rect 27252 45280 27304 45286
rect 27252 45222 27304 45228
rect 27172 44946 27200 45222
rect 27160 44940 27212 44946
rect 27160 44882 27212 44888
rect 26332 44804 26384 44810
rect 26332 44746 26384 44752
rect 26238 44296 26294 44305
rect 26238 44231 26294 44240
rect 25776 44092 26084 44112
rect 25776 44090 25782 44092
rect 25838 44090 25862 44092
rect 25918 44090 25942 44092
rect 25998 44090 26022 44092
rect 26078 44090 26084 44092
rect 25838 44038 25840 44090
rect 26020 44038 26022 44090
rect 25776 44036 25782 44038
rect 25838 44036 25862 44038
rect 25918 44036 25942 44038
rect 25998 44036 26022 44038
rect 26078 44036 26084 44038
rect 25776 44016 26084 44036
rect 25412 43852 25464 43858
rect 25412 43794 25464 43800
rect 25872 43852 25924 43858
rect 25872 43794 25924 43800
rect 25320 43444 25372 43450
rect 25320 43386 25372 43392
rect 25320 43308 25372 43314
rect 25320 43250 25372 43256
rect 25136 42832 25188 42838
rect 25136 42774 25188 42780
rect 25044 42764 25096 42770
rect 25044 42706 25096 42712
rect 24952 42628 25004 42634
rect 24952 42570 25004 42576
rect 24964 40633 24992 42570
rect 25044 42016 25096 42022
rect 25044 41958 25096 41964
rect 25056 41546 25084 41958
rect 25148 41682 25176 42774
rect 25332 42702 25360 43250
rect 25424 42838 25452 43794
rect 25884 43314 25912 43794
rect 26056 43784 26108 43790
rect 26056 43726 26108 43732
rect 25688 43308 25740 43314
rect 25688 43250 25740 43256
rect 25872 43308 25924 43314
rect 25872 43250 25924 43256
rect 25596 43240 25648 43246
rect 25596 43182 25648 43188
rect 25504 43104 25556 43110
rect 25504 43046 25556 43052
rect 25412 42832 25464 42838
rect 25412 42774 25464 42780
rect 25320 42696 25372 42702
rect 25320 42638 25372 42644
rect 25228 41744 25280 41750
rect 25228 41686 25280 41692
rect 25136 41676 25188 41682
rect 25136 41618 25188 41624
rect 25044 41540 25096 41546
rect 25044 41482 25096 41488
rect 25044 41064 25096 41070
rect 25044 41006 25096 41012
rect 24950 40624 25006 40633
rect 24950 40559 25006 40568
rect 24860 40384 24912 40390
rect 24860 40326 24912 40332
rect 24768 39840 24820 39846
rect 24768 39782 24820 39788
rect 24490 39672 24546 39681
rect 24490 39607 24546 39616
rect 24860 39636 24912 39642
rect 24860 39578 24912 39584
rect 24320 39494 24624 39522
rect 24596 39488 24624 39494
rect 24768 39500 24820 39506
rect 24596 39460 24768 39488
rect 24308 39432 24360 39438
rect 24308 39374 24360 39380
rect 24492 39432 24544 39438
rect 24544 39380 24624 39386
rect 24492 39374 24624 39380
rect 24216 39364 24268 39370
rect 24216 39306 24268 39312
rect 23664 39092 23716 39098
rect 23664 39034 23716 39040
rect 23756 39092 23808 39098
rect 23756 39034 23808 39040
rect 23768 38962 23796 39034
rect 23756 38956 23808 38962
rect 23756 38898 23808 38904
rect 24228 38894 24256 39306
rect 24320 38962 24348 39374
rect 24504 39358 24624 39374
rect 24308 38956 24360 38962
rect 24308 38898 24360 38904
rect 24400 38956 24452 38962
rect 24400 38898 24452 38904
rect 24216 38888 24268 38894
rect 24216 38830 24268 38836
rect 23584 38626 23704 38654
rect 23216 38168 23336 38196
rect 23480 38208 23532 38214
rect 23216 37398 23244 38168
rect 23480 38150 23532 38156
rect 23204 37392 23256 37398
rect 23204 37334 23256 37340
rect 23112 36100 23164 36106
rect 23112 36042 23164 36048
rect 23020 36032 23072 36038
rect 23020 35974 23072 35980
rect 22928 35828 22980 35834
rect 22928 35770 22980 35776
rect 22836 35488 22888 35494
rect 22836 35430 22888 35436
rect 22652 34740 22704 34746
rect 22652 34682 22704 34688
rect 22560 33856 22612 33862
rect 22560 33798 22612 33804
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22572 33590 22600 33798
rect 22560 33584 22612 33590
rect 22560 33526 22612 33532
rect 22756 33522 22784 33798
rect 22744 33516 22796 33522
rect 22744 33458 22796 33464
rect 22836 33516 22888 33522
rect 22836 33458 22888 33464
rect 22560 33448 22612 33454
rect 22560 33390 22612 33396
rect 22572 32366 22600 33390
rect 22848 32570 22876 33458
rect 22836 32564 22888 32570
rect 22836 32506 22888 32512
rect 22940 32450 22968 35770
rect 22756 32422 22968 32450
rect 22560 32360 22612 32366
rect 22560 32302 22612 32308
rect 22572 31686 22600 32302
rect 22560 31680 22612 31686
rect 22560 31622 22612 31628
rect 22572 31278 22600 31622
rect 22560 31272 22612 31278
rect 22560 31214 22612 31220
rect 22572 30734 22600 31214
rect 22560 30728 22612 30734
rect 22560 30670 22612 30676
rect 22572 29850 22600 30670
rect 22560 29844 22612 29850
rect 22560 29786 22612 29792
rect 22756 29510 22784 32422
rect 22928 31952 22980 31958
rect 22928 31894 22980 31900
rect 22836 31340 22888 31346
rect 22836 31282 22888 31288
rect 22848 30870 22876 31282
rect 22836 30864 22888 30870
rect 22836 30806 22888 30812
rect 22744 29504 22796 29510
rect 22744 29446 22796 29452
rect 22480 28172 22784 28200
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 22468 27872 22520 27878
rect 22468 27814 22520 27820
rect 21916 27124 21968 27130
rect 21916 27066 21968 27072
rect 22100 27124 22152 27130
rect 22100 27066 22152 27072
rect 22376 27124 22428 27130
rect 22376 27066 22428 27072
rect 21916 26920 21968 26926
rect 21916 26862 21968 26868
rect 21928 26586 21956 26862
rect 21916 26580 21968 26586
rect 21916 26522 21968 26528
rect 21928 25906 21956 26522
rect 21916 25900 21968 25906
rect 21916 25842 21968 25848
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21916 23316 21968 23322
rect 21968 23276 22048 23304
rect 21916 23258 21968 23264
rect 21640 23180 21692 23186
rect 21640 23122 21692 23128
rect 21652 22642 21680 23122
rect 21732 23112 21784 23118
rect 21732 23054 21784 23060
rect 21744 22658 21772 23054
rect 22020 22778 22048 23276
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 22112 22658 22140 27066
rect 22480 26994 22508 27814
rect 22572 27674 22600 28018
rect 22652 27872 22704 27878
rect 22652 27814 22704 27820
rect 22560 27668 22612 27674
rect 22560 27610 22612 27616
rect 22468 26988 22520 26994
rect 22468 26930 22520 26936
rect 22572 26382 22600 27610
rect 22664 26586 22692 27814
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 22560 26376 22612 26382
rect 22560 26318 22612 26324
rect 22664 25770 22692 26522
rect 22192 25764 22244 25770
rect 22192 25706 22244 25712
rect 22652 25764 22704 25770
rect 22652 25706 22704 25712
rect 22204 23798 22232 25706
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 22376 24744 22428 24750
rect 22376 24686 22428 24692
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 22296 24274 22324 24346
rect 22284 24268 22336 24274
rect 22284 24210 22336 24216
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22192 23792 22244 23798
rect 22192 23734 22244 23740
rect 22204 22710 22232 23734
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 21640 22636 21692 22642
rect 21744 22630 21864 22658
rect 21928 22642 22140 22658
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 21640 22578 21692 22584
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20824 22094 20852 22578
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 20732 22066 20852 22094
rect 20732 21486 20760 22066
rect 21272 21956 21324 21962
rect 21272 21898 21324 21904
rect 20811 21788 21119 21808
rect 20811 21786 20817 21788
rect 20873 21786 20897 21788
rect 20953 21786 20977 21788
rect 21033 21786 21057 21788
rect 21113 21786 21119 21788
rect 20873 21734 20875 21786
rect 21055 21734 21057 21786
rect 20811 21732 20817 21734
rect 20873 21732 20897 21734
rect 20953 21732 20977 21734
rect 21033 21732 21057 21734
rect 21113 21732 21119 21734
rect 20811 21712 21119 21732
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20810 21448 20866 21457
rect 20732 20942 20760 21422
rect 20810 21383 20866 21392
rect 20720 20936 20772 20942
rect 20626 20904 20682 20913
rect 20720 20878 20772 20884
rect 20626 20839 20628 20848
rect 20680 20839 20682 20848
rect 20628 20810 20680 20816
rect 20640 20779 20668 20810
rect 20824 20788 20852 21383
rect 20732 20760 20852 20788
rect 21180 20800 21232 20806
rect 20732 20482 20760 20760
rect 21180 20742 21232 20748
rect 20811 20700 21119 20720
rect 20811 20698 20817 20700
rect 20873 20698 20897 20700
rect 20953 20698 20977 20700
rect 21033 20698 21057 20700
rect 21113 20698 21119 20700
rect 20873 20646 20875 20698
rect 21055 20646 21057 20698
rect 20811 20644 20817 20646
rect 20873 20644 20897 20646
rect 20953 20644 20977 20646
rect 21033 20644 21057 20646
rect 21113 20644 21119 20646
rect 20811 20624 21119 20644
rect 21192 20534 21220 20742
rect 21284 20534 21312 21898
rect 21180 20528 21232 20534
rect 20628 20460 20680 20466
rect 20732 20454 21036 20482
rect 21180 20470 21232 20476
rect 21272 20528 21324 20534
rect 21272 20470 21324 20476
rect 20628 20402 20680 20408
rect 20640 20058 20668 20402
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20364 17864 20392 19654
rect 20548 19378 20576 19790
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20444 18692 20496 18698
rect 20444 18634 20496 18640
rect 20456 18426 20484 18634
rect 20640 18630 20668 19994
rect 21008 19854 21036 20454
rect 21192 19922 21220 20470
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 20812 19780 20864 19786
rect 20732 19740 20812 19768
rect 20732 19496 20760 19740
rect 20812 19722 20864 19728
rect 20811 19612 21119 19632
rect 20811 19610 20817 19612
rect 20873 19610 20897 19612
rect 20953 19610 20977 19612
rect 21033 19610 21057 19612
rect 21113 19610 21119 19612
rect 20873 19558 20875 19610
rect 21055 19558 21057 19610
rect 20811 19556 20817 19558
rect 20873 19556 20897 19558
rect 20953 19556 20977 19558
rect 21033 19556 21057 19558
rect 21113 19556 21119 19558
rect 20811 19536 21119 19556
rect 20732 19468 20852 19496
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20732 18902 20760 19314
rect 20720 18896 20772 18902
rect 20720 18838 20772 18844
rect 20824 18714 20852 19468
rect 21180 19440 21232 19446
rect 21180 19382 21232 19388
rect 20904 19236 20956 19242
rect 20904 19178 20956 19184
rect 20916 18834 20944 19178
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 20732 18686 20852 18714
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20628 17876 20680 17882
rect 20364 17836 20484 17864
rect 20350 17776 20406 17785
rect 20350 17711 20352 17720
rect 20404 17711 20406 17720
rect 20352 17682 20404 17688
rect 20456 17626 20484 17836
rect 20628 17818 20680 17824
rect 20640 17678 20668 17818
rect 20628 17672 20680 17678
rect 20534 17640 20590 17649
rect 20456 17598 20534 17626
rect 20628 17614 20680 17620
rect 20534 17575 20590 17584
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20364 16658 20392 16934
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20364 16250 20392 16390
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20364 15094 20392 16050
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20364 14006 20392 15030
rect 20352 14000 20404 14006
rect 20352 13942 20404 13948
rect 20456 13326 20484 15982
rect 20548 13394 20576 17575
rect 20640 14929 20668 17614
rect 20626 14920 20682 14929
rect 20626 14855 20682 14864
rect 20640 14618 20668 14855
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20364 12730 20392 13262
rect 20456 12968 20484 13262
rect 20456 12940 20576 12968
rect 20548 12900 20576 12940
rect 20628 12912 20680 12918
rect 20548 12872 20628 12900
rect 20628 12854 20680 12860
rect 20364 12702 20484 12730
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20364 11830 20392 12582
rect 20352 11824 20404 11830
rect 20352 11766 20404 11772
rect 20456 11778 20484 12702
rect 20628 12640 20680 12646
rect 20732 12617 20760 18686
rect 20811 18524 21119 18544
rect 20811 18522 20817 18524
rect 20873 18522 20897 18524
rect 20953 18522 20977 18524
rect 21033 18522 21057 18524
rect 21113 18522 21119 18524
rect 20873 18470 20875 18522
rect 21055 18470 21057 18522
rect 20811 18468 20817 18470
rect 20873 18468 20897 18470
rect 20953 18468 20977 18470
rect 21033 18468 21057 18470
rect 21113 18468 21119 18470
rect 20811 18448 21119 18468
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20824 17882 20852 18226
rect 21192 18086 21220 19382
rect 21284 18766 21312 19790
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21086 17912 21142 17921
rect 20812 17876 20864 17882
rect 21086 17847 21142 17856
rect 20812 17818 20864 17824
rect 21100 17814 21128 17847
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 21180 17808 21232 17814
rect 21284 17785 21312 18702
rect 21180 17750 21232 17756
rect 21270 17776 21326 17785
rect 20810 17640 20866 17649
rect 20810 17575 20812 17584
rect 20864 17575 20866 17584
rect 20812 17546 20864 17552
rect 20811 17436 21119 17456
rect 20811 17434 20817 17436
rect 20873 17434 20897 17436
rect 20953 17434 20977 17436
rect 21033 17434 21057 17436
rect 21113 17434 21119 17436
rect 20873 17382 20875 17434
rect 21055 17382 21057 17434
rect 20811 17380 20817 17382
rect 20873 17380 20897 17382
rect 20953 17380 20977 17382
rect 21033 17380 21057 17382
rect 21113 17380 21119 17382
rect 20811 17360 21119 17380
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20916 16998 20944 17138
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 21008 16658 21036 17138
rect 21192 17134 21220 17750
rect 21270 17711 21326 17720
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21192 16697 21220 17070
rect 21284 16833 21312 17478
rect 21270 16824 21326 16833
rect 21270 16759 21326 16768
rect 21178 16688 21234 16697
rect 20996 16652 21048 16658
rect 21178 16623 21234 16632
rect 20996 16594 21048 16600
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 20811 16348 21119 16368
rect 20811 16346 20817 16348
rect 20873 16346 20897 16348
rect 20953 16346 20977 16348
rect 21033 16346 21057 16348
rect 21113 16346 21119 16348
rect 20873 16294 20875 16346
rect 21055 16294 21057 16346
rect 20811 16292 20817 16294
rect 20873 16292 20897 16294
rect 20953 16292 20977 16294
rect 21033 16292 21057 16294
rect 21113 16292 21119 16294
rect 20811 16272 21119 16292
rect 21192 16182 21220 16458
rect 21180 16176 21232 16182
rect 21180 16118 21232 16124
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 20811 15260 21119 15280
rect 20811 15258 20817 15260
rect 20873 15258 20897 15260
rect 20953 15258 20977 15260
rect 21033 15258 21057 15260
rect 21113 15258 21119 15260
rect 20873 15206 20875 15258
rect 21055 15206 21057 15258
rect 20811 15204 20817 15206
rect 20873 15204 20897 15206
rect 20953 15204 20977 15206
rect 21033 15204 21057 15206
rect 21113 15204 21119 15206
rect 20811 15184 21119 15204
rect 21192 15094 21220 15846
rect 21284 15178 21312 16526
rect 21376 16046 21404 22374
rect 21456 22160 21508 22166
rect 21456 22102 21508 22108
rect 21468 21350 21496 22102
rect 21546 21448 21602 21457
rect 21546 21383 21602 21392
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 21468 20398 21496 21286
rect 21560 21010 21588 21383
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 21546 20904 21602 20913
rect 21744 20874 21772 21286
rect 21546 20839 21602 20848
rect 21732 20868 21784 20874
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21468 17746 21496 18022
rect 21560 17814 21588 20839
rect 21732 20810 21784 20816
rect 21744 20505 21772 20810
rect 21730 20496 21786 20505
rect 21730 20431 21786 20440
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 21548 17808 21600 17814
rect 21652 17785 21680 20198
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21744 19174 21772 19790
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21744 17882 21772 18906
rect 21836 17898 21864 22630
rect 21916 22636 22140 22642
rect 21968 22630 22140 22636
rect 21916 22578 21968 22584
rect 21914 22536 21970 22545
rect 21914 22471 21970 22480
rect 21928 22098 21956 22471
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 22020 22030 22048 22630
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 22020 21690 22048 21966
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 21916 21616 21968 21622
rect 21916 21558 21968 21564
rect 21928 20534 21956 21558
rect 22112 21418 22140 21830
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22100 21412 22152 21418
rect 22100 21354 22152 21360
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 21916 20528 21968 20534
rect 21916 20470 21968 20476
rect 22112 20466 22140 20878
rect 22204 20806 22232 21422
rect 22296 21010 22324 24006
rect 22284 21004 22336 21010
rect 22284 20946 22336 20952
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 21928 19378 21956 20334
rect 22112 19922 22140 20402
rect 22296 19990 22324 20402
rect 22284 19984 22336 19990
rect 22284 19926 22336 19932
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 22112 19802 22140 19858
rect 22112 19774 22232 19802
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22008 19508 22060 19514
rect 22008 19450 22060 19456
rect 22020 19417 22048 19450
rect 22006 19408 22062 19417
rect 21916 19372 21968 19378
rect 22112 19378 22140 19654
rect 22006 19343 22062 19352
rect 22100 19372 22152 19378
rect 21916 19314 21968 19320
rect 22100 19314 22152 19320
rect 21928 19258 21956 19314
rect 21928 19230 22140 19258
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22020 18426 22048 19110
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 21732 17876 21784 17882
rect 21836 17870 21956 17898
rect 21732 17818 21784 17824
rect 21548 17750 21600 17756
rect 21638 17776 21694 17785
rect 21456 17740 21508 17746
rect 21638 17711 21694 17720
rect 21456 17682 21508 17688
rect 21468 17202 21496 17682
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21454 16688 21510 16697
rect 21454 16623 21456 16632
rect 21508 16623 21510 16632
rect 21456 16594 21508 16600
rect 21468 16046 21496 16594
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21284 15150 21496 15178
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 20916 14822 20944 15030
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 21100 14414 21128 14894
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 20811 14172 21119 14192
rect 20811 14170 20817 14172
rect 20873 14170 20897 14172
rect 20953 14170 20977 14172
rect 21033 14170 21057 14172
rect 21113 14170 21119 14172
rect 20873 14118 20875 14170
rect 21055 14118 21057 14170
rect 20811 14116 20817 14118
rect 20873 14116 20897 14118
rect 20953 14116 20977 14118
rect 21033 14116 21057 14118
rect 21113 14116 21119 14118
rect 20811 14096 21119 14116
rect 21192 13258 21220 15030
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21284 14550 21312 14894
rect 21272 14544 21324 14550
rect 21272 14486 21324 14492
rect 21272 14408 21324 14414
rect 21270 14376 21272 14385
rect 21324 14376 21326 14385
rect 21270 14311 21326 14320
rect 21376 13326 21404 14962
rect 21468 13462 21496 15150
rect 21456 13456 21508 13462
rect 21456 13398 21508 13404
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 20811 13084 21119 13104
rect 20811 13082 20817 13084
rect 20873 13082 20897 13084
rect 20953 13082 20977 13084
rect 21033 13082 21057 13084
rect 21113 13082 21119 13084
rect 20873 13030 20875 13082
rect 21055 13030 21057 13082
rect 20811 13028 20817 13030
rect 20873 13028 20897 13030
rect 20953 13028 20977 13030
rect 21033 13028 21057 13030
rect 21113 13028 21119 13030
rect 20811 13008 21119 13028
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20628 12582 20680 12588
rect 20718 12608 20774 12617
rect 20640 12458 20668 12582
rect 20718 12543 20774 12552
rect 20640 12430 20760 12458
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20456 11750 20576 11778
rect 20442 10704 20498 10713
rect 20442 10639 20498 10648
rect 20456 10606 20484 10639
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20548 9217 20576 11750
rect 20640 11286 20668 12310
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20732 11150 20760 12430
rect 20916 12306 20944 12718
rect 21284 12594 21312 13126
rect 21192 12566 21312 12594
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20811 11996 21119 12016
rect 20811 11994 20817 11996
rect 20873 11994 20897 11996
rect 20953 11994 20977 11996
rect 21033 11994 21057 11996
rect 21113 11994 21119 11996
rect 20873 11942 20875 11994
rect 21055 11942 21057 11994
rect 20811 11940 20817 11942
rect 20873 11940 20897 11942
rect 20953 11940 20977 11942
rect 21033 11940 21057 11942
rect 21113 11940 21119 11942
rect 20811 11920 21119 11940
rect 20996 11756 21048 11762
rect 21192 11744 21220 12566
rect 21376 12424 21404 13262
rect 21468 12850 21496 13262
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21456 12708 21508 12714
rect 21456 12650 21508 12656
rect 21048 11716 21220 11744
rect 20996 11698 21048 11704
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20824 11218 20852 11630
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20640 10266 20668 10610
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20732 9466 20760 11086
rect 21192 11082 21220 11716
rect 21284 12396 21404 12424
rect 21284 11626 21312 12396
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21272 11620 21324 11626
rect 21272 11562 21324 11568
rect 21284 11150 21312 11562
rect 21376 11354 21404 12242
rect 21468 12220 21496 12650
rect 21560 12374 21588 17546
rect 21652 17338 21680 17614
rect 21744 17338 21772 17614
rect 21640 17332 21692 17338
rect 21640 17274 21692 17280
rect 21732 17332 21784 17338
rect 21732 17274 21784 17280
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21652 16590 21680 17002
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21548 12368 21600 12374
rect 21548 12310 21600 12316
rect 21468 12192 21588 12220
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21468 11762 21496 12038
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21456 11280 21508 11286
rect 21376 11228 21456 11234
rect 21376 11222 21508 11228
rect 21376 11206 21496 11222
rect 21272 11144 21324 11150
rect 21272 11086 21324 11092
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 20811 10908 21119 10928
rect 20811 10906 20817 10908
rect 20873 10906 20897 10908
rect 20953 10906 20977 10908
rect 21033 10906 21057 10908
rect 21113 10906 21119 10908
rect 20873 10854 20875 10906
rect 21055 10854 21057 10906
rect 20811 10852 20817 10854
rect 20873 10852 20897 10854
rect 20953 10852 20977 10854
rect 21033 10852 21057 10854
rect 21113 10852 21119 10854
rect 20811 10832 21119 10852
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 20811 9820 21119 9840
rect 20811 9818 20817 9820
rect 20873 9818 20897 9820
rect 20953 9818 20977 9820
rect 21033 9818 21057 9820
rect 21113 9818 21119 9820
rect 20873 9766 20875 9818
rect 21055 9766 21057 9818
rect 20811 9764 20817 9766
rect 20873 9764 20897 9766
rect 20953 9764 20977 9766
rect 21033 9764 21057 9766
rect 21113 9764 21119 9766
rect 20811 9744 21119 9764
rect 20732 9438 20852 9466
rect 20824 9382 20852 9438
rect 20628 9376 20680 9382
rect 20812 9376 20864 9382
rect 20680 9324 20760 9330
rect 20628 9318 20760 9324
rect 20812 9318 20864 9324
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20640 9302 20760 9318
rect 20534 9208 20590 9217
rect 20534 9143 20590 9152
rect 20548 8974 20576 9143
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20640 8430 20668 8842
rect 20732 8838 20760 9302
rect 20902 9072 20958 9081
rect 20902 9007 20958 9016
rect 20916 8974 20944 9007
rect 21008 8974 21036 9318
rect 21192 9081 21220 10066
rect 21284 10062 21312 11086
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21272 9920 21324 9926
rect 21376 9908 21404 11206
rect 21560 11150 21588 12192
rect 21548 11144 21600 11150
rect 21454 11112 21510 11121
rect 21548 11086 21600 11092
rect 21454 11047 21510 11056
rect 21468 10062 21496 11047
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21324 9880 21404 9908
rect 21272 9862 21324 9868
rect 21284 9518 21312 9862
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21272 9512 21324 9518
rect 21272 9454 21324 9460
rect 21376 9110 21404 9522
rect 21364 9104 21416 9110
rect 21178 9072 21234 9081
rect 21364 9046 21416 9052
rect 21178 9007 21234 9016
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20811 8732 21119 8752
rect 20811 8730 20817 8732
rect 20873 8730 20897 8732
rect 20953 8730 20977 8732
rect 21033 8730 21057 8732
rect 21113 8730 21119 8732
rect 20873 8678 20875 8730
rect 21055 8678 21057 8730
rect 20811 8676 20817 8678
rect 20873 8676 20897 8678
rect 20953 8676 20977 8678
rect 21033 8676 21057 8678
rect 21113 8676 21119 8678
rect 20811 8656 21119 8676
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20732 7410 20760 7822
rect 20811 7644 21119 7664
rect 20811 7642 20817 7644
rect 20873 7642 20897 7644
rect 20953 7642 20977 7644
rect 21033 7642 21057 7644
rect 21113 7642 21119 7644
rect 20873 7590 20875 7642
rect 21055 7590 21057 7642
rect 20811 7588 20817 7590
rect 20873 7588 20897 7590
rect 20953 7588 20977 7590
rect 21033 7588 21057 7590
rect 21113 7588 21119 7590
rect 20811 7568 21119 7588
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20456 7002 20484 7346
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20732 6934 20760 7346
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20720 6928 20772 6934
rect 20720 6870 20772 6876
rect 20824 6866 20852 7142
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 20088 5846 20116 6666
rect 20076 5840 20128 5846
rect 20076 5782 20128 5788
rect 19668 5664 19748 5692
rect 19800 5704 19852 5710
rect 19616 5646 19668 5652
rect 19800 5646 19852 5652
rect 19812 5302 19840 5646
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19800 5296 19852 5302
rect 19800 5238 19852 5244
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18892 3602 18920 3878
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 15200 3052 15252 3058
rect 15120 3012 15200 3040
rect 15200 2994 15252 3000
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15488 2990 15516 3130
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15846 2748 16154 2768
rect 15846 2746 15852 2748
rect 15908 2746 15932 2748
rect 15988 2746 16012 2748
rect 16068 2746 16092 2748
rect 16148 2746 16154 2748
rect 15908 2694 15910 2746
rect 16090 2694 16092 2746
rect 15846 2692 15852 2694
rect 15908 2692 15932 2694
rect 15988 2692 16012 2694
rect 16068 2692 16092 2694
rect 16148 2692 16154 2694
rect 15846 2672 16154 2692
rect 20180 2650 20208 6666
rect 20456 6322 20484 6734
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20732 4622 20760 6734
rect 20811 6556 21119 6576
rect 20811 6554 20817 6556
rect 20873 6554 20897 6556
rect 20953 6554 20977 6556
rect 21033 6554 21057 6556
rect 21113 6554 21119 6556
rect 20873 6502 20875 6554
rect 21055 6502 21057 6554
rect 20811 6500 20817 6502
rect 20873 6500 20897 6502
rect 20953 6500 20977 6502
rect 21033 6500 21057 6502
rect 21113 6500 21119 6502
rect 20811 6480 21119 6500
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 21192 5914 21220 6190
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 21192 5778 21220 5850
rect 21180 5772 21232 5778
rect 21180 5714 21232 5720
rect 20984 5704 21036 5710
rect 21036 5672 21050 5681
rect 20984 5646 20994 5652
rect 21284 5642 21312 8026
rect 21364 6180 21416 6186
rect 21364 6122 21416 6128
rect 21376 5817 21404 6122
rect 21362 5808 21418 5817
rect 21362 5743 21418 5752
rect 21364 5704 21416 5710
rect 21468 5681 21496 9998
rect 21560 7478 21588 11086
rect 21548 7472 21600 7478
rect 21548 7414 21600 7420
rect 21652 6458 21680 16050
rect 21744 13920 21772 16934
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21836 14278 21864 15370
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21928 14074 21956 17870
rect 22008 17808 22060 17814
rect 22008 17750 22060 17756
rect 22020 17678 22048 17750
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 22112 15502 22140 19230
rect 22204 18834 22232 19774
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22192 18828 22244 18834
rect 22192 18770 22244 18776
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22204 17678 22232 18022
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22296 16522 22324 19450
rect 22388 17882 22416 24686
rect 22480 24206 22508 25638
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 22664 24410 22692 24754
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22468 24200 22520 24206
rect 22468 24142 22520 24148
rect 22468 23112 22520 23118
rect 22468 23054 22520 23060
rect 22480 22166 22508 23054
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22468 22160 22520 22166
rect 22468 22102 22520 22108
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22480 21146 22508 21626
rect 22468 21140 22520 21146
rect 22468 21082 22520 21088
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22480 20398 22508 20878
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22480 19854 22508 20334
rect 22572 20330 22600 22578
rect 22756 21894 22784 28172
rect 22848 25906 22876 30806
rect 22940 29646 22968 31894
rect 23032 31142 23060 35974
rect 23216 35834 23244 37334
rect 23296 37324 23348 37330
rect 23296 37266 23348 37272
rect 23308 37126 23336 37266
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 23296 37120 23348 37126
rect 23296 37062 23348 37068
rect 23400 36938 23428 37198
rect 23308 36922 23428 36938
rect 23296 36916 23428 36922
rect 23348 36910 23428 36916
rect 23296 36858 23348 36864
rect 23492 36786 23520 38150
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23296 36304 23348 36310
rect 23296 36246 23348 36252
rect 23204 35828 23256 35834
rect 23204 35770 23256 35776
rect 23308 35034 23336 36246
rect 23388 35692 23440 35698
rect 23388 35634 23440 35640
rect 23400 35290 23428 35634
rect 23572 35488 23624 35494
rect 23572 35430 23624 35436
rect 23388 35284 23440 35290
rect 23388 35226 23440 35232
rect 23480 35080 23532 35086
rect 23308 35028 23480 35034
rect 23308 35022 23532 35028
rect 23308 35006 23520 35022
rect 23112 32836 23164 32842
rect 23112 32778 23164 32784
rect 23124 32026 23152 32778
rect 23204 32496 23256 32502
rect 23204 32438 23256 32444
rect 23112 32020 23164 32026
rect 23112 31962 23164 31968
rect 23216 31482 23244 32438
rect 23204 31476 23256 31482
rect 23204 31418 23256 31424
rect 23020 31136 23072 31142
rect 23020 31078 23072 31084
rect 22928 29640 22980 29646
rect 22928 29582 22980 29588
rect 22928 28756 22980 28762
rect 22928 28698 22980 28704
rect 22940 27878 22968 28698
rect 22928 27872 22980 27878
rect 22928 27814 22980 27820
rect 22836 25900 22888 25906
rect 22836 25842 22888 25848
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 23124 25498 23152 25842
rect 23308 25514 23336 35006
rect 23584 33522 23612 35430
rect 23676 34202 23704 38626
rect 23756 37868 23808 37874
rect 23756 37810 23808 37816
rect 23768 37466 23796 37810
rect 23940 37664 23992 37670
rect 23940 37606 23992 37612
rect 23756 37460 23808 37466
rect 23756 37402 23808 37408
rect 23952 37330 23980 37606
rect 23940 37324 23992 37330
rect 23940 37266 23992 37272
rect 23756 36032 23808 36038
rect 23756 35974 23808 35980
rect 23768 35698 23796 35974
rect 23756 35692 23808 35698
rect 23756 35634 23808 35640
rect 23848 35624 23900 35630
rect 23848 35566 23900 35572
rect 23860 34610 23888 35566
rect 24124 35012 24176 35018
rect 24124 34954 24176 34960
rect 23848 34604 23900 34610
rect 23848 34546 23900 34552
rect 24032 34604 24084 34610
rect 24032 34546 24084 34552
rect 23664 34196 23716 34202
rect 23664 34138 23716 34144
rect 23572 33516 23624 33522
rect 23572 33458 23624 33464
rect 23480 32904 23532 32910
rect 23480 32846 23532 32852
rect 23388 32768 23440 32774
rect 23388 32710 23440 32716
rect 23400 32434 23428 32710
rect 23492 32570 23520 32846
rect 23480 32564 23532 32570
rect 23480 32506 23532 32512
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 23400 31822 23428 32370
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 23584 31346 23612 33458
rect 23664 31816 23716 31822
rect 23664 31758 23716 31764
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23584 30734 23612 31282
rect 23676 30938 23704 31758
rect 24044 31278 24072 34546
rect 24032 31272 24084 31278
rect 24032 31214 24084 31220
rect 23664 30932 23716 30938
rect 23664 30874 23716 30880
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 23480 30660 23532 30666
rect 23480 30602 23532 30608
rect 23492 30054 23520 30602
rect 23480 30048 23532 30054
rect 23480 29990 23532 29996
rect 23388 29028 23440 29034
rect 23388 28970 23440 28976
rect 23400 28626 23428 28970
rect 23388 28620 23440 28626
rect 23388 28562 23440 28568
rect 23492 28082 23520 29990
rect 23676 29238 23704 30874
rect 23756 30320 23808 30326
rect 23756 30262 23808 30268
rect 23768 29510 23796 30262
rect 23848 30048 23900 30054
rect 23848 29990 23900 29996
rect 23860 29714 23888 29990
rect 23848 29708 23900 29714
rect 23848 29650 23900 29656
rect 23756 29504 23808 29510
rect 23756 29446 23808 29452
rect 23664 29232 23716 29238
rect 23664 29174 23716 29180
rect 23676 28558 23704 29174
rect 23664 28552 23716 28558
rect 23664 28494 23716 28500
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23572 28008 23624 28014
rect 23572 27950 23624 27956
rect 23584 27130 23612 27950
rect 23572 27124 23624 27130
rect 23572 27066 23624 27072
rect 23768 27062 23796 29446
rect 23860 28966 23888 29650
rect 23848 28960 23900 28966
rect 23848 28902 23900 28908
rect 23848 28416 23900 28422
rect 23848 28358 23900 28364
rect 23860 27470 23888 28358
rect 23940 27872 23992 27878
rect 23940 27814 23992 27820
rect 23952 27470 23980 27814
rect 23848 27464 23900 27470
rect 23848 27406 23900 27412
rect 23940 27464 23992 27470
rect 23940 27406 23992 27412
rect 23940 27328 23992 27334
rect 23940 27270 23992 27276
rect 23952 27130 23980 27270
rect 23940 27124 23992 27130
rect 23940 27066 23992 27072
rect 23756 27056 23808 27062
rect 23756 26998 23808 27004
rect 23664 26444 23716 26450
rect 23664 26386 23716 26392
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23480 26240 23532 26246
rect 23480 26182 23532 26188
rect 23112 25492 23164 25498
rect 23112 25434 23164 25440
rect 23216 25486 23336 25514
rect 23112 25220 23164 25226
rect 23112 25162 23164 25168
rect 22928 24608 22980 24614
rect 22928 24550 22980 24556
rect 22940 23730 22968 24550
rect 23124 23730 23152 25162
rect 23216 24274 23244 25486
rect 23296 25356 23348 25362
rect 23296 25298 23348 25304
rect 23308 24750 23336 25298
rect 23492 25294 23520 26182
rect 23584 26042 23612 26318
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23296 24744 23348 24750
rect 23296 24686 23348 24692
rect 23388 24744 23440 24750
rect 23388 24686 23440 24692
rect 23308 24274 23336 24686
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 22928 23724 22980 23730
rect 22928 23666 22980 23672
rect 23112 23724 23164 23730
rect 23112 23666 23164 23672
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 22848 23254 22876 23598
rect 23400 23322 23428 24686
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23492 24206 23520 24550
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 22836 23248 22888 23254
rect 22836 23190 22888 23196
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22652 21412 22704 21418
rect 22652 21354 22704 21360
rect 22664 21146 22692 21354
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22652 20868 22704 20874
rect 22652 20810 22704 20816
rect 22744 20868 22796 20874
rect 22744 20810 22796 20816
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22560 19916 22612 19922
rect 22560 19858 22612 19864
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22480 18290 22508 19790
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22388 17066 22416 17138
rect 22468 17128 22520 17134
rect 22468 17070 22520 17076
rect 22376 17060 22428 17066
rect 22376 17002 22428 17008
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22192 16108 22244 16114
rect 22296 16096 22324 16458
rect 22244 16068 22324 16096
rect 22192 16050 22244 16056
rect 22388 15910 22416 17002
rect 22376 15904 22428 15910
rect 22376 15846 22428 15852
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 22020 14618 22048 15302
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21744 13892 21956 13920
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21744 13394 21772 13738
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21364 5646 21416 5652
rect 21454 5672 21510 5681
rect 20994 5607 21050 5616
rect 21272 5636 21324 5642
rect 21272 5578 21324 5584
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 20811 5468 21119 5488
rect 20811 5466 20817 5468
rect 20873 5466 20897 5468
rect 20953 5466 20977 5468
rect 21033 5466 21057 5468
rect 21113 5466 21119 5468
rect 20873 5414 20875 5466
rect 21055 5414 21057 5466
rect 20811 5412 20817 5414
rect 20873 5412 20897 5414
rect 20953 5412 20977 5414
rect 21033 5412 21057 5414
rect 21113 5412 21119 5414
rect 20811 5392 21119 5412
rect 21192 5234 21220 5510
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21376 4826 21404 5646
rect 21454 5607 21510 5616
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20811 4380 21119 4400
rect 20811 4378 20817 4380
rect 20873 4378 20897 4380
rect 20953 4378 20977 4380
rect 21033 4378 21057 4380
rect 21113 4378 21119 4380
rect 20873 4326 20875 4378
rect 21055 4326 21057 4378
rect 20811 4324 20817 4326
rect 20873 4324 20897 4326
rect 20953 4324 20977 4326
rect 21033 4324 21057 4326
rect 21113 4324 21119 4326
rect 20811 4304 21119 4324
rect 21468 3398 21496 5607
rect 21548 5568 21600 5574
rect 21548 5510 21600 5516
rect 21560 4554 21588 5510
rect 21744 5234 21772 13330
rect 21824 13252 21876 13258
rect 21824 13194 21876 13200
rect 21836 12442 21864 13194
rect 21928 12832 21956 13892
rect 22112 13802 22140 15438
rect 22296 15026 22324 15506
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22192 14952 22244 14958
rect 22190 14920 22192 14929
rect 22244 14920 22246 14929
rect 22190 14855 22246 14864
rect 22100 13796 22152 13802
rect 22100 13738 22152 13744
rect 21928 12804 22048 12832
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 21824 12436 21876 12442
rect 21824 12378 21876 12384
rect 21822 11928 21878 11937
rect 21822 11863 21878 11872
rect 21836 11830 21864 11863
rect 21928 11830 21956 12582
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 21928 11150 21956 11766
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 21824 11076 21876 11082
rect 21824 11018 21876 11024
rect 21836 10130 21864 11018
rect 22020 10810 22048 12804
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 22112 11762 22140 12106
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22098 11656 22154 11665
rect 22098 11591 22154 11600
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 21836 8974 21864 10066
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21928 8498 21956 10542
rect 22112 9674 22140 11591
rect 22204 11218 22232 12718
rect 22296 12714 22324 14962
rect 22388 14822 22416 14962
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22284 12708 22336 12714
rect 22284 12650 22336 12656
rect 22284 12164 22336 12170
rect 22284 12106 22336 12112
rect 22296 11898 22324 12106
rect 22388 12102 22416 13874
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22388 11354 22416 11698
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 22204 10198 22232 11154
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22020 9646 22140 9674
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 21928 7818 21956 8434
rect 21916 7812 21968 7818
rect 21916 7754 21968 7760
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21836 5846 21864 6258
rect 21824 5840 21876 5846
rect 21824 5782 21876 5788
rect 21928 5710 21956 6598
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 22020 5234 22048 9646
rect 22296 9586 22324 9862
rect 22388 9654 22416 11086
rect 22376 9648 22428 9654
rect 22376 9590 22428 9596
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22112 8566 22140 9522
rect 22190 9208 22246 9217
rect 22246 9152 22324 9160
rect 22190 9143 22192 9152
rect 22244 9132 22324 9152
rect 22192 9114 22244 9120
rect 22190 9072 22246 9081
rect 22190 9007 22192 9016
rect 22244 9007 22246 9016
rect 22192 8978 22244 8984
rect 22100 8560 22152 8566
rect 22100 8502 22152 8508
rect 22112 7410 22140 8502
rect 22296 8022 22324 9132
rect 22388 8838 22416 9590
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22480 8566 22508 17070
rect 22572 8906 22600 19858
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 22468 8560 22520 8566
rect 22468 8502 22520 8508
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22284 8016 22336 8022
rect 22204 7976 22284 8004
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22112 6798 22140 7346
rect 22204 6798 22232 7976
rect 22284 7958 22336 7964
rect 22480 7818 22508 8366
rect 22376 7812 22428 7818
rect 22376 7754 22428 7760
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22112 6322 22140 6734
rect 22204 6662 22232 6734
rect 22296 6730 22324 7686
rect 22388 7002 22416 7754
rect 22376 6996 22428 7002
rect 22376 6938 22428 6944
rect 22284 6724 22336 6730
rect 22284 6666 22336 6672
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22284 6180 22336 6186
rect 22284 6122 22336 6128
rect 22296 5817 22324 6122
rect 22282 5808 22338 5817
rect 22282 5743 22338 5752
rect 22296 5710 22324 5743
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 22112 5234 22140 5510
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22572 5166 22600 5646
rect 22560 5160 22612 5166
rect 22560 5102 22612 5108
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22572 4622 22600 4966
rect 22664 4842 22692 20810
rect 22756 20330 22784 20810
rect 22744 20324 22796 20330
rect 22744 20266 22796 20272
rect 22756 19514 22784 20266
rect 22848 20262 22876 23190
rect 23388 23044 23440 23050
rect 23388 22986 23440 22992
rect 23400 22778 23428 22986
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23112 22500 23164 22506
rect 23112 22442 23164 22448
rect 23020 22432 23072 22438
rect 23020 22374 23072 22380
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 22940 20942 22968 21830
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 22928 20800 22980 20806
rect 22928 20742 22980 20748
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22756 17882 22784 18566
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22848 17814 22876 20198
rect 22836 17808 22888 17814
rect 22756 17756 22836 17762
rect 22756 17750 22888 17756
rect 22756 17734 22876 17750
rect 22756 16726 22784 17734
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 22744 16720 22796 16726
rect 22744 16662 22796 16668
rect 22744 16584 22796 16590
rect 22744 16526 22796 16532
rect 22756 13530 22784 16526
rect 22848 16250 22876 17614
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22836 15904 22888 15910
rect 22836 15846 22888 15852
rect 22848 15026 22876 15846
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22744 13524 22796 13530
rect 22744 13466 22796 13472
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22756 11150 22784 12174
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22744 8900 22796 8906
rect 22744 8842 22796 8848
rect 22756 6662 22784 8842
rect 22836 7948 22888 7954
rect 22836 7890 22888 7896
rect 22848 6798 22876 7890
rect 22940 7478 22968 20742
rect 23032 20466 23060 22374
rect 23124 22234 23152 22442
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 23124 20210 23152 22170
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23400 21690 23428 21966
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23204 21004 23256 21010
rect 23204 20946 23256 20952
rect 23216 20466 23244 20946
rect 23296 20936 23348 20942
rect 23296 20878 23348 20884
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 23032 20182 23152 20210
rect 23032 18630 23060 20182
rect 23112 20052 23164 20058
rect 23112 19994 23164 20000
rect 23124 19854 23152 19994
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 23124 18290 23152 19790
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23112 18284 23164 18290
rect 23112 18226 23164 18232
rect 23216 18222 23244 18770
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 23020 18148 23072 18154
rect 23020 18090 23072 18096
rect 23032 17134 23060 18090
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 23124 17202 23152 17478
rect 23216 17270 23244 18158
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 23032 15638 23060 17070
rect 23124 16794 23152 17138
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 23124 16250 23152 16526
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23020 15632 23072 15638
rect 23020 15574 23072 15580
rect 23216 15502 23244 17206
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 23020 15360 23072 15366
rect 23020 15302 23072 15308
rect 23032 11937 23060 15302
rect 23216 15178 23244 15438
rect 23124 15150 23244 15178
rect 23124 14958 23152 15150
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 23216 14385 23244 14962
rect 23202 14376 23258 14385
rect 23202 14311 23258 14320
rect 23216 13394 23244 14311
rect 23204 13388 23256 13394
rect 23204 13330 23256 13336
rect 23018 11928 23074 11937
rect 23018 11863 23074 11872
rect 23204 9444 23256 9450
rect 23204 9386 23256 9392
rect 23112 9104 23164 9110
rect 23112 9046 23164 9052
rect 23124 8537 23152 9046
rect 23216 8974 23244 9386
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23110 8528 23166 8537
rect 23020 8492 23072 8498
rect 23110 8463 23112 8472
rect 23020 8434 23072 8440
rect 23164 8463 23166 8472
rect 23112 8434 23164 8440
rect 23032 8106 23060 8434
rect 23032 8078 23152 8106
rect 23308 8090 23336 20878
rect 23400 20058 23428 21626
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23400 18834 23428 19790
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23400 17066 23428 18226
rect 23388 17060 23440 17066
rect 23388 17002 23440 17008
rect 23492 16794 23520 24006
rect 23584 17882 23612 25094
rect 23676 24818 23704 26386
rect 23756 25288 23808 25294
rect 23756 25230 23808 25236
rect 23664 24812 23716 24818
rect 23664 24754 23716 24760
rect 23768 24410 23796 25230
rect 23756 24404 23808 24410
rect 23756 24346 23808 24352
rect 23756 23316 23808 23322
rect 23756 23258 23808 23264
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23676 22778 23704 22918
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23768 22710 23796 23258
rect 23756 22704 23808 22710
rect 23756 22646 23808 22652
rect 23768 22166 23796 22646
rect 23756 22160 23808 22166
rect 23756 22102 23808 22108
rect 24044 22094 24072 31214
rect 24136 30258 24164 34954
rect 24320 34474 24348 38898
rect 24412 35222 24440 38898
rect 24492 38344 24544 38350
rect 24492 38286 24544 38292
rect 24504 37466 24532 38286
rect 24492 37460 24544 37466
rect 24492 37402 24544 37408
rect 24492 37256 24544 37262
rect 24490 37224 24492 37233
rect 24544 37224 24546 37233
rect 24490 37159 24546 37168
rect 24492 36916 24544 36922
rect 24492 36858 24544 36864
rect 24504 36174 24532 36858
rect 24596 36378 24624 39358
rect 24688 38962 24716 39460
rect 24768 39442 24820 39448
rect 24872 39370 24900 39578
rect 24860 39364 24912 39370
rect 24860 39306 24912 39312
rect 24676 38956 24728 38962
rect 24676 38898 24728 38904
rect 24676 38344 24728 38350
rect 24676 38286 24728 38292
rect 24584 36372 24636 36378
rect 24584 36314 24636 36320
rect 24492 36168 24544 36174
rect 24492 36110 24544 36116
rect 24400 35216 24452 35222
rect 24400 35158 24452 35164
rect 24308 34468 24360 34474
rect 24308 34410 24360 34416
rect 24412 33930 24440 35158
rect 24504 35018 24532 36110
rect 24492 35012 24544 35018
rect 24492 34954 24544 34960
rect 24688 34746 24716 38286
rect 24768 37868 24820 37874
rect 24768 37810 24820 37816
rect 24676 34740 24728 34746
rect 24676 34682 24728 34688
rect 24492 34604 24544 34610
rect 24492 34546 24544 34552
rect 24504 34202 24532 34546
rect 24676 34468 24728 34474
rect 24676 34410 24728 34416
rect 24492 34196 24544 34202
rect 24492 34138 24544 34144
rect 24400 33924 24452 33930
rect 24400 33866 24452 33872
rect 24688 33522 24716 34410
rect 24676 33516 24728 33522
rect 24676 33458 24728 33464
rect 24400 33312 24452 33318
rect 24400 33254 24452 33260
rect 24412 32366 24440 33254
rect 24780 33046 24808 37810
rect 24872 36854 24900 39306
rect 25056 39001 25084 41006
rect 25148 41002 25176 41618
rect 25136 40996 25188 41002
rect 25136 40938 25188 40944
rect 25136 40452 25188 40458
rect 25136 40394 25188 40400
rect 25148 39642 25176 40394
rect 25136 39636 25188 39642
rect 25136 39578 25188 39584
rect 25042 38992 25098 39001
rect 25042 38927 25098 38936
rect 24952 38752 25004 38758
rect 24952 38694 25004 38700
rect 24964 38350 24992 38694
rect 24952 38344 25004 38350
rect 24952 38286 25004 38292
rect 24952 37256 25004 37262
rect 24952 37198 25004 37204
rect 24860 36848 24912 36854
rect 24860 36790 24912 36796
rect 24860 36236 24912 36242
rect 24964 36224 24992 37198
rect 25056 36310 25084 38927
rect 25044 36304 25096 36310
rect 25044 36246 25096 36252
rect 24912 36196 24992 36224
rect 24860 36178 24912 36184
rect 24872 35154 24900 36178
rect 25136 35692 25188 35698
rect 25136 35634 25188 35640
rect 24952 35556 25004 35562
rect 24952 35498 25004 35504
rect 24860 35148 24912 35154
rect 24860 35090 24912 35096
rect 24964 35086 24992 35498
rect 25148 35290 25176 35634
rect 25136 35284 25188 35290
rect 25136 35226 25188 35232
rect 24952 35080 25004 35086
rect 24952 35022 25004 35028
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 24872 33998 24900 34546
rect 25240 34490 25268 41686
rect 25516 41614 25544 43046
rect 25608 42922 25636 43182
rect 25700 43110 25728 43250
rect 26068 43194 26096 43726
rect 26240 43716 26292 43722
rect 26240 43658 26292 43664
rect 26068 43166 26188 43194
rect 25688 43104 25740 43110
rect 25688 43046 25740 43052
rect 25776 43004 26084 43024
rect 25776 43002 25782 43004
rect 25838 43002 25862 43004
rect 25918 43002 25942 43004
rect 25998 43002 26022 43004
rect 26078 43002 26084 43004
rect 25838 42950 25840 43002
rect 26020 42950 26022 43002
rect 25776 42948 25782 42950
rect 25838 42948 25862 42950
rect 25918 42948 25942 42950
rect 25998 42948 26022 42950
rect 26078 42948 26084 42950
rect 25776 42928 26084 42948
rect 25608 42894 25728 42922
rect 25596 42696 25648 42702
rect 25596 42638 25648 42644
rect 25504 41608 25556 41614
rect 25502 41576 25504 41585
rect 25556 41576 25558 41585
rect 25502 41511 25558 41520
rect 25412 40656 25464 40662
rect 25412 40598 25464 40604
rect 25502 40624 25558 40633
rect 25320 39840 25372 39846
rect 25320 39782 25372 39788
rect 25332 39574 25360 39782
rect 25320 39568 25372 39574
rect 25320 39510 25372 39516
rect 25332 37618 25360 39510
rect 25424 39438 25452 40598
rect 25502 40559 25504 40568
rect 25556 40559 25558 40568
rect 25504 40530 25556 40536
rect 25608 39624 25636 42638
rect 25700 42566 25728 42894
rect 25872 42832 25924 42838
rect 25872 42774 25924 42780
rect 25884 42702 25912 42774
rect 25872 42696 25924 42702
rect 25872 42638 25924 42644
rect 26160 42634 26188 43166
rect 26252 42702 26280 43658
rect 26344 43450 26372 44746
rect 26792 44736 26844 44742
rect 26792 44678 26844 44684
rect 26608 43648 26660 43654
rect 26608 43590 26660 43596
rect 26332 43444 26384 43450
rect 26332 43386 26384 43392
rect 26516 43444 26568 43450
rect 26516 43386 26568 43392
rect 26332 43172 26384 43178
rect 26332 43114 26384 43120
rect 26240 42696 26292 42702
rect 26240 42638 26292 42644
rect 26148 42628 26200 42634
rect 26148 42570 26200 42576
rect 25688 42560 25740 42566
rect 25688 42502 25740 42508
rect 25700 41120 25728 42502
rect 25776 41916 26084 41936
rect 25776 41914 25782 41916
rect 25838 41914 25862 41916
rect 25918 41914 25942 41916
rect 25998 41914 26022 41916
rect 26078 41914 26084 41916
rect 25838 41862 25840 41914
rect 26020 41862 26022 41914
rect 25776 41860 25782 41862
rect 25838 41860 25862 41862
rect 25918 41860 25942 41862
rect 25998 41860 26022 41862
rect 26078 41860 26084 41862
rect 25776 41840 26084 41860
rect 26240 41540 26292 41546
rect 26240 41482 26292 41488
rect 26252 41274 26280 41482
rect 26240 41268 26292 41274
rect 26240 41210 26292 41216
rect 25780 41132 25832 41138
rect 25700 41092 25780 41120
rect 25780 41074 25832 41080
rect 25686 41032 25742 41041
rect 25686 40967 25742 40976
rect 25516 39596 25636 39624
rect 25412 39432 25464 39438
rect 25412 39374 25464 39380
rect 25516 39370 25544 39596
rect 25596 39500 25648 39506
rect 25700 39488 25728 40967
rect 25776 40828 26084 40848
rect 25776 40826 25782 40828
rect 25838 40826 25862 40828
rect 25918 40826 25942 40828
rect 25998 40826 26022 40828
rect 26078 40826 26084 40828
rect 25838 40774 25840 40826
rect 26020 40774 26022 40826
rect 25776 40772 25782 40774
rect 25838 40772 25862 40774
rect 25918 40772 25942 40774
rect 25998 40772 26022 40774
rect 26078 40772 26084 40774
rect 25776 40752 26084 40772
rect 25872 40520 25924 40526
rect 25872 40462 25924 40468
rect 25884 40186 25912 40462
rect 26240 40384 26292 40390
rect 26240 40326 26292 40332
rect 26252 40186 26280 40326
rect 25872 40180 25924 40186
rect 25872 40122 25924 40128
rect 26240 40180 26292 40186
rect 26240 40122 26292 40128
rect 26240 39840 26292 39846
rect 26240 39782 26292 39788
rect 25776 39740 26084 39760
rect 25776 39738 25782 39740
rect 25838 39738 25862 39740
rect 25918 39738 25942 39740
rect 25998 39738 26022 39740
rect 26078 39738 26084 39740
rect 25838 39686 25840 39738
rect 26020 39686 26022 39738
rect 25776 39684 25782 39686
rect 25838 39684 25862 39686
rect 25918 39684 25942 39686
rect 25998 39684 26022 39686
rect 26078 39684 26084 39686
rect 25776 39664 26084 39684
rect 25964 39568 26016 39574
rect 26252 39522 26280 39782
rect 25964 39510 26016 39516
rect 25700 39460 25820 39488
rect 25596 39442 25648 39448
rect 25504 39364 25556 39370
rect 25504 39306 25556 39312
rect 25504 38956 25556 38962
rect 25504 38898 25556 38904
rect 25412 38820 25464 38826
rect 25412 38762 25464 38768
rect 25424 37942 25452 38762
rect 25516 38350 25544 38898
rect 25608 38894 25636 39442
rect 25688 39364 25740 39370
rect 25688 39306 25740 39312
rect 25700 38962 25728 39306
rect 25792 38962 25820 39460
rect 25976 39438 26004 39510
rect 26068 39494 26280 39522
rect 25964 39432 26016 39438
rect 25964 39374 26016 39380
rect 26068 39302 26096 39494
rect 26148 39432 26200 39438
rect 26148 39374 26200 39380
rect 26160 39302 26188 39374
rect 26056 39296 26108 39302
rect 26056 39238 26108 39244
rect 26148 39296 26200 39302
rect 26148 39238 26200 39244
rect 26160 38962 26188 39238
rect 26344 39030 26372 43114
rect 26422 41304 26478 41313
rect 26422 41239 26424 41248
rect 26476 41239 26478 41248
rect 26424 41210 26476 41216
rect 26424 41064 26476 41070
rect 26424 41006 26476 41012
rect 26436 40526 26464 41006
rect 26528 40730 26556 43386
rect 26620 42566 26648 43590
rect 26804 43314 26832 44678
rect 27068 43784 27120 43790
rect 27068 43726 27120 43732
rect 27080 43314 27108 43726
rect 26792 43308 26844 43314
rect 26792 43250 26844 43256
rect 26976 43308 27028 43314
rect 26976 43250 27028 43256
rect 27068 43308 27120 43314
rect 27068 43250 27120 43256
rect 26700 42696 26752 42702
rect 26700 42638 26752 42644
rect 26608 42560 26660 42566
rect 26608 42502 26660 42508
rect 26712 42362 26740 42638
rect 26700 42356 26752 42362
rect 26700 42298 26752 42304
rect 26792 42356 26844 42362
rect 26792 42298 26844 42304
rect 26608 41132 26660 41138
rect 26608 41074 26660 41080
rect 26516 40724 26568 40730
rect 26516 40666 26568 40672
rect 26424 40520 26476 40526
rect 26424 40462 26476 40468
rect 26516 40452 26568 40458
rect 26516 40394 26568 40400
rect 26528 40202 26556 40394
rect 26436 40174 26556 40202
rect 26332 39024 26384 39030
rect 26332 38966 26384 38972
rect 25688 38956 25740 38962
rect 25688 38898 25740 38904
rect 25780 38956 25832 38962
rect 25780 38898 25832 38904
rect 26148 38956 26200 38962
rect 26148 38898 26200 38904
rect 25596 38888 25648 38894
rect 25596 38830 25648 38836
rect 25504 38344 25556 38350
rect 25504 38286 25556 38292
rect 25412 37936 25464 37942
rect 25412 37878 25464 37884
rect 25332 37590 25544 37618
rect 25148 34462 25268 34490
rect 24860 33992 24912 33998
rect 24860 33934 24912 33940
rect 24872 33318 24900 33934
rect 24952 33924 25004 33930
rect 24952 33866 25004 33872
rect 24860 33312 24912 33318
rect 24860 33254 24912 33260
rect 24768 33040 24820 33046
rect 24768 32982 24820 32988
rect 24400 32360 24452 32366
rect 24400 32302 24452 32308
rect 24412 31822 24440 32302
rect 24780 32230 24808 32982
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 24768 32224 24820 32230
rect 24688 32172 24768 32178
rect 24688 32166 24820 32172
rect 24688 32150 24808 32166
rect 24688 32026 24716 32150
rect 24872 32026 24900 32846
rect 24676 32020 24728 32026
rect 24676 31962 24728 31968
rect 24860 32020 24912 32026
rect 24860 31962 24912 31968
rect 24400 31816 24452 31822
rect 24400 31758 24452 31764
rect 24216 31272 24268 31278
rect 24216 31214 24268 31220
rect 24860 31272 24912 31278
rect 24860 31214 24912 31220
rect 24228 30258 24256 31214
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24124 30252 24176 30258
rect 24124 30194 24176 30200
rect 24216 30252 24268 30258
rect 24216 30194 24268 30200
rect 24596 29850 24624 30670
rect 24872 30258 24900 31214
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24768 30184 24820 30190
rect 24768 30126 24820 30132
rect 24584 29844 24636 29850
rect 24584 29786 24636 29792
rect 24780 29782 24808 30126
rect 24872 29782 24900 30194
rect 24768 29776 24820 29782
rect 24768 29718 24820 29724
rect 24860 29776 24912 29782
rect 24860 29718 24912 29724
rect 24676 29640 24728 29646
rect 24676 29582 24728 29588
rect 24492 29232 24544 29238
rect 24492 29174 24544 29180
rect 24216 29164 24268 29170
rect 24216 29106 24268 29112
rect 24124 28416 24176 28422
rect 24124 28358 24176 28364
rect 24136 28218 24164 28358
rect 24124 28212 24176 28218
rect 24124 28154 24176 28160
rect 24228 24682 24256 29106
rect 24504 28150 24532 29174
rect 24688 29170 24716 29582
rect 24676 29164 24728 29170
rect 24676 29106 24728 29112
rect 24780 29034 24808 29718
rect 24872 29102 24900 29718
rect 24964 29714 24992 33866
rect 25148 32978 25176 34462
rect 25228 34400 25280 34406
rect 25228 34342 25280 34348
rect 25240 34066 25268 34342
rect 25228 34060 25280 34066
rect 25228 34002 25280 34008
rect 25516 33522 25544 37590
rect 25608 36666 25636 38830
rect 25700 37874 25728 38898
rect 25792 38826 25820 38898
rect 25780 38820 25832 38826
rect 25780 38762 25832 38768
rect 25776 38652 26084 38672
rect 25776 38650 25782 38652
rect 25838 38650 25862 38652
rect 25918 38650 25942 38652
rect 25998 38650 26022 38652
rect 26078 38650 26084 38652
rect 25838 38598 25840 38650
rect 26020 38598 26022 38650
rect 25776 38596 25782 38598
rect 25838 38596 25862 38598
rect 25918 38596 25942 38598
rect 25998 38596 26022 38598
rect 26078 38596 26084 38598
rect 25776 38576 26084 38596
rect 25688 37868 25740 37874
rect 25688 37810 25740 37816
rect 25700 37244 25728 37810
rect 25776 37564 26084 37584
rect 25776 37562 25782 37564
rect 25838 37562 25862 37564
rect 25918 37562 25942 37564
rect 25998 37562 26022 37564
rect 26078 37562 26084 37564
rect 25838 37510 25840 37562
rect 26020 37510 26022 37562
rect 25776 37508 25782 37510
rect 25838 37508 25862 37510
rect 25918 37508 25942 37510
rect 25998 37508 26022 37510
rect 26078 37508 26084 37510
rect 25776 37488 26084 37508
rect 26160 37330 26188 38898
rect 26332 38820 26384 38826
rect 26332 38762 26384 38768
rect 26148 37324 26200 37330
rect 26148 37266 26200 37272
rect 25780 37256 25832 37262
rect 25700 37216 25780 37244
rect 25700 36786 25728 37216
rect 25780 37198 25832 37204
rect 25780 37120 25832 37126
rect 25780 37062 25832 37068
rect 25688 36780 25740 36786
rect 25688 36722 25740 36728
rect 25792 36718 25820 37062
rect 26056 36848 26108 36854
rect 26056 36790 26108 36796
rect 25780 36712 25832 36718
rect 25608 36660 25780 36666
rect 25608 36654 25832 36660
rect 26068 36666 26096 36790
rect 26160 36786 26188 37266
rect 26148 36780 26200 36786
rect 26148 36722 26200 36728
rect 25608 36638 25820 36654
rect 26068 36638 26280 36666
rect 25700 36242 25728 36638
rect 25776 36476 26084 36496
rect 25776 36474 25782 36476
rect 25838 36474 25862 36476
rect 25918 36474 25942 36476
rect 25998 36474 26022 36476
rect 26078 36474 26084 36476
rect 25838 36422 25840 36474
rect 26020 36422 26022 36474
rect 25776 36420 25782 36422
rect 25838 36420 25862 36422
rect 25918 36420 25942 36422
rect 25998 36420 26022 36422
rect 26078 36420 26084 36422
rect 25776 36400 26084 36420
rect 25688 36236 25740 36242
rect 25688 36178 25740 36184
rect 25776 35388 26084 35408
rect 25776 35386 25782 35388
rect 25838 35386 25862 35388
rect 25918 35386 25942 35388
rect 25998 35386 26022 35388
rect 26078 35386 26084 35388
rect 25838 35334 25840 35386
rect 26020 35334 26022 35386
rect 25776 35332 25782 35334
rect 25838 35332 25862 35334
rect 25918 35332 25942 35334
rect 25998 35332 26022 35334
rect 26078 35332 26084 35334
rect 25776 35312 26084 35332
rect 25776 34300 26084 34320
rect 25776 34298 25782 34300
rect 25838 34298 25862 34300
rect 25918 34298 25942 34300
rect 25998 34298 26022 34300
rect 26078 34298 26084 34300
rect 25838 34246 25840 34298
rect 26020 34246 26022 34298
rect 25776 34244 25782 34246
rect 25838 34244 25862 34246
rect 25918 34244 25942 34246
rect 25998 34244 26022 34246
rect 26078 34244 26084 34246
rect 25776 34224 26084 34244
rect 26148 33924 26200 33930
rect 26148 33866 26200 33872
rect 26160 33658 26188 33866
rect 26148 33652 26200 33658
rect 26148 33594 26200 33600
rect 25504 33516 25556 33522
rect 25504 33458 25556 33464
rect 25136 32972 25188 32978
rect 25136 32914 25188 32920
rect 25148 31754 25176 32914
rect 25228 32768 25280 32774
rect 25228 32710 25280 32716
rect 25056 31726 25176 31754
rect 24952 29708 25004 29714
rect 24952 29650 25004 29656
rect 25056 29594 25084 31726
rect 25136 30660 25188 30666
rect 25136 30602 25188 30608
rect 25148 30394 25176 30602
rect 25136 30388 25188 30394
rect 25136 30330 25188 30336
rect 24964 29578 25084 29594
rect 24952 29572 25084 29578
rect 25004 29566 25084 29572
rect 24952 29514 25004 29520
rect 24860 29096 24912 29102
rect 24860 29038 24912 29044
rect 24584 29028 24636 29034
rect 24584 28970 24636 28976
rect 24768 29028 24820 29034
rect 24768 28970 24820 28976
rect 24492 28144 24544 28150
rect 24492 28086 24544 28092
rect 24400 27328 24452 27334
rect 24400 27270 24452 27276
rect 24308 26988 24360 26994
rect 24308 26930 24360 26936
rect 24216 24676 24268 24682
rect 24216 24618 24268 24624
rect 23952 22066 24072 22094
rect 23952 21962 23980 22066
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 23940 21956 23992 21962
rect 23940 21898 23992 21904
rect 24228 21350 24256 21966
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 23756 21004 23808 21010
rect 23756 20946 23808 20952
rect 23768 20262 23796 20946
rect 24032 20936 24084 20942
rect 24032 20878 24084 20884
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23756 19916 23808 19922
rect 23756 19858 23808 19864
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23676 19310 23704 19382
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23676 18766 23704 19110
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23768 18222 23796 19858
rect 23940 19848 23992 19854
rect 23940 19790 23992 19796
rect 23952 19310 23980 19790
rect 23940 19304 23992 19310
rect 23940 19246 23992 19252
rect 23952 18630 23980 19246
rect 23940 18624 23992 18630
rect 23940 18566 23992 18572
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23480 16788 23532 16794
rect 23480 16730 23532 16736
rect 23388 16720 23440 16726
rect 23388 16662 23440 16668
rect 23400 16522 23428 16662
rect 23584 16658 23612 17682
rect 23664 17604 23716 17610
rect 23664 17546 23716 17552
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23400 15502 23428 16050
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23400 14278 23428 15438
rect 23492 15026 23520 15438
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23492 14006 23520 14350
rect 23584 14346 23612 15302
rect 23572 14340 23624 14346
rect 23572 14282 23624 14288
rect 23480 14000 23532 14006
rect 23480 13942 23532 13948
rect 23676 13530 23704 17546
rect 23756 17128 23808 17134
rect 23756 17070 23808 17076
rect 23768 16046 23796 17070
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 23768 15706 23796 15982
rect 23756 15700 23808 15706
rect 23756 15642 23808 15648
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23768 13938 23796 14758
rect 23756 13932 23808 13938
rect 23756 13874 23808 13880
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23492 8430 23520 8910
rect 23768 8430 23796 12106
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 22928 7472 22980 7478
rect 22928 7414 22980 7420
rect 23032 6798 23060 7482
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 23124 6730 23152 8078
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 23216 6798 23244 7822
rect 23480 7812 23532 7818
rect 23480 7754 23532 7760
rect 23492 7478 23520 7754
rect 23480 7472 23532 7478
rect 23480 7414 23532 7420
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23400 7002 23428 7346
rect 23388 6996 23440 7002
rect 23388 6938 23440 6944
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23112 6724 23164 6730
rect 23112 6666 23164 6672
rect 22744 6656 22796 6662
rect 22744 6598 22796 6604
rect 22928 6656 22980 6662
rect 22928 6598 22980 6604
rect 22744 6316 22796 6322
rect 22744 6258 22796 6264
rect 22756 5914 22784 6258
rect 22744 5908 22796 5914
rect 22744 5850 22796 5856
rect 22940 5642 22968 6598
rect 22928 5636 22980 5642
rect 22928 5578 22980 5584
rect 22664 4826 22784 4842
rect 22664 4820 22796 4826
rect 22664 4814 22744 4820
rect 22744 4762 22796 4768
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 21548 4548 21600 4554
rect 21548 4490 21600 4496
rect 23124 4486 23152 6666
rect 23216 5710 23244 6734
rect 23584 6118 23612 7822
rect 23768 7410 23796 8366
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 23204 5704 23256 5710
rect 23204 5646 23256 5652
rect 23860 5302 23888 18226
rect 23952 17921 23980 18226
rect 23938 17912 23994 17921
rect 23938 17847 23994 17856
rect 23938 17776 23994 17785
rect 23938 17711 23994 17720
rect 23952 15434 23980 17711
rect 23940 15428 23992 15434
rect 23940 15370 23992 15376
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 23952 11762 23980 13942
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23952 11218 23980 11698
rect 24044 11354 24072 20878
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24228 18426 24256 19314
rect 24216 18420 24268 18426
rect 24216 18362 24268 18368
rect 24216 17672 24268 17678
rect 24216 17614 24268 17620
rect 24124 16448 24176 16454
rect 24124 16390 24176 16396
rect 24136 16250 24164 16390
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 24136 15570 24164 16186
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24228 15162 24256 17614
rect 24320 16794 24348 26930
rect 24412 26042 24440 27270
rect 24492 26308 24544 26314
rect 24492 26250 24544 26256
rect 24400 26036 24452 26042
rect 24400 25978 24452 25984
rect 24400 25832 24452 25838
rect 24400 25774 24452 25780
rect 24412 21146 24440 25774
rect 24504 23866 24532 26250
rect 24596 24206 24624 28970
rect 24780 28558 24808 28970
rect 24872 28762 24900 29038
rect 24860 28756 24912 28762
rect 24860 28698 24912 28704
rect 24858 28656 24914 28665
rect 24858 28591 24914 28600
rect 24768 28552 24820 28558
rect 24768 28494 24820 28500
rect 24872 28082 24900 28591
rect 24964 28218 24992 29514
rect 25044 29504 25096 29510
rect 25044 29446 25096 29452
rect 25056 28422 25084 29446
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 24952 28212 25004 28218
rect 24952 28154 25004 28160
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 24872 27538 24900 28018
rect 24860 27532 24912 27538
rect 24860 27474 24912 27480
rect 25044 27464 25096 27470
rect 25044 27406 25096 27412
rect 24676 26852 24728 26858
rect 24676 26794 24728 26800
rect 24688 25838 24716 26794
rect 24676 25832 24728 25838
rect 24676 25774 24728 25780
rect 24688 25362 24716 25774
rect 25056 25770 25084 27406
rect 25136 27328 25188 27334
rect 25136 27270 25188 27276
rect 25148 27062 25176 27270
rect 25136 27056 25188 27062
rect 25136 26998 25188 27004
rect 25240 26382 25268 32710
rect 25516 32366 25544 33458
rect 25596 33312 25648 33318
rect 25596 33254 25648 33260
rect 25608 32434 25636 33254
rect 25776 33212 26084 33232
rect 25776 33210 25782 33212
rect 25838 33210 25862 33212
rect 25918 33210 25942 33212
rect 25998 33210 26022 33212
rect 26078 33210 26084 33212
rect 25838 33158 25840 33210
rect 26020 33158 26022 33210
rect 25776 33156 25782 33158
rect 25838 33156 25862 33158
rect 25918 33156 25942 33158
rect 25998 33156 26022 33158
rect 26078 33156 26084 33158
rect 25776 33136 26084 33156
rect 26252 32978 26280 36638
rect 26344 33930 26372 38762
rect 26436 38554 26464 40174
rect 26516 40112 26568 40118
rect 26516 40054 26568 40060
rect 26424 38548 26476 38554
rect 26424 38490 26476 38496
rect 26528 38350 26556 40054
rect 26620 39438 26648 41074
rect 26804 40186 26832 42298
rect 26988 42226 27016 43250
rect 27160 43104 27212 43110
rect 27160 43046 27212 43052
rect 27172 42770 27200 43046
rect 27160 42764 27212 42770
rect 27160 42706 27212 42712
rect 26976 42220 27028 42226
rect 26976 42162 27028 42168
rect 26976 42084 27028 42090
rect 26976 42026 27028 42032
rect 26988 41682 27016 42026
rect 26976 41676 27028 41682
rect 26976 41618 27028 41624
rect 27160 41540 27212 41546
rect 27160 41482 27212 41488
rect 26976 41472 27028 41478
rect 26976 41414 27028 41420
rect 26988 41206 27016 41414
rect 26976 41200 27028 41206
rect 26976 41142 27028 41148
rect 27172 40662 27200 41482
rect 27160 40656 27212 40662
rect 27160 40598 27212 40604
rect 26884 40520 26936 40526
rect 26884 40462 26936 40468
rect 26792 40180 26844 40186
rect 26792 40122 26844 40128
rect 26700 40112 26752 40118
rect 26700 40054 26752 40060
rect 26790 40080 26846 40089
rect 26608 39432 26660 39438
rect 26608 39374 26660 39380
rect 26712 39137 26740 40054
rect 26790 40015 26846 40024
rect 26804 39506 26832 40015
rect 26792 39500 26844 39506
rect 26792 39442 26844 39448
rect 26698 39128 26754 39137
rect 26698 39063 26754 39072
rect 26516 38344 26568 38350
rect 26516 38286 26568 38292
rect 26528 37874 26556 38286
rect 26896 38010 26924 40462
rect 27068 40384 27120 40390
rect 27068 40326 27120 40332
rect 26976 40044 27028 40050
rect 26976 39986 27028 39992
rect 26988 38554 27016 39986
rect 27080 38962 27108 40326
rect 27160 40180 27212 40186
rect 27160 40122 27212 40128
rect 27068 38956 27120 38962
rect 27068 38898 27120 38904
rect 27068 38752 27120 38758
rect 27068 38694 27120 38700
rect 26976 38548 27028 38554
rect 26976 38490 27028 38496
rect 27080 38350 27108 38694
rect 27172 38418 27200 40122
rect 27264 39846 27292 45222
rect 27448 44985 27476 45426
rect 27528 45416 27580 45422
rect 27526 45384 27528 45393
rect 27580 45384 27582 45393
rect 27526 45319 27582 45328
rect 27528 45280 27580 45286
rect 27528 45222 27580 45228
rect 27540 45082 27568 45222
rect 27528 45076 27580 45082
rect 27528 45018 27580 45024
rect 27434 44976 27490 44985
rect 27434 44911 27490 44920
rect 27528 44736 27580 44742
rect 27528 44678 27580 44684
rect 27540 44538 27568 44678
rect 27528 44532 27580 44538
rect 27528 44474 27580 44480
rect 27434 42800 27490 42809
rect 27434 42735 27436 42744
rect 27488 42735 27490 42744
rect 27436 42706 27488 42712
rect 27344 42696 27396 42702
rect 27344 42638 27396 42644
rect 27356 41818 27384 42638
rect 27528 42560 27580 42566
rect 27528 42502 27580 42508
rect 27436 42288 27488 42294
rect 27434 42256 27436 42265
rect 27488 42256 27490 42265
rect 27434 42191 27490 42200
rect 27344 41812 27396 41818
rect 27344 41754 27396 41760
rect 27540 41614 27568 42502
rect 27528 41608 27580 41614
rect 27434 41576 27490 41585
rect 27528 41550 27580 41556
rect 27434 41511 27490 41520
rect 27342 40352 27398 40361
rect 27342 40287 27398 40296
rect 27356 40186 27384 40287
rect 27344 40180 27396 40186
rect 27344 40122 27396 40128
rect 27252 39840 27304 39846
rect 27252 39782 27304 39788
rect 27252 39432 27304 39438
rect 27448 39386 27476 41511
rect 27632 39642 27660 45426
rect 27710 45384 27766 45393
rect 27710 45319 27712 45328
rect 27764 45319 27766 45328
rect 27712 45290 27764 45296
rect 27710 43208 27766 43217
rect 27816 43178 27844 47200
rect 27894 46880 27950 46889
rect 27894 46815 27950 46824
rect 27908 44470 27936 46815
rect 28552 45608 28580 47200
rect 28906 46064 28962 46073
rect 28906 45999 28962 46008
rect 28368 45580 28580 45608
rect 28264 45076 28316 45082
rect 28264 45018 28316 45024
rect 28080 44872 28132 44878
rect 28080 44814 28132 44820
rect 27896 44464 27948 44470
rect 27896 44406 27948 44412
rect 28092 44266 28120 44814
rect 28080 44260 28132 44266
rect 28080 44202 28132 44208
rect 28092 43790 28120 44202
rect 28276 44198 28304 45018
rect 28264 44192 28316 44198
rect 28264 44134 28316 44140
rect 28276 43994 28304 44134
rect 28264 43988 28316 43994
rect 28264 43930 28316 43936
rect 28080 43784 28132 43790
rect 28080 43726 28132 43732
rect 28092 43178 28120 43726
rect 27710 43143 27766 43152
rect 27804 43172 27856 43178
rect 27724 43110 27752 43143
rect 27804 43114 27856 43120
rect 28080 43172 28132 43178
rect 28080 43114 28132 43120
rect 27712 43104 27764 43110
rect 27712 43046 27764 43052
rect 27712 42288 27764 42294
rect 27988 42288 28040 42294
rect 27712 42230 27764 42236
rect 27908 42248 27988 42276
rect 27724 41478 27752 42230
rect 27712 41472 27764 41478
rect 27712 41414 27764 41420
rect 27908 40934 27936 42248
rect 27988 42230 28040 42236
rect 27988 41608 28040 41614
rect 27988 41550 28040 41556
rect 27896 40928 27948 40934
rect 27896 40870 27948 40876
rect 27620 39636 27672 39642
rect 27620 39578 27672 39584
rect 27528 39568 27580 39574
rect 27526 39536 27528 39545
rect 27580 39536 27582 39545
rect 27526 39471 27582 39480
rect 27304 39380 27476 39386
rect 27252 39374 27476 39380
rect 27264 39358 27476 39374
rect 27160 38412 27212 38418
rect 27160 38354 27212 38360
rect 27068 38344 27120 38350
rect 27068 38286 27120 38292
rect 26884 38004 26936 38010
rect 26884 37946 26936 37952
rect 26516 37868 26568 37874
rect 26516 37810 26568 37816
rect 26528 35834 26556 37810
rect 26700 37256 26752 37262
rect 26700 37198 26752 37204
rect 26712 36310 26740 37198
rect 26976 36712 27028 36718
rect 26976 36654 27028 36660
rect 26700 36304 26752 36310
rect 26700 36246 26752 36252
rect 26516 35828 26568 35834
rect 26516 35770 26568 35776
rect 26424 35488 26476 35494
rect 26424 35430 26476 35436
rect 26436 35086 26464 35430
rect 26424 35080 26476 35086
rect 26424 35022 26476 35028
rect 26608 34740 26660 34746
rect 26608 34682 26660 34688
rect 26620 34202 26648 34682
rect 26608 34196 26660 34202
rect 26608 34138 26660 34144
rect 26332 33924 26384 33930
rect 26332 33866 26384 33872
rect 26240 32972 26292 32978
rect 26240 32914 26292 32920
rect 26148 32904 26200 32910
rect 26148 32846 26200 32852
rect 26160 32434 26188 32846
rect 25596 32428 25648 32434
rect 25596 32370 25648 32376
rect 26148 32428 26200 32434
rect 26148 32370 26200 32376
rect 25504 32360 25556 32366
rect 25504 32302 25556 32308
rect 26240 32292 26292 32298
rect 26240 32234 26292 32240
rect 25688 32224 25740 32230
rect 25688 32166 25740 32172
rect 25700 31822 25728 32166
rect 25776 32124 26084 32144
rect 25776 32122 25782 32124
rect 25838 32122 25862 32124
rect 25918 32122 25942 32124
rect 25998 32122 26022 32124
rect 26078 32122 26084 32124
rect 25838 32070 25840 32122
rect 26020 32070 26022 32122
rect 25776 32068 25782 32070
rect 25838 32068 25862 32070
rect 25918 32068 25942 32070
rect 25998 32068 26022 32070
rect 26078 32068 26084 32070
rect 25776 32048 26084 32068
rect 26148 32020 26200 32026
rect 26148 31962 26200 31968
rect 25688 31816 25740 31822
rect 25688 31758 25740 31764
rect 26160 31754 26188 31962
rect 26068 31726 26188 31754
rect 26068 31278 26096 31726
rect 26148 31476 26200 31482
rect 26148 31418 26200 31424
rect 25688 31272 25740 31278
rect 25688 31214 25740 31220
rect 26056 31272 26108 31278
rect 26056 31214 26108 31220
rect 25700 30326 25728 31214
rect 25776 31036 26084 31056
rect 25776 31034 25782 31036
rect 25838 31034 25862 31036
rect 25918 31034 25942 31036
rect 25998 31034 26022 31036
rect 26078 31034 26084 31036
rect 25838 30982 25840 31034
rect 26020 30982 26022 31034
rect 25776 30980 25782 30982
rect 25838 30980 25862 30982
rect 25918 30980 25942 30982
rect 25998 30980 26022 30982
rect 26078 30980 26084 30982
rect 25776 30960 26084 30980
rect 26160 30938 26188 31418
rect 26148 30932 26200 30938
rect 26148 30874 26200 30880
rect 25688 30320 25740 30326
rect 25688 30262 25740 30268
rect 26160 30258 26188 30874
rect 26148 30252 26200 30258
rect 26148 30194 26200 30200
rect 25776 29948 26084 29968
rect 25776 29946 25782 29948
rect 25838 29946 25862 29948
rect 25918 29946 25942 29948
rect 25998 29946 26022 29948
rect 26078 29946 26084 29948
rect 25838 29894 25840 29946
rect 26020 29894 26022 29946
rect 25776 29892 25782 29894
rect 25838 29892 25862 29894
rect 25918 29892 25942 29894
rect 25998 29892 26022 29894
rect 26078 29892 26084 29894
rect 25776 29872 26084 29892
rect 25504 29572 25556 29578
rect 25504 29514 25556 29520
rect 25516 29306 25544 29514
rect 25504 29300 25556 29306
rect 25504 29242 25556 29248
rect 25776 28860 26084 28880
rect 25776 28858 25782 28860
rect 25838 28858 25862 28860
rect 25918 28858 25942 28860
rect 25998 28858 26022 28860
rect 26078 28858 26084 28860
rect 25838 28806 25840 28858
rect 26020 28806 26022 28858
rect 25776 28804 25782 28806
rect 25838 28804 25862 28806
rect 25918 28804 25942 28806
rect 25998 28804 26022 28806
rect 26078 28804 26084 28806
rect 25776 28784 26084 28804
rect 25776 27772 26084 27792
rect 25776 27770 25782 27772
rect 25838 27770 25862 27772
rect 25918 27770 25942 27772
rect 25998 27770 26022 27772
rect 26078 27770 26084 27772
rect 25838 27718 25840 27770
rect 26020 27718 26022 27770
rect 25776 27716 25782 27718
rect 25838 27716 25862 27718
rect 25918 27716 25942 27718
rect 25998 27716 26022 27718
rect 26078 27716 26084 27718
rect 25776 27696 26084 27716
rect 25688 27464 25740 27470
rect 25688 27406 25740 27412
rect 25320 27396 25372 27402
rect 25320 27338 25372 27344
rect 25228 26376 25280 26382
rect 25228 26318 25280 26324
rect 25332 25906 25360 27338
rect 25412 26920 25464 26926
rect 25412 26862 25464 26868
rect 25504 26920 25556 26926
rect 25504 26862 25556 26868
rect 25320 25900 25372 25906
rect 25320 25842 25372 25848
rect 25044 25764 25096 25770
rect 25044 25706 25096 25712
rect 25136 25424 25188 25430
rect 25136 25366 25188 25372
rect 24676 25356 24728 25362
rect 24676 25298 24728 25304
rect 24688 24970 24716 25298
rect 24688 24942 24900 24970
rect 24676 24812 24728 24818
rect 24676 24754 24728 24760
rect 24688 24410 24716 24754
rect 24872 24750 24900 24942
rect 24860 24744 24912 24750
rect 24860 24686 24912 24692
rect 25044 24608 25096 24614
rect 25044 24550 25096 24556
rect 24676 24404 24728 24410
rect 24676 24346 24728 24352
rect 24584 24200 24636 24206
rect 25056 24188 25084 24550
rect 25148 24342 25176 25366
rect 25332 25294 25360 25842
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25228 24948 25280 24954
rect 25228 24890 25280 24896
rect 25136 24336 25188 24342
rect 25136 24278 25188 24284
rect 25136 24200 25188 24206
rect 25056 24160 25136 24188
rect 24584 24142 24636 24148
rect 25136 24142 25188 24148
rect 24492 23860 24544 23866
rect 24492 23802 24544 23808
rect 24860 23724 24912 23730
rect 24860 23666 24912 23672
rect 24872 23322 24900 23666
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24492 23180 24544 23186
rect 24492 23122 24544 23128
rect 24400 21140 24452 21146
rect 24400 21082 24452 21088
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24412 19666 24440 20878
rect 24504 19854 24532 23122
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 24676 22976 24728 22982
rect 24676 22918 24728 22924
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24596 21146 24624 22578
rect 24584 21140 24636 21146
rect 24584 21082 24636 21088
rect 24688 20466 24716 22918
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24780 21486 24808 22646
rect 24860 22568 24912 22574
rect 24860 22510 24912 22516
rect 24768 21480 24820 21486
rect 24768 21422 24820 21428
rect 24780 21321 24808 21422
rect 24766 21312 24822 21321
rect 24766 21247 24822 21256
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24780 20602 24808 21082
rect 24872 21010 24900 22510
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24964 20942 24992 21626
rect 24952 20936 25004 20942
rect 24952 20878 25004 20884
rect 25056 20618 25084 23054
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 25148 20942 25176 22714
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 24964 20590 25084 20618
rect 24780 20466 24808 20538
rect 24676 20460 24728 20466
rect 24676 20402 24728 20408
rect 24768 20460 24820 20466
rect 24768 20402 24820 20408
rect 24584 20392 24636 20398
rect 24584 20334 24636 20340
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24412 19638 24532 19666
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24308 16652 24360 16658
rect 24308 16594 24360 16600
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24228 14074 24256 14962
rect 24216 14068 24268 14074
rect 24216 14010 24268 14016
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 24228 12238 24256 12854
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 23940 11212 23992 11218
rect 23940 11154 23992 11160
rect 23952 9926 23980 11154
rect 24228 10606 24256 12174
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23952 9586 23980 9862
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 23952 8498 23980 9522
rect 24044 9178 24072 9522
rect 24228 9382 24256 10542
rect 24216 9376 24268 9382
rect 24216 9318 24268 9324
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 24124 8900 24176 8906
rect 24124 8842 24176 8848
rect 24136 8634 24164 8842
rect 24216 8832 24268 8838
rect 24216 8774 24268 8780
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24228 8566 24256 8774
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23952 8022 23980 8434
rect 24320 8090 24348 16594
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24412 13326 24440 15438
rect 24504 14006 24532 19638
rect 24492 14000 24544 14006
rect 24492 13942 24544 13948
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24412 12918 24440 13262
rect 24400 12912 24452 12918
rect 24400 12854 24452 12860
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 24400 12368 24452 12374
rect 24400 12310 24452 12316
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 23940 8016 23992 8022
rect 23940 7958 23992 7964
rect 23952 6322 23980 7958
rect 24308 7880 24360 7886
rect 24308 7822 24360 7828
rect 24320 7546 24348 7822
rect 24308 7540 24360 7546
rect 24308 7482 24360 7488
rect 24412 7478 24440 12310
rect 24504 12170 24532 12786
rect 24492 12164 24544 12170
rect 24492 12106 24544 12112
rect 24596 10538 24624 20334
rect 24766 19816 24822 19825
rect 24766 19751 24768 19760
rect 24820 19751 24822 19760
rect 24768 19722 24820 19728
rect 24964 19514 24992 20590
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 24674 19408 24730 19417
rect 24674 19343 24730 19352
rect 24688 13938 24716 19343
rect 24860 18760 24912 18766
rect 24858 18728 24860 18737
rect 24912 18728 24914 18737
rect 24858 18663 24914 18672
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24766 18320 24822 18329
rect 24766 18255 24822 18264
rect 24780 15722 24808 18255
rect 24872 18086 24900 18566
rect 24964 18290 24992 19450
rect 25056 18970 25084 20402
rect 25044 18964 25096 18970
rect 25044 18906 25096 18912
rect 25148 18850 25176 20742
rect 25240 20602 25268 24890
rect 25332 24886 25360 25230
rect 25320 24880 25372 24886
rect 25320 24822 25372 24828
rect 25318 24304 25374 24313
rect 25318 24239 25320 24248
rect 25372 24239 25374 24248
rect 25320 24210 25372 24216
rect 25320 23520 25372 23526
rect 25320 23462 25372 23468
rect 25332 21962 25360 23462
rect 25424 23322 25452 26862
rect 25516 26450 25544 26862
rect 25700 26790 25728 27406
rect 26252 26994 26280 32234
rect 26344 31890 26372 33866
rect 26620 33522 26648 34138
rect 26608 33516 26660 33522
rect 26608 33458 26660 33464
rect 26516 32972 26568 32978
rect 26516 32914 26568 32920
rect 26424 32428 26476 32434
rect 26424 32370 26476 32376
rect 26332 31884 26384 31890
rect 26332 31826 26384 31832
rect 26436 31822 26464 32370
rect 26424 31816 26476 31822
rect 26424 31758 26476 31764
rect 26436 30258 26464 31758
rect 26528 31754 26556 32914
rect 26516 31748 26568 31754
rect 26516 31690 26568 31696
rect 26528 30666 26556 31690
rect 26712 31414 26740 36246
rect 26988 35290 27016 36654
rect 26976 35284 27028 35290
rect 26976 35226 27028 35232
rect 26976 34604 27028 34610
rect 26976 34546 27028 34552
rect 26884 34060 26936 34066
rect 26884 34002 26936 34008
rect 26896 33454 26924 34002
rect 26884 33448 26936 33454
rect 26884 33390 26936 33396
rect 26896 32502 26924 33390
rect 26988 33114 27016 34546
rect 27160 34400 27212 34406
rect 27160 34342 27212 34348
rect 27068 33992 27120 33998
rect 27068 33934 27120 33940
rect 26976 33108 27028 33114
rect 26976 33050 27028 33056
rect 26884 32496 26936 32502
rect 26884 32438 26936 32444
rect 27080 32434 27108 33934
rect 27172 32978 27200 34342
rect 27264 33561 27292 39358
rect 27804 39296 27856 39302
rect 27804 39238 27856 39244
rect 27816 39030 27844 39238
rect 27804 39024 27856 39030
rect 27804 38966 27856 38972
rect 27896 37868 27948 37874
rect 27896 37810 27948 37816
rect 27344 37256 27396 37262
rect 27342 37224 27344 37233
rect 27804 37256 27856 37262
rect 27396 37224 27398 37233
rect 27804 37198 27856 37204
rect 27342 37159 27398 37168
rect 27344 37120 27396 37126
rect 27344 37062 27396 37068
rect 27356 36106 27384 37062
rect 27344 36100 27396 36106
rect 27344 36042 27396 36048
rect 27712 36032 27764 36038
rect 27712 35974 27764 35980
rect 27724 35698 27752 35974
rect 27816 35834 27844 37198
rect 27908 35834 27936 37810
rect 28000 37398 28028 41550
rect 27988 37392 28040 37398
rect 27988 37334 28040 37340
rect 27988 37120 28040 37126
rect 27988 37062 28040 37068
rect 28000 36174 28028 37062
rect 27988 36168 28040 36174
rect 27988 36110 28040 36116
rect 27804 35828 27856 35834
rect 27804 35770 27856 35776
rect 27896 35828 27948 35834
rect 27896 35770 27948 35776
rect 27712 35692 27764 35698
rect 27712 35634 27764 35640
rect 27988 34944 28040 34950
rect 27988 34886 28040 34892
rect 28000 33998 28028 34886
rect 27988 33992 28040 33998
rect 27988 33934 28040 33940
rect 27436 33924 27488 33930
rect 27436 33866 27488 33872
rect 27448 33658 27476 33866
rect 27620 33856 27672 33862
rect 27620 33798 27672 33804
rect 27436 33652 27488 33658
rect 27436 33594 27488 33600
rect 27250 33552 27306 33561
rect 27250 33487 27306 33496
rect 27160 32972 27212 32978
rect 27160 32914 27212 32920
rect 27264 32858 27292 33487
rect 27172 32830 27292 32858
rect 27172 32434 27200 32830
rect 27252 32496 27304 32502
rect 27252 32438 27304 32444
rect 27068 32428 27120 32434
rect 27068 32370 27120 32376
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 26884 32292 26936 32298
rect 26884 32234 26936 32240
rect 26792 32224 26844 32230
rect 26792 32166 26844 32172
rect 26804 31958 26832 32166
rect 26896 32026 26924 32234
rect 27160 32224 27212 32230
rect 27160 32166 27212 32172
rect 26884 32020 26936 32026
rect 26884 31962 26936 31968
rect 26792 31952 26844 31958
rect 26792 31894 26844 31900
rect 26896 31890 26924 31962
rect 26884 31884 26936 31890
rect 26884 31826 26936 31832
rect 26792 31816 26844 31822
rect 26792 31758 26844 31764
rect 26700 31408 26752 31414
rect 26700 31350 26752 31356
rect 26516 30660 26568 30666
rect 26516 30602 26568 30608
rect 26424 30252 26476 30258
rect 26424 30194 26476 30200
rect 26436 30122 26464 30194
rect 26804 30190 26832 31758
rect 27068 31408 27120 31414
rect 27068 31350 27120 31356
rect 27080 30258 27108 31350
rect 27172 31346 27200 32166
rect 27264 31822 27292 32438
rect 27448 32366 27476 33594
rect 27632 32842 27660 33798
rect 27712 33652 27764 33658
rect 27712 33594 27764 33600
rect 27620 32836 27672 32842
rect 27620 32778 27672 32784
rect 27724 32502 27752 33594
rect 27804 33516 27856 33522
rect 27804 33458 27856 33464
rect 27816 32570 27844 33458
rect 27804 32564 27856 32570
rect 27804 32506 27856 32512
rect 27712 32496 27764 32502
rect 27712 32438 27764 32444
rect 27436 32360 27488 32366
rect 27436 32302 27488 32308
rect 27252 31816 27304 31822
rect 27252 31758 27304 31764
rect 27436 31680 27488 31686
rect 27436 31622 27488 31628
rect 27448 31414 27476 31622
rect 27436 31408 27488 31414
rect 27436 31350 27488 31356
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 27712 30660 27764 30666
rect 27712 30602 27764 30608
rect 27724 30326 27752 30602
rect 27712 30320 27764 30326
rect 27712 30262 27764 30268
rect 27068 30252 27120 30258
rect 27068 30194 27120 30200
rect 26792 30184 26844 30190
rect 26792 30126 26844 30132
rect 26424 30116 26476 30122
rect 26424 30058 26476 30064
rect 28092 30054 28120 43114
rect 28276 43110 28304 43930
rect 28264 43104 28316 43110
rect 28264 43046 28316 43052
rect 28276 42022 28304 43046
rect 28264 42016 28316 42022
rect 28264 41958 28316 41964
rect 28368 41721 28396 45580
rect 28446 45520 28502 45529
rect 28446 45455 28502 45464
rect 28540 45484 28592 45490
rect 28460 44538 28488 45455
rect 28540 45426 28592 45432
rect 28552 44538 28580 45426
rect 28448 44532 28500 44538
rect 28448 44474 28500 44480
rect 28540 44532 28592 44538
rect 28540 44474 28592 44480
rect 28920 43450 28948 45999
rect 29184 45484 29236 45490
rect 29184 45426 29236 45432
rect 29000 44260 29052 44266
rect 29000 44202 29052 44208
rect 29012 43790 29040 44202
rect 29092 43852 29144 43858
rect 29092 43794 29144 43800
rect 29000 43784 29052 43790
rect 29000 43726 29052 43732
rect 28908 43444 28960 43450
rect 28908 43386 28960 43392
rect 28448 42696 28500 42702
rect 28448 42638 28500 42644
rect 28908 42696 28960 42702
rect 28908 42638 28960 42644
rect 28354 41712 28410 41721
rect 28354 41647 28410 41656
rect 28356 41200 28408 41206
rect 28170 41168 28226 41177
rect 28356 41142 28408 41148
rect 28170 41103 28226 41112
rect 28184 41002 28212 41103
rect 28264 41064 28316 41070
rect 28264 41006 28316 41012
rect 28172 40996 28224 41002
rect 28172 40938 28224 40944
rect 28276 40225 28304 41006
rect 28368 40934 28396 41142
rect 28356 40928 28408 40934
rect 28356 40870 28408 40876
rect 28262 40216 28318 40225
rect 28262 40151 28318 40160
rect 28368 40089 28396 40870
rect 28460 40202 28488 42638
rect 28632 42560 28684 42566
rect 28632 42502 28684 42508
rect 28540 42220 28592 42226
rect 28540 42162 28592 42168
rect 28552 41750 28580 42162
rect 28644 42022 28672 42502
rect 28632 42016 28684 42022
rect 28632 41958 28684 41964
rect 28644 41818 28672 41958
rect 28632 41812 28684 41818
rect 28632 41754 28684 41760
rect 28816 41812 28868 41818
rect 28816 41754 28868 41760
rect 28540 41744 28592 41750
rect 28540 41686 28592 41692
rect 28552 41138 28580 41686
rect 28724 41472 28776 41478
rect 28724 41414 28776 41420
rect 28540 41132 28592 41138
rect 28540 41074 28592 41080
rect 28552 40662 28580 41074
rect 28540 40656 28592 40662
rect 28540 40598 28592 40604
rect 28632 40384 28684 40390
rect 28632 40326 28684 40332
rect 28460 40174 28580 40202
rect 28354 40080 28410 40089
rect 28354 40015 28410 40024
rect 28448 40044 28500 40050
rect 28448 39986 28500 39992
rect 28172 39840 28224 39846
rect 28172 39782 28224 39788
rect 28184 36174 28212 39782
rect 28356 39364 28408 39370
rect 28356 39306 28408 39312
rect 28368 38962 28396 39306
rect 28356 38956 28408 38962
rect 28356 38898 28408 38904
rect 28368 38554 28396 38898
rect 28356 38548 28408 38554
rect 28356 38490 28408 38496
rect 28264 37936 28316 37942
rect 28264 37878 28316 37884
rect 28276 37466 28304 37878
rect 28264 37460 28316 37466
rect 28264 37402 28316 37408
rect 28276 36378 28304 37402
rect 28460 36854 28488 39986
rect 28552 39574 28580 40174
rect 28540 39568 28592 39574
rect 28540 39510 28592 39516
rect 28540 39432 28592 39438
rect 28540 39374 28592 39380
rect 28552 39098 28580 39374
rect 28540 39092 28592 39098
rect 28540 39034 28592 39040
rect 28644 38350 28672 40326
rect 28736 39438 28764 41414
rect 28828 40730 28856 41754
rect 28816 40724 28868 40730
rect 28816 40666 28868 40672
rect 28920 40610 28948 42638
rect 29104 41818 29132 43794
rect 29196 42537 29224 45426
rect 29182 42528 29238 42537
rect 29182 42463 29238 42472
rect 29092 41812 29144 41818
rect 29092 41754 29144 41760
rect 29288 41414 29316 47200
rect 30024 45626 30052 47495
rect 30102 47200 30158 48000
rect 30838 47200 30894 48000
rect 31574 47200 31630 48000
rect 30012 45620 30064 45626
rect 30012 45562 30064 45568
rect 30012 44736 30064 44742
rect 30012 44678 30064 44684
rect 30024 44577 30052 44678
rect 30010 44568 30066 44577
rect 30010 44503 30066 44512
rect 29552 44396 29604 44402
rect 29552 44338 29604 44344
rect 29920 44396 29972 44402
rect 29920 44338 29972 44344
rect 29288 41386 29500 41414
rect 29184 40928 29236 40934
rect 29184 40870 29236 40876
rect 29196 40730 29224 40870
rect 29184 40724 29236 40730
rect 29184 40666 29236 40672
rect 28828 40582 28948 40610
rect 28828 40050 28856 40582
rect 28908 40520 28960 40526
rect 28908 40462 28960 40468
rect 29092 40520 29144 40526
rect 29092 40462 29144 40468
rect 28816 40044 28868 40050
rect 28816 39986 28868 39992
rect 28724 39432 28776 39438
rect 28724 39374 28776 39380
rect 28828 39284 28856 39986
rect 28920 39386 28948 40462
rect 29104 40118 29132 40462
rect 29092 40112 29144 40118
rect 29092 40054 29144 40060
rect 29196 39642 29224 40666
rect 29472 40186 29500 41386
rect 29564 41070 29592 44338
rect 29644 44192 29696 44198
rect 29644 44134 29696 44140
rect 29552 41064 29604 41070
rect 29552 41006 29604 41012
rect 29460 40180 29512 40186
rect 29460 40122 29512 40128
rect 29656 39982 29684 44134
rect 29736 42628 29788 42634
rect 29736 42570 29788 42576
rect 29748 41138 29776 42570
rect 29736 41132 29788 41138
rect 29736 41074 29788 41080
rect 29932 40497 29960 44338
rect 30116 44033 30144 47200
rect 30102 44024 30158 44033
rect 30852 43994 30880 47200
rect 31588 44130 31616 47200
rect 31576 44124 31628 44130
rect 31576 44066 31628 44072
rect 30102 43959 30158 43968
rect 30840 43988 30892 43994
rect 30840 43930 30892 43936
rect 30012 43920 30064 43926
rect 30010 43888 30012 43897
rect 30064 43888 30066 43897
rect 30010 43823 30066 43832
rect 30012 43104 30064 43110
rect 30010 43072 30012 43081
rect 30064 43072 30066 43081
rect 30010 43007 30066 43016
rect 30012 42560 30064 42566
rect 30012 42502 30064 42508
rect 30024 42401 30052 42502
rect 30010 42392 30066 42401
rect 30010 42327 30066 42336
rect 30012 42016 30064 42022
rect 30012 41958 30064 41964
rect 30024 41721 30052 41958
rect 30010 41712 30066 41721
rect 30010 41647 30066 41656
rect 30012 41472 30064 41478
rect 30012 41414 30064 41420
rect 30024 40905 30052 41414
rect 30104 40928 30156 40934
rect 30010 40896 30066 40905
rect 30104 40870 30156 40876
rect 30010 40831 30066 40840
rect 29918 40488 29974 40497
rect 29918 40423 29974 40432
rect 30012 40384 30064 40390
rect 30012 40326 30064 40332
rect 29644 39976 29696 39982
rect 29644 39918 29696 39924
rect 29368 39840 29420 39846
rect 29368 39782 29420 39788
rect 29184 39636 29236 39642
rect 29184 39578 29236 39584
rect 29092 39432 29144 39438
rect 28920 39358 29040 39386
rect 29092 39374 29144 39380
rect 28736 39256 28856 39284
rect 28908 39296 28960 39302
rect 28632 38344 28684 38350
rect 28632 38286 28684 38292
rect 28736 38196 28764 39256
rect 28908 39238 28960 39244
rect 28920 38729 28948 39238
rect 28906 38720 28962 38729
rect 28906 38655 28962 38664
rect 29012 38570 29040 39358
rect 29104 38826 29132 39374
rect 29092 38820 29144 38826
rect 29092 38762 29144 38768
rect 28644 38168 28764 38196
rect 28920 38542 29040 38570
rect 28540 37868 28592 37874
rect 28540 37810 28592 37816
rect 28448 36848 28500 36854
rect 28448 36790 28500 36796
rect 28264 36372 28316 36378
rect 28264 36314 28316 36320
rect 28172 36168 28224 36174
rect 28172 36110 28224 36116
rect 28552 35290 28580 37810
rect 28644 35698 28672 38168
rect 28724 37664 28776 37670
rect 28724 37606 28776 37612
rect 28632 35692 28684 35698
rect 28632 35634 28684 35640
rect 28356 35284 28408 35290
rect 28356 35226 28408 35232
rect 28540 35284 28592 35290
rect 28540 35226 28592 35232
rect 28264 35080 28316 35086
rect 28264 35022 28316 35028
rect 28172 34604 28224 34610
rect 28172 34546 28224 34552
rect 28184 32570 28212 34546
rect 28276 33114 28304 35022
rect 28368 34610 28396 35226
rect 28736 35086 28764 37606
rect 28920 37126 28948 38542
rect 29104 37806 29132 38762
rect 29380 38758 29408 39782
rect 30024 39409 30052 40326
rect 30116 40225 30144 40870
rect 30102 40216 30158 40225
rect 30102 40151 30158 40160
rect 30104 39840 30156 39846
rect 30104 39782 30156 39788
rect 30010 39400 30066 39409
rect 30010 39335 30066 39344
rect 29368 38752 29420 38758
rect 29368 38694 29420 38700
rect 29092 37800 29144 37806
rect 29092 37742 29144 37748
rect 29104 37330 29132 37742
rect 29380 37670 29408 38694
rect 30012 38208 30064 38214
rect 30012 38150 30064 38156
rect 29276 37664 29328 37670
rect 29276 37606 29328 37612
rect 29368 37664 29420 37670
rect 29368 37606 29420 37612
rect 29092 37324 29144 37330
rect 29092 37266 29144 37272
rect 28816 37120 28868 37126
rect 28816 37062 28868 37068
rect 28908 37120 28960 37126
rect 28908 37062 28960 37068
rect 28828 36922 28856 37062
rect 28816 36916 28868 36922
rect 28816 36858 28868 36864
rect 29092 36644 29144 36650
rect 29092 36586 29144 36592
rect 28906 36544 28962 36553
rect 28906 36479 28962 36488
rect 28920 36378 28948 36479
rect 28908 36372 28960 36378
rect 28908 36314 28960 36320
rect 29104 35698 29132 36586
rect 29288 36174 29316 37606
rect 29380 37466 29408 37606
rect 29368 37460 29420 37466
rect 29368 37402 29420 37408
rect 29380 36582 29408 37402
rect 30024 37233 30052 38150
rect 30116 37913 30144 39782
rect 30102 37904 30158 37913
rect 30102 37839 30158 37848
rect 30010 37224 30066 37233
rect 30010 37159 30066 37168
rect 29368 36576 29420 36582
rect 29368 36518 29420 36524
rect 29276 36168 29328 36174
rect 29276 36110 29328 36116
rect 30012 36032 30064 36038
rect 30012 35974 30064 35980
rect 30024 35737 30052 35974
rect 30010 35728 30066 35737
rect 29092 35692 29144 35698
rect 30010 35663 30066 35672
rect 29092 35634 29144 35640
rect 29104 35222 29132 35634
rect 29920 35488 29972 35494
rect 29920 35430 29972 35436
rect 29932 35290 29960 35430
rect 29920 35284 29972 35290
rect 29920 35226 29972 35232
rect 29092 35216 29144 35222
rect 29092 35158 29144 35164
rect 28724 35080 28776 35086
rect 28724 35022 28776 35028
rect 28906 35048 28962 35057
rect 28906 34983 28962 34992
rect 28920 34950 28948 34983
rect 28908 34944 28960 34950
rect 28908 34886 28960 34892
rect 29000 34944 29052 34950
rect 29000 34886 29052 34892
rect 29012 34746 29040 34886
rect 28448 34740 28500 34746
rect 28448 34682 28500 34688
rect 29000 34740 29052 34746
rect 29000 34682 29052 34688
rect 28356 34604 28408 34610
rect 28356 34546 28408 34552
rect 28460 34241 28488 34682
rect 28724 34672 28776 34678
rect 28724 34614 28776 34620
rect 28446 34232 28502 34241
rect 28446 34167 28502 34176
rect 28632 33924 28684 33930
rect 28632 33866 28684 33872
rect 28644 33658 28672 33866
rect 28736 33862 28764 34614
rect 29104 34610 29132 35158
rect 29460 35012 29512 35018
rect 29460 34954 29512 34960
rect 29472 34746 29500 34954
rect 29460 34740 29512 34746
rect 29460 34682 29512 34688
rect 29092 34604 29144 34610
rect 29092 34546 29144 34552
rect 29104 34134 29132 34546
rect 29828 34536 29880 34542
rect 29828 34478 29880 34484
rect 29276 34400 29328 34406
rect 29276 34342 29328 34348
rect 29288 34202 29316 34342
rect 29276 34196 29328 34202
rect 29276 34138 29328 34144
rect 29092 34128 29144 34134
rect 29092 34070 29144 34076
rect 28724 33856 28776 33862
rect 28724 33798 28776 33804
rect 28908 33856 28960 33862
rect 28908 33798 28960 33804
rect 28632 33652 28684 33658
rect 28632 33594 28684 33600
rect 28264 33108 28316 33114
rect 28264 33050 28316 33056
rect 28448 33108 28500 33114
rect 28448 33050 28500 33056
rect 28264 32904 28316 32910
rect 28264 32846 28316 32852
rect 28172 32564 28224 32570
rect 28172 32506 28224 32512
rect 28276 32026 28304 32846
rect 28460 32434 28488 33050
rect 28644 32502 28672 33594
rect 28736 33114 28764 33798
rect 28920 33561 28948 33798
rect 28906 33552 28962 33561
rect 28906 33487 28962 33496
rect 28724 33108 28776 33114
rect 28724 33050 28776 33056
rect 28632 32496 28684 32502
rect 28632 32438 28684 32444
rect 28724 32496 28776 32502
rect 28724 32438 28776 32444
rect 28448 32428 28500 32434
rect 28448 32370 28500 32376
rect 28264 32020 28316 32026
rect 28264 31962 28316 31968
rect 28736 31958 28764 32438
rect 29184 32428 29236 32434
rect 29184 32370 29236 32376
rect 28908 32292 28960 32298
rect 28908 32234 28960 32240
rect 28724 31952 28776 31958
rect 28724 31894 28776 31900
rect 28736 31482 28764 31894
rect 28724 31476 28776 31482
rect 28724 31418 28776 31424
rect 28920 31210 28948 32234
rect 29000 31816 29052 31822
rect 29000 31758 29052 31764
rect 29012 31482 29040 31758
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 28632 31204 28684 31210
rect 28632 31146 28684 31152
rect 28908 31204 28960 31210
rect 28908 31146 28960 31152
rect 28644 30734 28672 31146
rect 29092 31136 29144 31142
rect 29092 31078 29144 31084
rect 28356 30728 28408 30734
rect 28356 30670 28408 30676
rect 28632 30728 28684 30734
rect 28632 30670 28684 30676
rect 28172 30592 28224 30598
rect 28172 30534 28224 30540
rect 28184 30258 28212 30534
rect 28368 30394 28396 30670
rect 28448 30592 28500 30598
rect 28448 30534 28500 30540
rect 28356 30388 28408 30394
rect 28356 30330 28408 30336
rect 28460 30326 28488 30534
rect 28448 30320 28500 30326
rect 28448 30262 28500 30268
rect 28172 30252 28224 30258
rect 28172 30194 28224 30200
rect 28080 30048 28132 30054
rect 28080 29990 28132 29996
rect 27344 29844 27396 29850
rect 27344 29786 27396 29792
rect 27160 29640 27212 29646
rect 27160 29582 27212 29588
rect 26424 29504 26476 29510
rect 26424 29446 26476 29452
rect 26436 28490 26464 29446
rect 27172 29306 27200 29582
rect 27356 29578 27384 29786
rect 28644 29646 28672 30670
rect 29000 30252 29052 30258
rect 29000 30194 29052 30200
rect 29012 29850 29040 30194
rect 29000 29844 29052 29850
rect 29000 29786 29052 29792
rect 29104 29782 29132 31078
rect 29092 29776 29144 29782
rect 29092 29718 29144 29724
rect 28632 29640 28684 29646
rect 28632 29582 28684 29588
rect 27344 29572 27396 29578
rect 27344 29514 27396 29520
rect 27160 29300 27212 29306
rect 27160 29242 27212 29248
rect 27068 29164 27120 29170
rect 27068 29106 27120 29112
rect 26516 29028 26568 29034
rect 26516 28970 26568 28976
rect 26528 28558 26556 28970
rect 26516 28552 26568 28558
rect 26516 28494 26568 28500
rect 26424 28484 26476 28490
rect 26424 28426 26476 28432
rect 27080 28218 27108 29106
rect 27356 28762 27384 29514
rect 27436 29504 27488 29510
rect 27436 29446 27488 29452
rect 27448 29306 27476 29446
rect 27436 29300 27488 29306
rect 27436 29242 27488 29248
rect 27448 29102 27476 29242
rect 28644 29170 28672 29582
rect 28632 29164 28684 29170
rect 28632 29106 28684 29112
rect 27436 29096 27488 29102
rect 27436 29038 27488 29044
rect 27528 29096 27580 29102
rect 27528 29038 27580 29044
rect 27344 28756 27396 28762
rect 27344 28698 27396 28704
rect 27068 28212 27120 28218
rect 27068 28154 27120 28160
rect 27540 27606 27568 29038
rect 29104 28966 29132 29718
rect 29196 29306 29224 32370
rect 29288 32230 29316 34138
rect 29840 33522 29868 34478
rect 29932 34202 29960 35226
rect 30104 35148 30156 35154
rect 30104 35090 30156 35096
rect 30116 34202 30144 35090
rect 29920 34196 29972 34202
rect 29920 34138 29972 34144
rect 30104 34196 30156 34202
rect 30104 34138 30156 34144
rect 29828 33516 29880 33522
rect 29828 33458 29880 33464
rect 30012 33312 30064 33318
rect 30012 33254 30064 33260
rect 30024 32745 30052 33254
rect 30104 32768 30156 32774
rect 30010 32736 30066 32745
rect 30104 32710 30156 32716
rect 30010 32671 30066 32680
rect 29276 32224 29328 32230
rect 29276 32166 29328 32172
rect 29828 32224 29880 32230
rect 29828 32166 29880 32172
rect 29840 29646 29868 32166
rect 30116 32065 30144 32710
rect 30102 32056 30158 32065
rect 30102 31991 30158 32000
rect 30104 31748 30156 31754
rect 30104 31690 30156 31696
rect 30012 31680 30064 31686
rect 30012 31622 30064 31628
rect 30024 31385 30052 31622
rect 30010 31376 30066 31385
rect 30010 31311 30066 31320
rect 29920 31136 29972 31142
rect 29920 31078 29972 31084
rect 29932 30938 29960 31078
rect 30116 30938 30144 31690
rect 29920 30932 29972 30938
rect 29920 30874 29972 30880
rect 30104 30932 30156 30938
rect 30104 30874 30156 30880
rect 30102 30560 30158 30569
rect 30102 30495 30158 30504
rect 30012 30048 30064 30054
rect 30012 29990 30064 29996
rect 30024 29889 30052 29990
rect 30010 29880 30066 29889
rect 30116 29850 30144 30495
rect 30010 29815 30066 29824
rect 30104 29844 30156 29850
rect 30104 29786 30156 29792
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29184 29300 29236 29306
rect 29184 29242 29236 29248
rect 30010 29064 30066 29073
rect 30010 28999 30012 29008
rect 30064 28999 30066 29008
rect 30012 28970 30064 28976
rect 29092 28960 29144 28966
rect 29092 28902 29144 28908
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 27528 27600 27580 27606
rect 27528 27542 27580 27548
rect 29840 27538 29868 28494
rect 30012 28416 30064 28422
rect 30010 28384 30012 28393
rect 30064 28384 30066 28393
rect 30010 28319 30066 28328
rect 30012 27872 30064 27878
rect 30012 27814 30064 27820
rect 30024 27577 30052 27814
rect 30010 27568 30066 27577
rect 29828 27532 29880 27538
rect 30010 27503 30066 27512
rect 29828 27474 29880 27480
rect 26332 27464 26384 27470
rect 26332 27406 26384 27412
rect 26240 26988 26292 26994
rect 26240 26930 26292 26936
rect 25688 26784 25740 26790
rect 25688 26726 25740 26732
rect 25776 26684 26084 26704
rect 25776 26682 25782 26684
rect 25838 26682 25862 26684
rect 25918 26682 25942 26684
rect 25998 26682 26022 26684
rect 26078 26682 26084 26684
rect 25838 26630 25840 26682
rect 26020 26630 26022 26682
rect 25776 26628 25782 26630
rect 25838 26628 25862 26630
rect 25918 26628 25942 26630
rect 25998 26628 26022 26630
rect 26078 26628 26084 26630
rect 25776 26608 26084 26628
rect 26344 26586 26372 27406
rect 30010 26888 30066 26897
rect 30010 26823 30012 26832
rect 30064 26823 30066 26832
rect 30012 26794 30064 26800
rect 26332 26580 26384 26586
rect 26332 26522 26384 26528
rect 25504 26444 25556 26450
rect 25504 26386 25556 26392
rect 26792 26376 26844 26382
rect 26792 26318 26844 26324
rect 29828 26376 29880 26382
rect 29828 26318 29880 26324
rect 26700 25968 26752 25974
rect 26700 25910 26752 25916
rect 26332 25832 26384 25838
rect 26332 25774 26384 25780
rect 25776 25596 26084 25616
rect 25776 25594 25782 25596
rect 25838 25594 25862 25596
rect 25918 25594 25942 25596
rect 25998 25594 26022 25596
rect 26078 25594 26084 25596
rect 25838 25542 25840 25594
rect 26020 25542 26022 25594
rect 25776 25540 25782 25542
rect 25838 25540 25862 25542
rect 25918 25540 25942 25542
rect 25998 25540 26022 25542
rect 26078 25540 26084 25542
rect 25776 25520 26084 25540
rect 25688 25220 25740 25226
rect 25688 25162 25740 25168
rect 26240 25220 26292 25226
rect 26240 25162 26292 25168
rect 25596 24200 25648 24206
rect 25596 24142 25648 24148
rect 25608 23526 25636 24142
rect 25700 23633 25728 25162
rect 25964 25152 26016 25158
rect 25964 25094 26016 25100
rect 25976 24750 26004 25094
rect 25964 24744 26016 24750
rect 25964 24686 26016 24692
rect 25776 24508 26084 24528
rect 25776 24506 25782 24508
rect 25838 24506 25862 24508
rect 25918 24506 25942 24508
rect 25998 24506 26022 24508
rect 26078 24506 26084 24508
rect 25838 24454 25840 24506
rect 26020 24454 26022 24506
rect 25776 24452 25782 24454
rect 25838 24452 25862 24454
rect 25918 24452 25942 24454
rect 25998 24452 26022 24454
rect 26078 24452 26084 24454
rect 25776 24432 26084 24452
rect 26252 24410 26280 25162
rect 26240 24404 26292 24410
rect 26240 24346 26292 24352
rect 25780 24064 25832 24070
rect 25780 24006 25832 24012
rect 25792 23730 25820 24006
rect 26344 23866 26372 25774
rect 26608 24404 26660 24410
rect 26608 24346 26660 24352
rect 26620 24206 26648 24346
rect 26608 24200 26660 24206
rect 26608 24142 26660 24148
rect 26332 23860 26384 23866
rect 26332 23802 26384 23808
rect 25780 23724 25832 23730
rect 25780 23666 25832 23672
rect 25686 23624 25742 23633
rect 25686 23559 25742 23568
rect 25596 23520 25648 23526
rect 25596 23462 25648 23468
rect 25412 23316 25464 23322
rect 25412 23258 25464 23264
rect 25608 23254 25636 23462
rect 25596 23248 25648 23254
rect 25596 23190 25648 23196
rect 25504 23112 25556 23118
rect 25504 23054 25556 23060
rect 25516 22234 25544 23054
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25504 22228 25556 22234
rect 25504 22170 25556 22176
rect 25608 22166 25636 22510
rect 25700 22216 25728 23559
rect 25776 23420 26084 23440
rect 25776 23418 25782 23420
rect 25838 23418 25862 23420
rect 25918 23418 25942 23420
rect 25998 23418 26022 23420
rect 26078 23418 26084 23420
rect 25838 23366 25840 23418
rect 26020 23366 26022 23418
rect 25776 23364 25782 23366
rect 25838 23364 25862 23366
rect 25918 23364 25942 23366
rect 25998 23364 26022 23366
rect 26078 23364 26084 23366
rect 25776 23344 26084 23364
rect 26516 22976 26568 22982
rect 26516 22918 26568 22924
rect 26332 22432 26384 22438
rect 26332 22374 26384 22380
rect 25776 22332 26084 22352
rect 25776 22330 25782 22332
rect 25838 22330 25862 22332
rect 25918 22330 25942 22332
rect 25998 22330 26022 22332
rect 26078 22330 26084 22332
rect 25838 22278 25840 22330
rect 26020 22278 26022 22330
rect 25776 22276 25782 22278
rect 25838 22276 25862 22278
rect 25918 22276 25942 22278
rect 25998 22276 26022 22278
rect 26078 22276 26084 22278
rect 25776 22256 26084 22276
rect 25700 22188 25820 22216
rect 25596 22160 25648 22166
rect 25596 22102 25648 22108
rect 25688 22092 25740 22098
rect 25688 22034 25740 22040
rect 25412 22024 25464 22030
rect 25412 21966 25464 21972
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25320 21956 25372 21962
rect 25320 21898 25372 21904
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25332 18970 25360 20878
rect 25320 18964 25372 18970
rect 25320 18906 25372 18912
rect 25148 18822 25268 18850
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24872 16046 24900 18022
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24964 16590 24992 17478
rect 25056 17338 25084 17546
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 25148 16266 25176 18702
rect 25240 16402 25268 18822
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 25332 17882 25360 18702
rect 25320 17876 25372 17882
rect 25320 17818 25372 17824
rect 25240 16374 25360 16402
rect 25148 16238 25268 16266
rect 25136 16108 25188 16114
rect 25136 16050 25188 16056
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24780 15694 24900 15722
rect 25148 15706 25176 16050
rect 24872 15502 24900 15694
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24872 13530 24900 15438
rect 25136 14340 25188 14346
rect 25136 14282 25188 14288
rect 25148 13530 25176 14282
rect 25240 13530 25268 16238
rect 25332 15434 25360 16374
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 25228 13524 25280 13530
rect 25228 13466 25280 13472
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24688 12714 24716 13330
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24780 12918 24808 13262
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 25320 13184 25372 13190
rect 25320 13126 25372 13132
rect 24768 12912 24820 12918
rect 24768 12854 24820 12860
rect 24872 12850 24900 13126
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24676 12708 24728 12714
rect 24676 12650 24728 12656
rect 24688 12306 24716 12650
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24676 12300 24728 12306
rect 24676 12242 24728 12248
rect 24872 11830 24900 12582
rect 25136 12096 25188 12102
rect 25136 12038 25188 12044
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 25148 11150 25176 12038
rect 25332 11898 25360 13126
rect 25424 12918 25452 21966
rect 25608 19990 25636 21966
rect 25700 21690 25728 22034
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25792 21570 25820 22188
rect 25700 21542 25820 21570
rect 26148 21616 26200 21622
rect 26148 21558 26200 21564
rect 25596 19984 25648 19990
rect 25596 19926 25648 19932
rect 25596 19712 25648 19718
rect 25596 19654 25648 19660
rect 25504 18964 25556 18970
rect 25504 18906 25556 18912
rect 25516 18834 25544 18906
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 25516 17728 25544 18770
rect 25608 18766 25636 19654
rect 25700 19310 25728 21542
rect 25776 21244 26084 21264
rect 25776 21242 25782 21244
rect 25838 21242 25862 21244
rect 25918 21242 25942 21244
rect 25998 21242 26022 21244
rect 26078 21242 26084 21244
rect 25838 21190 25840 21242
rect 26020 21190 26022 21242
rect 25776 21188 25782 21190
rect 25838 21188 25862 21190
rect 25918 21188 25942 21190
rect 25998 21188 26022 21190
rect 26078 21188 26084 21190
rect 25776 21168 26084 21188
rect 25964 21004 26016 21010
rect 25964 20946 26016 20952
rect 25976 20398 26004 20946
rect 26160 20602 26188 21558
rect 26238 21040 26294 21049
rect 26238 20975 26294 20984
rect 26252 20602 26280 20975
rect 26344 20806 26372 22374
rect 26332 20800 26384 20806
rect 26332 20742 26384 20748
rect 26148 20596 26200 20602
rect 26148 20538 26200 20544
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26160 20398 26188 20538
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 25964 20392 26016 20398
rect 25964 20334 26016 20340
rect 26148 20392 26200 20398
rect 26148 20334 26200 20340
rect 25776 20156 26084 20176
rect 25776 20154 25782 20156
rect 25838 20154 25862 20156
rect 25918 20154 25942 20156
rect 25998 20154 26022 20156
rect 26078 20154 26084 20156
rect 25838 20102 25840 20154
rect 26020 20102 26022 20154
rect 25776 20100 25782 20102
rect 25838 20100 25862 20102
rect 25918 20100 25942 20102
rect 25998 20100 26022 20102
rect 26078 20100 26084 20102
rect 25776 20080 26084 20100
rect 26160 20058 26188 20334
rect 26148 20052 26200 20058
rect 26148 19994 26200 20000
rect 26056 19984 26108 19990
rect 26056 19926 26108 19932
rect 25688 19304 25740 19310
rect 25688 19246 25740 19252
rect 25700 18850 25728 19246
rect 26068 19156 26096 19926
rect 26252 19514 26280 20402
rect 26528 19854 26556 22918
rect 26712 20448 26740 25910
rect 26804 25226 26832 26318
rect 29840 26042 29868 26318
rect 30012 26240 30064 26246
rect 30010 26208 30012 26217
rect 30064 26208 30066 26217
rect 30010 26143 30066 26152
rect 29828 26036 29880 26042
rect 29828 25978 29880 25984
rect 27620 25764 27672 25770
rect 27620 25706 27672 25712
rect 27528 25424 27580 25430
rect 27528 25366 27580 25372
rect 26792 25220 26844 25226
rect 26792 25162 26844 25168
rect 26884 25152 26936 25158
rect 26884 25094 26936 25100
rect 26896 24313 26924 25094
rect 26882 24304 26938 24313
rect 26882 24239 26938 24248
rect 26896 24206 26924 24239
rect 26884 24200 26936 24206
rect 26884 24142 26936 24148
rect 27160 24200 27212 24206
rect 27160 24142 27212 24148
rect 26896 22574 26924 24142
rect 27068 24064 27120 24070
rect 27068 24006 27120 24012
rect 26884 22568 26936 22574
rect 26884 22510 26936 22516
rect 27080 22094 27108 24006
rect 27172 23254 27200 24142
rect 27344 24064 27396 24070
rect 27344 24006 27396 24012
rect 27436 24064 27488 24070
rect 27436 24006 27488 24012
rect 27160 23248 27212 23254
rect 27160 23190 27212 23196
rect 27356 23118 27384 24006
rect 27344 23112 27396 23118
rect 27344 23054 27396 23060
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27080 22066 27292 22094
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 26792 21956 26844 21962
rect 26792 21898 26844 21904
rect 26804 21010 26832 21898
rect 27068 21888 27120 21894
rect 27068 21830 27120 21836
rect 26792 21004 26844 21010
rect 26792 20946 26844 20952
rect 26804 20516 26832 20946
rect 26804 20488 27016 20516
rect 26712 20420 26924 20448
rect 26608 20256 26660 20262
rect 26608 20198 26660 20204
rect 26516 19848 26568 19854
rect 26516 19790 26568 19796
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26068 19128 26188 19156
rect 25776 19068 26084 19088
rect 25776 19066 25782 19068
rect 25838 19066 25862 19068
rect 25918 19066 25942 19068
rect 25998 19066 26022 19068
rect 26078 19066 26084 19068
rect 25838 19014 25840 19066
rect 26020 19014 26022 19066
rect 25776 19012 25782 19014
rect 25838 19012 25862 19014
rect 25918 19012 25942 19014
rect 25998 19012 26022 19014
rect 26078 19012 26084 19014
rect 25776 18992 26084 19012
rect 25700 18822 25912 18850
rect 25884 18766 25912 18822
rect 25596 18760 25648 18766
rect 25596 18702 25648 18708
rect 25872 18760 25924 18766
rect 25872 18702 25924 18708
rect 25594 18048 25650 18057
rect 25594 17983 25650 17992
rect 25608 17864 25636 17983
rect 25776 17980 26084 18000
rect 25776 17978 25782 17980
rect 25838 17978 25862 17980
rect 25918 17978 25942 17980
rect 25998 17978 26022 17980
rect 26078 17978 26084 17980
rect 25838 17926 25840 17978
rect 26020 17926 26022 17978
rect 25776 17924 25782 17926
rect 25838 17924 25862 17926
rect 25918 17924 25942 17926
rect 25998 17924 26022 17926
rect 26078 17924 26084 17926
rect 25776 17904 26084 17924
rect 25688 17876 25740 17882
rect 25608 17836 25688 17864
rect 25688 17818 25740 17824
rect 26054 17776 26110 17785
rect 25596 17740 25648 17746
rect 25516 17700 25596 17728
rect 26054 17711 26110 17720
rect 25596 17682 25648 17688
rect 26068 17678 26096 17711
rect 26056 17672 26108 17678
rect 26056 17614 26108 17620
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 25516 15094 25544 17138
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 25700 16590 25728 16934
rect 25776 16892 26084 16912
rect 25776 16890 25782 16892
rect 25838 16890 25862 16892
rect 25918 16890 25942 16892
rect 25998 16890 26022 16892
rect 26078 16890 26084 16892
rect 25838 16838 25840 16890
rect 26020 16838 26022 16890
rect 25776 16836 25782 16838
rect 25838 16836 25862 16838
rect 25918 16836 25942 16838
rect 25998 16836 26022 16838
rect 26078 16836 26084 16838
rect 25776 16816 26084 16836
rect 25688 16584 25740 16590
rect 25688 16526 25740 16532
rect 26160 16046 26188 19128
rect 26252 18698 26280 19314
rect 26332 19236 26384 19242
rect 26332 19178 26384 19184
rect 26240 18692 26292 18698
rect 26240 18634 26292 18640
rect 26252 17338 26280 18634
rect 26344 18154 26372 19178
rect 26516 18964 26568 18970
rect 26516 18906 26568 18912
rect 26424 18828 26476 18834
rect 26424 18770 26476 18776
rect 26332 18148 26384 18154
rect 26332 18090 26384 18096
rect 26436 17649 26464 18770
rect 26422 17640 26478 17649
rect 26422 17575 26478 17584
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26148 15904 26200 15910
rect 26148 15846 26200 15852
rect 25776 15804 26084 15824
rect 25776 15802 25782 15804
rect 25838 15802 25862 15804
rect 25918 15802 25942 15804
rect 25998 15802 26022 15804
rect 26078 15802 26084 15804
rect 25838 15750 25840 15802
rect 26020 15750 26022 15802
rect 25776 15748 25782 15750
rect 25838 15748 25862 15750
rect 25918 15748 25942 15750
rect 25998 15748 26022 15750
rect 26078 15748 26084 15750
rect 25776 15728 26084 15748
rect 26160 15570 26188 15846
rect 26148 15564 26200 15570
rect 26148 15506 26200 15512
rect 26160 15094 26188 15506
rect 25504 15088 25556 15094
rect 25504 15030 25556 15036
rect 26148 15088 26200 15094
rect 26148 15030 26200 15036
rect 25412 12912 25464 12918
rect 25412 12854 25464 12860
rect 25412 12776 25464 12782
rect 25412 12718 25464 12724
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 24584 10532 24636 10538
rect 24584 10474 24636 10480
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 24964 8294 24992 8978
rect 25136 8900 25188 8906
rect 25136 8842 25188 8848
rect 24952 8288 25004 8294
rect 24952 8230 25004 8236
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24964 6798 24992 8230
rect 25148 7886 25176 8842
rect 25240 8537 25268 9998
rect 25320 8968 25372 8974
rect 25424 8956 25452 12718
rect 25516 11830 25544 15030
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25608 13938 25636 14962
rect 26344 14890 26372 17478
rect 26436 16522 26464 17478
rect 26424 16516 26476 16522
rect 26424 16458 26476 16464
rect 26528 15162 26556 18906
rect 26516 15156 26568 15162
rect 26516 15098 26568 15104
rect 26516 15020 26568 15026
rect 26516 14962 26568 14968
rect 26332 14884 26384 14890
rect 26332 14826 26384 14832
rect 26424 14884 26476 14890
rect 26424 14826 26476 14832
rect 25776 14716 26084 14736
rect 25776 14714 25782 14716
rect 25838 14714 25862 14716
rect 25918 14714 25942 14716
rect 25998 14714 26022 14716
rect 26078 14714 26084 14716
rect 25838 14662 25840 14714
rect 26020 14662 26022 14714
rect 25776 14660 25782 14662
rect 25838 14660 25862 14662
rect 25918 14660 25942 14662
rect 25998 14660 26022 14662
rect 26078 14660 26084 14662
rect 25776 14640 26084 14660
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25700 13938 25728 14214
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25688 13932 25740 13938
rect 25688 13874 25740 13880
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 25608 13258 25636 13874
rect 25700 13326 25728 13874
rect 25776 13628 26084 13648
rect 25776 13626 25782 13628
rect 25838 13626 25862 13628
rect 25918 13626 25942 13628
rect 25998 13626 26022 13628
rect 26078 13626 26084 13628
rect 25838 13574 25840 13626
rect 26020 13574 26022 13626
rect 25776 13572 25782 13574
rect 25838 13572 25862 13574
rect 25918 13572 25942 13574
rect 25998 13572 26022 13574
rect 26078 13572 26084 13574
rect 25776 13552 26084 13572
rect 26344 13326 26372 13874
rect 25688 13320 25740 13326
rect 25688 13262 25740 13268
rect 26332 13320 26384 13326
rect 26332 13262 26384 13268
rect 25596 13252 25648 13258
rect 25596 13194 25648 13200
rect 25608 12850 25636 13194
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25776 12540 26084 12560
rect 25776 12538 25782 12540
rect 25838 12538 25862 12540
rect 25918 12538 25942 12540
rect 25998 12538 26022 12540
rect 26078 12538 26084 12540
rect 25838 12486 25840 12538
rect 26020 12486 26022 12538
rect 25776 12484 25782 12486
rect 25838 12484 25862 12486
rect 25918 12484 25942 12486
rect 25998 12484 26022 12486
rect 26078 12484 26084 12486
rect 25776 12464 26084 12484
rect 26252 12238 26280 12922
rect 26436 12434 26464 14826
rect 26528 13938 26556 14962
rect 26516 13932 26568 13938
rect 26516 13874 26568 13880
rect 26620 13818 26648 20198
rect 26700 19984 26752 19990
rect 26700 19926 26752 19932
rect 26344 12406 26464 12434
rect 26528 13790 26648 13818
rect 26240 12232 26292 12238
rect 26240 12174 26292 12180
rect 25688 12164 25740 12170
rect 25688 12106 25740 12112
rect 25504 11824 25556 11830
rect 25504 11766 25556 11772
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 25608 11150 25636 11494
rect 25700 11354 25728 12106
rect 26148 12096 26200 12102
rect 26148 12038 26200 12044
rect 25776 11452 26084 11472
rect 25776 11450 25782 11452
rect 25838 11450 25862 11452
rect 25918 11450 25942 11452
rect 25998 11450 26022 11452
rect 26078 11450 26084 11452
rect 25838 11398 25840 11450
rect 26020 11398 26022 11450
rect 25776 11396 25782 11398
rect 25838 11396 25862 11398
rect 25918 11396 25942 11398
rect 25998 11396 26022 11398
rect 26078 11396 26084 11398
rect 25776 11376 26084 11396
rect 25688 11348 25740 11354
rect 25688 11290 25740 11296
rect 25596 11144 25648 11150
rect 25596 11086 25648 11092
rect 25608 10674 25636 11086
rect 25596 10668 25648 10674
rect 25596 10610 25648 10616
rect 25688 10668 25740 10674
rect 25688 10610 25740 10616
rect 25372 8928 25452 8956
rect 25320 8910 25372 8916
rect 25226 8528 25282 8537
rect 25226 8463 25282 8472
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25240 6848 25268 8463
rect 25332 8362 25360 8910
rect 25320 8356 25372 8362
rect 25320 8298 25372 8304
rect 25320 6860 25372 6866
rect 25240 6820 25320 6848
rect 25320 6802 25372 6808
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 23952 5778 23980 6258
rect 23940 5772 23992 5778
rect 23940 5714 23992 5720
rect 23848 5296 23900 5302
rect 23848 5238 23900 5244
rect 24964 5234 24992 6734
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 24952 5228 25004 5234
rect 24952 5170 25004 5176
rect 23216 4826 23244 5170
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 24964 4622 24992 5170
rect 25332 5166 25360 6802
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 25424 6390 25452 6734
rect 25700 6458 25728 10610
rect 26056 10600 26108 10606
rect 26160 10588 26188 12038
rect 26108 10560 26188 10588
rect 26056 10542 26108 10548
rect 25776 10364 26084 10384
rect 25776 10362 25782 10364
rect 25838 10362 25862 10364
rect 25918 10362 25942 10364
rect 25998 10362 26022 10364
rect 26078 10362 26084 10364
rect 25838 10310 25840 10362
rect 26020 10310 26022 10362
rect 25776 10308 25782 10310
rect 25838 10308 25862 10310
rect 25918 10308 25942 10310
rect 25998 10308 26022 10310
rect 26078 10308 26084 10310
rect 25776 10288 26084 10308
rect 26160 9586 26188 10560
rect 26148 9580 26200 9586
rect 26148 9522 26200 9528
rect 25776 9276 26084 9296
rect 25776 9274 25782 9276
rect 25838 9274 25862 9276
rect 25918 9274 25942 9276
rect 25998 9274 26022 9276
rect 26078 9274 26084 9276
rect 25838 9222 25840 9274
rect 26020 9222 26022 9274
rect 25776 9220 25782 9222
rect 25838 9220 25862 9222
rect 25918 9220 25942 9222
rect 25998 9220 26022 9222
rect 26078 9220 26084 9222
rect 25776 9200 26084 9220
rect 26160 8974 26188 9522
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 26148 8492 26200 8498
rect 26148 8434 26200 8440
rect 25776 8188 26084 8208
rect 25776 8186 25782 8188
rect 25838 8186 25862 8188
rect 25918 8186 25942 8188
rect 25998 8186 26022 8188
rect 26078 8186 26084 8188
rect 25838 8134 25840 8186
rect 26020 8134 26022 8186
rect 25776 8132 25782 8134
rect 25838 8132 25862 8134
rect 25918 8132 25942 8134
rect 25998 8132 26022 8134
rect 26078 8132 26084 8134
rect 25776 8112 26084 8132
rect 25776 7100 26084 7120
rect 25776 7098 25782 7100
rect 25838 7098 25862 7100
rect 25918 7098 25942 7100
rect 25998 7098 26022 7100
rect 26078 7098 26084 7100
rect 25838 7046 25840 7098
rect 26020 7046 26022 7098
rect 25776 7044 25782 7046
rect 25838 7044 25862 7046
rect 25918 7044 25942 7046
rect 25998 7044 26022 7046
rect 26078 7044 26084 7046
rect 25776 7024 26084 7044
rect 26160 6866 26188 8434
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 26252 7342 26280 8366
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26148 6860 26200 6866
rect 26148 6802 26200 6808
rect 25688 6452 25740 6458
rect 25688 6394 25740 6400
rect 25412 6384 25464 6390
rect 25412 6326 25464 6332
rect 25596 6316 25648 6322
rect 25596 6258 25648 6264
rect 25608 5370 25636 6258
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 25700 5234 25728 6394
rect 26160 6186 26188 6802
rect 26344 6798 26372 12406
rect 26528 12374 26556 13790
rect 26608 13728 26660 13734
rect 26608 13670 26660 13676
rect 26516 12368 26568 12374
rect 26516 12310 26568 12316
rect 26620 11234 26648 13670
rect 26712 11286 26740 19926
rect 26792 15156 26844 15162
rect 26792 15098 26844 15104
rect 26804 14414 26832 15098
rect 26792 14408 26844 14414
rect 26792 14350 26844 14356
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26804 12850 26832 13262
rect 26792 12844 26844 12850
rect 26792 12786 26844 12792
rect 26804 12238 26832 12786
rect 26896 12434 26924 20420
rect 26988 19990 27016 20488
rect 26976 19984 27028 19990
rect 26976 19926 27028 19932
rect 26988 19718 27016 19926
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 26988 17746 27016 19654
rect 26976 17740 27028 17746
rect 26976 17682 27028 17688
rect 26974 17640 27030 17649
rect 26974 17575 27030 17584
rect 26988 14618 27016 17575
rect 26976 14612 27028 14618
rect 26976 14554 27028 14560
rect 26976 14340 27028 14346
rect 26976 14282 27028 14288
rect 26988 13734 27016 14282
rect 26976 13728 27028 13734
rect 26976 13670 27028 13676
rect 26988 13326 27016 13670
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 26896 12406 27016 12434
rect 26792 12232 26844 12238
rect 26792 12174 26844 12180
rect 26884 11620 26936 11626
rect 26884 11562 26936 11568
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 26528 11218 26648 11234
rect 26700 11280 26752 11286
rect 26700 11222 26752 11228
rect 26516 11212 26648 11218
rect 26568 11206 26648 11212
rect 26516 11154 26568 11160
rect 26528 10810 26556 11154
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26516 10804 26568 10810
rect 26516 10746 26568 10752
rect 26528 10674 26556 10746
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26148 6180 26200 6186
rect 26148 6122 26200 6128
rect 25776 6012 26084 6032
rect 25776 6010 25782 6012
rect 25838 6010 25862 6012
rect 25918 6010 25942 6012
rect 25998 6010 26022 6012
rect 26078 6010 26084 6012
rect 25838 5958 25840 6010
rect 26020 5958 26022 6010
rect 25776 5956 25782 5958
rect 25838 5956 25862 5958
rect 25918 5956 25942 5958
rect 25998 5956 26022 5958
rect 26078 5956 26084 5958
rect 25776 5936 26084 5956
rect 26160 5794 26188 6122
rect 26344 5846 26372 6734
rect 26620 5914 26648 11086
rect 26804 10606 26832 11290
rect 26896 11082 26924 11562
rect 26884 11076 26936 11082
rect 26884 11018 26936 11024
rect 26792 10600 26844 10606
rect 26792 10542 26844 10548
rect 26896 10062 26924 11018
rect 26988 10130 27016 12406
rect 27080 10606 27108 21830
rect 27172 21622 27200 21966
rect 27264 21894 27292 22066
rect 27356 21962 27384 22578
rect 27448 22098 27476 24006
rect 27540 22710 27568 25366
rect 27632 25226 27660 25706
rect 30012 25696 30064 25702
rect 30012 25638 30064 25644
rect 30024 25401 30052 25638
rect 30010 25392 30066 25401
rect 30010 25327 30066 25336
rect 28908 25288 28960 25294
rect 28908 25230 28960 25236
rect 27620 25220 27672 25226
rect 27620 25162 27672 25168
rect 28632 25220 28684 25226
rect 28632 25162 28684 25168
rect 27528 22704 27580 22710
rect 27528 22646 27580 22652
rect 27632 22438 27660 25162
rect 28356 24812 28408 24818
rect 28356 24754 28408 24760
rect 28540 24812 28592 24818
rect 28540 24754 28592 24760
rect 28080 24268 28132 24274
rect 28080 24210 28132 24216
rect 27804 24200 27856 24206
rect 27804 24142 27856 24148
rect 27712 23860 27764 23866
rect 27712 23802 27764 23808
rect 27620 22432 27672 22438
rect 27620 22374 27672 22380
rect 27620 22228 27672 22234
rect 27620 22170 27672 22176
rect 27436 22092 27488 22098
rect 27436 22034 27488 22040
rect 27344 21956 27396 21962
rect 27344 21898 27396 21904
rect 27252 21888 27304 21894
rect 27252 21830 27304 21836
rect 27160 21616 27212 21622
rect 27160 21558 27212 21564
rect 27252 21548 27304 21554
rect 27356 21536 27384 21898
rect 27304 21508 27384 21536
rect 27252 21490 27304 21496
rect 27264 20466 27292 21490
rect 27344 21072 27396 21078
rect 27632 21026 27660 22170
rect 27344 21014 27396 21020
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 27252 19848 27304 19854
rect 27172 19808 27252 19836
rect 27172 18766 27200 19808
rect 27252 19790 27304 19796
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 27172 17202 27200 18702
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 27264 17338 27292 18226
rect 27252 17332 27304 17338
rect 27252 17274 27304 17280
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 27172 16590 27200 17138
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27252 16584 27304 16590
rect 27356 16572 27384 21014
rect 27540 20998 27660 21026
rect 27436 20800 27488 20806
rect 27436 20742 27488 20748
rect 27448 20534 27476 20742
rect 27436 20528 27488 20534
rect 27436 20470 27488 20476
rect 27540 20482 27568 20998
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27632 20602 27660 20878
rect 27620 20596 27672 20602
rect 27620 20538 27672 20544
rect 27540 20454 27660 20482
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 27436 19984 27488 19990
rect 27436 19926 27488 19932
rect 27448 17134 27476 19926
rect 27540 19310 27568 20198
rect 27528 19304 27580 19310
rect 27528 19246 27580 19252
rect 27632 18850 27660 20454
rect 27724 20330 27752 23802
rect 27816 23526 27844 24142
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 27804 23520 27856 23526
rect 27804 23462 27856 23468
rect 27816 22642 27844 23462
rect 28000 22778 28028 23666
rect 28092 23186 28120 24210
rect 28264 24200 28316 24206
rect 28264 24142 28316 24148
rect 28172 24064 28224 24070
rect 28172 24006 28224 24012
rect 28080 23180 28132 23186
rect 28080 23122 28132 23128
rect 27988 22772 28040 22778
rect 27988 22714 28040 22720
rect 27804 22636 27856 22642
rect 27804 22578 27856 22584
rect 28092 22574 28120 23122
rect 28080 22568 28132 22574
rect 28080 22510 28132 22516
rect 27988 22500 28040 22506
rect 27988 22442 28040 22448
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 27816 21010 27844 22374
rect 27894 22128 27950 22137
rect 27894 22063 27950 22072
rect 27908 21554 27936 22063
rect 28000 21554 28028 22442
rect 28092 22137 28120 22510
rect 28078 22128 28134 22137
rect 28078 22063 28134 22072
rect 28080 22024 28132 22030
rect 28080 21966 28132 21972
rect 27896 21548 27948 21554
rect 27896 21490 27948 21496
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 27804 21004 27856 21010
rect 27804 20946 27856 20952
rect 27712 20324 27764 20330
rect 27712 20266 27764 20272
rect 27712 19848 27764 19854
rect 27712 19790 27764 19796
rect 27540 18822 27660 18850
rect 27540 17746 27568 18822
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27632 18358 27660 18702
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 27724 18193 27752 19790
rect 27710 18184 27766 18193
rect 27710 18119 27766 18128
rect 27620 17808 27672 17814
rect 27618 17776 27620 17785
rect 27672 17776 27674 17785
rect 27528 17740 27580 17746
rect 27618 17711 27674 17720
rect 27528 17682 27580 17688
rect 27436 17128 27488 17134
rect 27436 17070 27488 17076
rect 27448 16726 27476 17070
rect 27540 16794 27568 17682
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 27528 16788 27580 16794
rect 27528 16730 27580 16736
rect 27436 16720 27488 16726
rect 27436 16662 27488 16668
rect 27304 16544 27384 16572
rect 27252 16526 27304 16532
rect 27172 16250 27200 16526
rect 27344 16448 27396 16454
rect 27344 16390 27396 16396
rect 27160 16244 27212 16250
rect 27160 16186 27212 16192
rect 27172 13938 27200 16186
rect 27356 16182 27384 16390
rect 27344 16176 27396 16182
rect 27344 16118 27396 16124
rect 27252 15904 27304 15910
rect 27252 15846 27304 15852
rect 27264 15366 27292 15846
rect 27252 15360 27304 15366
rect 27252 15302 27304 15308
rect 27264 14414 27292 15302
rect 27252 14408 27304 14414
rect 27252 14350 27304 14356
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27068 10600 27120 10606
rect 27068 10542 27120 10548
rect 26976 10124 27028 10130
rect 26976 10066 27028 10072
rect 26884 10056 26936 10062
rect 26884 9998 26936 10004
rect 26988 9654 27016 10066
rect 26976 9648 27028 9654
rect 26976 9590 27028 9596
rect 26988 8974 27016 9590
rect 26976 8968 27028 8974
rect 26976 8910 27028 8916
rect 27172 8566 27200 10610
rect 27356 9042 27384 16118
rect 27448 15094 27476 16662
rect 27540 16114 27568 16730
rect 27632 16726 27660 17614
rect 27620 16720 27672 16726
rect 27620 16662 27672 16668
rect 27816 16640 27844 20946
rect 27908 20466 27936 21490
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 28092 20058 28120 21966
rect 28184 21622 28212 24006
rect 28172 21616 28224 21622
rect 28172 21558 28224 21564
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28184 20942 28212 21422
rect 28172 20936 28224 20942
rect 28172 20878 28224 20884
rect 28184 20398 28212 20878
rect 28172 20392 28224 20398
rect 28172 20334 28224 20340
rect 28184 20074 28212 20334
rect 28276 20233 28304 24142
rect 28368 23225 28396 24754
rect 28448 23792 28500 23798
rect 28448 23734 28500 23740
rect 28354 23216 28410 23225
rect 28354 23151 28410 23160
rect 28356 23044 28408 23050
rect 28356 22986 28408 22992
rect 28368 22234 28396 22986
rect 28460 22642 28488 23734
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28356 22228 28408 22234
rect 28356 22170 28408 22176
rect 28356 21956 28408 21962
rect 28356 21898 28408 21904
rect 28368 20942 28396 21898
rect 28460 21554 28488 22578
rect 28448 21548 28500 21554
rect 28448 21490 28500 21496
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28460 20466 28488 21490
rect 28552 21049 28580 24754
rect 28644 22234 28672 25162
rect 28816 25152 28868 25158
rect 28816 25094 28868 25100
rect 28724 24608 28776 24614
rect 28724 24550 28776 24556
rect 28632 22228 28684 22234
rect 28632 22170 28684 22176
rect 28630 22128 28686 22137
rect 28736 22098 28764 24550
rect 28828 24342 28856 25094
rect 28816 24336 28868 24342
rect 28816 24278 28868 24284
rect 28816 23724 28868 23730
rect 28816 23666 28868 23672
rect 28630 22063 28686 22072
rect 28724 22092 28776 22098
rect 28644 22030 28672 22063
rect 28724 22034 28776 22040
rect 28632 22024 28684 22030
rect 28632 21966 28684 21972
rect 28538 21040 28594 21049
rect 28538 20975 28594 20984
rect 28448 20460 28500 20466
rect 28448 20402 28500 20408
rect 28262 20224 28318 20233
rect 28262 20159 28318 20168
rect 28080 20052 28132 20058
rect 28184 20046 28304 20074
rect 28080 19994 28132 20000
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 28000 18358 28028 19790
rect 28172 19508 28224 19514
rect 28172 19450 28224 19456
rect 27988 18352 28040 18358
rect 27988 18294 28040 18300
rect 28000 17746 28028 18294
rect 28080 18080 28132 18086
rect 28080 18022 28132 18028
rect 27988 17740 28040 17746
rect 27988 17682 28040 17688
rect 27896 17536 27948 17542
rect 27896 17478 27948 17484
rect 27724 16612 27844 16640
rect 27620 16176 27672 16182
rect 27620 16118 27672 16124
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27436 15088 27488 15094
rect 27436 15030 27488 15036
rect 27448 14482 27476 15030
rect 27632 14618 27660 16118
rect 27724 14890 27752 16612
rect 27712 14884 27764 14890
rect 27712 14826 27764 14832
rect 27620 14612 27672 14618
rect 27620 14554 27672 14560
rect 27724 14482 27752 14826
rect 27436 14476 27488 14482
rect 27436 14418 27488 14424
rect 27712 14476 27764 14482
rect 27712 14418 27764 14424
rect 27448 13818 27476 14418
rect 27908 13938 27936 17478
rect 28000 17134 28028 17682
rect 28092 17202 28120 18022
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 27988 17128 28040 17134
rect 27988 17070 28040 17076
rect 28000 16658 28028 17070
rect 28080 16720 28132 16726
rect 28080 16662 28132 16668
rect 27988 16652 28040 16658
rect 27988 16594 28040 16600
rect 27988 16040 28040 16046
rect 27988 15982 28040 15988
rect 28000 14346 28028 15982
rect 28092 15978 28120 16662
rect 28080 15972 28132 15978
rect 28080 15914 28132 15920
rect 28184 15706 28212 19450
rect 28276 18222 28304 20046
rect 28356 19712 28408 19718
rect 28356 19654 28408 19660
rect 28368 18290 28396 19654
rect 28460 19378 28488 20402
rect 28540 19780 28592 19786
rect 28540 19722 28592 19728
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 28460 19242 28488 19314
rect 28448 19236 28500 19242
rect 28448 19178 28500 19184
rect 28460 18766 28488 19178
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28264 18216 28316 18222
rect 28264 18158 28316 18164
rect 28276 16726 28304 18158
rect 28356 17604 28408 17610
rect 28356 17546 28408 17552
rect 28264 16720 28316 16726
rect 28264 16662 28316 16668
rect 28264 16584 28316 16590
rect 28264 16526 28316 16532
rect 28276 16250 28304 16526
rect 28264 16244 28316 16250
rect 28264 16186 28316 16192
rect 28264 15972 28316 15978
rect 28264 15914 28316 15920
rect 28172 15700 28224 15706
rect 28172 15642 28224 15648
rect 28080 15632 28132 15638
rect 28080 15574 28132 15580
rect 27988 14340 28040 14346
rect 27988 14282 28040 14288
rect 27896 13932 27948 13938
rect 27896 13874 27948 13880
rect 27528 13864 27580 13870
rect 27448 13812 27528 13818
rect 27448 13806 27580 13812
rect 27448 13790 27568 13806
rect 28000 13802 28028 14282
rect 28092 13938 28120 15574
rect 28172 15428 28224 15434
rect 28172 15370 28224 15376
rect 28184 14074 28212 15370
rect 28172 14068 28224 14074
rect 28172 14010 28224 14016
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 28276 13818 28304 15914
rect 28184 13802 28304 13818
rect 27620 13796 27672 13802
rect 27620 13738 27672 13744
rect 27988 13796 28040 13802
rect 27988 13738 28040 13744
rect 28172 13796 28304 13802
rect 28224 13790 28304 13796
rect 28172 13738 28224 13744
rect 27632 13682 27660 13738
rect 27540 13654 27660 13682
rect 27712 13728 27764 13734
rect 27712 13670 27764 13676
rect 27540 13512 27568 13654
rect 27448 13484 27568 13512
rect 27448 13326 27476 13484
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 27632 12986 27660 13262
rect 27620 12980 27672 12986
rect 27620 12922 27672 12928
rect 27724 12238 27752 13670
rect 27896 13252 27948 13258
rect 27896 13194 27948 13200
rect 27804 13184 27856 13190
rect 27804 13126 27856 13132
rect 27816 12850 27844 13126
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 27804 12368 27856 12374
rect 27804 12310 27856 12316
rect 27712 12232 27764 12238
rect 27712 12174 27764 12180
rect 27712 12096 27764 12102
rect 27712 12038 27764 12044
rect 27724 11762 27752 12038
rect 27712 11756 27764 11762
rect 27712 11698 27764 11704
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27528 9988 27580 9994
rect 27528 9930 27580 9936
rect 27344 9036 27396 9042
rect 27344 8978 27396 8984
rect 27160 8560 27212 8566
rect 27160 8502 27212 8508
rect 27172 8090 27200 8502
rect 27356 8430 27384 8978
rect 27344 8424 27396 8430
rect 27344 8366 27396 8372
rect 27540 8090 27568 9930
rect 27632 9586 27660 11630
rect 27816 11506 27844 12310
rect 27724 11478 27844 11506
rect 27620 9580 27672 9586
rect 27620 9522 27672 9528
rect 27160 8084 27212 8090
rect 27160 8026 27212 8032
rect 27528 8084 27580 8090
rect 27528 8026 27580 8032
rect 27632 8022 27660 9522
rect 27724 8514 27752 11478
rect 27802 11384 27858 11393
rect 27802 11319 27858 11328
rect 27816 11150 27844 11319
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27724 8486 27844 8514
rect 27712 8424 27764 8430
rect 27712 8366 27764 8372
rect 27620 8016 27672 8022
rect 27620 7958 27672 7964
rect 27632 7886 27660 7958
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27620 7744 27672 7750
rect 27620 7686 27672 7692
rect 27252 7404 27304 7410
rect 27252 7346 27304 7352
rect 27264 7002 27292 7346
rect 27252 6996 27304 7002
rect 27252 6938 27304 6944
rect 26700 6792 26752 6798
rect 26700 6734 26752 6740
rect 26712 6254 26740 6734
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 26700 6248 26752 6254
rect 26700 6190 26752 6196
rect 26608 5908 26660 5914
rect 26608 5850 26660 5856
rect 26068 5766 26188 5794
rect 26332 5840 26384 5846
rect 26332 5782 26384 5788
rect 25688 5228 25740 5234
rect 25688 5170 25740 5176
rect 26068 5166 26096 5766
rect 26148 5636 26200 5642
rect 26148 5578 26200 5584
rect 25320 5160 25372 5166
rect 25780 5160 25832 5166
rect 25320 5102 25372 5108
rect 25700 5108 25780 5114
rect 25700 5102 25832 5108
rect 26056 5160 26108 5166
rect 26056 5102 26108 5108
rect 24952 4616 25004 4622
rect 24952 4558 25004 4564
rect 25332 4554 25360 5102
rect 25700 5086 25820 5102
rect 25700 4706 25728 5086
rect 25776 4924 26084 4944
rect 25776 4922 25782 4924
rect 25838 4922 25862 4924
rect 25918 4922 25942 4924
rect 25998 4922 26022 4924
rect 26078 4922 26084 4924
rect 25838 4870 25840 4922
rect 26020 4870 26022 4922
rect 25776 4868 25782 4870
rect 25838 4868 25862 4870
rect 25918 4868 25942 4870
rect 25998 4868 26022 4870
rect 26078 4868 26084 4870
rect 25776 4848 26084 4868
rect 26160 4826 26188 5578
rect 26148 4820 26200 4826
rect 26148 4762 26200 4768
rect 25700 4690 25820 4706
rect 25700 4684 25832 4690
rect 25700 4678 25780 4684
rect 25780 4626 25832 4632
rect 26620 4622 26648 5850
rect 27356 5642 27384 6598
rect 27632 6322 27660 7686
rect 27724 7206 27752 8366
rect 27712 7200 27764 7206
rect 27712 7142 27764 7148
rect 27724 6798 27752 7142
rect 27712 6792 27764 6798
rect 27712 6734 27764 6740
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 27436 6248 27488 6254
rect 27488 6196 27660 6202
rect 27436 6190 27660 6196
rect 27448 6186 27660 6190
rect 27448 6180 27672 6186
rect 27448 6174 27620 6180
rect 27620 6122 27672 6128
rect 27724 5710 27752 6734
rect 27816 6662 27844 8486
rect 27908 7546 27936 13194
rect 28000 13190 28028 13738
rect 28264 13728 28316 13734
rect 28264 13670 28316 13676
rect 28172 13524 28224 13530
rect 28172 13466 28224 13472
rect 27988 13184 28040 13190
rect 27988 13126 28040 13132
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 28092 11014 28120 11698
rect 28080 11008 28132 11014
rect 28080 10950 28132 10956
rect 28092 10810 28120 10950
rect 28080 10804 28132 10810
rect 28080 10746 28132 10752
rect 28080 9444 28132 9450
rect 28080 9386 28132 9392
rect 27988 9036 28040 9042
rect 27988 8978 28040 8984
rect 28000 7886 28028 8978
rect 27988 7880 28040 7886
rect 27988 7822 28040 7828
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 27908 7002 27936 7482
rect 28000 7274 28028 7822
rect 28092 7818 28120 9386
rect 28184 9178 28212 13466
rect 28276 13326 28304 13670
rect 28264 13320 28316 13326
rect 28368 13308 28396 17546
rect 28460 17202 28488 18702
rect 28552 18154 28580 19722
rect 28828 19553 28856 23666
rect 28920 22409 28948 25230
rect 30010 24712 30066 24721
rect 29828 24676 29880 24682
rect 30010 24647 30012 24656
rect 29828 24618 29880 24624
rect 30064 24647 30066 24656
rect 30012 24618 30064 24624
rect 29840 24206 29868 24618
rect 29828 24200 29880 24206
rect 29828 24142 29880 24148
rect 30012 24064 30064 24070
rect 30012 24006 30064 24012
rect 30024 23905 30052 24006
rect 30010 23896 30066 23905
rect 30010 23831 30066 23840
rect 30104 23724 30156 23730
rect 30104 23666 30156 23672
rect 29828 23520 29880 23526
rect 29828 23462 29880 23468
rect 29000 22636 29052 22642
rect 29000 22578 29052 22584
rect 28906 22400 28962 22409
rect 28906 22335 28962 22344
rect 28908 22228 28960 22234
rect 28908 22170 28960 22176
rect 28920 21729 28948 22170
rect 29012 22098 29040 22578
rect 29552 22432 29604 22438
rect 29552 22374 29604 22380
rect 29000 22092 29052 22098
rect 29000 22034 29052 22040
rect 29564 22030 29592 22374
rect 29552 22024 29604 22030
rect 29552 21966 29604 21972
rect 28906 21720 28962 21729
rect 28906 21655 28962 21664
rect 29092 20936 29144 20942
rect 29092 20878 29144 20884
rect 28814 19544 28870 19553
rect 28814 19479 28870 19488
rect 29000 19372 29052 19378
rect 29000 19314 29052 19320
rect 28724 19236 28776 19242
rect 28724 19178 28776 19184
rect 28632 18760 28684 18766
rect 28632 18702 28684 18708
rect 28540 18148 28592 18154
rect 28540 18090 28592 18096
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 28460 16114 28488 17138
rect 28448 16108 28500 16114
rect 28448 16050 28500 16056
rect 28460 15502 28488 16050
rect 28448 15496 28500 15502
rect 28448 15438 28500 15444
rect 28460 15026 28488 15438
rect 28552 15065 28580 17614
rect 28538 15056 28594 15065
rect 28448 15020 28500 15026
rect 28538 14991 28594 15000
rect 28448 14962 28500 14968
rect 28540 14408 28592 14414
rect 28644 14385 28672 18702
rect 28736 18290 28764 19178
rect 29012 18834 29040 19314
rect 29000 18828 29052 18834
rect 29000 18770 29052 18776
rect 29104 18442 29132 20878
rect 29460 19848 29512 19854
rect 29512 19808 29592 19836
rect 29460 19790 29512 19796
rect 29184 19508 29236 19514
rect 29184 19450 29236 19456
rect 29012 18414 29132 18442
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 29012 17954 29040 18414
rect 29092 18352 29144 18358
rect 29092 18294 29144 18300
rect 29104 18154 29132 18294
rect 29092 18148 29144 18154
rect 29092 18090 29144 18096
rect 28920 17926 29040 17954
rect 28816 17740 28868 17746
rect 28816 17682 28868 17688
rect 28724 17196 28776 17202
rect 28724 17138 28776 17144
rect 28736 16794 28764 17138
rect 28724 16788 28776 16794
rect 28724 16730 28776 16736
rect 28540 14350 28592 14356
rect 28630 14376 28686 14385
rect 28552 13530 28580 14350
rect 28630 14311 28686 14320
rect 28724 13864 28776 13870
rect 28724 13806 28776 13812
rect 28632 13796 28684 13802
rect 28632 13738 28684 13744
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 28448 13320 28500 13326
rect 28368 13280 28448 13308
rect 28264 13262 28316 13268
rect 28448 13262 28500 13268
rect 28276 12850 28304 13262
rect 28264 12844 28316 12850
rect 28264 12786 28316 12792
rect 28552 12782 28580 13466
rect 28644 13462 28672 13738
rect 28632 13456 28684 13462
rect 28632 13398 28684 13404
rect 28736 12918 28764 13806
rect 28828 13569 28856 17682
rect 28920 15881 28948 17926
rect 29196 16980 29224 19450
rect 29368 18828 29420 18834
rect 29368 18770 29420 18776
rect 29276 16992 29328 16998
rect 29196 16952 29276 16980
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 28906 15872 28962 15881
rect 28906 15807 28962 15816
rect 29012 15722 29040 16594
rect 29196 16590 29224 16952
rect 29276 16934 29328 16940
rect 29380 16794 29408 18770
rect 29460 18624 29512 18630
rect 29460 18566 29512 18572
rect 29472 18290 29500 18566
rect 29460 18284 29512 18290
rect 29460 18226 29512 18232
rect 29472 17814 29500 18226
rect 29460 17808 29512 17814
rect 29460 17750 29512 17756
rect 29564 16998 29592 19808
rect 29736 18692 29788 18698
rect 29736 18634 29788 18640
rect 29748 18426 29776 18634
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 29552 16992 29604 16998
rect 29552 16934 29604 16940
rect 29368 16788 29420 16794
rect 29368 16730 29420 16736
rect 29184 16584 29236 16590
rect 29184 16526 29236 16532
rect 29564 16454 29592 16934
rect 29840 16522 29868 23462
rect 30116 18057 30144 23666
rect 30102 18048 30158 18057
rect 30102 17983 30158 17992
rect 29828 16516 29880 16522
rect 29828 16458 29880 16464
rect 29552 16448 29604 16454
rect 29552 16390 29604 16396
rect 29644 16448 29696 16454
rect 29644 16390 29696 16396
rect 29656 16182 29684 16390
rect 29644 16176 29696 16182
rect 29644 16118 29696 16124
rect 28920 15694 29040 15722
rect 28920 15638 28948 15694
rect 28908 15632 28960 15638
rect 28908 15574 28960 15580
rect 28908 15496 28960 15502
rect 28908 15438 28960 15444
rect 28814 13560 28870 13569
rect 28814 13495 28870 13504
rect 28816 13184 28868 13190
rect 28816 13126 28868 13132
rect 28828 12918 28856 13126
rect 28724 12912 28776 12918
rect 28724 12854 28776 12860
rect 28816 12912 28868 12918
rect 28920 12889 28948 15438
rect 29092 15428 29144 15434
rect 29092 15370 29144 15376
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 29012 13530 29040 14962
rect 29104 14822 29132 15370
rect 29184 15360 29236 15366
rect 29184 15302 29236 15308
rect 29092 14816 29144 14822
rect 29092 14758 29144 14764
rect 29000 13524 29052 13530
rect 29000 13466 29052 13472
rect 29104 13326 29132 14758
rect 29092 13320 29144 13326
rect 29092 13262 29144 13268
rect 28816 12854 28868 12860
rect 28906 12880 28962 12889
rect 28540 12776 28592 12782
rect 28540 12718 28592 12724
rect 28264 12232 28316 12238
rect 28264 12174 28316 12180
rect 28276 11150 28304 12174
rect 28552 11830 28580 12718
rect 28540 11824 28592 11830
rect 28540 11766 28592 11772
rect 28552 11218 28580 11766
rect 28736 11694 28764 12854
rect 29196 12850 29224 15302
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 29920 14000 29972 14006
rect 29920 13942 29972 13948
rect 29736 13932 29788 13938
rect 29736 13874 29788 13880
rect 29552 13320 29604 13326
rect 29552 13262 29604 13268
rect 29564 12986 29592 13262
rect 29748 12986 29776 13874
rect 29552 12980 29604 12986
rect 29552 12922 29604 12928
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 28906 12815 28962 12824
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 29184 12232 29236 12238
rect 29184 12174 29236 12180
rect 28908 12096 28960 12102
rect 28814 12064 28870 12073
rect 28908 12038 28960 12044
rect 28814 11999 28870 12008
rect 28724 11688 28776 11694
rect 28724 11630 28776 11636
rect 28632 11620 28684 11626
rect 28632 11562 28684 11568
rect 28540 11212 28592 11218
rect 28540 11154 28592 11160
rect 28644 11150 28672 11562
rect 28736 11354 28764 11630
rect 28724 11348 28776 11354
rect 28724 11290 28776 11296
rect 28264 11144 28316 11150
rect 28264 11086 28316 11092
rect 28632 11144 28684 11150
rect 28632 11086 28684 11092
rect 28540 10600 28592 10606
rect 28540 10542 28592 10548
rect 28552 10266 28580 10542
rect 28540 10260 28592 10266
rect 28540 10202 28592 10208
rect 28172 9172 28224 9178
rect 28172 9114 28224 9120
rect 28552 7886 28580 10202
rect 28644 9042 28672 11086
rect 28736 10606 28764 11290
rect 28724 10600 28776 10606
rect 28724 10542 28776 10548
rect 28736 10062 28764 10542
rect 28724 10056 28776 10062
rect 28724 9998 28776 10004
rect 28736 9518 28764 9998
rect 28724 9512 28776 9518
rect 28724 9454 28776 9460
rect 28632 9036 28684 9042
rect 28632 8978 28684 8984
rect 28736 8430 28764 9454
rect 28828 8974 28856 11999
rect 28816 8968 28868 8974
rect 28816 8910 28868 8916
rect 28816 8832 28868 8838
rect 28816 8774 28868 8780
rect 28724 8424 28776 8430
rect 28724 8366 28776 8372
rect 28724 8016 28776 8022
rect 28724 7958 28776 7964
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28080 7812 28132 7818
rect 28080 7754 28132 7760
rect 28092 7342 28120 7754
rect 28736 7410 28764 7958
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 28724 7404 28776 7410
rect 28724 7346 28776 7352
rect 28080 7336 28132 7342
rect 28080 7278 28132 7284
rect 27988 7268 28040 7274
rect 27988 7210 28040 7216
rect 27896 6996 27948 7002
rect 27896 6938 27948 6944
rect 27896 6724 27948 6730
rect 27896 6666 27948 6672
rect 27804 6656 27856 6662
rect 27804 6598 27856 6604
rect 27816 6322 27844 6598
rect 27908 6458 27936 6666
rect 27896 6452 27948 6458
rect 27896 6394 27948 6400
rect 28368 6322 28396 7346
rect 28632 7336 28684 7342
rect 28632 7278 28684 7284
rect 27804 6316 27856 6322
rect 27804 6258 27856 6264
rect 28356 6316 28408 6322
rect 28356 6258 28408 6264
rect 28368 6118 28396 6258
rect 28644 6254 28672 7278
rect 28724 7268 28776 7274
rect 28724 7210 28776 7216
rect 28736 6254 28764 7210
rect 28828 6322 28856 8774
rect 28920 7954 28948 12038
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29012 11286 29040 11698
rect 29092 11552 29144 11558
rect 29092 11494 29144 11500
rect 29000 11280 29052 11286
rect 29000 11222 29052 11228
rect 29104 10742 29132 11494
rect 29092 10736 29144 10742
rect 29196 10713 29224 12174
rect 29092 10678 29144 10684
rect 29182 10704 29238 10713
rect 29182 10639 29238 10648
rect 29276 9920 29328 9926
rect 29276 9862 29328 9868
rect 29000 8492 29052 8498
rect 29000 8434 29052 8440
rect 28908 7948 28960 7954
rect 28908 7890 28960 7896
rect 29012 6458 29040 8434
rect 29092 7472 29144 7478
rect 29092 7414 29144 7420
rect 29000 6452 29052 6458
rect 29000 6394 29052 6400
rect 28816 6316 28868 6322
rect 28816 6258 28868 6264
rect 28632 6248 28684 6254
rect 28632 6190 28684 6196
rect 28724 6248 28776 6254
rect 28724 6190 28776 6196
rect 28356 6112 28408 6118
rect 28356 6054 28408 6060
rect 27712 5704 27764 5710
rect 27712 5646 27764 5652
rect 27344 5636 27396 5642
rect 27344 5578 27396 5584
rect 29000 5092 29052 5098
rect 29000 5034 29052 5040
rect 26608 4616 26660 4622
rect 26608 4558 26660 4564
rect 25320 4548 25372 4554
rect 25320 4490 25372 4496
rect 23112 4480 23164 4486
rect 23112 4422 23164 4428
rect 25776 3836 26084 3856
rect 25776 3834 25782 3836
rect 25838 3834 25862 3836
rect 25918 3834 25942 3836
rect 25998 3834 26022 3836
rect 26078 3834 26084 3836
rect 25838 3782 25840 3834
rect 26020 3782 26022 3834
rect 25776 3780 25782 3782
rect 25838 3780 25862 3782
rect 25918 3780 25942 3782
rect 25998 3780 26022 3782
rect 26078 3780 26084 3782
rect 25776 3760 26084 3780
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 20811 3292 21119 3312
rect 20811 3290 20817 3292
rect 20873 3290 20897 3292
rect 20953 3290 20977 3292
rect 21033 3290 21057 3292
rect 21113 3290 21119 3292
rect 20873 3238 20875 3290
rect 21055 3238 21057 3290
rect 20811 3236 20817 3238
rect 20873 3236 20897 3238
rect 20953 3236 20977 3238
rect 21033 3236 21057 3238
rect 21113 3236 21119 3238
rect 20811 3216 21119 3236
rect 25776 2748 26084 2768
rect 25776 2746 25782 2748
rect 25838 2746 25862 2748
rect 25918 2746 25942 2748
rect 25998 2746 26022 2748
rect 26078 2746 26084 2748
rect 25838 2694 25840 2746
rect 26020 2694 26022 2746
rect 25776 2692 25782 2694
rect 25838 2692 25862 2694
rect 25918 2692 25942 2694
rect 25998 2692 26022 2694
rect 26078 2692 26084 2694
rect 25776 2672 26084 2692
rect 29012 2650 29040 5034
rect 29104 3194 29132 7414
rect 29288 7410 29316 9862
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29564 7546 29592 9522
rect 29932 8634 29960 13942
rect 30116 13734 30144 14350
rect 30104 13728 30156 13734
rect 30104 13670 30156 13676
rect 30116 12850 30144 13670
rect 30104 12844 30156 12850
rect 30104 12786 30156 12792
rect 30012 12640 30064 12646
rect 30012 12582 30064 12588
rect 30024 9450 30052 12582
rect 30196 12232 30248 12238
rect 30196 12174 30248 12180
rect 30104 11552 30156 11558
rect 30104 11494 30156 11500
rect 30116 11218 30144 11494
rect 30104 11212 30156 11218
rect 30104 11154 30156 11160
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 30012 9444 30064 9450
rect 30012 9386 30064 9392
rect 29920 8628 29972 8634
rect 29920 8570 29972 8576
rect 29552 7540 29604 7546
rect 29552 7482 29604 7488
rect 29276 7404 29328 7410
rect 29276 7346 29328 7352
rect 29932 6322 29960 8570
rect 30024 7410 30052 9386
rect 30116 9217 30144 9998
rect 30208 9897 30236 12174
rect 30194 9888 30250 9897
rect 30194 9823 30250 9832
rect 30102 9208 30158 9217
rect 30102 9143 30158 9152
rect 30104 8968 30156 8974
rect 30104 8910 30156 8916
rect 30116 8401 30144 8910
rect 30102 8392 30158 8401
rect 30102 8327 30158 8336
rect 30104 7880 30156 7886
rect 30104 7822 30156 7828
rect 30116 7721 30144 7822
rect 30102 7712 30158 7721
rect 30102 7647 30158 7656
rect 30012 7404 30064 7410
rect 30012 7346 30064 7352
rect 30102 6896 30158 6905
rect 30102 6831 30158 6840
rect 30116 6798 30144 6831
rect 30104 6792 30156 6798
rect 30104 6734 30156 6740
rect 29920 6316 29972 6322
rect 29920 6258 29972 6264
rect 30104 6316 30156 6322
rect 30104 6258 30156 6264
rect 30116 6225 30144 6258
rect 30102 6216 30158 6225
rect 30102 6151 30158 6160
rect 29920 5636 29972 5642
rect 29920 5578 29972 5584
rect 29184 5568 29236 5574
rect 29932 5545 29960 5578
rect 30012 5568 30064 5574
rect 29184 5510 29236 5516
rect 29918 5536 29974 5545
rect 29196 4010 29224 5510
rect 30012 5510 30064 5516
rect 29918 5471 29974 5480
rect 30024 5302 30052 5510
rect 30012 5296 30064 5302
rect 30012 5238 30064 5244
rect 29920 5228 29972 5234
rect 29920 5170 29972 5176
rect 29932 4729 29960 5170
rect 30012 5024 30064 5030
rect 30012 4966 30064 4972
rect 30024 4758 30052 4966
rect 30012 4752 30064 4758
rect 29918 4720 29974 4729
rect 30012 4694 30064 4700
rect 29918 4655 29974 4664
rect 29920 4548 29972 4554
rect 29920 4490 29972 4496
rect 29932 4049 29960 4490
rect 30012 4140 30064 4146
rect 30012 4082 30064 4088
rect 29918 4040 29974 4049
rect 29184 4004 29236 4010
rect 29918 3975 29974 3984
rect 29184 3946 29236 3952
rect 29828 3528 29880 3534
rect 29828 3470 29880 3476
rect 29092 3188 29144 3194
rect 29092 3130 29144 3136
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 29840 2553 29868 3470
rect 30024 3233 30052 4082
rect 30010 3224 30066 3233
rect 30010 3159 30066 3168
rect 29920 3052 29972 3058
rect 29920 2994 29972 3000
rect 29826 2544 29882 2553
rect 29826 2479 29882 2488
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1596 1057 1624 2246
rect 10880 2204 11188 2224
rect 10880 2202 10886 2204
rect 10942 2202 10966 2204
rect 11022 2202 11046 2204
rect 11102 2202 11126 2204
rect 11182 2202 11188 2204
rect 10942 2150 10944 2202
rect 11124 2150 11126 2202
rect 10880 2148 10886 2150
rect 10942 2148 10966 2150
rect 11022 2148 11046 2150
rect 11102 2148 11126 2150
rect 11182 2148 11188 2150
rect 10880 2128 11188 2148
rect 20811 2204 21119 2224
rect 20811 2202 20817 2204
rect 20873 2202 20897 2204
rect 20953 2202 20977 2204
rect 21033 2202 21057 2204
rect 21113 2202 21119 2204
rect 20873 2150 20875 2202
rect 21055 2150 21057 2202
rect 20811 2148 20817 2150
rect 20873 2148 20897 2150
rect 20953 2148 20977 2150
rect 21033 2148 21057 2150
rect 21113 2148 21119 2150
rect 20811 2128 21119 2148
rect 28736 1057 28764 2382
rect 29736 2372 29788 2378
rect 29736 2314 29788 2320
rect 1582 1048 1638 1057
rect 1582 983 1638 992
rect 28722 1048 28778 1057
rect 28722 983 28778 992
rect 29748 377 29776 2314
rect 29932 1737 29960 2994
rect 29918 1728 29974 1737
rect 29918 1663 29974 1672
rect 29734 368 29790 377
rect 29734 303 29790 312
<< via2 >>
rect 1582 44920 1638 44976
rect 2778 46960 2834 47016
rect 1582 42880 1638 42936
rect 1582 40976 1638 41032
rect 1582 38936 1638 38992
rect 1582 36896 1638 36952
rect 1582 35028 1584 35048
rect 1584 35028 1636 35048
rect 1636 35028 1638 35048
rect 1582 34992 1638 35028
rect 1582 32952 1638 33008
rect 1398 30912 1454 30968
rect 1582 28872 1638 28928
rect 1582 26968 1638 27024
rect 1582 24928 1638 24984
rect 1582 22924 1584 22944
rect 1584 22924 1636 22944
rect 1636 22924 1638 22944
rect 1582 22888 1638 22924
rect 1582 20984 1638 21040
rect 1582 18944 1638 19000
rect 1582 16940 1584 16960
rect 1584 16940 1636 16960
rect 1636 16940 1638 16960
rect 1582 16904 1638 16940
rect 1582 14884 1638 14920
rect 1582 14864 1584 14884
rect 1584 14864 1636 14884
rect 1636 14864 1638 14884
rect 1582 12960 1638 13016
rect 1582 10956 1584 10976
rect 1584 10956 1636 10976
rect 1636 10956 1638 10976
rect 1582 10920 1638 10956
rect 1582 8880 1638 8936
rect 1582 6976 1638 7032
rect 1582 4972 1584 4992
rect 1584 4972 1636 4992
rect 1636 4972 1638 4992
rect 1582 4936 1638 4972
rect 5921 45178 5977 45180
rect 6001 45178 6057 45180
rect 6081 45178 6137 45180
rect 6161 45178 6217 45180
rect 5921 45126 5967 45178
rect 5967 45126 5977 45178
rect 6001 45126 6031 45178
rect 6031 45126 6043 45178
rect 6043 45126 6057 45178
rect 6081 45126 6095 45178
rect 6095 45126 6107 45178
rect 6107 45126 6137 45178
rect 6161 45126 6171 45178
rect 6171 45126 6217 45178
rect 5921 45124 5977 45126
rect 6001 45124 6057 45126
rect 6081 45124 6137 45126
rect 6161 45124 6217 45126
rect 5921 44090 5977 44092
rect 6001 44090 6057 44092
rect 6081 44090 6137 44092
rect 6161 44090 6217 44092
rect 5921 44038 5967 44090
rect 5967 44038 5977 44090
rect 6001 44038 6031 44090
rect 6031 44038 6043 44090
rect 6043 44038 6057 44090
rect 6081 44038 6095 44090
rect 6095 44038 6107 44090
rect 6107 44038 6137 44090
rect 6161 44038 6171 44090
rect 6171 44038 6217 44090
rect 5921 44036 5977 44038
rect 6001 44036 6057 44038
rect 6081 44036 6137 44038
rect 6161 44036 6217 44038
rect 5921 43002 5977 43004
rect 6001 43002 6057 43004
rect 6081 43002 6137 43004
rect 6161 43002 6217 43004
rect 5921 42950 5967 43002
rect 5967 42950 5977 43002
rect 6001 42950 6031 43002
rect 6031 42950 6043 43002
rect 6043 42950 6057 43002
rect 6081 42950 6095 43002
rect 6095 42950 6107 43002
rect 6107 42950 6137 43002
rect 6161 42950 6171 43002
rect 6171 42950 6217 43002
rect 5921 42948 5977 42950
rect 6001 42948 6057 42950
rect 6081 42948 6137 42950
rect 6161 42948 6217 42950
rect 5921 41914 5977 41916
rect 6001 41914 6057 41916
rect 6081 41914 6137 41916
rect 6161 41914 6217 41916
rect 5921 41862 5967 41914
rect 5967 41862 5977 41914
rect 6001 41862 6031 41914
rect 6031 41862 6043 41914
rect 6043 41862 6057 41914
rect 6081 41862 6095 41914
rect 6095 41862 6107 41914
rect 6107 41862 6137 41914
rect 6161 41862 6171 41914
rect 6171 41862 6217 41914
rect 5921 41860 5977 41862
rect 6001 41860 6057 41862
rect 6081 41860 6137 41862
rect 6161 41860 6217 41862
rect 5921 40826 5977 40828
rect 6001 40826 6057 40828
rect 6081 40826 6137 40828
rect 6161 40826 6217 40828
rect 5921 40774 5967 40826
rect 5967 40774 5977 40826
rect 6001 40774 6031 40826
rect 6031 40774 6043 40826
rect 6043 40774 6057 40826
rect 6081 40774 6095 40826
rect 6095 40774 6107 40826
rect 6107 40774 6137 40826
rect 6161 40774 6171 40826
rect 6171 40774 6217 40826
rect 5921 40772 5977 40774
rect 6001 40772 6057 40774
rect 6081 40772 6137 40774
rect 6161 40772 6217 40774
rect 5921 39738 5977 39740
rect 6001 39738 6057 39740
rect 6081 39738 6137 39740
rect 6161 39738 6217 39740
rect 5921 39686 5967 39738
rect 5967 39686 5977 39738
rect 6001 39686 6031 39738
rect 6031 39686 6043 39738
rect 6043 39686 6057 39738
rect 6081 39686 6095 39738
rect 6095 39686 6107 39738
rect 6107 39686 6137 39738
rect 6161 39686 6171 39738
rect 6171 39686 6217 39738
rect 5921 39684 5977 39686
rect 6001 39684 6057 39686
rect 6081 39684 6137 39686
rect 6161 39684 6217 39686
rect 5921 38650 5977 38652
rect 6001 38650 6057 38652
rect 6081 38650 6137 38652
rect 6161 38650 6217 38652
rect 5921 38598 5967 38650
rect 5967 38598 5977 38650
rect 6001 38598 6031 38650
rect 6031 38598 6043 38650
rect 6043 38598 6057 38650
rect 6081 38598 6095 38650
rect 6095 38598 6107 38650
rect 6107 38598 6137 38650
rect 6161 38598 6171 38650
rect 6171 38598 6217 38650
rect 5921 38596 5977 38598
rect 6001 38596 6057 38598
rect 6081 38596 6137 38598
rect 6161 38596 6217 38598
rect 5921 37562 5977 37564
rect 6001 37562 6057 37564
rect 6081 37562 6137 37564
rect 6161 37562 6217 37564
rect 5921 37510 5967 37562
rect 5967 37510 5977 37562
rect 6001 37510 6031 37562
rect 6031 37510 6043 37562
rect 6043 37510 6057 37562
rect 6081 37510 6095 37562
rect 6095 37510 6107 37562
rect 6107 37510 6137 37562
rect 6161 37510 6171 37562
rect 6171 37510 6217 37562
rect 5921 37508 5977 37510
rect 6001 37508 6057 37510
rect 6081 37508 6137 37510
rect 6161 37508 6217 37510
rect 5921 36474 5977 36476
rect 6001 36474 6057 36476
rect 6081 36474 6137 36476
rect 6161 36474 6217 36476
rect 5921 36422 5967 36474
rect 5967 36422 5977 36474
rect 6001 36422 6031 36474
rect 6031 36422 6043 36474
rect 6043 36422 6057 36474
rect 6081 36422 6095 36474
rect 6095 36422 6107 36474
rect 6107 36422 6137 36474
rect 6161 36422 6171 36474
rect 6171 36422 6217 36474
rect 5921 36420 5977 36422
rect 6001 36420 6057 36422
rect 6081 36420 6137 36422
rect 6161 36420 6217 36422
rect 5921 35386 5977 35388
rect 6001 35386 6057 35388
rect 6081 35386 6137 35388
rect 6161 35386 6217 35388
rect 5921 35334 5967 35386
rect 5967 35334 5977 35386
rect 6001 35334 6031 35386
rect 6031 35334 6043 35386
rect 6043 35334 6057 35386
rect 6081 35334 6095 35386
rect 6095 35334 6107 35386
rect 6107 35334 6137 35386
rect 6161 35334 6171 35386
rect 6171 35334 6217 35386
rect 5921 35332 5977 35334
rect 6001 35332 6057 35334
rect 6081 35332 6137 35334
rect 6161 35332 6217 35334
rect 5921 34298 5977 34300
rect 6001 34298 6057 34300
rect 6081 34298 6137 34300
rect 6161 34298 6217 34300
rect 5921 34246 5967 34298
rect 5967 34246 5977 34298
rect 6001 34246 6031 34298
rect 6031 34246 6043 34298
rect 6043 34246 6057 34298
rect 6081 34246 6095 34298
rect 6095 34246 6107 34298
rect 6107 34246 6137 34298
rect 6161 34246 6171 34298
rect 6171 34246 6217 34298
rect 5921 34244 5977 34246
rect 6001 34244 6057 34246
rect 6081 34244 6137 34246
rect 6161 34244 6217 34246
rect 5921 33210 5977 33212
rect 6001 33210 6057 33212
rect 6081 33210 6137 33212
rect 6161 33210 6217 33212
rect 5921 33158 5967 33210
rect 5967 33158 5977 33210
rect 6001 33158 6031 33210
rect 6031 33158 6043 33210
rect 6043 33158 6057 33210
rect 6081 33158 6095 33210
rect 6095 33158 6107 33210
rect 6107 33158 6137 33210
rect 6161 33158 6171 33210
rect 6171 33158 6217 33210
rect 5921 33156 5977 33158
rect 6001 33156 6057 33158
rect 6081 33156 6137 33158
rect 6161 33156 6217 33158
rect 5921 32122 5977 32124
rect 6001 32122 6057 32124
rect 6081 32122 6137 32124
rect 6161 32122 6217 32124
rect 5921 32070 5967 32122
rect 5967 32070 5977 32122
rect 6001 32070 6031 32122
rect 6031 32070 6043 32122
rect 6043 32070 6057 32122
rect 6081 32070 6095 32122
rect 6095 32070 6107 32122
rect 6107 32070 6137 32122
rect 6161 32070 6171 32122
rect 6171 32070 6217 32122
rect 5921 32068 5977 32070
rect 6001 32068 6057 32070
rect 6081 32068 6137 32070
rect 6161 32068 6217 32070
rect 5921 31034 5977 31036
rect 6001 31034 6057 31036
rect 6081 31034 6137 31036
rect 6161 31034 6217 31036
rect 5921 30982 5967 31034
rect 5967 30982 5977 31034
rect 6001 30982 6031 31034
rect 6031 30982 6043 31034
rect 6043 30982 6057 31034
rect 6081 30982 6095 31034
rect 6095 30982 6107 31034
rect 6107 30982 6137 31034
rect 6161 30982 6171 31034
rect 6171 30982 6217 31034
rect 5921 30980 5977 30982
rect 6001 30980 6057 30982
rect 6081 30980 6137 30982
rect 6161 30980 6217 30982
rect 5921 29946 5977 29948
rect 6001 29946 6057 29948
rect 6081 29946 6137 29948
rect 6161 29946 6217 29948
rect 5921 29894 5967 29946
rect 5967 29894 5977 29946
rect 6001 29894 6031 29946
rect 6031 29894 6043 29946
rect 6043 29894 6057 29946
rect 6081 29894 6095 29946
rect 6095 29894 6107 29946
rect 6107 29894 6137 29946
rect 6161 29894 6171 29946
rect 6171 29894 6217 29946
rect 5921 29892 5977 29894
rect 6001 29892 6057 29894
rect 6081 29892 6137 29894
rect 6161 29892 6217 29894
rect 5921 28858 5977 28860
rect 6001 28858 6057 28860
rect 6081 28858 6137 28860
rect 6161 28858 6217 28860
rect 5921 28806 5967 28858
rect 5967 28806 5977 28858
rect 6001 28806 6031 28858
rect 6031 28806 6043 28858
rect 6043 28806 6057 28858
rect 6081 28806 6095 28858
rect 6095 28806 6107 28858
rect 6107 28806 6137 28858
rect 6161 28806 6171 28858
rect 6171 28806 6217 28858
rect 5921 28804 5977 28806
rect 6001 28804 6057 28806
rect 6081 28804 6137 28806
rect 6161 28804 6217 28806
rect 10886 45722 10942 45724
rect 10966 45722 11022 45724
rect 11046 45722 11102 45724
rect 11126 45722 11182 45724
rect 10886 45670 10932 45722
rect 10932 45670 10942 45722
rect 10966 45670 10996 45722
rect 10996 45670 11008 45722
rect 11008 45670 11022 45722
rect 11046 45670 11060 45722
rect 11060 45670 11072 45722
rect 11072 45670 11102 45722
rect 11126 45670 11136 45722
rect 11136 45670 11182 45722
rect 10886 45668 10942 45670
rect 10966 45668 11022 45670
rect 11046 45668 11102 45670
rect 11126 45668 11182 45670
rect 10886 44634 10942 44636
rect 10966 44634 11022 44636
rect 11046 44634 11102 44636
rect 11126 44634 11182 44636
rect 10886 44582 10932 44634
rect 10932 44582 10942 44634
rect 10966 44582 10996 44634
rect 10996 44582 11008 44634
rect 11008 44582 11022 44634
rect 11046 44582 11060 44634
rect 11060 44582 11072 44634
rect 11072 44582 11102 44634
rect 11126 44582 11136 44634
rect 11136 44582 11182 44634
rect 10886 44580 10942 44582
rect 10966 44580 11022 44582
rect 11046 44580 11102 44582
rect 11126 44580 11182 44582
rect 10886 43546 10942 43548
rect 10966 43546 11022 43548
rect 11046 43546 11102 43548
rect 11126 43546 11182 43548
rect 10886 43494 10932 43546
rect 10932 43494 10942 43546
rect 10966 43494 10996 43546
rect 10996 43494 11008 43546
rect 11008 43494 11022 43546
rect 11046 43494 11060 43546
rect 11060 43494 11072 43546
rect 11072 43494 11102 43546
rect 11126 43494 11136 43546
rect 11136 43494 11182 43546
rect 10886 43492 10942 43494
rect 10966 43492 11022 43494
rect 11046 43492 11102 43494
rect 11126 43492 11182 43494
rect 10886 42458 10942 42460
rect 10966 42458 11022 42460
rect 11046 42458 11102 42460
rect 11126 42458 11182 42460
rect 10886 42406 10932 42458
rect 10932 42406 10942 42458
rect 10966 42406 10996 42458
rect 10996 42406 11008 42458
rect 11008 42406 11022 42458
rect 11046 42406 11060 42458
rect 11060 42406 11072 42458
rect 11072 42406 11102 42458
rect 11126 42406 11136 42458
rect 11136 42406 11182 42458
rect 10886 42404 10942 42406
rect 10966 42404 11022 42406
rect 11046 42404 11102 42406
rect 11126 42404 11182 42406
rect 10886 41370 10942 41372
rect 10966 41370 11022 41372
rect 11046 41370 11102 41372
rect 11126 41370 11182 41372
rect 10886 41318 10932 41370
rect 10932 41318 10942 41370
rect 10966 41318 10996 41370
rect 10996 41318 11008 41370
rect 11008 41318 11022 41370
rect 11046 41318 11060 41370
rect 11060 41318 11072 41370
rect 11072 41318 11102 41370
rect 11126 41318 11136 41370
rect 11136 41318 11182 41370
rect 10886 41316 10942 41318
rect 10966 41316 11022 41318
rect 11046 41316 11102 41318
rect 11126 41316 11182 41318
rect 10886 40282 10942 40284
rect 10966 40282 11022 40284
rect 11046 40282 11102 40284
rect 11126 40282 11182 40284
rect 10886 40230 10932 40282
rect 10932 40230 10942 40282
rect 10966 40230 10996 40282
rect 10996 40230 11008 40282
rect 11008 40230 11022 40282
rect 11046 40230 11060 40282
rect 11060 40230 11072 40282
rect 11072 40230 11102 40282
rect 11126 40230 11136 40282
rect 11136 40230 11182 40282
rect 10886 40228 10942 40230
rect 10966 40228 11022 40230
rect 11046 40228 11102 40230
rect 11126 40228 11182 40230
rect 10886 39194 10942 39196
rect 10966 39194 11022 39196
rect 11046 39194 11102 39196
rect 11126 39194 11182 39196
rect 10886 39142 10932 39194
rect 10932 39142 10942 39194
rect 10966 39142 10996 39194
rect 10996 39142 11008 39194
rect 11008 39142 11022 39194
rect 11046 39142 11060 39194
rect 11060 39142 11072 39194
rect 11072 39142 11102 39194
rect 11126 39142 11136 39194
rect 11136 39142 11182 39194
rect 10886 39140 10942 39142
rect 10966 39140 11022 39142
rect 11046 39140 11102 39142
rect 11126 39140 11182 39142
rect 10886 38106 10942 38108
rect 10966 38106 11022 38108
rect 11046 38106 11102 38108
rect 11126 38106 11182 38108
rect 10886 38054 10932 38106
rect 10932 38054 10942 38106
rect 10966 38054 10996 38106
rect 10996 38054 11008 38106
rect 11008 38054 11022 38106
rect 11046 38054 11060 38106
rect 11060 38054 11072 38106
rect 11072 38054 11102 38106
rect 11126 38054 11136 38106
rect 11136 38054 11182 38106
rect 10886 38052 10942 38054
rect 10966 38052 11022 38054
rect 11046 38052 11102 38054
rect 11126 38052 11182 38054
rect 9954 30096 10010 30152
rect 5921 27770 5977 27772
rect 6001 27770 6057 27772
rect 6081 27770 6137 27772
rect 6161 27770 6217 27772
rect 5921 27718 5967 27770
rect 5967 27718 5977 27770
rect 6001 27718 6031 27770
rect 6031 27718 6043 27770
rect 6043 27718 6057 27770
rect 6081 27718 6095 27770
rect 6095 27718 6107 27770
rect 6107 27718 6137 27770
rect 6161 27718 6171 27770
rect 6171 27718 6217 27770
rect 5921 27716 5977 27718
rect 6001 27716 6057 27718
rect 6081 27716 6137 27718
rect 6161 27716 6217 27718
rect 5921 26682 5977 26684
rect 6001 26682 6057 26684
rect 6081 26682 6137 26684
rect 6161 26682 6217 26684
rect 5921 26630 5967 26682
rect 5967 26630 5977 26682
rect 6001 26630 6031 26682
rect 6031 26630 6043 26682
rect 6043 26630 6057 26682
rect 6081 26630 6095 26682
rect 6095 26630 6107 26682
rect 6107 26630 6137 26682
rect 6161 26630 6171 26682
rect 6171 26630 6217 26682
rect 5921 26628 5977 26630
rect 6001 26628 6057 26630
rect 6081 26628 6137 26630
rect 6161 26628 6217 26630
rect 5921 25594 5977 25596
rect 6001 25594 6057 25596
rect 6081 25594 6137 25596
rect 6161 25594 6217 25596
rect 5921 25542 5967 25594
rect 5967 25542 5977 25594
rect 6001 25542 6031 25594
rect 6031 25542 6043 25594
rect 6043 25542 6057 25594
rect 6081 25542 6095 25594
rect 6095 25542 6107 25594
rect 6107 25542 6137 25594
rect 6161 25542 6171 25594
rect 6171 25542 6217 25594
rect 5921 25540 5977 25542
rect 6001 25540 6057 25542
rect 6081 25540 6137 25542
rect 6161 25540 6217 25542
rect 5921 24506 5977 24508
rect 6001 24506 6057 24508
rect 6081 24506 6137 24508
rect 6161 24506 6217 24508
rect 5921 24454 5967 24506
rect 5967 24454 5977 24506
rect 6001 24454 6031 24506
rect 6031 24454 6043 24506
rect 6043 24454 6057 24506
rect 6081 24454 6095 24506
rect 6095 24454 6107 24506
rect 6107 24454 6137 24506
rect 6161 24454 6171 24506
rect 6171 24454 6217 24506
rect 5921 24452 5977 24454
rect 6001 24452 6057 24454
rect 6081 24452 6137 24454
rect 6161 24452 6217 24454
rect 5921 23418 5977 23420
rect 6001 23418 6057 23420
rect 6081 23418 6137 23420
rect 6161 23418 6217 23420
rect 5921 23366 5967 23418
rect 5967 23366 5977 23418
rect 6001 23366 6031 23418
rect 6031 23366 6043 23418
rect 6043 23366 6057 23418
rect 6081 23366 6095 23418
rect 6095 23366 6107 23418
rect 6107 23366 6137 23418
rect 6161 23366 6171 23418
rect 6171 23366 6217 23418
rect 5921 23364 5977 23366
rect 6001 23364 6057 23366
rect 6081 23364 6137 23366
rect 6161 23364 6217 23366
rect 5921 22330 5977 22332
rect 6001 22330 6057 22332
rect 6081 22330 6137 22332
rect 6161 22330 6217 22332
rect 5921 22278 5967 22330
rect 5967 22278 5977 22330
rect 6001 22278 6031 22330
rect 6031 22278 6043 22330
rect 6043 22278 6057 22330
rect 6081 22278 6095 22330
rect 6095 22278 6107 22330
rect 6107 22278 6137 22330
rect 6161 22278 6171 22330
rect 6171 22278 6217 22330
rect 5921 22276 5977 22278
rect 6001 22276 6057 22278
rect 6081 22276 6137 22278
rect 6161 22276 6217 22278
rect 5921 21242 5977 21244
rect 6001 21242 6057 21244
rect 6081 21242 6137 21244
rect 6161 21242 6217 21244
rect 5921 21190 5967 21242
rect 5967 21190 5977 21242
rect 6001 21190 6031 21242
rect 6031 21190 6043 21242
rect 6043 21190 6057 21242
rect 6081 21190 6095 21242
rect 6095 21190 6107 21242
rect 6107 21190 6137 21242
rect 6161 21190 6171 21242
rect 6171 21190 6217 21242
rect 5921 21188 5977 21190
rect 6001 21188 6057 21190
rect 6081 21188 6137 21190
rect 6161 21188 6217 21190
rect 5921 20154 5977 20156
rect 6001 20154 6057 20156
rect 6081 20154 6137 20156
rect 6161 20154 6217 20156
rect 5921 20102 5967 20154
rect 5967 20102 5977 20154
rect 6001 20102 6031 20154
rect 6031 20102 6043 20154
rect 6043 20102 6057 20154
rect 6081 20102 6095 20154
rect 6095 20102 6107 20154
rect 6107 20102 6137 20154
rect 6161 20102 6171 20154
rect 6171 20102 6217 20154
rect 5921 20100 5977 20102
rect 6001 20100 6057 20102
rect 6081 20100 6137 20102
rect 6161 20100 6217 20102
rect 5921 19066 5977 19068
rect 6001 19066 6057 19068
rect 6081 19066 6137 19068
rect 6161 19066 6217 19068
rect 5921 19014 5967 19066
rect 5967 19014 5977 19066
rect 6001 19014 6031 19066
rect 6031 19014 6043 19066
rect 6043 19014 6057 19066
rect 6081 19014 6095 19066
rect 6095 19014 6107 19066
rect 6107 19014 6137 19066
rect 6161 19014 6171 19066
rect 6171 19014 6217 19066
rect 5921 19012 5977 19014
rect 6001 19012 6057 19014
rect 6081 19012 6137 19014
rect 6161 19012 6217 19014
rect 10230 33940 10232 33960
rect 10232 33940 10284 33960
rect 10284 33940 10286 33960
rect 10230 33904 10286 33940
rect 10414 33904 10470 33960
rect 10886 37018 10942 37020
rect 10966 37018 11022 37020
rect 11046 37018 11102 37020
rect 11126 37018 11182 37020
rect 10886 36966 10932 37018
rect 10932 36966 10942 37018
rect 10966 36966 10996 37018
rect 10996 36966 11008 37018
rect 11008 36966 11022 37018
rect 11046 36966 11060 37018
rect 11060 36966 11072 37018
rect 11072 36966 11102 37018
rect 11126 36966 11136 37018
rect 11136 36966 11182 37018
rect 10886 36964 10942 36966
rect 10966 36964 11022 36966
rect 11046 36964 11102 36966
rect 11126 36964 11182 36966
rect 10886 35930 10942 35932
rect 10966 35930 11022 35932
rect 11046 35930 11102 35932
rect 11126 35930 11182 35932
rect 10886 35878 10932 35930
rect 10932 35878 10942 35930
rect 10966 35878 10996 35930
rect 10996 35878 11008 35930
rect 11008 35878 11022 35930
rect 11046 35878 11060 35930
rect 11060 35878 11072 35930
rect 11072 35878 11102 35930
rect 11126 35878 11136 35930
rect 11136 35878 11182 35930
rect 10886 35876 10942 35878
rect 10966 35876 11022 35878
rect 11046 35876 11102 35878
rect 11126 35876 11182 35878
rect 10886 34842 10942 34844
rect 10966 34842 11022 34844
rect 11046 34842 11102 34844
rect 11126 34842 11182 34844
rect 10886 34790 10932 34842
rect 10932 34790 10942 34842
rect 10966 34790 10996 34842
rect 10996 34790 11008 34842
rect 11008 34790 11022 34842
rect 11046 34790 11060 34842
rect 11060 34790 11072 34842
rect 11072 34790 11102 34842
rect 11126 34790 11136 34842
rect 11136 34790 11182 34842
rect 10886 34788 10942 34790
rect 10966 34788 11022 34790
rect 11046 34788 11102 34790
rect 11126 34788 11182 34790
rect 13542 44240 13598 44296
rect 14002 43832 14058 43888
rect 14278 44920 14334 44976
rect 14186 44140 14188 44160
rect 14188 44140 14240 44160
rect 14240 44140 14242 44160
rect 14186 44104 14242 44140
rect 14646 44804 14702 44840
rect 14646 44784 14648 44804
rect 14648 44784 14700 44804
rect 14700 44784 14702 44804
rect 10886 33754 10942 33756
rect 10966 33754 11022 33756
rect 11046 33754 11102 33756
rect 11126 33754 11182 33756
rect 10886 33702 10932 33754
rect 10932 33702 10942 33754
rect 10966 33702 10996 33754
rect 10996 33702 11008 33754
rect 11008 33702 11022 33754
rect 11046 33702 11060 33754
rect 11060 33702 11072 33754
rect 11072 33702 11102 33754
rect 11126 33702 11136 33754
rect 11136 33702 11182 33754
rect 10886 33700 10942 33702
rect 10966 33700 11022 33702
rect 11046 33700 11102 33702
rect 11126 33700 11182 33702
rect 10230 29552 10286 29608
rect 10886 32666 10942 32668
rect 10966 32666 11022 32668
rect 11046 32666 11102 32668
rect 11126 32666 11182 32668
rect 10886 32614 10932 32666
rect 10932 32614 10942 32666
rect 10966 32614 10996 32666
rect 10996 32614 11008 32666
rect 11008 32614 11022 32666
rect 11046 32614 11060 32666
rect 11060 32614 11072 32666
rect 11072 32614 11102 32666
rect 11126 32614 11136 32666
rect 11136 32614 11182 32666
rect 10886 32612 10942 32614
rect 10966 32612 11022 32614
rect 11046 32612 11102 32614
rect 11126 32612 11182 32614
rect 10886 31578 10942 31580
rect 10966 31578 11022 31580
rect 11046 31578 11102 31580
rect 11126 31578 11182 31580
rect 10886 31526 10932 31578
rect 10932 31526 10942 31578
rect 10966 31526 10996 31578
rect 10996 31526 11008 31578
rect 11008 31526 11022 31578
rect 11046 31526 11060 31578
rect 11060 31526 11072 31578
rect 11072 31526 11102 31578
rect 11126 31526 11136 31578
rect 11136 31526 11182 31578
rect 10886 31524 10942 31526
rect 10966 31524 11022 31526
rect 11046 31524 11102 31526
rect 11126 31524 11182 31526
rect 10886 30490 10942 30492
rect 10966 30490 11022 30492
rect 11046 30490 11102 30492
rect 11126 30490 11182 30492
rect 10886 30438 10932 30490
rect 10932 30438 10942 30490
rect 10966 30438 10996 30490
rect 10996 30438 11008 30490
rect 11008 30438 11022 30490
rect 11046 30438 11060 30490
rect 11060 30438 11072 30490
rect 11072 30438 11102 30490
rect 11126 30438 11136 30490
rect 11136 30438 11182 30490
rect 10886 30436 10942 30438
rect 10966 30436 11022 30438
rect 11046 30436 11102 30438
rect 11126 30436 11182 30438
rect 10886 29402 10942 29404
rect 10966 29402 11022 29404
rect 11046 29402 11102 29404
rect 11126 29402 11182 29404
rect 10886 29350 10932 29402
rect 10932 29350 10942 29402
rect 10966 29350 10996 29402
rect 10996 29350 11008 29402
rect 11008 29350 11022 29402
rect 11046 29350 11060 29402
rect 11060 29350 11072 29402
rect 11072 29350 11102 29402
rect 11126 29350 11136 29402
rect 11136 29350 11182 29402
rect 10886 29348 10942 29350
rect 10966 29348 11022 29350
rect 11046 29348 11102 29350
rect 11126 29348 11182 29350
rect 11150 29144 11206 29200
rect 10138 24656 10194 24712
rect 9678 23160 9734 23216
rect 10046 23160 10102 23216
rect 5921 17978 5977 17980
rect 6001 17978 6057 17980
rect 6081 17978 6137 17980
rect 6161 17978 6217 17980
rect 5921 17926 5967 17978
rect 5967 17926 5977 17978
rect 6001 17926 6031 17978
rect 6031 17926 6043 17978
rect 6043 17926 6057 17978
rect 6081 17926 6095 17978
rect 6095 17926 6107 17978
rect 6107 17926 6137 17978
rect 6161 17926 6171 17978
rect 6171 17926 6217 17978
rect 5921 17924 5977 17926
rect 6001 17924 6057 17926
rect 6081 17924 6137 17926
rect 6161 17924 6217 17926
rect 10046 21392 10102 21448
rect 9954 18808 10010 18864
rect 5921 16890 5977 16892
rect 6001 16890 6057 16892
rect 6081 16890 6137 16892
rect 6161 16890 6217 16892
rect 5921 16838 5967 16890
rect 5967 16838 5977 16890
rect 6001 16838 6031 16890
rect 6031 16838 6043 16890
rect 6043 16838 6057 16890
rect 6081 16838 6095 16890
rect 6095 16838 6107 16890
rect 6107 16838 6137 16890
rect 6161 16838 6171 16890
rect 6171 16838 6217 16890
rect 5921 16836 5977 16838
rect 6001 16836 6057 16838
rect 6081 16836 6137 16838
rect 6161 16836 6217 16838
rect 5921 15802 5977 15804
rect 6001 15802 6057 15804
rect 6081 15802 6137 15804
rect 6161 15802 6217 15804
rect 5921 15750 5967 15802
rect 5967 15750 5977 15802
rect 6001 15750 6031 15802
rect 6031 15750 6043 15802
rect 6043 15750 6057 15802
rect 6081 15750 6095 15802
rect 6095 15750 6107 15802
rect 6107 15750 6137 15802
rect 6161 15750 6171 15802
rect 6171 15750 6217 15802
rect 5921 15748 5977 15750
rect 6001 15748 6057 15750
rect 6081 15748 6137 15750
rect 6161 15748 6217 15750
rect 5921 14714 5977 14716
rect 6001 14714 6057 14716
rect 6081 14714 6137 14716
rect 6161 14714 6217 14716
rect 5921 14662 5967 14714
rect 5967 14662 5977 14714
rect 6001 14662 6031 14714
rect 6031 14662 6043 14714
rect 6043 14662 6057 14714
rect 6081 14662 6095 14714
rect 6095 14662 6107 14714
rect 6107 14662 6137 14714
rect 6161 14662 6171 14714
rect 6171 14662 6217 14714
rect 5921 14660 5977 14662
rect 6001 14660 6057 14662
rect 6081 14660 6137 14662
rect 6161 14660 6217 14662
rect 5921 13626 5977 13628
rect 6001 13626 6057 13628
rect 6081 13626 6137 13628
rect 6161 13626 6217 13628
rect 5921 13574 5967 13626
rect 5967 13574 5977 13626
rect 6001 13574 6031 13626
rect 6031 13574 6043 13626
rect 6043 13574 6057 13626
rect 6081 13574 6095 13626
rect 6095 13574 6107 13626
rect 6107 13574 6137 13626
rect 6161 13574 6171 13626
rect 6171 13574 6217 13626
rect 5921 13572 5977 13574
rect 6001 13572 6057 13574
rect 6081 13572 6137 13574
rect 6161 13572 6217 13574
rect 5921 12538 5977 12540
rect 6001 12538 6057 12540
rect 6081 12538 6137 12540
rect 6161 12538 6217 12540
rect 5921 12486 5967 12538
rect 5967 12486 5977 12538
rect 6001 12486 6031 12538
rect 6031 12486 6043 12538
rect 6043 12486 6057 12538
rect 6081 12486 6095 12538
rect 6095 12486 6107 12538
rect 6107 12486 6137 12538
rect 6161 12486 6171 12538
rect 6171 12486 6217 12538
rect 5921 12484 5977 12486
rect 6001 12484 6057 12486
rect 6081 12484 6137 12486
rect 6161 12484 6217 12486
rect 5921 11450 5977 11452
rect 6001 11450 6057 11452
rect 6081 11450 6137 11452
rect 6161 11450 6217 11452
rect 5921 11398 5967 11450
rect 5967 11398 5977 11450
rect 6001 11398 6031 11450
rect 6031 11398 6043 11450
rect 6043 11398 6057 11450
rect 6081 11398 6095 11450
rect 6095 11398 6107 11450
rect 6107 11398 6137 11450
rect 6161 11398 6171 11450
rect 6171 11398 6217 11450
rect 5921 11396 5977 11398
rect 6001 11396 6057 11398
rect 6081 11396 6137 11398
rect 6161 11396 6217 11398
rect 5921 10362 5977 10364
rect 6001 10362 6057 10364
rect 6081 10362 6137 10364
rect 6161 10362 6217 10364
rect 5921 10310 5967 10362
rect 5967 10310 5977 10362
rect 6001 10310 6031 10362
rect 6031 10310 6043 10362
rect 6043 10310 6057 10362
rect 6081 10310 6095 10362
rect 6095 10310 6107 10362
rect 6107 10310 6137 10362
rect 6161 10310 6171 10362
rect 6171 10310 6217 10362
rect 5921 10308 5977 10310
rect 6001 10308 6057 10310
rect 6081 10308 6137 10310
rect 6161 10308 6217 10310
rect 5921 9274 5977 9276
rect 6001 9274 6057 9276
rect 6081 9274 6137 9276
rect 6161 9274 6217 9276
rect 5921 9222 5967 9274
rect 5967 9222 5977 9274
rect 6001 9222 6031 9274
rect 6031 9222 6043 9274
rect 6043 9222 6057 9274
rect 6081 9222 6095 9274
rect 6095 9222 6107 9274
rect 6107 9222 6137 9274
rect 6161 9222 6171 9274
rect 6171 9222 6217 9274
rect 5921 9220 5977 9222
rect 6001 9220 6057 9222
rect 6081 9220 6137 9222
rect 6161 9220 6217 9222
rect 5921 8186 5977 8188
rect 6001 8186 6057 8188
rect 6081 8186 6137 8188
rect 6161 8186 6217 8188
rect 5921 8134 5967 8186
rect 5967 8134 5977 8186
rect 6001 8134 6031 8186
rect 6031 8134 6043 8186
rect 6043 8134 6057 8186
rect 6081 8134 6095 8186
rect 6095 8134 6107 8186
rect 6107 8134 6137 8186
rect 6161 8134 6171 8186
rect 6171 8134 6217 8186
rect 5921 8132 5977 8134
rect 6001 8132 6057 8134
rect 6081 8132 6137 8134
rect 6161 8132 6217 8134
rect 5921 7098 5977 7100
rect 6001 7098 6057 7100
rect 6081 7098 6137 7100
rect 6161 7098 6217 7100
rect 5921 7046 5967 7098
rect 5967 7046 5977 7098
rect 6001 7046 6031 7098
rect 6031 7046 6043 7098
rect 6043 7046 6057 7098
rect 6081 7046 6095 7098
rect 6095 7046 6107 7098
rect 6107 7046 6137 7098
rect 6161 7046 6171 7098
rect 6171 7046 6217 7098
rect 5921 7044 5977 7046
rect 6001 7044 6057 7046
rect 6081 7044 6137 7046
rect 6161 7044 6217 7046
rect 5921 6010 5977 6012
rect 6001 6010 6057 6012
rect 6081 6010 6137 6012
rect 6161 6010 6217 6012
rect 5921 5958 5967 6010
rect 5967 5958 5977 6010
rect 6001 5958 6031 6010
rect 6031 5958 6043 6010
rect 6043 5958 6057 6010
rect 6081 5958 6095 6010
rect 6095 5958 6107 6010
rect 6107 5958 6137 6010
rect 6161 5958 6171 6010
rect 6171 5958 6217 6010
rect 5921 5956 5977 5958
rect 6001 5956 6057 5958
rect 6081 5956 6137 5958
rect 6161 5956 6217 5958
rect 5921 4922 5977 4924
rect 6001 4922 6057 4924
rect 6081 4922 6137 4924
rect 6161 4922 6217 4924
rect 5921 4870 5967 4922
rect 5967 4870 5977 4922
rect 6001 4870 6031 4922
rect 6031 4870 6043 4922
rect 6043 4870 6057 4922
rect 6081 4870 6095 4922
rect 6095 4870 6107 4922
rect 6107 4870 6137 4922
rect 6161 4870 6171 4922
rect 6171 4870 6217 4922
rect 5921 4868 5977 4870
rect 6001 4868 6057 4870
rect 6081 4868 6137 4870
rect 6161 4868 6217 4870
rect 5921 3834 5977 3836
rect 6001 3834 6057 3836
rect 6081 3834 6137 3836
rect 6161 3834 6217 3836
rect 5921 3782 5967 3834
rect 5967 3782 5977 3834
rect 6001 3782 6031 3834
rect 6031 3782 6043 3834
rect 6043 3782 6057 3834
rect 6081 3782 6095 3834
rect 6095 3782 6107 3834
rect 6107 3782 6137 3834
rect 6161 3782 6171 3834
rect 6171 3782 6217 3834
rect 5921 3780 5977 3782
rect 6001 3780 6057 3782
rect 6081 3780 6137 3782
rect 6161 3780 6217 3782
rect 1582 2916 1638 2952
rect 1582 2896 1584 2916
rect 1584 2896 1636 2916
rect 1636 2896 1638 2916
rect 5921 2746 5977 2748
rect 6001 2746 6057 2748
rect 6081 2746 6137 2748
rect 6161 2746 6217 2748
rect 5921 2694 5967 2746
rect 5967 2694 5977 2746
rect 6001 2694 6031 2746
rect 6031 2694 6043 2746
rect 6043 2694 6057 2746
rect 6081 2694 6095 2746
rect 6095 2694 6107 2746
rect 6107 2694 6137 2746
rect 6161 2694 6171 2746
rect 6171 2694 6217 2746
rect 5921 2692 5977 2694
rect 6001 2692 6057 2694
rect 6081 2692 6137 2694
rect 6161 2692 6217 2694
rect 10886 28314 10942 28316
rect 10966 28314 11022 28316
rect 11046 28314 11102 28316
rect 11126 28314 11182 28316
rect 10886 28262 10932 28314
rect 10932 28262 10942 28314
rect 10966 28262 10996 28314
rect 10996 28262 11008 28314
rect 11008 28262 11022 28314
rect 11046 28262 11060 28314
rect 11060 28262 11072 28314
rect 11072 28262 11102 28314
rect 11126 28262 11136 28314
rect 11136 28262 11182 28314
rect 10886 28260 10942 28262
rect 10966 28260 11022 28262
rect 11046 28260 11102 28262
rect 11126 28260 11182 28262
rect 10886 27226 10942 27228
rect 10966 27226 11022 27228
rect 11046 27226 11102 27228
rect 11126 27226 11182 27228
rect 10886 27174 10932 27226
rect 10932 27174 10942 27226
rect 10966 27174 10996 27226
rect 10996 27174 11008 27226
rect 11008 27174 11022 27226
rect 11046 27174 11060 27226
rect 11060 27174 11072 27226
rect 11072 27174 11102 27226
rect 11126 27174 11136 27226
rect 11136 27174 11182 27226
rect 10886 27172 10942 27174
rect 10966 27172 11022 27174
rect 11046 27172 11102 27174
rect 11126 27172 11182 27174
rect 10886 26138 10942 26140
rect 10966 26138 11022 26140
rect 11046 26138 11102 26140
rect 11126 26138 11182 26140
rect 10886 26086 10932 26138
rect 10932 26086 10942 26138
rect 10966 26086 10996 26138
rect 10996 26086 11008 26138
rect 11008 26086 11022 26138
rect 11046 26086 11060 26138
rect 11060 26086 11072 26138
rect 11072 26086 11102 26138
rect 11126 26086 11136 26138
rect 11136 26086 11182 26138
rect 10886 26084 10942 26086
rect 10966 26084 11022 26086
rect 11046 26084 11102 26086
rect 11126 26084 11182 26086
rect 10598 24656 10654 24712
rect 10886 25050 10942 25052
rect 10966 25050 11022 25052
rect 11046 25050 11102 25052
rect 11126 25050 11182 25052
rect 10886 24998 10932 25050
rect 10932 24998 10942 25050
rect 10966 24998 10996 25050
rect 10996 24998 11008 25050
rect 11008 24998 11022 25050
rect 11046 24998 11060 25050
rect 11060 24998 11072 25050
rect 11072 24998 11102 25050
rect 11126 24998 11136 25050
rect 11136 24998 11182 25050
rect 10886 24996 10942 24998
rect 10966 24996 11022 24998
rect 11046 24996 11102 24998
rect 11126 24996 11182 24998
rect 11334 24268 11390 24304
rect 11334 24248 11336 24268
rect 11336 24248 11388 24268
rect 11388 24248 11390 24268
rect 10886 23962 10942 23964
rect 10966 23962 11022 23964
rect 11046 23962 11102 23964
rect 11126 23962 11182 23964
rect 10886 23910 10932 23962
rect 10932 23910 10942 23962
rect 10966 23910 10996 23962
rect 10996 23910 11008 23962
rect 11008 23910 11022 23962
rect 11046 23910 11060 23962
rect 11060 23910 11072 23962
rect 11072 23910 11102 23962
rect 11126 23910 11136 23962
rect 11136 23910 11182 23962
rect 10886 23908 10942 23910
rect 10966 23908 11022 23910
rect 11046 23908 11102 23910
rect 11126 23908 11182 23910
rect 11242 23704 11298 23760
rect 10886 22874 10942 22876
rect 10966 22874 11022 22876
rect 11046 22874 11102 22876
rect 11126 22874 11182 22876
rect 10886 22822 10932 22874
rect 10932 22822 10942 22874
rect 10966 22822 10996 22874
rect 10996 22822 11008 22874
rect 11008 22822 11022 22874
rect 11046 22822 11060 22874
rect 11060 22822 11072 22874
rect 11072 22822 11102 22874
rect 11126 22822 11136 22874
rect 11136 22822 11182 22874
rect 10886 22820 10942 22822
rect 10966 22820 11022 22822
rect 11046 22820 11102 22822
rect 11126 22820 11182 22822
rect 11334 22344 11390 22400
rect 10886 21786 10942 21788
rect 10966 21786 11022 21788
rect 11046 21786 11102 21788
rect 11126 21786 11182 21788
rect 10886 21734 10932 21786
rect 10932 21734 10942 21786
rect 10966 21734 10996 21786
rect 10996 21734 11008 21786
rect 11008 21734 11022 21786
rect 11046 21734 11060 21786
rect 11060 21734 11072 21786
rect 11072 21734 11102 21786
rect 11126 21734 11136 21786
rect 11136 21734 11182 21786
rect 10886 21732 10942 21734
rect 10966 21732 11022 21734
rect 11046 21732 11102 21734
rect 11126 21732 11182 21734
rect 11058 21528 11114 21584
rect 10886 20698 10942 20700
rect 10966 20698 11022 20700
rect 11046 20698 11102 20700
rect 11126 20698 11182 20700
rect 10886 20646 10932 20698
rect 10932 20646 10942 20698
rect 10966 20646 10996 20698
rect 10996 20646 11008 20698
rect 11008 20646 11022 20698
rect 11046 20646 11060 20698
rect 11060 20646 11072 20698
rect 11072 20646 11102 20698
rect 11126 20646 11136 20698
rect 11136 20646 11182 20698
rect 10886 20644 10942 20646
rect 10966 20644 11022 20646
rect 11046 20644 11102 20646
rect 11126 20644 11182 20646
rect 10886 19610 10942 19612
rect 10966 19610 11022 19612
rect 11046 19610 11102 19612
rect 11126 19610 11182 19612
rect 10886 19558 10932 19610
rect 10932 19558 10942 19610
rect 10966 19558 10996 19610
rect 10996 19558 11008 19610
rect 11008 19558 11022 19610
rect 11046 19558 11060 19610
rect 11060 19558 11072 19610
rect 11072 19558 11102 19610
rect 11126 19558 11136 19610
rect 11136 19558 11182 19610
rect 10886 19556 10942 19558
rect 10966 19556 11022 19558
rect 11046 19556 11102 19558
rect 11126 19556 11182 19558
rect 10886 18522 10942 18524
rect 10966 18522 11022 18524
rect 11046 18522 11102 18524
rect 11126 18522 11182 18524
rect 10886 18470 10932 18522
rect 10932 18470 10942 18522
rect 10966 18470 10996 18522
rect 10996 18470 11008 18522
rect 11008 18470 11022 18522
rect 11046 18470 11060 18522
rect 11060 18470 11072 18522
rect 11072 18470 11102 18522
rect 11126 18470 11136 18522
rect 11136 18470 11182 18522
rect 10886 18468 10942 18470
rect 10966 18468 11022 18470
rect 11046 18468 11102 18470
rect 11126 18468 11182 18470
rect 11426 21292 11428 21312
rect 11428 21292 11480 21312
rect 11480 21292 11482 21312
rect 11426 21256 11482 21292
rect 11518 21120 11574 21176
rect 10886 17434 10942 17436
rect 10966 17434 11022 17436
rect 11046 17434 11102 17436
rect 11126 17434 11182 17436
rect 10886 17382 10932 17434
rect 10932 17382 10942 17434
rect 10966 17382 10996 17434
rect 10996 17382 11008 17434
rect 11008 17382 11022 17434
rect 11046 17382 11060 17434
rect 11060 17382 11072 17434
rect 11072 17382 11102 17434
rect 11126 17382 11136 17434
rect 11136 17382 11182 17434
rect 10886 17380 10942 17382
rect 10966 17380 11022 17382
rect 11046 17380 11102 17382
rect 11126 17380 11182 17382
rect 10886 16346 10942 16348
rect 10966 16346 11022 16348
rect 11046 16346 11102 16348
rect 11126 16346 11182 16348
rect 10886 16294 10932 16346
rect 10932 16294 10942 16346
rect 10966 16294 10996 16346
rect 10996 16294 11008 16346
rect 11008 16294 11022 16346
rect 11046 16294 11060 16346
rect 11060 16294 11072 16346
rect 11072 16294 11102 16346
rect 11126 16294 11136 16346
rect 11136 16294 11182 16346
rect 10886 16292 10942 16294
rect 10966 16292 11022 16294
rect 11046 16292 11102 16294
rect 11126 16292 11182 16294
rect 10886 15258 10942 15260
rect 10966 15258 11022 15260
rect 11046 15258 11102 15260
rect 11126 15258 11182 15260
rect 10886 15206 10932 15258
rect 10932 15206 10942 15258
rect 10966 15206 10996 15258
rect 10996 15206 11008 15258
rect 11008 15206 11022 15258
rect 11046 15206 11060 15258
rect 11060 15206 11072 15258
rect 11072 15206 11102 15258
rect 11126 15206 11136 15258
rect 11136 15206 11182 15258
rect 10886 15204 10942 15206
rect 10966 15204 11022 15206
rect 11046 15204 11102 15206
rect 11126 15204 11182 15206
rect 10886 14170 10942 14172
rect 10966 14170 11022 14172
rect 11046 14170 11102 14172
rect 11126 14170 11182 14172
rect 10886 14118 10932 14170
rect 10932 14118 10942 14170
rect 10966 14118 10996 14170
rect 10996 14118 11008 14170
rect 11008 14118 11022 14170
rect 11046 14118 11060 14170
rect 11060 14118 11072 14170
rect 11072 14118 11102 14170
rect 11126 14118 11136 14170
rect 11136 14118 11182 14170
rect 10886 14116 10942 14118
rect 10966 14116 11022 14118
rect 11046 14116 11102 14118
rect 11126 14116 11182 14118
rect 10886 13082 10942 13084
rect 10966 13082 11022 13084
rect 11046 13082 11102 13084
rect 11126 13082 11182 13084
rect 10886 13030 10932 13082
rect 10932 13030 10942 13082
rect 10966 13030 10996 13082
rect 10996 13030 11008 13082
rect 11008 13030 11022 13082
rect 11046 13030 11060 13082
rect 11060 13030 11072 13082
rect 11072 13030 11102 13082
rect 11126 13030 11136 13082
rect 11136 13030 11182 13082
rect 10886 13028 10942 13030
rect 10966 13028 11022 13030
rect 11046 13028 11102 13030
rect 11126 13028 11182 13030
rect 10886 11994 10942 11996
rect 10966 11994 11022 11996
rect 11046 11994 11102 11996
rect 11126 11994 11182 11996
rect 10886 11942 10932 11994
rect 10932 11942 10942 11994
rect 10966 11942 10996 11994
rect 10996 11942 11008 11994
rect 11008 11942 11022 11994
rect 11046 11942 11060 11994
rect 11060 11942 11072 11994
rect 11072 11942 11102 11994
rect 11126 11942 11136 11994
rect 11136 11942 11182 11994
rect 10886 11940 10942 11942
rect 10966 11940 11022 11942
rect 11046 11940 11102 11942
rect 11126 11940 11182 11942
rect 12806 29280 12862 29336
rect 13266 29416 13322 29472
rect 12898 29144 12954 29200
rect 12346 22344 12402 22400
rect 12438 22072 12494 22128
rect 12254 21428 12256 21448
rect 12256 21428 12308 21448
rect 12308 21428 12310 21448
rect 12254 21392 12310 21428
rect 12530 21120 12586 21176
rect 12254 18808 12310 18864
rect 13358 25744 13414 25800
rect 13358 25064 13414 25120
rect 15198 45328 15254 45384
rect 15852 45178 15908 45180
rect 15932 45178 15988 45180
rect 16012 45178 16068 45180
rect 16092 45178 16148 45180
rect 15852 45126 15898 45178
rect 15898 45126 15908 45178
rect 15932 45126 15962 45178
rect 15962 45126 15974 45178
rect 15974 45126 15988 45178
rect 16012 45126 16026 45178
rect 16026 45126 16038 45178
rect 16038 45126 16068 45178
rect 16092 45126 16102 45178
rect 16102 45126 16148 45178
rect 15852 45124 15908 45126
rect 15932 45124 15988 45126
rect 16012 45124 16068 45126
rect 16092 45124 16148 45126
rect 15290 44104 15346 44160
rect 15852 44090 15908 44092
rect 15932 44090 15988 44092
rect 16012 44090 16068 44092
rect 16092 44090 16148 44092
rect 15852 44038 15898 44090
rect 15898 44038 15908 44090
rect 15932 44038 15962 44090
rect 15962 44038 15974 44090
rect 15974 44038 15988 44090
rect 16012 44038 16026 44090
rect 16026 44038 16038 44090
rect 16038 44038 16068 44090
rect 16092 44038 16102 44090
rect 16102 44038 16148 44090
rect 15852 44036 15908 44038
rect 15932 44036 15988 44038
rect 16012 44036 16068 44038
rect 16092 44036 16148 44038
rect 17038 45328 17094 45384
rect 14002 25744 14058 25800
rect 12990 21256 13046 21312
rect 13082 18300 13084 18320
rect 13084 18300 13136 18320
rect 13136 18300 13138 18320
rect 13082 18264 13138 18300
rect 13358 17740 13414 17776
rect 13358 17720 13360 17740
rect 13360 17720 13412 17740
rect 13412 17720 13414 17740
rect 10886 10906 10942 10908
rect 10966 10906 11022 10908
rect 11046 10906 11102 10908
rect 11126 10906 11182 10908
rect 10886 10854 10932 10906
rect 10932 10854 10942 10906
rect 10966 10854 10996 10906
rect 10996 10854 11008 10906
rect 11008 10854 11022 10906
rect 11046 10854 11060 10906
rect 11060 10854 11072 10906
rect 11072 10854 11102 10906
rect 11126 10854 11136 10906
rect 11136 10854 11182 10906
rect 10886 10852 10942 10854
rect 10966 10852 11022 10854
rect 11046 10852 11102 10854
rect 11126 10852 11182 10854
rect 10886 9818 10942 9820
rect 10966 9818 11022 9820
rect 11046 9818 11102 9820
rect 11126 9818 11182 9820
rect 10886 9766 10932 9818
rect 10932 9766 10942 9818
rect 10966 9766 10996 9818
rect 10996 9766 11008 9818
rect 11008 9766 11022 9818
rect 11046 9766 11060 9818
rect 11060 9766 11072 9818
rect 11072 9766 11102 9818
rect 11126 9766 11136 9818
rect 11136 9766 11182 9818
rect 10886 9764 10942 9766
rect 10966 9764 11022 9766
rect 11046 9764 11102 9766
rect 11126 9764 11182 9766
rect 10886 8730 10942 8732
rect 10966 8730 11022 8732
rect 11046 8730 11102 8732
rect 11126 8730 11182 8732
rect 10886 8678 10932 8730
rect 10932 8678 10942 8730
rect 10966 8678 10996 8730
rect 10996 8678 11008 8730
rect 11008 8678 11022 8730
rect 11046 8678 11060 8730
rect 11060 8678 11072 8730
rect 11072 8678 11102 8730
rect 11126 8678 11136 8730
rect 11136 8678 11182 8730
rect 10886 8676 10942 8678
rect 10966 8676 11022 8678
rect 11046 8676 11102 8678
rect 11126 8676 11182 8678
rect 10886 7642 10942 7644
rect 10966 7642 11022 7644
rect 11046 7642 11102 7644
rect 11126 7642 11182 7644
rect 10886 7590 10932 7642
rect 10932 7590 10942 7642
rect 10966 7590 10996 7642
rect 10996 7590 11008 7642
rect 11008 7590 11022 7642
rect 11046 7590 11060 7642
rect 11060 7590 11072 7642
rect 11072 7590 11102 7642
rect 11126 7590 11136 7642
rect 11136 7590 11182 7642
rect 10886 7588 10942 7590
rect 10966 7588 11022 7590
rect 11046 7588 11102 7590
rect 11126 7588 11182 7590
rect 10886 6554 10942 6556
rect 10966 6554 11022 6556
rect 11046 6554 11102 6556
rect 11126 6554 11182 6556
rect 10886 6502 10932 6554
rect 10932 6502 10942 6554
rect 10966 6502 10996 6554
rect 10996 6502 11008 6554
rect 11008 6502 11022 6554
rect 11046 6502 11060 6554
rect 11060 6502 11072 6554
rect 11072 6502 11102 6554
rect 11126 6502 11136 6554
rect 11136 6502 11182 6554
rect 10886 6500 10942 6502
rect 10966 6500 11022 6502
rect 11046 6500 11102 6502
rect 11126 6500 11182 6502
rect 10886 5466 10942 5468
rect 10966 5466 11022 5468
rect 11046 5466 11102 5468
rect 11126 5466 11182 5468
rect 10886 5414 10932 5466
rect 10932 5414 10942 5466
rect 10966 5414 10996 5466
rect 10996 5414 11008 5466
rect 11008 5414 11022 5466
rect 11046 5414 11060 5466
rect 11060 5414 11072 5466
rect 11072 5414 11102 5466
rect 11126 5414 11136 5466
rect 11136 5414 11182 5466
rect 10886 5412 10942 5414
rect 10966 5412 11022 5414
rect 11046 5412 11102 5414
rect 11126 5412 11182 5414
rect 10886 4378 10942 4380
rect 10966 4378 11022 4380
rect 11046 4378 11102 4380
rect 11126 4378 11182 4380
rect 10886 4326 10932 4378
rect 10932 4326 10942 4378
rect 10966 4326 10996 4378
rect 10996 4326 11008 4378
rect 11008 4326 11022 4378
rect 11046 4326 11060 4378
rect 11060 4326 11072 4378
rect 11072 4326 11102 4378
rect 11126 4326 11136 4378
rect 11136 4326 11182 4378
rect 10886 4324 10942 4326
rect 10966 4324 11022 4326
rect 11046 4324 11102 4326
rect 11126 4324 11182 4326
rect 10886 3290 10942 3292
rect 10966 3290 11022 3292
rect 11046 3290 11102 3292
rect 11126 3290 11182 3292
rect 10886 3238 10932 3290
rect 10932 3238 10942 3290
rect 10966 3238 10996 3290
rect 10996 3238 11008 3290
rect 11008 3238 11022 3290
rect 11046 3238 11060 3290
rect 11060 3238 11072 3290
rect 11072 3238 11102 3290
rect 11126 3238 11136 3290
rect 11136 3238 11182 3290
rect 10886 3236 10942 3238
rect 10966 3236 11022 3238
rect 11046 3236 11102 3238
rect 11126 3236 11182 3238
rect 13818 19116 13820 19136
rect 13820 19116 13872 19136
rect 13872 19116 13874 19136
rect 13818 19080 13874 19116
rect 14094 23196 14096 23216
rect 14096 23196 14148 23216
rect 14148 23196 14150 23216
rect 14094 23160 14150 23196
rect 15852 43002 15908 43004
rect 15932 43002 15988 43004
rect 16012 43002 16068 43004
rect 16092 43002 16148 43004
rect 15852 42950 15898 43002
rect 15898 42950 15908 43002
rect 15932 42950 15962 43002
rect 15962 42950 15974 43002
rect 15974 42950 15988 43002
rect 16012 42950 16026 43002
rect 16026 42950 16038 43002
rect 16038 42950 16068 43002
rect 16092 42950 16102 43002
rect 16102 42950 16148 43002
rect 15852 42948 15908 42950
rect 15932 42948 15988 42950
rect 16012 42948 16068 42950
rect 16092 42948 16148 42950
rect 15852 41914 15908 41916
rect 15932 41914 15988 41916
rect 16012 41914 16068 41916
rect 16092 41914 16148 41916
rect 15852 41862 15898 41914
rect 15898 41862 15908 41914
rect 15932 41862 15962 41914
rect 15962 41862 15974 41914
rect 15974 41862 15988 41914
rect 16012 41862 16026 41914
rect 16026 41862 16038 41914
rect 16038 41862 16068 41914
rect 16092 41862 16102 41914
rect 16102 41862 16148 41914
rect 15852 41860 15908 41862
rect 15932 41860 15988 41862
rect 16012 41860 16068 41862
rect 16092 41860 16148 41862
rect 15852 40826 15908 40828
rect 15932 40826 15988 40828
rect 16012 40826 16068 40828
rect 16092 40826 16148 40828
rect 15852 40774 15898 40826
rect 15898 40774 15908 40826
rect 15932 40774 15962 40826
rect 15962 40774 15974 40826
rect 15974 40774 15988 40826
rect 16012 40774 16026 40826
rect 16026 40774 16038 40826
rect 16038 40774 16068 40826
rect 16092 40774 16102 40826
rect 16102 40774 16148 40826
rect 15852 40772 15908 40774
rect 15932 40772 15988 40774
rect 16012 40772 16068 40774
rect 16092 40772 16148 40774
rect 15852 39738 15908 39740
rect 15932 39738 15988 39740
rect 16012 39738 16068 39740
rect 16092 39738 16148 39740
rect 15852 39686 15898 39738
rect 15898 39686 15908 39738
rect 15932 39686 15962 39738
rect 15962 39686 15974 39738
rect 15974 39686 15988 39738
rect 16012 39686 16026 39738
rect 16026 39686 16038 39738
rect 16038 39686 16068 39738
rect 16092 39686 16102 39738
rect 16102 39686 16148 39738
rect 15852 39684 15908 39686
rect 15932 39684 15988 39686
rect 16012 39684 16068 39686
rect 16092 39684 16148 39686
rect 15852 38650 15908 38652
rect 15932 38650 15988 38652
rect 16012 38650 16068 38652
rect 16092 38650 16148 38652
rect 15852 38598 15898 38650
rect 15898 38598 15908 38650
rect 15932 38598 15962 38650
rect 15962 38598 15974 38650
rect 15974 38598 15988 38650
rect 16012 38598 16026 38650
rect 16026 38598 16038 38650
rect 16038 38598 16068 38650
rect 16092 38598 16102 38650
rect 16102 38598 16148 38650
rect 15852 38596 15908 38598
rect 15932 38596 15988 38598
rect 16012 38596 16068 38598
rect 16092 38596 16148 38598
rect 15852 37562 15908 37564
rect 15932 37562 15988 37564
rect 16012 37562 16068 37564
rect 16092 37562 16148 37564
rect 15852 37510 15898 37562
rect 15898 37510 15908 37562
rect 15932 37510 15962 37562
rect 15962 37510 15974 37562
rect 15974 37510 15988 37562
rect 16012 37510 16026 37562
rect 16026 37510 16038 37562
rect 16038 37510 16068 37562
rect 16092 37510 16102 37562
rect 16102 37510 16148 37562
rect 15852 37508 15908 37510
rect 15932 37508 15988 37510
rect 16012 37508 16068 37510
rect 16092 37508 16148 37510
rect 15852 36474 15908 36476
rect 15932 36474 15988 36476
rect 16012 36474 16068 36476
rect 16092 36474 16148 36476
rect 15852 36422 15898 36474
rect 15898 36422 15908 36474
rect 15932 36422 15962 36474
rect 15962 36422 15974 36474
rect 15974 36422 15988 36474
rect 16012 36422 16026 36474
rect 16026 36422 16038 36474
rect 16038 36422 16068 36474
rect 16092 36422 16102 36474
rect 16102 36422 16148 36474
rect 15852 36420 15908 36422
rect 15932 36420 15988 36422
rect 16012 36420 16068 36422
rect 16092 36420 16148 36422
rect 15852 35386 15908 35388
rect 15932 35386 15988 35388
rect 16012 35386 16068 35388
rect 16092 35386 16148 35388
rect 15852 35334 15898 35386
rect 15898 35334 15908 35386
rect 15932 35334 15962 35386
rect 15962 35334 15974 35386
rect 15974 35334 15988 35386
rect 16012 35334 16026 35386
rect 16026 35334 16038 35386
rect 16038 35334 16068 35386
rect 16092 35334 16102 35386
rect 16102 35334 16148 35386
rect 15852 35332 15908 35334
rect 15932 35332 15988 35334
rect 16012 35332 16068 35334
rect 16092 35332 16148 35334
rect 15852 34298 15908 34300
rect 15932 34298 15988 34300
rect 16012 34298 16068 34300
rect 16092 34298 16148 34300
rect 15852 34246 15898 34298
rect 15898 34246 15908 34298
rect 15932 34246 15962 34298
rect 15962 34246 15974 34298
rect 15974 34246 15988 34298
rect 16012 34246 16026 34298
rect 16026 34246 16038 34298
rect 16038 34246 16068 34298
rect 16092 34246 16102 34298
rect 16102 34246 16148 34298
rect 15852 34244 15908 34246
rect 15932 34244 15988 34246
rect 16012 34244 16068 34246
rect 16092 34244 16148 34246
rect 15658 31728 15714 31784
rect 15382 31456 15438 31512
rect 14462 23704 14518 23760
rect 14370 18808 14426 18864
rect 14738 18808 14794 18864
rect 15852 33210 15908 33212
rect 15932 33210 15988 33212
rect 16012 33210 16068 33212
rect 16092 33210 16148 33212
rect 15852 33158 15898 33210
rect 15898 33158 15908 33210
rect 15932 33158 15962 33210
rect 15962 33158 15974 33210
rect 15974 33158 15988 33210
rect 16012 33158 16026 33210
rect 16026 33158 16038 33210
rect 16038 33158 16068 33210
rect 16092 33158 16102 33210
rect 16102 33158 16148 33210
rect 15852 33156 15908 33158
rect 15932 33156 15988 33158
rect 16012 33156 16068 33158
rect 16092 33156 16148 33158
rect 15852 32122 15908 32124
rect 15932 32122 15988 32124
rect 16012 32122 16068 32124
rect 16092 32122 16148 32124
rect 15852 32070 15898 32122
rect 15898 32070 15908 32122
rect 15932 32070 15962 32122
rect 15962 32070 15974 32122
rect 15974 32070 15988 32122
rect 16012 32070 16026 32122
rect 16026 32070 16038 32122
rect 16038 32070 16068 32122
rect 16092 32070 16102 32122
rect 16102 32070 16148 32122
rect 15852 32068 15908 32070
rect 15932 32068 15988 32070
rect 16012 32068 16068 32070
rect 16092 32068 16148 32070
rect 15852 31034 15908 31036
rect 15932 31034 15988 31036
rect 16012 31034 16068 31036
rect 16092 31034 16148 31036
rect 15852 30982 15898 31034
rect 15898 30982 15908 31034
rect 15932 30982 15962 31034
rect 15962 30982 15974 31034
rect 15974 30982 15988 31034
rect 16012 30982 16026 31034
rect 16026 30982 16038 31034
rect 16038 30982 16068 31034
rect 16092 30982 16102 31034
rect 16102 30982 16148 31034
rect 15852 30980 15908 30982
rect 15932 30980 15988 30982
rect 16012 30980 16068 30982
rect 16092 30980 16148 30982
rect 15852 29946 15908 29948
rect 15932 29946 15988 29948
rect 16012 29946 16068 29948
rect 16092 29946 16148 29948
rect 15852 29894 15898 29946
rect 15898 29894 15908 29946
rect 15932 29894 15962 29946
rect 15962 29894 15974 29946
rect 15974 29894 15988 29946
rect 16012 29894 16026 29946
rect 16026 29894 16038 29946
rect 16038 29894 16068 29946
rect 16092 29894 16102 29946
rect 16102 29894 16148 29946
rect 15852 29892 15908 29894
rect 15932 29892 15988 29894
rect 16012 29892 16068 29894
rect 16092 29892 16148 29894
rect 16026 29144 16082 29200
rect 15852 28858 15908 28860
rect 15932 28858 15988 28860
rect 16012 28858 16068 28860
rect 16092 28858 16148 28860
rect 15852 28806 15898 28858
rect 15898 28806 15908 28858
rect 15932 28806 15962 28858
rect 15962 28806 15974 28858
rect 15974 28806 15988 28858
rect 16012 28806 16026 28858
rect 16026 28806 16038 28858
rect 16038 28806 16068 28858
rect 16092 28806 16102 28858
rect 16102 28806 16148 28858
rect 15852 28804 15908 28806
rect 15932 28804 15988 28806
rect 16012 28804 16068 28806
rect 16092 28804 16148 28806
rect 15852 27770 15908 27772
rect 15932 27770 15988 27772
rect 16012 27770 16068 27772
rect 16092 27770 16148 27772
rect 15852 27718 15898 27770
rect 15898 27718 15908 27770
rect 15932 27718 15962 27770
rect 15962 27718 15974 27770
rect 15974 27718 15988 27770
rect 16012 27718 16026 27770
rect 16026 27718 16038 27770
rect 16038 27718 16068 27770
rect 16092 27718 16102 27770
rect 16102 27718 16148 27770
rect 15852 27716 15908 27718
rect 15932 27716 15988 27718
rect 16012 27716 16068 27718
rect 16092 27716 16148 27718
rect 15852 26682 15908 26684
rect 15932 26682 15988 26684
rect 16012 26682 16068 26684
rect 16092 26682 16148 26684
rect 15852 26630 15898 26682
rect 15898 26630 15908 26682
rect 15932 26630 15962 26682
rect 15962 26630 15974 26682
rect 15974 26630 15988 26682
rect 16012 26630 16026 26682
rect 16026 26630 16038 26682
rect 16038 26630 16068 26682
rect 16092 26630 16102 26682
rect 16102 26630 16148 26682
rect 15852 26628 15908 26630
rect 15932 26628 15988 26630
rect 16012 26628 16068 26630
rect 16092 26628 16148 26630
rect 16210 25880 16266 25936
rect 15852 25594 15908 25596
rect 15932 25594 15988 25596
rect 16012 25594 16068 25596
rect 16092 25594 16148 25596
rect 15852 25542 15898 25594
rect 15898 25542 15908 25594
rect 15932 25542 15962 25594
rect 15962 25542 15974 25594
rect 15974 25542 15988 25594
rect 16012 25542 16026 25594
rect 16026 25542 16038 25594
rect 16038 25542 16068 25594
rect 16092 25542 16102 25594
rect 16102 25542 16148 25594
rect 15852 25540 15908 25542
rect 15932 25540 15988 25542
rect 16012 25540 16068 25542
rect 16092 25540 16148 25542
rect 15014 20576 15070 20632
rect 15014 19080 15070 19136
rect 15852 24506 15908 24508
rect 15932 24506 15988 24508
rect 16012 24506 16068 24508
rect 16092 24506 16148 24508
rect 15852 24454 15898 24506
rect 15898 24454 15908 24506
rect 15932 24454 15962 24506
rect 15962 24454 15974 24506
rect 15974 24454 15988 24506
rect 16012 24454 16026 24506
rect 16026 24454 16038 24506
rect 16038 24454 16068 24506
rect 16092 24454 16102 24506
rect 16102 24454 16148 24506
rect 15852 24452 15908 24454
rect 15932 24452 15988 24454
rect 16012 24452 16068 24454
rect 16092 24452 16148 24454
rect 17314 44920 17370 44976
rect 17222 44784 17278 44840
rect 17222 44240 17278 44296
rect 16578 30912 16634 30968
rect 16578 30776 16634 30832
rect 16302 25100 16304 25120
rect 16304 25100 16356 25120
rect 16356 25100 16358 25120
rect 16302 25064 16358 25100
rect 16302 24248 16358 24304
rect 15852 23418 15908 23420
rect 15932 23418 15988 23420
rect 16012 23418 16068 23420
rect 16092 23418 16148 23420
rect 15852 23366 15898 23418
rect 15898 23366 15908 23418
rect 15932 23366 15962 23418
rect 15962 23366 15974 23418
rect 15974 23366 15988 23418
rect 16012 23366 16026 23418
rect 16026 23366 16038 23418
rect 16038 23366 16068 23418
rect 16092 23366 16102 23418
rect 16102 23366 16148 23418
rect 15852 23364 15908 23366
rect 15932 23364 15988 23366
rect 16012 23364 16068 23366
rect 16092 23364 16148 23366
rect 15934 23196 15936 23216
rect 15936 23196 15988 23216
rect 15988 23196 15990 23216
rect 15934 23160 15990 23196
rect 15852 22330 15908 22332
rect 15932 22330 15988 22332
rect 16012 22330 16068 22332
rect 16092 22330 16148 22332
rect 15852 22278 15898 22330
rect 15898 22278 15908 22330
rect 15932 22278 15962 22330
rect 15962 22278 15974 22330
rect 15974 22278 15988 22330
rect 16012 22278 16026 22330
rect 16026 22278 16038 22330
rect 16038 22278 16068 22330
rect 16092 22278 16102 22330
rect 16102 22278 16148 22330
rect 15852 22276 15908 22278
rect 15932 22276 15988 22278
rect 16012 22276 16068 22278
rect 16092 22276 16148 22278
rect 15852 21242 15908 21244
rect 15932 21242 15988 21244
rect 16012 21242 16068 21244
rect 16092 21242 16148 21244
rect 15852 21190 15898 21242
rect 15898 21190 15908 21242
rect 15932 21190 15962 21242
rect 15962 21190 15974 21242
rect 15974 21190 15988 21242
rect 16012 21190 16026 21242
rect 16026 21190 16038 21242
rect 16038 21190 16068 21242
rect 16092 21190 16102 21242
rect 16102 21190 16148 21242
rect 15852 21188 15908 21190
rect 15932 21188 15988 21190
rect 16012 21188 16068 21190
rect 16092 21188 16148 21190
rect 15852 20154 15908 20156
rect 15932 20154 15988 20156
rect 16012 20154 16068 20156
rect 16092 20154 16148 20156
rect 15852 20102 15898 20154
rect 15898 20102 15908 20154
rect 15932 20102 15962 20154
rect 15962 20102 15974 20154
rect 15974 20102 15988 20154
rect 16012 20102 16026 20154
rect 16026 20102 16038 20154
rect 16038 20102 16068 20154
rect 16092 20102 16102 20154
rect 16102 20102 16148 20154
rect 15852 20100 15908 20102
rect 15932 20100 15988 20102
rect 16012 20100 16068 20102
rect 16092 20100 16148 20102
rect 15852 19066 15908 19068
rect 15932 19066 15988 19068
rect 16012 19066 16068 19068
rect 16092 19066 16148 19068
rect 15852 19014 15898 19066
rect 15898 19014 15908 19066
rect 15932 19014 15962 19066
rect 15962 19014 15974 19066
rect 15974 19014 15988 19066
rect 16012 19014 16026 19066
rect 16026 19014 16038 19066
rect 16038 19014 16068 19066
rect 16092 19014 16102 19066
rect 16102 19014 16148 19066
rect 15852 19012 15908 19014
rect 15932 19012 15988 19014
rect 16012 19012 16068 19014
rect 16092 19012 16148 19014
rect 15852 17978 15908 17980
rect 15932 17978 15988 17980
rect 16012 17978 16068 17980
rect 16092 17978 16148 17980
rect 15852 17926 15898 17978
rect 15898 17926 15908 17978
rect 15932 17926 15962 17978
rect 15962 17926 15974 17978
rect 15974 17926 15988 17978
rect 16012 17926 16026 17978
rect 16026 17926 16038 17978
rect 16038 17926 16068 17978
rect 16092 17926 16102 17978
rect 16102 17926 16148 17978
rect 15852 17924 15908 17926
rect 15932 17924 15988 17926
rect 16012 17924 16068 17926
rect 16092 17924 16148 17926
rect 18510 43052 18512 43072
rect 18512 43052 18564 43072
rect 18564 43052 18566 43072
rect 18510 43016 18566 43052
rect 16854 30368 16910 30424
rect 17222 34584 17278 34640
rect 16762 22480 16818 22536
rect 17222 29452 17224 29472
rect 17224 29452 17276 29472
rect 17276 29452 17278 29472
rect 17222 29416 17278 29452
rect 17314 28212 17370 28248
rect 17314 28192 17316 28212
rect 17316 28192 17368 28212
rect 17368 28192 17370 28212
rect 17590 33904 17646 33960
rect 17682 31864 17738 31920
rect 17590 30096 17646 30152
rect 17498 29688 17554 29744
rect 17866 27956 17868 27976
rect 17868 27956 17920 27976
rect 17920 27956 17922 27976
rect 17866 27920 17922 27956
rect 18326 33768 18382 33824
rect 18234 31456 18290 31512
rect 18142 30368 18198 30424
rect 18142 29688 18198 29744
rect 16302 17720 16358 17776
rect 16670 18300 16672 18320
rect 16672 18300 16724 18320
rect 16724 18300 16726 18320
rect 16670 18264 16726 18300
rect 15750 17040 15806 17096
rect 15934 17060 15990 17096
rect 15934 17040 15936 17060
rect 15936 17040 15988 17060
rect 15988 17040 15990 17060
rect 15852 16890 15908 16892
rect 15932 16890 15988 16892
rect 16012 16890 16068 16892
rect 16092 16890 16148 16892
rect 15852 16838 15898 16890
rect 15898 16838 15908 16890
rect 15932 16838 15962 16890
rect 15962 16838 15974 16890
rect 15974 16838 15988 16890
rect 16012 16838 16026 16890
rect 16026 16838 16038 16890
rect 16038 16838 16068 16890
rect 16092 16838 16102 16890
rect 16102 16838 16148 16890
rect 15852 16836 15908 16838
rect 15932 16836 15988 16838
rect 16012 16836 16068 16838
rect 16092 16836 16148 16838
rect 15852 15802 15908 15804
rect 15932 15802 15988 15804
rect 16012 15802 16068 15804
rect 16092 15802 16148 15804
rect 15852 15750 15898 15802
rect 15898 15750 15908 15802
rect 15932 15750 15962 15802
rect 15962 15750 15974 15802
rect 15974 15750 15988 15802
rect 16012 15750 16026 15802
rect 16026 15750 16038 15802
rect 16038 15750 16068 15802
rect 16092 15750 16102 15802
rect 16102 15750 16148 15802
rect 15852 15748 15908 15750
rect 15932 15748 15988 15750
rect 16012 15748 16068 15750
rect 16092 15748 16148 15750
rect 15852 14714 15908 14716
rect 15932 14714 15988 14716
rect 16012 14714 16068 14716
rect 16092 14714 16148 14716
rect 15852 14662 15898 14714
rect 15898 14662 15908 14714
rect 15932 14662 15962 14714
rect 15962 14662 15974 14714
rect 15974 14662 15988 14714
rect 16012 14662 16026 14714
rect 16026 14662 16038 14714
rect 16038 14662 16068 14714
rect 16092 14662 16102 14714
rect 16102 14662 16148 14714
rect 15852 14660 15908 14662
rect 15932 14660 15988 14662
rect 16012 14660 16068 14662
rect 16092 14660 16148 14662
rect 15852 13626 15908 13628
rect 15932 13626 15988 13628
rect 16012 13626 16068 13628
rect 16092 13626 16148 13628
rect 15852 13574 15898 13626
rect 15898 13574 15908 13626
rect 15932 13574 15962 13626
rect 15962 13574 15974 13626
rect 15974 13574 15988 13626
rect 16012 13574 16026 13626
rect 16026 13574 16038 13626
rect 16038 13574 16068 13626
rect 16092 13574 16102 13626
rect 16102 13574 16148 13626
rect 15852 13572 15908 13574
rect 15932 13572 15988 13574
rect 16012 13572 16068 13574
rect 16092 13572 16148 13574
rect 15852 12538 15908 12540
rect 15932 12538 15988 12540
rect 16012 12538 16068 12540
rect 16092 12538 16148 12540
rect 15852 12486 15898 12538
rect 15898 12486 15908 12538
rect 15932 12486 15962 12538
rect 15962 12486 15974 12538
rect 15974 12486 15988 12538
rect 16012 12486 16026 12538
rect 16026 12486 16038 12538
rect 16038 12486 16068 12538
rect 16092 12486 16102 12538
rect 16102 12486 16148 12538
rect 15852 12484 15908 12486
rect 15932 12484 15988 12486
rect 16012 12484 16068 12486
rect 16092 12484 16148 12486
rect 15852 11450 15908 11452
rect 15932 11450 15988 11452
rect 16012 11450 16068 11452
rect 16092 11450 16148 11452
rect 15852 11398 15898 11450
rect 15898 11398 15908 11450
rect 15932 11398 15962 11450
rect 15962 11398 15974 11450
rect 15974 11398 15988 11450
rect 16012 11398 16026 11450
rect 16026 11398 16038 11450
rect 16038 11398 16068 11450
rect 16092 11398 16102 11450
rect 16102 11398 16148 11450
rect 15852 11396 15908 11398
rect 15932 11396 15988 11398
rect 16012 11396 16068 11398
rect 16092 11396 16148 11398
rect 15852 10362 15908 10364
rect 15932 10362 15988 10364
rect 16012 10362 16068 10364
rect 16092 10362 16148 10364
rect 15852 10310 15898 10362
rect 15898 10310 15908 10362
rect 15932 10310 15962 10362
rect 15962 10310 15974 10362
rect 15974 10310 15988 10362
rect 16012 10310 16026 10362
rect 16026 10310 16038 10362
rect 16038 10310 16068 10362
rect 16092 10310 16102 10362
rect 16102 10310 16148 10362
rect 15852 10308 15908 10310
rect 15932 10308 15988 10310
rect 16012 10308 16068 10310
rect 16092 10308 16148 10310
rect 15852 9274 15908 9276
rect 15932 9274 15988 9276
rect 16012 9274 16068 9276
rect 16092 9274 16148 9276
rect 15852 9222 15898 9274
rect 15898 9222 15908 9274
rect 15932 9222 15962 9274
rect 15962 9222 15974 9274
rect 15974 9222 15988 9274
rect 16012 9222 16026 9274
rect 16026 9222 16038 9274
rect 16038 9222 16068 9274
rect 16092 9222 16102 9274
rect 16102 9222 16148 9274
rect 15852 9220 15908 9222
rect 15932 9220 15988 9222
rect 16012 9220 16068 9222
rect 16092 9220 16148 9222
rect 17130 22344 17186 22400
rect 17406 22208 17462 22264
rect 18050 25900 18106 25936
rect 18050 25880 18052 25900
rect 18052 25880 18104 25900
rect 18104 25880 18106 25900
rect 17866 21664 17922 21720
rect 18602 36216 18658 36272
rect 18510 35128 18566 35184
rect 19338 42336 19394 42392
rect 19430 42236 19432 42256
rect 19432 42236 19484 42256
rect 19484 42236 19486 42256
rect 19430 42200 19486 42236
rect 19890 42336 19946 42392
rect 19798 41112 19854 41168
rect 19614 40432 19670 40488
rect 19614 39636 19670 39672
rect 19614 39616 19616 39636
rect 19616 39616 19668 39636
rect 19668 39616 19670 39636
rect 18970 35128 19026 35184
rect 19062 35028 19064 35048
rect 19064 35028 19116 35048
rect 19116 35028 19118 35048
rect 19062 34992 19118 35028
rect 18970 34448 19026 34504
rect 18786 31864 18842 31920
rect 18510 30096 18566 30152
rect 18510 28056 18566 28112
rect 18878 30504 18934 30560
rect 18694 30096 18750 30152
rect 20817 45722 20873 45724
rect 20897 45722 20953 45724
rect 20977 45722 21033 45724
rect 21057 45722 21113 45724
rect 20817 45670 20863 45722
rect 20863 45670 20873 45722
rect 20897 45670 20927 45722
rect 20927 45670 20939 45722
rect 20939 45670 20953 45722
rect 20977 45670 20991 45722
rect 20991 45670 21003 45722
rect 21003 45670 21033 45722
rect 21057 45670 21067 45722
rect 21067 45670 21113 45722
rect 20817 45668 20873 45670
rect 20897 45668 20953 45670
rect 20977 45668 21033 45670
rect 21057 45668 21113 45670
rect 20350 38936 20406 38992
rect 20994 45328 21050 45384
rect 20994 44820 20996 44840
rect 20996 44820 21048 44840
rect 21048 44820 21050 44840
rect 20994 44784 21050 44820
rect 21454 45500 21456 45520
rect 21456 45500 21508 45520
rect 21508 45500 21510 45520
rect 21454 45464 21510 45500
rect 21454 44940 21510 44976
rect 21454 44920 21456 44940
rect 21456 44920 21508 44940
rect 21508 44920 21510 44940
rect 22006 44920 22062 44976
rect 22190 44956 22192 44976
rect 22192 44956 22244 44976
rect 22244 44956 22246 44976
rect 22190 44920 22246 44956
rect 20817 44634 20873 44636
rect 20897 44634 20953 44636
rect 20977 44634 21033 44636
rect 21057 44634 21113 44636
rect 20817 44582 20863 44634
rect 20863 44582 20873 44634
rect 20897 44582 20927 44634
rect 20927 44582 20939 44634
rect 20939 44582 20953 44634
rect 20977 44582 20991 44634
rect 20991 44582 21003 44634
rect 21003 44582 21033 44634
rect 21057 44582 21067 44634
rect 21067 44582 21113 44634
rect 20817 44580 20873 44582
rect 20897 44580 20953 44582
rect 20977 44580 21033 44582
rect 21057 44580 21113 44582
rect 20718 44240 20774 44296
rect 20817 43546 20873 43548
rect 20897 43546 20953 43548
rect 20977 43546 21033 43548
rect 21057 43546 21113 43548
rect 20817 43494 20863 43546
rect 20863 43494 20873 43546
rect 20897 43494 20927 43546
rect 20927 43494 20939 43546
rect 20939 43494 20953 43546
rect 20977 43494 20991 43546
rect 20991 43494 21003 43546
rect 21003 43494 21033 43546
rect 21057 43494 21067 43546
rect 21067 43494 21113 43546
rect 20817 43492 20873 43494
rect 20897 43492 20953 43494
rect 20977 43492 21033 43494
rect 21057 43492 21113 43494
rect 20817 42458 20873 42460
rect 20897 42458 20953 42460
rect 20977 42458 21033 42460
rect 21057 42458 21113 42460
rect 20817 42406 20863 42458
rect 20863 42406 20873 42458
rect 20897 42406 20927 42458
rect 20927 42406 20939 42458
rect 20939 42406 20953 42458
rect 20977 42406 20991 42458
rect 20991 42406 21003 42458
rect 21003 42406 21033 42458
rect 21057 42406 21067 42458
rect 21067 42406 21113 42458
rect 20817 42404 20873 42406
rect 20897 42404 20953 42406
rect 20977 42404 21033 42406
rect 21057 42404 21113 42406
rect 20626 42220 20682 42256
rect 20626 42200 20628 42220
rect 20628 42200 20680 42220
rect 20680 42200 20682 42220
rect 21178 42200 21234 42256
rect 20626 42064 20682 42120
rect 20817 41370 20873 41372
rect 20897 41370 20953 41372
rect 20977 41370 21033 41372
rect 21057 41370 21113 41372
rect 20817 41318 20863 41370
rect 20863 41318 20873 41370
rect 20897 41318 20927 41370
rect 20927 41318 20939 41370
rect 20939 41318 20953 41370
rect 20977 41318 20991 41370
rect 20991 41318 21003 41370
rect 21003 41318 21033 41370
rect 21057 41318 21067 41370
rect 21067 41318 21113 41370
rect 20817 41316 20873 41318
rect 20897 41316 20953 41318
rect 20977 41316 21033 41318
rect 21057 41316 21113 41318
rect 20817 40282 20873 40284
rect 20897 40282 20953 40284
rect 20977 40282 21033 40284
rect 21057 40282 21113 40284
rect 20817 40230 20863 40282
rect 20863 40230 20873 40282
rect 20897 40230 20927 40282
rect 20927 40230 20939 40282
rect 20939 40230 20953 40282
rect 20977 40230 20991 40282
rect 20991 40230 21003 40282
rect 21003 40230 21033 40282
rect 21057 40230 21067 40282
rect 21067 40230 21113 40282
rect 20817 40228 20873 40230
rect 20897 40228 20953 40230
rect 20977 40228 21033 40230
rect 21057 40228 21113 40230
rect 20817 39194 20873 39196
rect 20897 39194 20953 39196
rect 20977 39194 21033 39196
rect 21057 39194 21113 39196
rect 20817 39142 20863 39194
rect 20863 39142 20873 39194
rect 20897 39142 20927 39194
rect 20927 39142 20939 39194
rect 20939 39142 20953 39194
rect 20977 39142 20991 39194
rect 20991 39142 21003 39194
rect 21003 39142 21033 39194
rect 21057 39142 21067 39194
rect 21067 39142 21113 39194
rect 20817 39140 20873 39142
rect 20897 39140 20953 39142
rect 20977 39140 21033 39142
rect 21057 39140 21113 39142
rect 21454 44376 21510 44432
rect 21546 44104 21602 44160
rect 21546 42200 21602 42256
rect 21454 42064 21510 42120
rect 19982 35708 19984 35728
rect 19984 35708 20036 35728
rect 20036 35708 20038 35728
rect 19982 35672 20038 35708
rect 19614 34992 19670 35048
rect 19338 30676 19340 30696
rect 19340 30676 19392 30696
rect 19392 30676 19394 30696
rect 19338 30640 19394 30676
rect 19154 29280 19210 29336
rect 19154 28600 19210 28656
rect 19338 28600 19394 28656
rect 18970 28328 19026 28384
rect 19062 28192 19118 28248
rect 19338 28364 19340 28384
rect 19340 28364 19392 28384
rect 19392 28364 19394 28384
rect 19338 28328 19394 28364
rect 19062 28076 19118 28112
rect 19062 28056 19064 28076
rect 19064 28056 19116 28076
rect 19116 28056 19118 28076
rect 19338 28056 19394 28112
rect 18970 27784 19026 27840
rect 19246 27648 19302 27704
rect 19154 27124 19210 27160
rect 19154 27104 19156 27124
rect 19156 27104 19208 27124
rect 19208 27104 19210 27124
rect 18786 22480 18842 22536
rect 20442 35128 20498 35184
rect 20626 37188 20682 37224
rect 20626 37168 20628 37188
rect 20628 37168 20680 37188
rect 20680 37168 20682 37188
rect 21454 40180 21510 40216
rect 21454 40160 21456 40180
rect 21456 40160 21508 40180
rect 21508 40160 21510 40180
rect 20817 38106 20873 38108
rect 20897 38106 20953 38108
rect 20977 38106 21033 38108
rect 21057 38106 21113 38108
rect 20817 38054 20863 38106
rect 20863 38054 20873 38106
rect 20897 38054 20927 38106
rect 20927 38054 20939 38106
rect 20939 38054 20953 38106
rect 20977 38054 20991 38106
rect 20991 38054 21003 38106
rect 21003 38054 21033 38106
rect 21057 38054 21067 38106
rect 21067 38054 21113 38106
rect 20817 38052 20873 38054
rect 20897 38052 20953 38054
rect 20977 38052 21033 38054
rect 21057 38052 21113 38054
rect 21362 37168 21418 37224
rect 20817 37018 20873 37020
rect 20897 37018 20953 37020
rect 20977 37018 21033 37020
rect 21057 37018 21113 37020
rect 20817 36966 20863 37018
rect 20863 36966 20873 37018
rect 20897 36966 20927 37018
rect 20927 36966 20939 37018
rect 20939 36966 20953 37018
rect 20977 36966 20991 37018
rect 20991 36966 21003 37018
rect 21003 36966 21033 37018
rect 21057 36966 21067 37018
rect 21067 36966 21113 37018
rect 20817 36964 20873 36966
rect 20897 36964 20953 36966
rect 20977 36964 21033 36966
rect 21057 36964 21113 36966
rect 20817 35930 20873 35932
rect 20897 35930 20953 35932
rect 20977 35930 21033 35932
rect 21057 35930 21113 35932
rect 20817 35878 20863 35930
rect 20863 35878 20873 35930
rect 20897 35878 20927 35930
rect 20927 35878 20939 35930
rect 20939 35878 20953 35930
rect 20977 35878 20991 35930
rect 20991 35878 21003 35930
rect 21003 35878 21033 35930
rect 21057 35878 21067 35930
rect 21067 35878 21113 35930
rect 20817 35876 20873 35878
rect 20897 35876 20953 35878
rect 20977 35876 21033 35878
rect 21057 35876 21113 35878
rect 20810 35708 20812 35728
rect 20812 35708 20864 35728
rect 20864 35708 20866 35728
rect 20810 35672 20866 35708
rect 20902 35128 20958 35184
rect 20718 34992 20774 35048
rect 20817 34842 20873 34844
rect 20897 34842 20953 34844
rect 20977 34842 21033 34844
rect 21057 34842 21113 34844
rect 20817 34790 20863 34842
rect 20863 34790 20873 34842
rect 20897 34790 20927 34842
rect 20927 34790 20939 34842
rect 20939 34790 20953 34842
rect 20977 34790 20991 34842
rect 20991 34790 21003 34842
rect 21003 34790 21033 34842
rect 21057 34790 21067 34842
rect 21067 34790 21113 34842
rect 20817 34788 20873 34790
rect 20897 34788 20953 34790
rect 20977 34788 21033 34790
rect 21057 34788 21113 34790
rect 20817 33754 20873 33756
rect 20897 33754 20953 33756
rect 20977 33754 21033 33756
rect 21057 33754 21113 33756
rect 20817 33702 20863 33754
rect 20863 33702 20873 33754
rect 20897 33702 20927 33754
rect 20927 33702 20939 33754
rect 20939 33702 20953 33754
rect 20977 33702 20991 33754
rect 20991 33702 21003 33754
rect 21003 33702 21033 33754
rect 21057 33702 21067 33754
rect 21067 33702 21113 33754
rect 20817 33700 20873 33702
rect 20897 33700 20953 33702
rect 20977 33700 21033 33702
rect 21057 33700 21113 33702
rect 20810 33516 20866 33552
rect 20810 33496 20812 33516
rect 20812 33496 20864 33516
rect 20864 33496 20866 33516
rect 20817 32666 20873 32668
rect 20897 32666 20953 32668
rect 20977 32666 21033 32668
rect 21057 32666 21113 32668
rect 20817 32614 20863 32666
rect 20863 32614 20873 32666
rect 20897 32614 20927 32666
rect 20927 32614 20939 32666
rect 20939 32614 20953 32666
rect 20977 32614 20991 32666
rect 20991 32614 21003 32666
rect 21003 32614 21033 32666
rect 21057 32614 21067 32666
rect 21067 32614 21113 32666
rect 20817 32612 20873 32614
rect 20897 32612 20953 32614
rect 20977 32612 21033 32614
rect 21057 32612 21113 32614
rect 20817 31578 20873 31580
rect 20897 31578 20953 31580
rect 20977 31578 21033 31580
rect 21057 31578 21113 31580
rect 20817 31526 20863 31578
rect 20863 31526 20873 31578
rect 20897 31526 20927 31578
rect 20927 31526 20939 31578
rect 20939 31526 20953 31578
rect 20977 31526 20991 31578
rect 20991 31526 21003 31578
rect 21003 31526 21033 31578
rect 21057 31526 21067 31578
rect 21067 31526 21113 31578
rect 20817 31524 20873 31526
rect 20897 31524 20953 31526
rect 20977 31524 21033 31526
rect 21057 31524 21113 31526
rect 20817 30490 20873 30492
rect 20897 30490 20953 30492
rect 20977 30490 21033 30492
rect 21057 30490 21113 30492
rect 20817 30438 20863 30490
rect 20863 30438 20873 30490
rect 20897 30438 20927 30490
rect 20927 30438 20939 30490
rect 20939 30438 20953 30490
rect 20977 30438 20991 30490
rect 20991 30438 21003 30490
rect 21003 30438 21033 30490
rect 21057 30438 21067 30490
rect 21067 30438 21113 30490
rect 20817 30436 20873 30438
rect 20897 30436 20953 30438
rect 20977 30436 21033 30438
rect 21057 30436 21113 30438
rect 20166 28328 20222 28384
rect 19982 28056 20038 28112
rect 19062 22072 19118 22128
rect 18694 21664 18750 21720
rect 18970 21528 19026 21584
rect 15852 8186 15908 8188
rect 15932 8186 15988 8188
rect 16012 8186 16068 8188
rect 16092 8186 16148 8188
rect 15852 8134 15898 8186
rect 15898 8134 15908 8186
rect 15932 8134 15962 8186
rect 15962 8134 15974 8186
rect 15974 8134 15988 8186
rect 16012 8134 16026 8186
rect 16026 8134 16038 8186
rect 16038 8134 16068 8186
rect 16092 8134 16102 8186
rect 16102 8134 16148 8186
rect 15852 8132 15908 8134
rect 15932 8132 15988 8134
rect 16012 8132 16068 8134
rect 16092 8132 16148 8134
rect 15852 7098 15908 7100
rect 15932 7098 15988 7100
rect 16012 7098 16068 7100
rect 16092 7098 16148 7100
rect 15852 7046 15898 7098
rect 15898 7046 15908 7098
rect 15932 7046 15962 7098
rect 15962 7046 15974 7098
rect 15974 7046 15988 7098
rect 16012 7046 16026 7098
rect 16026 7046 16038 7098
rect 16038 7046 16068 7098
rect 16092 7046 16102 7098
rect 16102 7046 16148 7098
rect 15852 7044 15908 7046
rect 15932 7044 15988 7046
rect 16012 7044 16068 7046
rect 16092 7044 16148 7046
rect 15852 6010 15908 6012
rect 15932 6010 15988 6012
rect 16012 6010 16068 6012
rect 16092 6010 16148 6012
rect 15852 5958 15898 6010
rect 15898 5958 15908 6010
rect 15932 5958 15962 6010
rect 15962 5958 15974 6010
rect 15974 5958 15988 6010
rect 16012 5958 16026 6010
rect 16026 5958 16038 6010
rect 16038 5958 16068 6010
rect 16092 5958 16102 6010
rect 16102 5958 16148 6010
rect 15852 5956 15908 5958
rect 15932 5956 15988 5958
rect 16012 5956 16068 5958
rect 16092 5956 16148 5958
rect 15852 4922 15908 4924
rect 15932 4922 15988 4924
rect 16012 4922 16068 4924
rect 16092 4922 16148 4924
rect 15852 4870 15898 4922
rect 15898 4870 15908 4922
rect 15932 4870 15962 4922
rect 15962 4870 15974 4922
rect 15974 4870 15988 4922
rect 16012 4870 16026 4922
rect 16026 4870 16038 4922
rect 16038 4870 16068 4922
rect 16092 4870 16102 4922
rect 16102 4870 16148 4922
rect 15852 4868 15908 4870
rect 15932 4868 15988 4870
rect 16012 4868 16068 4870
rect 16092 4868 16148 4870
rect 19982 24248 20038 24304
rect 19614 20984 19670 21040
rect 19430 19760 19486 19816
rect 19522 18128 19578 18184
rect 19430 17992 19486 18048
rect 19798 17312 19854 17368
rect 20817 29402 20873 29404
rect 20897 29402 20953 29404
rect 20977 29402 21033 29404
rect 21057 29402 21113 29404
rect 20817 29350 20863 29402
rect 20863 29350 20873 29402
rect 20897 29350 20927 29402
rect 20927 29350 20939 29402
rect 20939 29350 20953 29402
rect 20977 29350 20991 29402
rect 20991 29350 21003 29402
rect 21003 29350 21033 29402
rect 21057 29350 21067 29402
rect 21067 29350 21113 29402
rect 20817 29348 20873 29350
rect 20897 29348 20953 29350
rect 20977 29348 21033 29350
rect 21057 29348 21113 29350
rect 20817 28314 20873 28316
rect 20897 28314 20953 28316
rect 20977 28314 21033 28316
rect 21057 28314 21113 28316
rect 20817 28262 20863 28314
rect 20863 28262 20873 28314
rect 20897 28262 20927 28314
rect 20927 28262 20939 28314
rect 20939 28262 20953 28314
rect 20977 28262 20991 28314
rect 20991 28262 21003 28314
rect 21003 28262 21033 28314
rect 21057 28262 21067 28314
rect 21067 28262 21113 28314
rect 20817 28260 20873 28262
rect 20897 28260 20953 28262
rect 20977 28260 21033 28262
rect 21057 28260 21113 28262
rect 20817 27226 20873 27228
rect 20897 27226 20953 27228
rect 20977 27226 21033 27228
rect 21057 27226 21113 27228
rect 20817 27174 20863 27226
rect 20863 27174 20873 27226
rect 20897 27174 20927 27226
rect 20927 27174 20939 27226
rect 20939 27174 20953 27226
rect 20977 27174 20991 27226
rect 20991 27174 21003 27226
rect 21003 27174 21033 27226
rect 21057 27174 21067 27226
rect 21067 27174 21113 27226
rect 20817 27172 20873 27174
rect 20897 27172 20953 27174
rect 20977 27172 21033 27174
rect 21057 27172 21113 27174
rect 20817 26138 20873 26140
rect 20897 26138 20953 26140
rect 20977 26138 21033 26140
rect 21057 26138 21113 26140
rect 20817 26086 20863 26138
rect 20863 26086 20873 26138
rect 20897 26086 20927 26138
rect 20927 26086 20939 26138
rect 20939 26086 20953 26138
rect 20977 26086 20991 26138
rect 20991 26086 21003 26138
rect 21003 26086 21033 26138
rect 21057 26086 21067 26138
rect 21067 26086 21113 26138
rect 20817 26084 20873 26086
rect 20897 26084 20953 26086
rect 20977 26084 21033 26086
rect 21057 26084 21113 26086
rect 21914 43188 21916 43208
rect 21916 43188 21968 43208
rect 21968 43188 21970 43208
rect 21914 43152 21970 43188
rect 21822 40568 21878 40624
rect 22190 44240 22246 44296
rect 22098 42744 22154 42800
rect 22282 43152 22338 43208
rect 21822 35264 21878 35320
rect 21638 28600 21694 28656
rect 20817 25050 20873 25052
rect 20897 25050 20953 25052
rect 20977 25050 21033 25052
rect 21057 25050 21113 25052
rect 20817 24998 20863 25050
rect 20863 24998 20873 25050
rect 20897 24998 20927 25050
rect 20927 24998 20939 25050
rect 20939 24998 20953 25050
rect 20977 24998 20991 25050
rect 20991 24998 21003 25050
rect 21003 24998 21033 25050
rect 21057 24998 21067 25050
rect 21067 24998 21113 25050
rect 20817 24996 20873 24998
rect 20897 24996 20953 24998
rect 20977 24996 21033 24998
rect 21057 24996 21113 24998
rect 20817 23962 20873 23964
rect 20897 23962 20953 23964
rect 20977 23962 21033 23964
rect 21057 23962 21113 23964
rect 20817 23910 20863 23962
rect 20863 23910 20873 23962
rect 20897 23910 20927 23962
rect 20927 23910 20939 23962
rect 20939 23910 20953 23962
rect 20977 23910 20991 23962
rect 20991 23910 21003 23962
rect 21003 23910 21033 23962
rect 21057 23910 21067 23962
rect 21067 23910 21113 23962
rect 20817 23908 20873 23910
rect 20897 23908 20953 23910
rect 20977 23908 21033 23910
rect 21057 23908 21113 23910
rect 20166 21256 20222 21312
rect 20074 20476 20076 20496
rect 20076 20476 20128 20496
rect 20128 20476 20130 20496
rect 20074 20440 20130 20476
rect 19982 18264 20038 18320
rect 15852 3834 15908 3836
rect 15932 3834 15988 3836
rect 16012 3834 16068 3836
rect 16092 3834 16148 3836
rect 15852 3782 15898 3834
rect 15898 3782 15908 3834
rect 15932 3782 15962 3834
rect 15962 3782 15974 3834
rect 15974 3782 15988 3834
rect 16012 3782 16026 3834
rect 16026 3782 16038 3834
rect 16038 3782 16068 3834
rect 16092 3782 16102 3834
rect 16102 3782 16148 3834
rect 15852 3780 15908 3782
rect 15932 3780 15988 3782
rect 16012 3780 16068 3782
rect 16092 3780 16148 3782
rect 20817 22874 20873 22876
rect 20897 22874 20953 22876
rect 20977 22874 21033 22876
rect 21057 22874 21113 22876
rect 20817 22822 20863 22874
rect 20863 22822 20873 22874
rect 20897 22822 20927 22874
rect 20927 22822 20939 22874
rect 20939 22822 20953 22874
rect 20977 22822 20991 22874
rect 20991 22822 21003 22874
rect 21003 22822 21033 22874
rect 21057 22822 21067 22874
rect 21067 22822 21113 22874
rect 20817 22820 20873 22822
rect 20897 22820 20953 22822
rect 20977 22820 21033 22822
rect 21057 22820 21113 22822
rect 22374 28464 22430 28520
rect 23846 45620 23902 45656
rect 23846 45600 23848 45620
rect 23848 45600 23900 45620
rect 23900 45600 23902 45620
rect 23386 44276 23388 44296
rect 23388 44276 23440 44296
rect 23440 44276 23442 44296
rect 23386 44240 23442 44276
rect 23386 44104 23442 44160
rect 23570 43732 23572 43752
rect 23572 43732 23624 43752
rect 23624 43732 23626 43752
rect 23570 43696 23626 43732
rect 30010 47504 30066 47560
rect 26146 45600 26202 45656
rect 25782 45178 25838 45180
rect 25862 45178 25918 45180
rect 25942 45178 25998 45180
rect 26022 45178 26078 45180
rect 25782 45126 25828 45178
rect 25828 45126 25838 45178
rect 25862 45126 25892 45178
rect 25892 45126 25904 45178
rect 25904 45126 25918 45178
rect 25942 45126 25956 45178
rect 25956 45126 25968 45178
rect 25968 45126 25998 45178
rect 26022 45126 26032 45178
rect 26032 45126 26078 45178
rect 25782 45124 25838 45126
rect 25862 45124 25918 45126
rect 25942 45124 25998 45126
rect 26022 45124 26078 45126
rect 24674 43732 24676 43752
rect 24676 43732 24728 43752
rect 24728 43732 24730 43752
rect 23386 43172 23442 43208
rect 23386 43152 23388 43172
rect 23388 43152 23440 43172
rect 23440 43152 23442 43172
rect 24674 43696 24730 43732
rect 23294 43016 23350 43072
rect 23846 42200 23902 42256
rect 23846 41676 23902 41712
rect 23846 41656 23848 41676
rect 23848 41656 23900 41676
rect 23900 41656 23902 41676
rect 23018 41248 23074 41304
rect 22834 40976 22890 41032
rect 23018 39092 23074 39128
rect 23018 39072 23020 39092
rect 23020 39072 23072 39092
rect 23072 39072 23074 39092
rect 23202 40296 23258 40352
rect 23478 39500 23534 39536
rect 23478 39480 23480 39500
rect 23480 39480 23532 39500
rect 23532 39480 23534 39500
rect 24674 42508 24676 42528
rect 24676 42508 24728 42528
rect 24728 42508 24730 42528
rect 24674 42472 24730 42508
rect 25226 44240 25282 44296
rect 25686 44396 25742 44432
rect 25686 44376 25688 44396
rect 25688 44376 25740 44396
rect 25740 44376 25742 44396
rect 26238 44240 26294 44296
rect 25782 44090 25838 44092
rect 25862 44090 25918 44092
rect 25942 44090 25998 44092
rect 26022 44090 26078 44092
rect 25782 44038 25828 44090
rect 25828 44038 25838 44090
rect 25862 44038 25892 44090
rect 25892 44038 25904 44090
rect 25904 44038 25918 44090
rect 25942 44038 25956 44090
rect 25956 44038 25968 44090
rect 25968 44038 25998 44090
rect 26022 44038 26032 44090
rect 26032 44038 26078 44090
rect 25782 44036 25838 44038
rect 25862 44036 25918 44038
rect 25942 44036 25998 44038
rect 26022 44036 26078 44038
rect 24950 40568 25006 40624
rect 24490 39616 24546 39672
rect 20817 21786 20873 21788
rect 20897 21786 20953 21788
rect 20977 21786 21033 21788
rect 21057 21786 21113 21788
rect 20817 21734 20863 21786
rect 20863 21734 20873 21786
rect 20897 21734 20927 21786
rect 20927 21734 20939 21786
rect 20939 21734 20953 21786
rect 20977 21734 20991 21786
rect 20991 21734 21003 21786
rect 21003 21734 21033 21786
rect 21057 21734 21067 21786
rect 21067 21734 21113 21786
rect 20817 21732 20873 21734
rect 20897 21732 20953 21734
rect 20977 21732 21033 21734
rect 21057 21732 21113 21734
rect 20810 21392 20866 21448
rect 20626 20868 20682 20904
rect 20626 20848 20628 20868
rect 20628 20848 20680 20868
rect 20680 20848 20682 20868
rect 20817 20698 20873 20700
rect 20897 20698 20953 20700
rect 20977 20698 21033 20700
rect 21057 20698 21113 20700
rect 20817 20646 20863 20698
rect 20863 20646 20873 20698
rect 20897 20646 20927 20698
rect 20927 20646 20939 20698
rect 20939 20646 20953 20698
rect 20977 20646 20991 20698
rect 20991 20646 21003 20698
rect 21003 20646 21033 20698
rect 21057 20646 21067 20698
rect 21067 20646 21113 20698
rect 20817 20644 20873 20646
rect 20897 20644 20953 20646
rect 20977 20644 21033 20646
rect 21057 20644 21113 20646
rect 20817 19610 20873 19612
rect 20897 19610 20953 19612
rect 20977 19610 21033 19612
rect 21057 19610 21113 19612
rect 20817 19558 20863 19610
rect 20863 19558 20873 19610
rect 20897 19558 20927 19610
rect 20927 19558 20939 19610
rect 20939 19558 20953 19610
rect 20977 19558 20991 19610
rect 20991 19558 21003 19610
rect 21003 19558 21033 19610
rect 21057 19558 21067 19610
rect 21067 19558 21113 19610
rect 20817 19556 20873 19558
rect 20897 19556 20953 19558
rect 20977 19556 21033 19558
rect 21057 19556 21113 19558
rect 20350 17740 20406 17776
rect 20350 17720 20352 17740
rect 20352 17720 20404 17740
rect 20404 17720 20406 17740
rect 20534 17584 20590 17640
rect 20626 14864 20682 14920
rect 20817 18522 20873 18524
rect 20897 18522 20953 18524
rect 20977 18522 21033 18524
rect 21057 18522 21113 18524
rect 20817 18470 20863 18522
rect 20863 18470 20873 18522
rect 20897 18470 20927 18522
rect 20927 18470 20939 18522
rect 20939 18470 20953 18522
rect 20977 18470 20991 18522
rect 20991 18470 21003 18522
rect 21003 18470 21033 18522
rect 21057 18470 21067 18522
rect 21067 18470 21113 18522
rect 20817 18468 20873 18470
rect 20897 18468 20953 18470
rect 20977 18468 21033 18470
rect 21057 18468 21113 18470
rect 21086 17856 21142 17912
rect 20810 17604 20866 17640
rect 20810 17584 20812 17604
rect 20812 17584 20864 17604
rect 20864 17584 20866 17604
rect 20817 17434 20873 17436
rect 20897 17434 20953 17436
rect 20977 17434 21033 17436
rect 21057 17434 21113 17436
rect 20817 17382 20863 17434
rect 20863 17382 20873 17434
rect 20897 17382 20927 17434
rect 20927 17382 20939 17434
rect 20939 17382 20953 17434
rect 20977 17382 20991 17434
rect 20991 17382 21003 17434
rect 21003 17382 21033 17434
rect 21057 17382 21067 17434
rect 21067 17382 21113 17434
rect 20817 17380 20873 17382
rect 20897 17380 20953 17382
rect 20977 17380 21033 17382
rect 21057 17380 21113 17382
rect 21270 17720 21326 17776
rect 21270 16768 21326 16824
rect 21178 16632 21234 16688
rect 20817 16346 20873 16348
rect 20897 16346 20953 16348
rect 20977 16346 21033 16348
rect 21057 16346 21113 16348
rect 20817 16294 20863 16346
rect 20863 16294 20873 16346
rect 20897 16294 20927 16346
rect 20927 16294 20939 16346
rect 20939 16294 20953 16346
rect 20977 16294 20991 16346
rect 20991 16294 21003 16346
rect 21003 16294 21033 16346
rect 21057 16294 21067 16346
rect 21067 16294 21113 16346
rect 20817 16292 20873 16294
rect 20897 16292 20953 16294
rect 20977 16292 21033 16294
rect 21057 16292 21113 16294
rect 20817 15258 20873 15260
rect 20897 15258 20953 15260
rect 20977 15258 21033 15260
rect 21057 15258 21113 15260
rect 20817 15206 20863 15258
rect 20863 15206 20873 15258
rect 20897 15206 20927 15258
rect 20927 15206 20939 15258
rect 20939 15206 20953 15258
rect 20977 15206 20991 15258
rect 20991 15206 21003 15258
rect 21003 15206 21033 15258
rect 21057 15206 21067 15258
rect 21067 15206 21113 15258
rect 20817 15204 20873 15206
rect 20897 15204 20953 15206
rect 20977 15204 21033 15206
rect 21057 15204 21113 15206
rect 21546 21392 21602 21448
rect 21546 20848 21602 20904
rect 21730 20440 21786 20496
rect 21914 22480 21970 22536
rect 22006 19352 22062 19408
rect 21638 17720 21694 17776
rect 21454 16652 21510 16688
rect 21454 16632 21456 16652
rect 21456 16632 21508 16652
rect 21508 16632 21510 16652
rect 20817 14170 20873 14172
rect 20897 14170 20953 14172
rect 20977 14170 21033 14172
rect 21057 14170 21113 14172
rect 20817 14118 20863 14170
rect 20863 14118 20873 14170
rect 20897 14118 20927 14170
rect 20927 14118 20939 14170
rect 20939 14118 20953 14170
rect 20977 14118 20991 14170
rect 20991 14118 21003 14170
rect 21003 14118 21033 14170
rect 21057 14118 21067 14170
rect 21067 14118 21113 14170
rect 20817 14116 20873 14118
rect 20897 14116 20953 14118
rect 20977 14116 21033 14118
rect 21057 14116 21113 14118
rect 21270 14356 21272 14376
rect 21272 14356 21324 14376
rect 21324 14356 21326 14376
rect 21270 14320 21326 14356
rect 20817 13082 20873 13084
rect 20897 13082 20953 13084
rect 20977 13082 21033 13084
rect 21057 13082 21113 13084
rect 20817 13030 20863 13082
rect 20863 13030 20873 13082
rect 20897 13030 20927 13082
rect 20927 13030 20939 13082
rect 20939 13030 20953 13082
rect 20977 13030 20991 13082
rect 20991 13030 21003 13082
rect 21003 13030 21033 13082
rect 21057 13030 21067 13082
rect 21067 13030 21113 13082
rect 20817 13028 20873 13030
rect 20897 13028 20953 13030
rect 20977 13028 21033 13030
rect 21057 13028 21113 13030
rect 20718 12552 20774 12608
rect 20442 10648 20498 10704
rect 20817 11994 20873 11996
rect 20897 11994 20953 11996
rect 20977 11994 21033 11996
rect 21057 11994 21113 11996
rect 20817 11942 20863 11994
rect 20863 11942 20873 11994
rect 20897 11942 20927 11994
rect 20927 11942 20939 11994
rect 20939 11942 20953 11994
rect 20977 11942 20991 11994
rect 20991 11942 21003 11994
rect 21003 11942 21033 11994
rect 21057 11942 21067 11994
rect 21067 11942 21113 11994
rect 20817 11940 20873 11942
rect 20897 11940 20953 11942
rect 20977 11940 21033 11942
rect 21057 11940 21113 11942
rect 20817 10906 20873 10908
rect 20897 10906 20953 10908
rect 20977 10906 21033 10908
rect 21057 10906 21113 10908
rect 20817 10854 20863 10906
rect 20863 10854 20873 10906
rect 20897 10854 20927 10906
rect 20927 10854 20939 10906
rect 20939 10854 20953 10906
rect 20977 10854 20991 10906
rect 20991 10854 21003 10906
rect 21003 10854 21033 10906
rect 21057 10854 21067 10906
rect 21067 10854 21113 10906
rect 20817 10852 20873 10854
rect 20897 10852 20953 10854
rect 20977 10852 21033 10854
rect 21057 10852 21113 10854
rect 20817 9818 20873 9820
rect 20897 9818 20953 9820
rect 20977 9818 21033 9820
rect 21057 9818 21113 9820
rect 20817 9766 20863 9818
rect 20863 9766 20873 9818
rect 20897 9766 20927 9818
rect 20927 9766 20939 9818
rect 20939 9766 20953 9818
rect 20977 9766 20991 9818
rect 20991 9766 21003 9818
rect 21003 9766 21033 9818
rect 21057 9766 21067 9818
rect 21067 9766 21113 9818
rect 20817 9764 20873 9766
rect 20897 9764 20953 9766
rect 20977 9764 21033 9766
rect 21057 9764 21113 9766
rect 20534 9152 20590 9208
rect 20902 9016 20958 9072
rect 21454 11056 21510 11112
rect 21178 9016 21234 9072
rect 20817 8730 20873 8732
rect 20897 8730 20953 8732
rect 20977 8730 21033 8732
rect 21057 8730 21113 8732
rect 20817 8678 20863 8730
rect 20863 8678 20873 8730
rect 20897 8678 20927 8730
rect 20927 8678 20939 8730
rect 20939 8678 20953 8730
rect 20977 8678 20991 8730
rect 20991 8678 21003 8730
rect 21003 8678 21033 8730
rect 21057 8678 21067 8730
rect 21067 8678 21113 8730
rect 20817 8676 20873 8678
rect 20897 8676 20953 8678
rect 20977 8676 21033 8678
rect 21057 8676 21113 8678
rect 20817 7642 20873 7644
rect 20897 7642 20953 7644
rect 20977 7642 21033 7644
rect 21057 7642 21113 7644
rect 20817 7590 20863 7642
rect 20863 7590 20873 7642
rect 20897 7590 20927 7642
rect 20927 7590 20939 7642
rect 20939 7590 20953 7642
rect 20977 7590 20991 7642
rect 20991 7590 21003 7642
rect 21003 7590 21033 7642
rect 21057 7590 21067 7642
rect 21067 7590 21113 7642
rect 20817 7588 20873 7590
rect 20897 7588 20953 7590
rect 20977 7588 21033 7590
rect 21057 7588 21113 7590
rect 15852 2746 15908 2748
rect 15932 2746 15988 2748
rect 16012 2746 16068 2748
rect 16092 2746 16148 2748
rect 15852 2694 15898 2746
rect 15898 2694 15908 2746
rect 15932 2694 15962 2746
rect 15962 2694 15974 2746
rect 15974 2694 15988 2746
rect 16012 2694 16026 2746
rect 16026 2694 16038 2746
rect 16038 2694 16068 2746
rect 16092 2694 16102 2746
rect 16102 2694 16148 2746
rect 15852 2692 15908 2694
rect 15932 2692 15988 2694
rect 16012 2692 16068 2694
rect 16092 2692 16148 2694
rect 20817 6554 20873 6556
rect 20897 6554 20953 6556
rect 20977 6554 21033 6556
rect 21057 6554 21113 6556
rect 20817 6502 20863 6554
rect 20863 6502 20873 6554
rect 20897 6502 20927 6554
rect 20927 6502 20939 6554
rect 20939 6502 20953 6554
rect 20977 6502 20991 6554
rect 20991 6502 21003 6554
rect 21003 6502 21033 6554
rect 21057 6502 21067 6554
rect 21067 6502 21113 6554
rect 20817 6500 20873 6502
rect 20897 6500 20953 6502
rect 20977 6500 21033 6502
rect 21057 6500 21113 6502
rect 20994 5652 21036 5672
rect 21036 5652 21050 5672
rect 20994 5616 21050 5652
rect 21362 5752 21418 5808
rect 20817 5466 20873 5468
rect 20897 5466 20953 5468
rect 20977 5466 21033 5468
rect 21057 5466 21113 5468
rect 20817 5414 20863 5466
rect 20863 5414 20873 5466
rect 20897 5414 20927 5466
rect 20927 5414 20939 5466
rect 20939 5414 20953 5466
rect 20977 5414 20991 5466
rect 20991 5414 21003 5466
rect 21003 5414 21033 5466
rect 21057 5414 21067 5466
rect 21067 5414 21113 5466
rect 20817 5412 20873 5414
rect 20897 5412 20953 5414
rect 20977 5412 21033 5414
rect 21057 5412 21113 5414
rect 21454 5616 21510 5672
rect 20817 4378 20873 4380
rect 20897 4378 20953 4380
rect 20977 4378 21033 4380
rect 21057 4378 21113 4380
rect 20817 4326 20863 4378
rect 20863 4326 20873 4378
rect 20897 4326 20927 4378
rect 20927 4326 20939 4378
rect 20939 4326 20953 4378
rect 20977 4326 20991 4378
rect 20991 4326 21003 4378
rect 21003 4326 21033 4378
rect 21057 4326 21067 4378
rect 21067 4326 21113 4378
rect 20817 4324 20873 4326
rect 20897 4324 20953 4326
rect 20977 4324 21033 4326
rect 21057 4324 21113 4326
rect 22190 14900 22192 14920
rect 22192 14900 22244 14920
rect 22244 14900 22246 14920
rect 22190 14864 22246 14900
rect 21822 11872 21878 11928
rect 22098 11600 22154 11656
rect 22190 9172 22246 9208
rect 22190 9152 22192 9172
rect 22192 9152 22244 9172
rect 22244 9152 22246 9172
rect 22190 9036 22246 9072
rect 22190 9016 22192 9036
rect 22192 9016 22244 9036
rect 22244 9016 22246 9036
rect 22282 5752 22338 5808
rect 23202 14320 23258 14376
rect 23018 11872 23074 11928
rect 23110 8492 23166 8528
rect 23110 8472 23112 8492
rect 23112 8472 23164 8492
rect 23164 8472 23166 8492
rect 24490 37204 24492 37224
rect 24492 37204 24544 37224
rect 24544 37204 24546 37224
rect 24490 37168 24546 37204
rect 25042 38936 25098 38992
rect 25782 43002 25838 43004
rect 25862 43002 25918 43004
rect 25942 43002 25998 43004
rect 26022 43002 26078 43004
rect 25782 42950 25828 43002
rect 25828 42950 25838 43002
rect 25862 42950 25892 43002
rect 25892 42950 25904 43002
rect 25904 42950 25918 43002
rect 25942 42950 25956 43002
rect 25956 42950 25968 43002
rect 25968 42950 25998 43002
rect 26022 42950 26032 43002
rect 26032 42950 26078 43002
rect 25782 42948 25838 42950
rect 25862 42948 25918 42950
rect 25942 42948 25998 42950
rect 26022 42948 26078 42950
rect 25502 41556 25504 41576
rect 25504 41556 25556 41576
rect 25556 41556 25558 41576
rect 25502 41520 25558 41556
rect 25502 40588 25558 40624
rect 25502 40568 25504 40588
rect 25504 40568 25556 40588
rect 25556 40568 25558 40588
rect 25782 41914 25838 41916
rect 25862 41914 25918 41916
rect 25942 41914 25998 41916
rect 26022 41914 26078 41916
rect 25782 41862 25828 41914
rect 25828 41862 25838 41914
rect 25862 41862 25892 41914
rect 25892 41862 25904 41914
rect 25904 41862 25918 41914
rect 25942 41862 25956 41914
rect 25956 41862 25968 41914
rect 25968 41862 25998 41914
rect 26022 41862 26032 41914
rect 26032 41862 26078 41914
rect 25782 41860 25838 41862
rect 25862 41860 25918 41862
rect 25942 41860 25998 41862
rect 26022 41860 26078 41862
rect 25686 40976 25742 41032
rect 25782 40826 25838 40828
rect 25862 40826 25918 40828
rect 25942 40826 25998 40828
rect 26022 40826 26078 40828
rect 25782 40774 25828 40826
rect 25828 40774 25838 40826
rect 25862 40774 25892 40826
rect 25892 40774 25904 40826
rect 25904 40774 25918 40826
rect 25942 40774 25956 40826
rect 25956 40774 25968 40826
rect 25968 40774 25998 40826
rect 26022 40774 26032 40826
rect 26032 40774 26078 40826
rect 25782 40772 25838 40774
rect 25862 40772 25918 40774
rect 25942 40772 25998 40774
rect 26022 40772 26078 40774
rect 25782 39738 25838 39740
rect 25862 39738 25918 39740
rect 25942 39738 25998 39740
rect 26022 39738 26078 39740
rect 25782 39686 25828 39738
rect 25828 39686 25838 39738
rect 25862 39686 25892 39738
rect 25892 39686 25904 39738
rect 25904 39686 25918 39738
rect 25942 39686 25956 39738
rect 25956 39686 25968 39738
rect 25968 39686 25998 39738
rect 26022 39686 26032 39738
rect 26032 39686 26078 39738
rect 25782 39684 25838 39686
rect 25862 39684 25918 39686
rect 25942 39684 25998 39686
rect 26022 39684 26078 39686
rect 26422 41268 26478 41304
rect 26422 41248 26424 41268
rect 26424 41248 26476 41268
rect 26476 41248 26478 41268
rect 25782 38650 25838 38652
rect 25862 38650 25918 38652
rect 25942 38650 25998 38652
rect 26022 38650 26078 38652
rect 25782 38598 25828 38650
rect 25828 38598 25838 38650
rect 25862 38598 25892 38650
rect 25892 38598 25904 38650
rect 25904 38598 25918 38650
rect 25942 38598 25956 38650
rect 25956 38598 25968 38650
rect 25968 38598 25998 38650
rect 26022 38598 26032 38650
rect 26032 38598 26078 38650
rect 25782 38596 25838 38598
rect 25862 38596 25918 38598
rect 25942 38596 25998 38598
rect 26022 38596 26078 38598
rect 25782 37562 25838 37564
rect 25862 37562 25918 37564
rect 25942 37562 25998 37564
rect 26022 37562 26078 37564
rect 25782 37510 25828 37562
rect 25828 37510 25838 37562
rect 25862 37510 25892 37562
rect 25892 37510 25904 37562
rect 25904 37510 25918 37562
rect 25942 37510 25956 37562
rect 25956 37510 25968 37562
rect 25968 37510 25998 37562
rect 26022 37510 26032 37562
rect 26032 37510 26078 37562
rect 25782 37508 25838 37510
rect 25862 37508 25918 37510
rect 25942 37508 25998 37510
rect 26022 37508 26078 37510
rect 25782 36474 25838 36476
rect 25862 36474 25918 36476
rect 25942 36474 25998 36476
rect 26022 36474 26078 36476
rect 25782 36422 25828 36474
rect 25828 36422 25838 36474
rect 25862 36422 25892 36474
rect 25892 36422 25904 36474
rect 25904 36422 25918 36474
rect 25942 36422 25956 36474
rect 25956 36422 25968 36474
rect 25968 36422 25998 36474
rect 26022 36422 26032 36474
rect 26032 36422 26078 36474
rect 25782 36420 25838 36422
rect 25862 36420 25918 36422
rect 25942 36420 25998 36422
rect 26022 36420 26078 36422
rect 25782 35386 25838 35388
rect 25862 35386 25918 35388
rect 25942 35386 25998 35388
rect 26022 35386 26078 35388
rect 25782 35334 25828 35386
rect 25828 35334 25838 35386
rect 25862 35334 25892 35386
rect 25892 35334 25904 35386
rect 25904 35334 25918 35386
rect 25942 35334 25956 35386
rect 25956 35334 25968 35386
rect 25968 35334 25998 35386
rect 26022 35334 26032 35386
rect 26032 35334 26078 35386
rect 25782 35332 25838 35334
rect 25862 35332 25918 35334
rect 25942 35332 25998 35334
rect 26022 35332 26078 35334
rect 25782 34298 25838 34300
rect 25862 34298 25918 34300
rect 25942 34298 25998 34300
rect 26022 34298 26078 34300
rect 25782 34246 25828 34298
rect 25828 34246 25838 34298
rect 25862 34246 25892 34298
rect 25892 34246 25904 34298
rect 25904 34246 25918 34298
rect 25942 34246 25956 34298
rect 25956 34246 25968 34298
rect 25968 34246 25998 34298
rect 26022 34246 26032 34298
rect 26032 34246 26078 34298
rect 25782 34244 25838 34246
rect 25862 34244 25918 34246
rect 25942 34244 25998 34246
rect 26022 34244 26078 34246
rect 23938 17856 23994 17912
rect 23938 17720 23994 17776
rect 24858 28600 24914 28656
rect 25782 33210 25838 33212
rect 25862 33210 25918 33212
rect 25942 33210 25998 33212
rect 26022 33210 26078 33212
rect 25782 33158 25828 33210
rect 25828 33158 25838 33210
rect 25862 33158 25892 33210
rect 25892 33158 25904 33210
rect 25904 33158 25918 33210
rect 25942 33158 25956 33210
rect 25956 33158 25968 33210
rect 25968 33158 25998 33210
rect 26022 33158 26032 33210
rect 26032 33158 26078 33210
rect 25782 33156 25838 33158
rect 25862 33156 25918 33158
rect 25942 33156 25998 33158
rect 26022 33156 26078 33158
rect 26790 40024 26846 40080
rect 26698 39072 26754 39128
rect 27526 45364 27528 45384
rect 27528 45364 27580 45384
rect 27580 45364 27582 45384
rect 27526 45328 27582 45364
rect 27434 44920 27490 44976
rect 27434 42764 27490 42800
rect 27434 42744 27436 42764
rect 27436 42744 27488 42764
rect 27488 42744 27490 42764
rect 27434 42236 27436 42256
rect 27436 42236 27488 42256
rect 27488 42236 27490 42256
rect 27434 42200 27490 42236
rect 27434 41520 27490 41576
rect 27342 40296 27398 40352
rect 27710 45348 27766 45384
rect 27710 45328 27712 45348
rect 27712 45328 27764 45348
rect 27764 45328 27766 45348
rect 27710 43152 27766 43208
rect 27894 46824 27950 46880
rect 28906 46008 28962 46064
rect 27526 39516 27528 39536
rect 27528 39516 27580 39536
rect 27580 39516 27582 39536
rect 27526 39480 27582 39516
rect 25782 32122 25838 32124
rect 25862 32122 25918 32124
rect 25942 32122 25998 32124
rect 26022 32122 26078 32124
rect 25782 32070 25828 32122
rect 25828 32070 25838 32122
rect 25862 32070 25892 32122
rect 25892 32070 25904 32122
rect 25904 32070 25918 32122
rect 25942 32070 25956 32122
rect 25956 32070 25968 32122
rect 25968 32070 25998 32122
rect 26022 32070 26032 32122
rect 26032 32070 26078 32122
rect 25782 32068 25838 32070
rect 25862 32068 25918 32070
rect 25942 32068 25998 32070
rect 26022 32068 26078 32070
rect 25782 31034 25838 31036
rect 25862 31034 25918 31036
rect 25942 31034 25998 31036
rect 26022 31034 26078 31036
rect 25782 30982 25828 31034
rect 25828 30982 25838 31034
rect 25862 30982 25892 31034
rect 25892 30982 25904 31034
rect 25904 30982 25918 31034
rect 25942 30982 25956 31034
rect 25956 30982 25968 31034
rect 25968 30982 25998 31034
rect 26022 30982 26032 31034
rect 26032 30982 26078 31034
rect 25782 30980 25838 30982
rect 25862 30980 25918 30982
rect 25942 30980 25998 30982
rect 26022 30980 26078 30982
rect 25782 29946 25838 29948
rect 25862 29946 25918 29948
rect 25942 29946 25998 29948
rect 26022 29946 26078 29948
rect 25782 29894 25828 29946
rect 25828 29894 25838 29946
rect 25862 29894 25892 29946
rect 25892 29894 25904 29946
rect 25904 29894 25918 29946
rect 25942 29894 25956 29946
rect 25956 29894 25968 29946
rect 25968 29894 25998 29946
rect 26022 29894 26032 29946
rect 26032 29894 26078 29946
rect 25782 29892 25838 29894
rect 25862 29892 25918 29894
rect 25942 29892 25998 29894
rect 26022 29892 26078 29894
rect 25782 28858 25838 28860
rect 25862 28858 25918 28860
rect 25942 28858 25998 28860
rect 26022 28858 26078 28860
rect 25782 28806 25828 28858
rect 25828 28806 25838 28858
rect 25862 28806 25892 28858
rect 25892 28806 25904 28858
rect 25904 28806 25918 28858
rect 25942 28806 25956 28858
rect 25956 28806 25968 28858
rect 25968 28806 25998 28858
rect 26022 28806 26032 28858
rect 26032 28806 26078 28858
rect 25782 28804 25838 28806
rect 25862 28804 25918 28806
rect 25942 28804 25998 28806
rect 26022 28804 26078 28806
rect 25782 27770 25838 27772
rect 25862 27770 25918 27772
rect 25942 27770 25998 27772
rect 26022 27770 26078 27772
rect 25782 27718 25828 27770
rect 25828 27718 25838 27770
rect 25862 27718 25892 27770
rect 25892 27718 25904 27770
rect 25904 27718 25918 27770
rect 25942 27718 25956 27770
rect 25956 27718 25968 27770
rect 25968 27718 25998 27770
rect 26022 27718 26032 27770
rect 26032 27718 26078 27770
rect 25782 27716 25838 27718
rect 25862 27716 25918 27718
rect 25942 27716 25998 27718
rect 26022 27716 26078 27718
rect 24766 21256 24822 21312
rect 24766 19780 24822 19816
rect 24766 19760 24768 19780
rect 24768 19760 24820 19780
rect 24820 19760 24822 19780
rect 24674 19352 24730 19408
rect 24858 18708 24860 18728
rect 24860 18708 24912 18728
rect 24912 18708 24914 18728
rect 24858 18672 24914 18708
rect 24766 18264 24822 18320
rect 25318 24268 25374 24304
rect 25318 24248 25320 24268
rect 25320 24248 25372 24268
rect 25372 24248 25374 24268
rect 27342 37204 27344 37224
rect 27344 37204 27396 37224
rect 27396 37204 27398 37224
rect 27342 37168 27398 37204
rect 27250 33496 27306 33552
rect 28446 45464 28502 45520
rect 28354 41656 28410 41712
rect 28170 41112 28226 41168
rect 28262 40160 28318 40216
rect 28354 40024 28410 40080
rect 29182 42472 29238 42528
rect 30010 44512 30066 44568
rect 30102 43968 30158 44024
rect 30010 43868 30012 43888
rect 30012 43868 30064 43888
rect 30064 43868 30066 43888
rect 30010 43832 30066 43868
rect 30010 43052 30012 43072
rect 30012 43052 30064 43072
rect 30064 43052 30066 43072
rect 30010 43016 30066 43052
rect 30010 42336 30066 42392
rect 30010 41656 30066 41712
rect 30010 40840 30066 40896
rect 29918 40432 29974 40488
rect 28906 38664 28962 38720
rect 30102 40160 30158 40216
rect 30010 39344 30066 39400
rect 28906 36488 28962 36544
rect 30102 37848 30158 37904
rect 30010 37168 30066 37224
rect 30010 35672 30066 35728
rect 28906 34992 28962 35048
rect 28446 34176 28502 34232
rect 28906 33496 28962 33552
rect 30010 32680 30066 32736
rect 30102 32000 30158 32056
rect 30010 31320 30066 31376
rect 30102 30504 30158 30560
rect 30010 29824 30066 29880
rect 30010 29028 30066 29064
rect 30010 29008 30012 29028
rect 30012 29008 30064 29028
rect 30064 29008 30066 29028
rect 30010 28364 30012 28384
rect 30012 28364 30064 28384
rect 30064 28364 30066 28384
rect 30010 28328 30066 28364
rect 30010 27512 30066 27568
rect 25782 26682 25838 26684
rect 25862 26682 25918 26684
rect 25942 26682 25998 26684
rect 26022 26682 26078 26684
rect 25782 26630 25828 26682
rect 25828 26630 25838 26682
rect 25862 26630 25892 26682
rect 25892 26630 25904 26682
rect 25904 26630 25918 26682
rect 25942 26630 25956 26682
rect 25956 26630 25968 26682
rect 25968 26630 25998 26682
rect 26022 26630 26032 26682
rect 26032 26630 26078 26682
rect 25782 26628 25838 26630
rect 25862 26628 25918 26630
rect 25942 26628 25998 26630
rect 26022 26628 26078 26630
rect 30010 26852 30066 26888
rect 30010 26832 30012 26852
rect 30012 26832 30064 26852
rect 30064 26832 30066 26852
rect 25782 25594 25838 25596
rect 25862 25594 25918 25596
rect 25942 25594 25998 25596
rect 26022 25594 26078 25596
rect 25782 25542 25828 25594
rect 25828 25542 25838 25594
rect 25862 25542 25892 25594
rect 25892 25542 25904 25594
rect 25904 25542 25918 25594
rect 25942 25542 25956 25594
rect 25956 25542 25968 25594
rect 25968 25542 25998 25594
rect 26022 25542 26032 25594
rect 26032 25542 26078 25594
rect 25782 25540 25838 25542
rect 25862 25540 25918 25542
rect 25942 25540 25998 25542
rect 26022 25540 26078 25542
rect 25782 24506 25838 24508
rect 25862 24506 25918 24508
rect 25942 24506 25998 24508
rect 26022 24506 26078 24508
rect 25782 24454 25828 24506
rect 25828 24454 25838 24506
rect 25862 24454 25892 24506
rect 25892 24454 25904 24506
rect 25904 24454 25918 24506
rect 25942 24454 25956 24506
rect 25956 24454 25968 24506
rect 25968 24454 25998 24506
rect 26022 24454 26032 24506
rect 26032 24454 26078 24506
rect 25782 24452 25838 24454
rect 25862 24452 25918 24454
rect 25942 24452 25998 24454
rect 26022 24452 26078 24454
rect 25686 23568 25742 23624
rect 25782 23418 25838 23420
rect 25862 23418 25918 23420
rect 25942 23418 25998 23420
rect 26022 23418 26078 23420
rect 25782 23366 25828 23418
rect 25828 23366 25838 23418
rect 25862 23366 25892 23418
rect 25892 23366 25904 23418
rect 25904 23366 25918 23418
rect 25942 23366 25956 23418
rect 25956 23366 25968 23418
rect 25968 23366 25998 23418
rect 26022 23366 26032 23418
rect 26032 23366 26078 23418
rect 25782 23364 25838 23366
rect 25862 23364 25918 23366
rect 25942 23364 25998 23366
rect 26022 23364 26078 23366
rect 25782 22330 25838 22332
rect 25862 22330 25918 22332
rect 25942 22330 25998 22332
rect 26022 22330 26078 22332
rect 25782 22278 25828 22330
rect 25828 22278 25838 22330
rect 25862 22278 25892 22330
rect 25892 22278 25904 22330
rect 25904 22278 25918 22330
rect 25942 22278 25956 22330
rect 25956 22278 25968 22330
rect 25968 22278 25998 22330
rect 26022 22278 26032 22330
rect 26032 22278 26078 22330
rect 25782 22276 25838 22278
rect 25862 22276 25918 22278
rect 25942 22276 25998 22278
rect 26022 22276 26078 22278
rect 25782 21242 25838 21244
rect 25862 21242 25918 21244
rect 25942 21242 25998 21244
rect 26022 21242 26078 21244
rect 25782 21190 25828 21242
rect 25828 21190 25838 21242
rect 25862 21190 25892 21242
rect 25892 21190 25904 21242
rect 25904 21190 25918 21242
rect 25942 21190 25956 21242
rect 25956 21190 25968 21242
rect 25968 21190 25998 21242
rect 26022 21190 26032 21242
rect 26032 21190 26078 21242
rect 25782 21188 25838 21190
rect 25862 21188 25918 21190
rect 25942 21188 25998 21190
rect 26022 21188 26078 21190
rect 26238 20984 26294 21040
rect 25782 20154 25838 20156
rect 25862 20154 25918 20156
rect 25942 20154 25998 20156
rect 26022 20154 26078 20156
rect 25782 20102 25828 20154
rect 25828 20102 25838 20154
rect 25862 20102 25892 20154
rect 25892 20102 25904 20154
rect 25904 20102 25918 20154
rect 25942 20102 25956 20154
rect 25956 20102 25968 20154
rect 25968 20102 25998 20154
rect 26022 20102 26032 20154
rect 26032 20102 26078 20154
rect 25782 20100 25838 20102
rect 25862 20100 25918 20102
rect 25942 20100 25998 20102
rect 26022 20100 26078 20102
rect 30010 26188 30012 26208
rect 30012 26188 30064 26208
rect 30064 26188 30066 26208
rect 30010 26152 30066 26188
rect 26882 24248 26938 24304
rect 25782 19066 25838 19068
rect 25862 19066 25918 19068
rect 25942 19066 25998 19068
rect 26022 19066 26078 19068
rect 25782 19014 25828 19066
rect 25828 19014 25838 19066
rect 25862 19014 25892 19066
rect 25892 19014 25904 19066
rect 25904 19014 25918 19066
rect 25942 19014 25956 19066
rect 25956 19014 25968 19066
rect 25968 19014 25998 19066
rect 26022 19014 26032 19066
rect 26032 19014 26078 19066
rect 25782 19012 25838 19014
rect 25862 19012 25918 19014
rect 25942 19012 25998 19014
rect 26022 19012 26078 19014
rect 25594 17992 25650 18048
rect 25782 17978 25838 17980
rect 25862 17978 25918 17980
rect 25942 17978 25998 17980
rect 26022 17978 26078 17980
rect 25782 17926 25828 17978
rect 25828 17926 25838 17978
rect 25862 17926 25892 17978
rect 25892 17926 25904 17978
rect 25904 17926 25918 17978
rect 25942 17926 25956 17978
rect 25956 17926 25968 17978
rect 25968 17926 25998 17978
rect 26022 17926 26032 17978
rect 26032 17926 26078 17978
rect 25782 17924 25838 17926
rect 25862 17924 25918 17926
rect 25942 17924 25998 17926
rect 26022 17924 26078 17926
rect 26054 17720 26110 17776
rect 25782 16890 25838 16892
rect 25862 16890 25918 16892
rect 25942 16890 25998 16892
rect 26022 16890 26078 16892
rect 25782 16838 25828 16890
rect 25828 16838 25838 16890
rect 25862 16838 25892 16890
rect 25892 16838 25904 16890
rect 25904 16838 25918 16890
rect 25942 16838 25956 16890
rect 25956 16838 25968 16890
rect 25968 16838 25998 16890
rect 26022 16838 26032 16890
rect 26032 16838 26078 16890
rect 25782 16836 25838 16838
rect 25862 16836 25918 16838
rect 25942 16836 25998 16838
rect 26022 16836 26078 16838
rect 26422 17584 26478 17640
rect 25782 15802 25838 15804
rect 25862 15802 25918 15804
rect 25942 15802 25998 15804
rect 26022 15802 26078 15804
rect 25782 15750 25828 15802
rect 25828 15750 25838 15802
rect 25862 15750 25892 15802
rect 25892 15750 25904 15802
rect 25904 15750 25918 15802
rect 25942 15750 25956 15802
rect 25956 15750 25968 15802
rect 25968 15750 25998 15802
rect 26022 15750 26032 15802
rect 26032 15750 26078 15802
rect 25782 15748 25838 15750
rect 25862 15748 25918 15750
rect 25942 15748 25998 15750
rect 26022 15748 26078 15750
rect 25782 14714 25838 14716
rect 25862 14714 25918 14716
rect 25942 14714 25998 14716
rect 26022 14714 26078 14716
rect 25782 14662 25828 14714
rect 25828 14662 25838 14714
rect 25862 14662 25892 14714
rect 25892 14662 25904 14714
rect 25904 14662 25918 14714
rect 25942 14662 25956 14714
rect 25956 14662 25968 14714
rect 25968 14662 25998 14714
rect 26022 14662 26032 14714
rect 26032 14662 26078 14714
rect 25782 14660 25838 14662
rect 25862 14660 25918 14662
rect 25942 14660 25998 14662
rect 26022 14660 26078 14662
rect 25782 13626 25838 13628
rect 25862 13626 25918 13628
rect 25942 13626 25998 13628
rect 26022 13626 26078 13628
rect 25782 13574 25828 13626
rect 25828 13574 25838 13626
rect 25862 13574 25892 13626
rect 25892 13574 25904 13626
rect 25904 13574 25918 13626
rect 25942 13574 25956 13626
rect 25956 13574 25968 13626
rect 25968 13574 25998 13626
rect 26022 13574 26032 13626
rect 26032 13574 26078 13626
rect 25782 13572 25838 13574
rect 25862 13572 25918 13574
rect 25942 13572 25998 13574
rect 26022 13572 26078 13574
rect 25782 12538 25838 12540
rect 25862 12538 25918 12540
rect 25942 12538 25998 12540
rect 26022 12538 26078 12540
rect 25782 12486 25828 12538
rect 25828 12486 25838 12538
rect 25862 12486 25892 12538
rect 25892 12486 25904 12538
rect 25904 12486 25918 12538
rect 25942 12486 25956 12538
rect 25956 12486 25968 12538
rect 25968 12486 25998 12538
rect 26022 12486 26032 12538
rect 26032 12486 26078 12538
rect 25782 12484 25838 12486
rect 25862 12484 25918 12486
rect 25942 12484 25998 12486
rect 26022 12484 26078 12486
rect 25782 11450 25838 11452
rect 25862 11450 25918 11452
rect 25942 11450 25998 11452
rect 26022 11450 26078 11452
rect 25782 11398 25828 11450
rect 25828 11398 25838 11450
rect 25862 11398 25892 11450
rect 25892 11398 25904 11450
rect 25904 11398 25918 11450
rect 25942 11398 25956 11450
rect 25956 11398 25968 11450
rect 25968 11398 25998 11450
rect 26022 11398 26032 11450
rect 26032 11398 26078 11450
rect 25782 11396 25838 11398
rect 25862 11396 25918 11398
rect 25942 11396 25998 11398
rect 26022 11396 26078 11398
rect 25226 8472 25282 8528
rect 25782 10362 25838 10364
rect 25862 10362 25918 10364
rect 25942 10362 25998 10364
rect 26022 10362 26078 10364
rect 25782 10310 25828 10362
rect 25828 10310 25838 10362
rect 25862 10310 25892 10362
rect 25892 10310 25904 10362
rect 25904 10310 25918 10362
rect 25942 10310 25956 10362
rect 25956 10310 25968 10362
rect 25968 10310 25998 10362
rect 26022 10310 26032 10362
rect 26032 10310 26078 10362
rect 25782 10308 25838 10310
rect 25862 10308 25918 10310
rect 25942 10308 25998 10310
rect 26022 10308 26078 10310
rect 25782 9274 25838 9276
rect 25862 9274 25918 9276
rect 25942 9274 25998 9276
rect 26022 9274 26078 9276
rect 25782 9222 25828 9274
rect 25828 9222 25838 9274
rect 25862 9222 25892 9274
rect 25892 9222 25904 9274
rect 25904 9222 25918 9274
rect 25942 9222 25956 9274
rect 25956 9222 25968 9274
rect 25968 9222 25998 9274
rect 26022 9222 26032 9274
rect 26032 9222 26078 9274
rect 25782 9220 25838 9222
rect 25862 9220 25918 9222
rect 25942 9220 25998 9222
rect 26022 9220 26078 9222
rect 25782 8186 25838 8188
rect 25862 8186 25918 8188
rect 25942 8186 25998 8188
rect 26022 8186 26078 8188
rect 25782 8134 25828 8186
rect 25828 8134 25838 8186
rect 25862 8134 25892 8186
rect 25892 8134 25904 8186
rect 25904 8134 25918 8186
rect 25942 8134 25956 8186
rect 25956 8134 25968 8186
rect 25968 8134 25998 8186
rect 26022 8134 26032 8186
rect 26032 8134 26078 8186
rect 25782 8132 25838 8134
rect 25862 8132 25918 8134
rect 25942 8132 25998 8134
rect 26022 8132 26078 8134
rect 25782 7098 25838 7100
rect 25862 7098 25918 7100
rect 25942 7098 25998 7100
rect 26022 7098 26078 7100
rect 25782 7046 25828 7098
rect 25828 7046 25838 7098
rect 25862 7046 25892 7098
rect 25892 7046 25904 7098
rect 25904 7046 25918 7098
rect 25942 7046 25956 7098
rect 25956 7046 25968 7098
rect 25968 7046 25998 7098
rect 26022 7046 26032 7098
rect 26032 7046 26078 7098
rect 25782 7044 25838 7046
rect 25862 7044 25918 7046
rect 25942 7044 25998 7046
rect 26022 7044 26078 7046
rect 26974 17584 27030 17640
rect 25782 6010 25838 6012
rect 25862 6010 25918 6012
rect 25942 6010 25998 6012
rect 26022 6010 26078 6012
rect 25782 5958 25828 6010
rect 25828 5958 25838 6010
rect 25862 5958 25892 6010
rect 25892 5958 25904 6010
rect 25904 5958 25918 6010
rect 25942 5958 25956 6010
rect 25956 5958 25968 6010
rect 25968 5958 25998 6010
rect 26022 5958 26032 6010
rect 26032 5958 26078 6010
rect 25782 5956 25838 5958
rect 25862 5956 25918 5958
rect 25942 5956 25998 5958
rect 26022 5956 26078 5958
rect 30010 25336 30066 25392
rect 27894 22072 27950 22128
rect 28078 22072 28134 22128
rect 27710 18128 27766 18184
rect 27618 17756 27620 17776
rect 27620 17756 27672 17776
rect 27672 17756 27674 17776
rect 27618 17720 27674 17756
rect 28354 23160 28410 23216
rect 28630 22072 28686 22128
rect 28538 20984 28594 21040
rect 28262 20168 28318 20224
rect 27802 11328 27858 11384
rect 25782 4922 25838 4924
rect 25862 4922 25918 4924
rect 25942 4922 25998 4924
rect 26022 4922 26078 4924
rect 25782 4870 25828 4922
rect 25828 4870 25838 4922
rect 25862 4870 25892 4922
rect 25892 4870 25904 4922
rect 25904 4870 25918 4922
rect 25942 4870 25956 4922
rect 25956 4870 25968 4922
rect 25968 4870 25998 4922
rect 26022 4870 26032 4922
rect 26032 4870 26078 4922
rect 25782 4868 25838 4870
rect 25862 4868 25918 4870
rect 25942 4868 25998 4870
rect 26022 4868 26078 4870
rect 30010 24676 30066 24712
rect 30010 24656 30012 24676
rect 30012 24656 30064 24676
rect 30064 24656 30066 24676
rect 30010 23840 30066 23896
rect 28906 22344 28962 22400
rect 28906 21664 28962 21720
rect 28814 19488 28870 19544
rect 28538 15000 28594 15056
rect 28630 14320 28686 14376
rect 28906 15816 28962 15872
rect 30102 17992 30158 18048
rect 28814 13504 28870 13560
rect 28906 12824 28962 12880
rect 28814 12008 28870 12064
rect 29182 10648 29238 10704
rect 25782 3834 25838 3836
rect 25862 3834 25918 3836
rect 25942 3834 25998 3836
rect 26022 3834 26078 3836
rect 25782 3782 25828 3834
rect 25828 3782 25838 3834
rect 25862 3782 25892 3834
rect 25892 3782 25904 3834
rect 25904 3782 25918 3834
rect 25942 3782 25956 3834
rect 25956 3782 25968 3834
rect 25968 3782 25998 3834
rect 26022 3782 26032 3834
rect 26032 3782 26078 3834
rect 25782 3780 25838 3782
rect 25862 3780 25918 3782
rect 25942 3780 25998 3782
rect 26022 3780 26078 3782
rect 20817 3290 20873 3292
rect 20897 3290 20953 3292
rect 20977 3290 21033 3292
rect 21057 3290 21113 3292
rect 20817 3238 20863 3290
rect 20863 3238 20873 3290
rect 20897 3238 20927 3290
rect 20927 3238 20939 3290
rect 20939 3238 20953 3290
rect 20977 3238 20991 3290
rect 20991 3238 21003 3290
rect 21003 3238 21033 3290
rect 21057 3238 21067 3290
rect 21067 3238 21113 3290
rect 20817 3236 20873 3238
rect 20897 3236 20953 3238
rect 20977 3236 21033 3238
rect 21057 3236 21113 3238
rect 25782 2746 25838 2748
rect 25862 2746 25918 2748
rect 25942 2746 25998 2748
rect 26022 2746 26078 2748
rect 25782 2694 25828 2746
rect 25828 2694 25838 2746
rect 25862 2694 25892 2746
rect 25892 2694 25904 2746
rect 25904 2694 25918 2746
rect 25942 2694 25956 2746
rect 25956 2694 25968 2746
rect 25968 2694 25998 2746
rect 26022 2694 26032 2746
rect 26032 2694 26078 2746
rect 25782 2692 25838 2694
rect 25862 2692 25918 2694
rect 25942 2692 25998 2694
rect 26022 2692 26078 2694
rect 30194 9832 30250 9888
rect 30102 9152 30158 9208
rect 30102 8336 30158 8392
rect 30102 7656 30158 7712
rect 30102 6840 30158 6896
rect 30102 6160 30158 6216
rect 29918 5480 29974 5536
rect 29918 4664 29974 4720
rect 29918 3984 29974 4040
rect 30010 3168 30066 3224
rect 29826 2488 29882 2544
rect 10886 2202 10942 2204
rect 10966 2202 11022 2204
rect 11046 2202 11102 2204
rect 11126 2202 11182 2204
rect 10886 2150 10932 2202
rect 10932 2150 10942 2202
rect 10966 2150 10996 2202
rect 10996 2150 11008 2202
rect 11008 2150 11022 2202
rect 11046 2150 11060 2202
rect 11060 2150 11072 2202
rect 11072 2150 11102 2202
rect 11126 2150 11136 2202
rect 11136 2150 11182 2202
rect 10886 2148 10942 2150
rect 10966 2148 11022 2150
rect 11046 2148 11102 2150
rect 11126 2148 11182 2150
rect 20817 2202 20873 2204
rect 20897 2202 20953 2204
rect 20977 2202 21033 2204
rect 21057 2202 21113 2204
rect 20817 2150 20863 2202
rect 20863 2150 20873 2202
rect 20897 2150 20927 2202
rect 20927 2150 20939 2202
rect 20939 2150 20953 2202
rect 20977 2150 20991 2202
rect 20991 2150 21003 2202
rect 21003 2150 21033 2202
rect 21057 2150 21067 2202
rect 21067 2150 21113 2202
rect 20817 2148 20873 2150
rect 20897 2148 20953 2150
rect 20977 2148 21033 2150
rect 21057 2148 21113 2150
rect 1582 992 1638 1048
rect 28722 992 28778 1048
rect 29918 1672 29974 1728
rect 29734 312 29790 368
<< metal3 >>
rect 30005 47562 30071 47565
rect 31200 47562 32000 47592
rect 30005 47560 32000 47562
rect 30005 47504 30010 47560
rect 30066 47504 32000 47560
rect 30005 47502 32000 47504
rect 30005 47499 30071 47502
rect 31200 47472 32000 47502
rect 0 47018 800 47048
rect 2773 47018 2839 47021
rect 0 47016 2839 47018
rect 0 46960 2778 47016
rect 2834 46960 2839 47016
rect 0 46958 2839 46960
rect 0 46928 800 46958
rect 2773 46955 2839 46958
rect 27889 46882 27955 46885
rect 31200 46882 32000 46912
rect 27889 46880 32000 46882
rect 27889 46824 27894 46880
rect 27950 46824 32000 46880
rect 27889 46822 32000 46824
rect 27889 46819 27955 46822
rect 31200 46792 32000 46822
rect 28901 46066 28967 46069
rect 31200 46066 32000 46096
rect 28901 46064 32000 46066
rect 28901 46008 28906 46064
rect 28962 46008 32000 46064
rect 28901 46006 32000 46008
rect 28901 46003 28967 46006
rect 31200 45976 32000 46006
rect 10874 45728 11194 45729
rect 10874 45664 10882 45728
rect 10946 45664 10962 45728
rect 11026 45664 11042 45728
rect 11106 45664 11122 45728
rect 11186 45664 11194 45728
rect 10874 45663 11194 45664
rect 20805 45728 21125 45729
rect 20805 45664 20813 45728
rect 20877 45664 20893 45728
rect 20957 45664 20973 45728
rect 21037 45664 21053 45728
rect 21117 45664 21125 45728
rect 20805 45663 21125 45664
rect 23841 45658 23907 45661
rect 26141 45658 26207 45661
rect 23841 45656 26207 45658
rect 23841 45600 23846 45656
rect 23902 45600 26146 45656
rect 26202 45600 26207 45656
rect 23841 45598 26207 45600
rect 23841 45595 23907 45598
rect 26141 45595 26207 45598
rect 21449 45522 21515 45525
rect 28441 45522 28507 45525
rect 21449 45520 28507 45522
rect 21449 45464 21454 45520
rect 21510 45464 28446 45520
rect 28502 45464 28507 45520
rect 21449 45462 28507 45464
rect 21449 45459 21515 45462
rect 28441 45459 28507 45462
rect 15193 45386 15259 45389
rect 17033 45386 17099 45389
rect 15193 45384 17099 45386
rect 15193 45328 15198 45384
rect 15254 45328 17038 45384
rect 17094 45328 17099 45384
rect 15193 45326 17099 45328
rect 15193 45323 15259 45326
rect 17033 45323 17099 45326
rect 20989 45386 21055 45389
rect 27521 45386 27587 45389
rect 20989 45384 27587 45386
rect 20989 45328 20994 45384
rect 21050 45328 27526 45384
rect 27582 45328 27587 45384
rect 20989 45326 27587 45328
rect 20989 45323 21055 45326
rect 27521 45323 27587 45326
rect 27705 45386 27771 45389
rect 31200 45386 32000 45416
rect 27705 45384 32000 45386
rect 27705 45328 27710 45384
rect 27766 45328 32000 45384
rect 27705 45326 32000 45328
rect 27705 45323 27771 45326
rect 31200 45296 32000 45326
rect 5909 45184 6229 45185
rect 5909 45120 5917 45184
rect 5981 45120 5997 45184
rect 6061 45120 6077 45184
rect 6141 45120 6157 45184
rect 6221 45120 6229 45184
rect 5909 45119 6229 45120
rect 15840 45184 16160 45185
rect 15840 45120 15848 45184
rect 15912 45120 15928 45184
rect 15992 45120 16008 45184
rect 16072 45120 16088 45184
rect 16152 45120 16160 45184
rect 15840 45119 16160 45120
rect 25770 45184 26090 45185
rect 25770 45120 25778 45184
rect 25842 45120 25858 45184
rect 25922 45120 25938 45184
rect 26002 45120 26018 45184
rect 26082 45120 26090 45184
rect 25770 45119 26090 45120
rect 0 44978 800 45008
rect 1577 44978 1643 44981
rect 0 44976 1643 44978
rect 0 44920 1582 44976
rect 1638 44920 1643 44976
rect 0 44918 1643 44920
rect 0 44888 800 44918
rect 1577 44915 1643 44918
rect 14273 44978 14339 44981
rect 17309 44978 17375 44981
rect 14273 44976 17375 44978
rect 14273 44920 14278 44976
rect 14334 44920 17314 44976
rect 17370 44920 17375 44976
rect 14273 44918 17375 44920
rect 14273 44915 14339 44918
rect 17309 44915 17375 44918
rect 21449 44978 21515 44981
rect 22001 44978 22067 44981
rect 21449 44976 22067 44978
rect 21449 44920 21454 44976
rect 21510 44920 22006 44976
rect 22062 44920 22067 44976
rect 21449 44918 22067 44920
rect 21449 44915 21515 44918
rect 22001 44915 22067 44918
rect 22185 44978 22251 44981
rect 27429 44978 27495 44981
rect 22185 44976 27495 44978
rect 22185 44920 22190 44976
rect 22246 44920 27434 44976
rect 27490 44920 27495 44976
rect 22185 44918 27495 44920
rect 22185 44915 22251 44918
rect 27429 44915 27495 44918
rect 14641 44842 14707 44845
rect 17217 44842 17283 44845
rect 14641 44840 17283 44842
rect 14641 44784 14646 44840
rect 14702 44784 17222 44840
rect 17278 44784 17283 44840
rect 14641 44782 17283 44784
rect 14641 44779 14707 44782
rect 17217 44779 17283 44782
rect 20989 44842 21055 44845
rect 21214 44842 21220 44844
rect 20989 44840 21220 44842
rect 20989 44784 20994 44840
rect 21050 44784 21220 44840
rect 20989 44782 21220 44784
rect 20989 44779 21055 44782
rect 21214 44780 21220 44782
rect 21284 44780 21290 44844
rect 10874 44640 11194 44641
rect 10874 44576 10882 44640
rect 10946 44576 10962 44640
rect 11026 44576 11042 44640
rect 11106 44576 11122 44640
rect 11186 44576 11194 44640
rect 10874 44575 11194 44576
rect 20805 44640 21125 44641
rect 20805 44576 20813 44640
rect 20877 44576 20893 44640
rect 20957 44576 20973 44640
rect 21037 44576 21053 44640
rect 21117 44576 21125 44640
rect 20805 44575 21125 44576
rect 30005 44570 30071 44573
rect 31200 44570 32000 44600
rect 30005 44568 32000 44570
rect 30005 44512 30010 44568
rect 30066 44512 32000 44568
rect 30005 44510 32000 44512
rect 30005 44507 30071 44510
rect 31200 44480 32000 44510
rect 21449 44434 21515 44437
rect 25681 44434 25747 44437
rect 21449 44432 25747 44434
rect 21449 44376 21454 44432
rect 21510 44376 25686 44432
rect 25742 44376 25747 44432
rect 21449 44374 25747 44376
rect 21449 44371 21515 44374
rect 25681 44371 25747 44374
rect 13537 44298 13603 44301
rect 17217 44298 17283 44301
rect 13537 44296 17283 44298
rect 13537 44240 13542 44296
rect 13598 44240 17222 44296
rect 17278 44240 17283 44296
rect 13537 44238 17283 44240
rect 13537 44235 13603 44238
rect 17217 44235 17283 44238
rect 20713 44298 20779 44301
rect 22185 44298 22251 44301
rect 20713 44296 22251 44298
rect 20713 44240 20718 44296
rect 20774 44240 22190 44296
rect 22246 44240 22251 44296
rect 20713 44238 22251 44240
rect 20713 44235 20779 44238
rect 21590 44165 21650 44238
rect 22185 44235 22251 44238
rect 23381 44298 23447 44301
rect 25221 44298 25287 44301
rect 26233 44298 26299 44301
rect 23381 44296 25287 44298
rect 23381 44240 23386 44296
rect 23442 44240 25226 44296
rect 25282 44240 25287 44296
rect 23381 44238 25287 44240
rect 23381 44235 23447 44238
rect 25221 44235 25287 44238
rect 25454 44296 26299 44298
rect 25454 44240 26238 44296
rect 26294 44240 26299 44296
rect 25454 44238 26299 44240
rect 14181 44162 14247 44165
rect 15285 44162 15351 44165
rect 14181 44160 15351 44162
rect 14181 44104 14186 44160
rect 14242 44104 15290 44160
rect 15346 44104 15351 44160
rect 14181 44102 15351 44104
rect 14181 44099 14247 44102
rect 15285 44099 15351 44102
rect 21541 44160 21650 44165
rect 21541 44104 21546 44160
rect 21602 44104 21650 44160
rect 21541 44102 21650 44104
rect 23381 44162 23447 44165
rect 25454 44162 25514 44238
rect 26233 44235 26299 44238
rect 23381 44160 25514 44162
rect 23381 44104 23386 44160
rect 23442 44104 25514 44160
rect 23381 44102 25514 44104
rect 21541 44099 21607 44102
rect 23381 44099 23447 44102
rect 5909 44096 6229 44097
rect 5909 44032 5917 44096
rect 5981 44032 5997 44096
rect 6061 44032 6077 44096
rect 6141 44032 6157 44096
rect 6221 44032 6229 44096
rect 5909 44031 6229 44032
rect 15840 44096 16160 44097
rect 15840 44032 15848 44096
rect 15912 44032 15928 44096
rect 15992 44032 16008 44096
rect 16072 44032 16088 44096
rect 16152 44032 16160 44096
rect 15840 44031 16160 44032
rect 25770 44096 26090 44097
rect 25770 44032 25778 44096
rect 25842 44032 25858 44096
rect 25922 44032 25938 44096
rect 26002 44032 26018 44096
rect 26082 44032 26090 44096
rect 25770 44031 26090 44032
rect 30097 44026 30163 44029
rect 26190 44024 30163 44026
rect 26190 43968 30102 44024
rect 30158 43968 30163 44024
rect 26190 43966 30163 43968
rect 13997 43890 14063 43893
rect 26190 43890 26250 43966
rect 30097 43963 30163 43966
rect 13997 43888 26250 43890
rect 13997 43832 14002 43888
rect 14058 43832 26250 43888
rect 13997 43830 26250 43832
rect 30005 43890 30071 43893
rect 31200 43890 32000 43920
rect 30005 43888 32000 43890
rect 30005 43832 30010 43888
rect 30066 43832 32000 43888
rect 30005 43830 32000 43832
rect 13997 43827 14063 43830
rect 30005 43827 30071 43830
rect 31200 43800 32000 43830
rect 23565 43754 23631 43757
rect 24669 43754 24735 43757
rect 23565 43752 24735 43754
rect 23565 43696 23570 43752
rect 23626 43696 24674 43752
rect 24730 43696 24735 43752
rect 23565 43694 24735 43696
rect 23565 43691 23631 43694
rect 24669 43691 24735 43694
rect 10874 43552 11194 43553
rect 10874 43488 10882 43552
rect 10946 43488 10962 43552
rect 11026 43488 11042 43552
rect 11106 43488 11122 43552
rect 11186 43488 11194 43552
rect 10874 43487 11194 43488
rect 20805 43552 21125 43553
rect 20805 43488 20813 43552
rect 20877 43488 20893 43552
rect 20957 43488 20973 43552
rect 21037 43488 21053 43552
rect 21117 43488 21125 43552
rect 20805 43487 21125 43488
rect 21909 43210 21975 43213
rect 22277 43210 22343 43213
rect 21909 43208 22343 43210
rect 21909 43152 21914 43208
rect 21970 43152 22282 43208
rect 22338 43152 22343 43208
rect 21909 43150 22343 43152
rect 21909 43147 21975 43150
rect 22277 43147 22343 43150
rect 23381 43210 23447 43213
rect 27705 43210 27771 43213
rect 23381 43208 27771 43210
rect 23381 43152 23386 43208
rect 23442 43152 27710 43208
rect 27766 43152 27771 43208
rect 23381 43150 27771 43152
rect 23381 43147 23447 43150
rect 27705 43147 27771 43150
rect 18505 43074 18571 43077
rect 23289 43074 23355 43077
rect 18505 43072 23355 43074
rect 18505 43016 18510 43072
rect 18566 43016 23294 43072
rect 23350 43016 23355 43072
rect 18505 43014 23355 43016
rect 18505 43011 18571 43014
rect 23289 43011 23355 43014
rect 30005 43074 30071 43077
rect 31200 43074 32000 43104
rect 30005 43072 32000 43074
rect 30005 43016 30010 43072
rect 30066 43016 32000 43072
rect 30005 43014 32000 43016
rect 30005 43011 30071 43014
rect 5909 43008 6229 43009
rect 0 42938 800 42968
rect 5909 42944 5917 43008
rect 5981 42944 5997 43008
rect 6061 42944 6077 43008
rect 6141 42944 6157 43008
rect 6221 42944 6229 43008
rect 5909 42943 6229 42944
rect 15840 43008 16160 43009
rect 15840 42944 15848 43008
rect 15912 42944 15928 43008
rect 15992 42944 16008 43008
rect 16072 42944 16088 43008
rect 16152 42944 16160 43008
rect 15840 42943 16160 42944
rect 25770 43008 26090 43009
rect 25770 42944 25778 43008
rect 25842 42944 25858 43008
rect 25922 42944 25938 43008
rect 26002 42944 26018 43008
rect 26082 42944 26090 43008
rect 31200 42984 32000 43014
rect 25770 42943 26090 42944
rect 1577 42938 1643 42941
rect 0 42936 1643 42938
rect 0 42880 1582 42936
rect 1638 42880 1643 42936
rect 0 42878 1643 42880
rect 0 42848 800 42878
rect 1577 42875 1643 42878
rect 22093 42802 22159 42805
rect 27429 42802 27495 42805
rect 22093 42800 27495 42802
rect 22093 42744 22098 42800
rect 22154 42744 27434 42800
rect 27490 42744 27495 42800
rect 22093 42742 27495 42744
rect 22093 42739 22159 42742
rect 27429 42739 27495 42742
rect 24669 42530 24735 42533
rect 29177 42530 29243 42533
rect 24669 42528 29243 42530
rect 24669 42472 24674 42528
rect 24730 42472 29182 42528
rect 29238 42472 29243 42528
rect 24669 42470 29243 42472
rect 24669 42467 24735 42470
rect 29177 42467 29243 42470
rect 10874 42464 11194 42465
rect 10874 42400 10882 42464
rect 10946 42400 10962 42464
rect 11026 42400 11042 42464
rect 11106 42400 11122 42464
rect 11186 42400 11194 42464
rect 10874 42399 11194 42400
rect 20805 42464 21125 42465
rect 20805 42400 20813 42464
rect 20877 42400 20893 42464
rect 20957 42400 20973 42464
rect 21037 42400 21053 42464
rect 21117 42400 21125 42464
rect 20805 42399 21125 42400
rect 19333 42394 19399 42397
rect 19885 42394 19951 42397
rect 19333 42392 19951 42394
rect 19333 42336 19338 42392
rect 19394 42336 19890 42392
rect 19946 42336 19951 42392
rect 19333 42334 19951 42336
rect 19333 42331 19399 42334
rect 19885 42331 19951 42334
rect 30005 42394 30071 42397
rect 31200 42394 32000 42424
rect 30005 42392 32000 42394
rect 30005 42336 30010 42392
rect 30066 42336 32000 42392
rect 30005 42334 32000 42336
rect 30005 42331 30071 42334
rect 31200 42304 32000 42334
rect 19425 42258 19491 42261
rect 20621 42258 20687 42261
rect 19425 42256 20687 42258
rect 19425 42200 19430 42256
rect 19486 42200 20626 42256
rect 20682 42200 20687 42256
rect 19425 42198 20687 42200
rect 19425 42195 19491 42198
rect 20621 42195 20687 42198
rect 21173 42258 21239 42261
rect 21541 42258 21607 42261
rect 21173 42256 21607 42258
rect 21173 42200 21178 42256
rect 21234 42200 21546 42256
rect 21602 42200 21607 42256
rect 21173 42198 21607 42200
rect 21173 42195 21239 42198
rect 21541 42195 21607 42198
rect 23841 42258 23907 42261
rect 27429 42258 27495 42261
rect 23841 42256 27495 42258
rect 23841 42200 23846 42256
rect 23902 42200 27434 42256
rect 27490 42200 27495 42256
rect 23841 42198 27495 42200
rect 23841 42195 23907 42198
rect 27429 42195 27495 42198
rect 20621 42122 20687 42125
rect 21449 42122 21515 42125
rect 20621 42120 21515 42122
rect 20621 42064 20626 42120
rect 20682 42064 21454 42120
rect 21510 42064 21515 42120
rect 20621 42062 21515 42064
rect 20621 42059 20687 42062
rect 21449 42059 21515 42062
rect 5909 41920 6229 41921
rect 5909 41856 5917 41920
rect 5981 41856 5997 41920
rect 6061 41856 6077 41920
rect 6141 41856 6157 41920
rect 6221 41856 6229 41920
rect 5909 41855 6229 41856
rect 15840 41920 16160 41921
rect 15840 41856 15848 41920
rect 15912 41856 15928 41920
rect 15992 41856 16008 41920
rect 16072 41856 16088 41920
rect 16152 41856 16160 41920
rect 15840 41855 16160 41856
rect 25770 41920 26090 41921
rect 25770 41856 25778 41920
rect 25842 41856 25858 41920
rect 25922 41856 25938 41920
rect 26002 41856 26018 41920
rect 26082 41856 26090 41920
rect 25770 41855 26090 41856
rect 23841 41714 23907 41717
rect 28349 41714 28415 41717
rect 23841 41712 28415 41714
rect 23841 41656 23846 41712
rect 23902 41656 28354 41712
rect 28410 41656 28415 41712
rect 23841 41654 28415 41656
rect 23841 41651 23907 41654
rect 28349 41651 28415 41654
rect 30005 41714 30071 41717
rect 31200 41714 32000 41744
rect 30005 41712 32000 41714
rect 30005 41656 30010 41712
rect 30066 41656 32000 41712
rect 30005 41654 32000 41656
rect 30005 41651 30071 41654
rect 31200 41624 32000 41654
rect 25497 41578 25563 41581
rect 27429 41578 27495 41581
rect 25497 41576 27495 41578
rect 25497 41520 25502 41576
rect 25558 41520 27434 41576
rect 27490 41520 27495 41576
rect 25497 41518 27495 41520
rect 25497 41515 25563 41518
rect 27429 41515 27495 41518
rect 10874 41376 11194 41377
rect 10874 41312 10882 41376
rect 10946 41312 10962 41376
rect 11026 41312 11042 41376
rect 11106 41312 11122 41376
rect 11186 41312 11194 41376
rect 10874 41311 11194 41312
rect 20805 41376 21125 41377
rect 20805 41312 20813 41376
rect 20877 41312 20893 41376
rect 20957 41312 20973 41376
rect 21037 41312 21053 41376
rect 21117 41312 21125 41376
rect 20805 41311 21125 41312
rect 23013 41306 23079 41309
rect 26417 41306 26483 41309
rect 23013 41304 26483 41306
rect 23013 41248 23018 41304
rect 23074 41248 26422 41304
rect 26478 41248 26483 41304
rect 23013 41246 26483 41248
rect 23013 41243 23079 41246
rect 26417 41243 26483 41246
rect 19793 41170 19859 41173
rect 28165 41170 28231 41173
rect 19793 41168 28231 41170
rect 19793 41112 19798 41168
rect 19854 41112 28170 41168
rect 28226 41112 28231 41168
rect 19793 41110 28231 41112
rect 19793 41107 19859 41110
rect 28165 41107 28231 41110
rect 0 41034 800 41064
rect 1577 41034 1643 41037
rect 0 41032 1643 41034
rect 0 40976 1582 41032
rect 1638 40976 1643 41032
rect 0 40974 1643 40976
rect 0 40944 800 40974
rect 1577 40971 1643 40974
rect 22829 41034 22895 41037
rect 25681 41034 25747 41037
rect 22829 41032 25747 41034
rect 22829 40976 22834 41032
rect 22890 40976 25686 41032
rect 25742 40976 25747 41032
rect 22829 40974 25747 40976
rect 22829 40971 22895 40974
rect 25681 40971 25747 40974
rect 30005 40898 30071 40901
rect 31200 40898 32000 40928
rect 30005 40896 32000 40898
rect 30005 40840 30010 40896
rect 30066 40840 32000 40896
rect 30005 40838 32000 40840
rect 30005 40835 30071 40838
rect 5909 40832 6229 40833
rect 5909 40768 5917 40832
rect 5981 40768 5997 40832
rect 6061 40768 6077 40832
rect 6141 40768 6157 40832
rect 6221 40768 6229 40832
rect 5909 40767 6229 40768
rect 15840 40832 16160 40833
rect 15840 40768 15848 40832
rect 15912 40768 15928 40832
rect 15992 40768 16008 40832
rect 16072 40768 16088 40832
rect 16152 40768 16160 40832
rect 15840 40767 16160 40768
rect 25770 40832 26090 40833
rect 25770 40768 25778 40832
rect 25842 40768 25858 40832
rect 25922 40768 25938 40832
rect 26002 40768 26018 40832
rect 26082 40768 26090 40832
rect 31200 40808 32000 40838
rect 25770 40767 26090 40768
rect 21214 40564 21220 40628
rect 21284 40626 21290 40628
rect 21817 40626 21883 40629
rect 21284 40624 21883 40626
rect 21284 40568 21822 40624
rect 21878 40568 21883 40624
rect 21284 40566 21883 40568
rect 21284 40564 21290 40566
rect 21817 40563 21883 40566
rect 24945 40626 25011 40629
rect 25497 40626 25563 40629
rect 24945 40624 25563 40626
rect 24945 40568 24950 40624
rect 25006 40568 25502 40624
rect 25558 40568 25563 40624
rect 24945 40566 25563 40568
rect 24945 40563 25011 40566
rect 25497 40563 25563 40566
rect 19609 40490 19675 40493
rect 29913 40490 29979 40493
rect 19609 40488 29979 40490
rect 19609 40432 19614 40488
rect 19670 40432 29918 40488
rect 29974 40432 29979 40488
rect 19609 40430 29979 40432
rect 19609 40427 19675 40430
rect 29913 40427 29979 40430
rect 23197 40354 23263 40357
rect 27337 40354 27403 40357
rect 23197 40352 27403 40354
rect 23197 40296 23202 40352
rect 23258 40296 27342 40352
rect 27398 40296 27403 40352
rect 23197 40294 27403 40296
rect 23197 40291 23263 40294
rect 27337 40291 27403 40294
rect 10874 40288 11194 40289
rect 10874 40224 10882 40288
rect 10946 40224 10962 40288
rect 11026 40224 11042 40288
rect 11106 40224 11122 40288
rect 11186 40224 11194 40288
rect 10874 40223 11194 40224
rect 20805 40288 21125 40289
rect 20805 40224 20813 40288
rect 20877 40224 20893 40288
rect 20957 40224 20973 40288
rect 21037 40224 21053 40288
rect 21117 40224 21125 40288
rect 20805 40223 21125 40224
rect 21449 40218 21515 40221
rect 28257 40218 28323 40221
rect 21449 40216 28323 40218
rect 21449 40160 21454 40216
rect 21510 40160 28262 40216
rect 28318 40160 28323 40216
rect 21449 40158 28323 40160
rect 21449 40155 21515 40158
rect 28257 40155 28323 40158
rect 30097 40218 30163 40221
rect 31200 40218 32000 40248
rect 30097 40216 32000 40218
rect 30097 40160 30102 40216
rect 30158 40160 32000 40216
rect 30097 40158 32000 40160
rect 30097 40155 30163 40158
rect 31200 40128 32000 40158
rect 26785 40082 26851 40085
rect 28349 40082 28415 40085
rect 26785 40080 28415 40082
rect 26785 40024 26790 40080
rect 26846 40024 28354 40080
rect 28410 40024 28415 40080
rect 26785 40022 28415 40024
rect 26785 40019 26851 40022
rect 28349 40019 28415 40022
rect 5909 39744 6229 39745
rect 5909 39680 5917 39744
rect 5981 39680 5997 39744
rect 6061 39680 6077 39744
rect 6141 39680 6157 39744
rect 6221 39680 6229 39744
rect 5909 39679 6229 39680
rect 15840 39744 16160 39745
rect 15840 39680 15848 39744
rect 15912 39680 15928 39744
rect 15992 39680 16008 39744
rect 16072 39680 16088 39744
rect 16152 39680 16160 39744
rect 15840 39679 16160 39680
rect 25770 39744 26090 39745
rect 25770 39680 25778 39744
rect 25842 39680 25858 39744
rect 25922 39680 25938 39744
rect 26002 39680 26018 39744
rect 26082 39680 26090 39744
rect 25770 39679 26090 39680
rect 19609 39674 19675 39677
rect 24485 39674 24551 39677
rect 19609 39672 24551 39674
rect 19609 39616 19614 39672
rect 19670 39616 24490 39672
rect 24546 39616 24551 39672
rect 19609 39614 24551 39616
rect 19609 39611 19675 39614
rect 24485 39611 24551 39614
rect 23473 39538 23539 39541
rect 27521 39538 27587 39541
rect 23473 39536 27587 39538
rect 23473 39480 23478 39536
rect 23534 39480 27526 39536
rect 27582 39480 27587 39536
rect 23473 39478 27587 39480
rect 23473 39475 23539 39478
rect 27521 39475 27587 39478
rect 30005 39402 30071 39405
rect 31200 39402 32000 39432
rect 30005 39400 32000 39402
rect 30005 39344 30010 39400
rect 30066 39344 32000 39400
rect 30005 39342 32000 39344
rect 30005 39339 30071 39342
rect 31200 39312 32000 39342
rect 10874 39200 11194 39201
rect 10874 39136 10882 39200
rect 10946 39136 10962 39200
rect 11026 39136 11042 39200
rect 11106 39136 11122 39200
rect 11186 39136 11194 39200
rect 10874 39135 11194 39136
rect 20805 39200 21125 39201
rect 20805 39136 20813 39200
rect 20877 39136 20893 39200
rect 20957 39136 20973 39200
rect 21037 39136 21053 39200
rect 21117 39136 21125 39200
rect 20805 39135 21125 39136
rect 23013 39130 23079 39133
rect 26693 39130 26759 39133
rect 23013 39128 26759 39130
rect 23013 39072 23018 39128
rect 23074 39072 26698 39128
rect 26754 39072 26759 39128
rect 23013 39070 26759 39072
rect 23013 39067 23079 39070
rect 26693 39067 26759 39070
rect 0 38994 800 39024
rect 1577 38994 1643 38997
rect 0 38992 1643 38994
rect 0 38936 1582 38992
rect 1638 38936 1643 38992
rect 0 38934 1643 38936
rect 0 38904 800 38934
rect 1577 38931 1643 38934
rect 20345 38994 20411 38997
rect 25037 38994 25103 38997
rect 20345 38992 25103 38994
rect 20345 38936 20350 38992
rect 20406 38936 25042 38992
rect 25098 38936 25103 38992
rect 20345 38934 25103 38936
rect 20345 38931 20411 38934
rect 25037 38931 25103 38934
rect 28901 38722 28967 38725
rect 31200 38722 32000 38752
rect 28901 38720 32000 38722
rect 28901 38664 28906 38720
rect 28962 38664 32000 38720
rect 28901 38662 32000 38664
rect 28901 38659 28967 38662
rect 5909 38656 6229 38657
rect 5909 38592 5917 38656
rect 5981 38592 5997 38656
rect 6061 38592 6077 38656
rect 6141 38592 6157 38656
rect 6221 38592 6229 38656
rect 5909 38591 6229 38592
rect 15840 38656 16160 38657
rect 15840 38592 15848 38656
rect 15912 38592 15928 38656
rect 15992 38592 16008 38656
rect 16072 38592 16088 38656
rect 16152 38592 16160 38656
rect 15840 38591 16160 38592
rect 25770 38656 26090 38657
rect 25770 38592 25778 38656
rect 25842 38592 25858 38656
rect 25922 38592 25938 38656
rect 26002 38592 26018 38656
rect 26082 38592 26090 38656
rect 31200 38632 32000 38662
rect 25770 38591 26090 38592
rect 10874 38112 11194 38113
rect 10874 38048 10882 38112
rect 10946 38048 10962 38112
rect 11026 38048 11042 38112
rect 11106 38048 11122 38112
rect 11186 38048 11194 38112
rect 10874 38047 11194 38048
rect 20805 38112 21125 38113
rect 20805 38048 20813 38112
rect 20877 38048 20893 38112
rect 20957 38048 20973 38112
rect 21037 38048 21053 38112
rect 21117 38048 21125 38112
rect 20805 38047 21125 38048
rect 30097 37906 30163 37909
rect 31200 37906 32000 37936
rect 30097 37904 32000 37906
rect 30097 37848 30102 37904
rect 30158 37848 32000 37904
rect 30097 37846 32000 37848
rect 30097 37843 30163 37846
rect 31200 37816 32000 37846
rect 5909 37568 6229 37569
rect 5909 37504 5917 37568
rect 5981 37504 5997 37568
rect 6061 37504 6077 37568
rect 6141 37504 6157 37568
rect 6221 37504 6229 37568
rect 5909 37503 6229 37504
rect 15840 37568 16160 37569
rect 15840 37504 15848 37568
rect 15912 37504 15928 37568
rect 15992 37504 16008 37568
rect 16072 37504 16088 37568
rect 16152 37504 16160 37568
rect 15840 37503 16160 37504
rect 25770 37568 26090 37569
rect 25770 37504 25778 37568
rect 25842 37504 25858 37568
rect 25922 37504 25938 37568
rect 26002 37504 26018 37568
rect 26082 37504 26090 37568
rect 25770 37503 26090 37504
rect 20621 37226 20687 37229
rect 21357 37226 21423 37229
rect 20621 37224 21423 37226
rect 20621 37168 20626 37224
rect 20682 37168 21362 37224
rect 21418 37168 21423 37224
rect 20621 37166 21423 37168
rect 20621 37163 20687 37166
rect 21357 37163 21423 37166
rect 24485 37226 24551 37229
rect 27337 37226 27403 37229
rect 24485 37224 27403 37226
rect 24485 37168 24490 37224
rect 24546 37168 27342 37224
rect 27398 37168 27403 37224
rect 24485 37166 27403 37168
rect 24485 37163 24551 37166
rect 27337 37163 27403 37166
rect 30005 37226 30071 37229
rect 31200 37226 32000 37256
rect 30005 37224 32000 37226
rect 30005 37168 30010 37224
rect 30066 37168 32000 37224
rect 30005 37166 32000 37168
rect 30005 37163 30071 37166
rect 31200 37136 32000 37166
rect 10874 37024 11194 37025
rect 0 36954 800 36984
rect 10874 36960 10882 37024
rect 10946 36960 10962 37024
rect 11026 36960 11042 37024
rect 11106 36960 11122 37024
rect 11186 36960 11194 37024
rect 10874 36959 11194 36960
rect 20805 37024 21125 37025
rect 20805 36960 20813 37024
rect 20877 36960 20893 37024
rect 20957 36960 20973 37024
rect 21037 36960 21053 37024
rect 21117 36960 21125 37024
rect 20805 36959 21125 36960
rect 1577 36954 1643 36957
rect 0 36952 1643 36954
rect 0 36896 1582 36952
rect 1638 36896 1643 36952
rect 0 36894 1643 36896
rect 0 36864 800 36894
rect 1577 36891 1643 36894
rect 28901 36546 28967 36549
rect 31200 36546 32000 36576
rect 28901 36544 32000 36546
rect 28901 36488 28906 36544
rect 28962 36488 32000 36544
rect 28901 36486 32000 36488
rect 28901 36483 28967 36486
rect 5909 36480 6229 36481
rect 5909 36416 5917 36480
rect 5981 36416 5997 36480
rect 6061 36416 6077 36480
rect 6141 36416 6157 36480
rect 6221 36416 6229 36480
rect 5909 36415 6229 36416
rect 15840 36480 16160 36481
rect 15840 36416 15848 36480
rect 15912 36416 15928 36480
rect 15992 36416 16008 36480
rect 16072 36416 16088 36480
rect 16152 36416 16160 36480
rect 15840 36415 16160 36416
rect 25770 36480 26090 36481
rect 25770 36416 25778 36480
rect 25842 36416 25858 36480
rect 25922 36416 25938 36480
rect 26002 36416 26018 36480
rect 26082 36416 26090 36480
rect 31200 36456 32000 36486
rect 25770 36415 26090 36416
rect 18597 36276 18663 36277
rect 18597 36274 18644 36276
rect 18552 36272 18644 36274
rect 18552 36216 18602 36272
rect 18552 36214 18644 36216
rect 18597 36212 18644 36214
rect 18708 36212 18714 36276
rect 18597 36211 18663 36212
rect 10874 35936 11194 35937
rect 10874 35872 10882 35936
rect 10946 35872 10962 35936
rect 11026 35872 11042 35936
rect 11106 35872 11122 35936
rect 11186 35872 11194 35936
rect 10874 35871 11194 35872
rect 20805 35936 21125 35937
rect 20805 35872 20813 35936
rect 20877 35872 20893 35936
rect 20957 35872 20973 35936
rect 21037 35872 21053 35936
rect 21117 35872 21125 35936
rect 20805 35871 21125 35872
rect 19977 35730 20043 35733
rect 20805 35730 20871 35733
rect 19977 35728 20871 35730
rect 19977 35672 19982 35728
rect 20038 35672 20810 35728
rect 20866 35672 20871 35728
rect 19977 35670 20871 35672
rect 19977 35667 20043 35670
rect 20805 35667 20871 35670
rect 30005 35730 30071 35733
rect 31200 35730 32000 35760
rect 30005 35728 32000 35730
rect 30005 35672 30010 35728
rect 30066 35672 32000 35728
rect 30005 35670 32000 35672
rect 30005 35667 30071 35670
rect 31200 35640 32000 35670
rect 5909 35392 6229 35393
rect 5909 35328 5917 35392
rect 5981 35328 5997 35392
rect 6061 35328 6077 35392
rect 6141 35328 6157 35392
rect 6221 35328 6229 35392
rect 5909 35327 6229 35328
rect 15840 35392 16160 35393
rect 15840 35328 15848 35392
rect 15912 35328 15928 35392
rect 15992 35328 16008 35392
rect 16072 35328 16088 35392
rect 16152 35328 16160 35392
rect 15840 35327 16160 35328
rect 25770 35392 26090 35393
rect 25770 35328 25778 35392
rect 25842 35328 25858 35392
rect 25922 35328 25938 35392
rect 26002 35328 26018 35392
rect 26082 35328 26090 35392
rect 25770 35327 26090 35328
rect 21817 35322 21883 35325
rect 18508 35320 21883 35322
rect 18508 35264 21822 35320
rect 21878 35264 21883 35320
rect 18508 35262 21883 35264
rect 18508 35189 18568 35262
rect 21817 35259 21883 35262
rect 18505 35184 18571 35189
rect 18965 35186 19031 35189
rect 18505 35128 18510 35184
rect 18566 35128 18571 35184
rect 18505 35123 18571 35128
rect 18830 35184 19031 35186
rect 18830 35128 18970 35184
rect 19026 35128 19031 35184
rect 18830 35126 19031 35128
rect 0 35050 800 35080
rect 1577 35050 1643 35053
rect 0 35048 1643 35050
rect 0 34992 1582 35048
rect 1638 34992 1643 35048
rect 0 34990 1643 34992
rect 0 34960 800 34990
rect 1577 34987 1643 34990
rect 18830 34914 18890 35126
rect 18965 35123 19031 35126
rect 20437 35186 20503 35189
rect 20897 35186 20963 35189
rect 20437 35184 20963 35186
rect 20437 35128 20442 35184
rect 20498 35128 20902 35184
rect 20958 35128 20963 35184
rect 20437 35126 20963 35128
rect 20437 35123 20503 35126
rect 20897 35123 20963 35126
rect 19057 35052 19123 35053
rect 19006 34988 19012 35052
rect 19076 35050 19123 35052
rect 19609 35050 19675 35053
rect 20713 35050 20779 35053
rect 19076 35048 19168 35050
rect 19118 34992 19168 35048
rect 19076 34990 19168 34992
rect 19609 35048 20779 35050
rect 19609 34992 19614 35048
rect 19670 34992 20718 35048
rect 20774 34992 20779 35048
rect 19609 34990 20779 34992
rect 19076 34988 19123 34990
rect 19057 34987 19123 34988
rect 19609 34987 19675 34990
rect 20713 34987 20779 34990
rect 28901 35050 28967 35053
rect 31200 35050 32000 35080
rect 28901 35048 32000 35050
rect 28901 34992 28906 35048
rect 28962 34992 32000 35048
rect 28901 34990 32000 34992
rect 28901 34987 28967 34990
rect 31200 34960 32000 34990
rect 18830 34854 19074 34914
rect 10874 34848 11194 34849
rect 10874 34784 10882 34848
rect 10946 34784 10962 34848
rect 11026 34784 11042 34848
rect 11106 34784 11122 34848
rect 11186 34784 11194 34848
rect 10874 34783 11194 34784
rect 17217 34642 17283 34645
rect 17350 34642 17356 34644
rect 17217 34640 17356 34642
rect 17217 34584 17222 34640
rect 17278 34584 17356 34640
rect 17217 34582 17356 34584
rect 17217 34579 17283 34582
rect 17350 34580 17356 34582
rect 17420 34580 17426 34644
rect 19014 34509 19074 34854
rect 20805 34848 21125 34849
rect 20805 34784 20813 34848
rect 20877 34784 20893 34848
rect 20957 34784 20973 34848
rect 21037 34784 21053 34848
rect 21117 34784 21125 34848
rect 20805 34783 21125 34784
rect 18965 34504 19074 34509
rect 18965 34448 18970 34504
rect 19026 34448 19074 34504
rect 18965 34446 19074 34448
rect 18965 34443 19031 34446
rect 5909 34304 6229 34305
rect 5909 34240 5917 34304
rect 5981 34240 5997 34304
rect 6061 34240 6077 34304
rect 6141 34240 6157 34304
rect 6221 34240 6229 34304
rect 5909 34239 6229 34240
rect 15840 34304 16160 34305
rect 15840 34240 15848 34304
rect 15912 34240 15928 34304
rect 15992 34240 16008 34304
rect 16072 34240 16088 34304
rect 16152 34240 16160 34304
rect 15840 34239 16160 34240
rect 25770 34304 26090 34305
rect 25770 34240 25778 34304
rect 25842 34240 25858 34304
rect 25922 34240 25938 34304
rect 26002 34240 26018 34304
rect 26082 34240 26090 34304
rect 25770 34239 26090 34240
rect 28441 34234 28507 34237
rect 31200 34234 32000 34264
rect 28441 34232 32000 34234
rect 28441 34176 28446 34232
rect 28502 34176 32000 34232
rect 28441 34174 32000 34176
rect 28441 34171 28507 34174
rect 31200 34144 32000 34174
rect 10225 33962 10291 33965
rect 10409 33962 10475 33965
rect 10225 33960 10475 33962
rect 10225 33904 10230 33960
rect 10286 33904 10414 33960
rect 10470 33904 10475 33960
rect 10225 33902 10475 33904
rect 10225 33899 10291 33902
rect 10409 33899 10475 33902
rect 16614 33900 16620 33964
rect 16684 33962 16690 33964
rect 17585 33962 17651 33965
rect 16684 33960 17651 33962
rect 16684 33904 17590 33960
rect 17646 33904 17651 33960
rect 16684 33902 17651 33904
rect 16684 33900 16690 33902
rect 17585 33899 17651 33902
rect 18321 33826 18387 33829
rect 19006 33826 19012 33828
rect 18321 33824 19012 33826
rect 18321 33768 18326 33824
rect 18382 33768 19012 33824
rect 18321 33766 19012 33768
rect 18321 33763 18387 33766
rect 19006 33764 19012 33766
rect 19076 33764 19082 33828
rect 10874 33760 11194 33761
rect 10874 33696 10882 33760
rect 10946 33696 10962 33760
rect 11026 33696 11042 33760
rect 11106 33696 11122 33760
rect 11186 33696 11194 33760
rect 10874 33695 11194 33696
rect 20805 33760 21125 33761
rect 20805 33696 20813 33760
rect 20877 33696 20893 33760
rect 20957 33696 20973 33760
rect 21037 33696 21053 33760
rect 21117 33696 21125 33760
rect 20805 33695 21125 33696
rect 20805 33554 20871 33557
rect 27245 33554 27311 33557
rect 20805 33552 27311 33554
rect 20805 33496 20810 33552
rect 20866 33496 27250 33552
rect 27306 33496 27311 33552
rect 20805 33494 27311 33496
rect 20805 33491 20871 33494
rect 27245 33491 27311 33494
rect 28901 33554 28967 33557
rect 31200 33554 32000 33584
rect 28901 33552 32000 33554
rect 28901 33496 28906 33552
rect 28962 33496 32000 33552
rect 28901 33494 32000 33496
rect 28901 33491 28967 33494
rect 31200 33464 32000 33494
rect 5909 33216 6229 33217
rect 5909 33152 5917 33216
rect 5981 33152 5997 33216
rect 6061 33152 6077 33216
rect 6141 33152 6157 33216
rect 6221 33152 6229 33216
rect 5909 33151 6229 33152
rect 15840 33216 16160 33217
rect 15840 33152 15848 33216
rect 15912 33152 15928 33216
rect 15992 33152 16008 33216
rect 16072 33152 16088 33216
rect 16152 33152 16160 33216
rect 15840 33151 16160 33152
rect 25770 33216 26090 33217
rect 25770 33152 25778 33216
rect 25842 33152 25858 33216
rect 25922 33152 25938 33216
rect 26002 33152 26018 33216
rect 26082 33152 26090 33216
rect 25770 33151 26090 33152
rect 0 33010 800 33040
rect 1577 33010 1643 33013
rect 0 33008 1643 33010
rect 0 32952 1582 33008
rect 1638 32952 1643 33008
rect 0 32950 1643 32952
rect 0 32920 800 32950
rect 1577 32947 1643 32950
rect 30005 32738 30071 32741
rect 31200 32738 32000 32768
rect 30005 32736 32000 32738
rect 30005 32680 30010 32736
rect 30066 32680 32000 32736
rect 30005 32678 32000 32680
rect 30005 32675 30071 32678
rect 10874 32672 11194 32673
rect 10874 32608 10882 32672
rect 10946 32608 10962 32672
rect 11026 32608 11042 32672
rect 11106 32608 11122 32672
rect 11186 32608 11194 32672
rect 10874 32607 11194 32608
rect 20805 32672 21125 32673
rect 20805 32608 20813 32672
rect 20877 32608 20893 32672
rect 20957 32608 20973 32672
rect 21037 32608 21053 32672
rect 21117 32608 21125 32672
rect 31200 32648 32000 32678
rect 20805 32607 21125 32608
rect 5909 32128 6229 32129
rect 5909 32064 5917 32128
rect 5981 32064 5997 32128
rect 6061 32064 6077 32128
rect 6141 32064 6157 32128
rect 6221 32064 6229 32128
rect 5909 32063 6229 32064
rect 15840 32128 16160 32129
rect 15840 32064 15848 32128
rect 15912 32064 15928 32128
rect 15992 32064 16008 32128
rect 16072 32064 16088 32128
rect 16152 32064 16160 32128
rect 15840 32063 16160 32064
rect 25770 32128 26090 32129
rect 25770 32064 25778 32128
rect 25842 32064 25858 32128
rect 25922 32064 25938 32128
rect 26002 32064 26018 32128
rect 26082 32064 26090 32128
rect 25770 32063 26090 32064
rect 30097 32058 30163 32061
rect 31200 32058 32000 32088
rect 30097 32056 32000 32058
rect 30097 32000 30102 32056
rect 30158 32000 32000 32056
rect 30097 31998 32000 32000
rect 30097 31995 30163 31998
rect 31200 31968 32000 31998
rect 17534 31860 17540 31924
rect 17604 31922 17610 31924
rect 17677 31922 17743 31925
rect 18781 31922 18847 31925
rect 17604 31920 17743 31922
rect 17604 31864 17682 31920
rect 17738 31864 17743 31920
rect 17604 31862 17743 31864
rect 17604 31860 17610 31862
rect 17677 31859 17743 31862
rect 18278 31920 18847 31922
rect 18278 31864 18786 31920
rect 18842 31864 18847 31920
rect 18278 31862 18847 31864
rect 15653 31786 15719 31789
rect 18278 31786 18338 31862
rect 18781 31859 18847 31862
rect 15653 31784 18338 31786
rect 15653 31728 15658 31784
rect 15714 31728 18338 31784
rect 15653 31726 18338 31728
rect 15653 31723 15719 31726
rect 10874 31584 11194 31585
rect 10874 31520 10882 31584
rect 10946 31520 10962 31584
rect 11026 31520 11042 31584
rect 11106 31520 11122 31584
rect 11186 31520 11194 31584
rect 10874 31519 11194 31520
rect 20805 31584 21125 31585
rect 20805 31520 20813 31584
rect 20877 31520 20893 31584
rect 20957 31520 20973 31584
rect 21037 31520 21053 31584
rect 21117 31520 21125 31584
rect 20805 31519 21125 31520
rect 15377 31514 15443 31517
rect 18229 31514 18295 31517
rect 15377 31512 18295 31514
rect 15377 31456 15382 31512
rect 15438 31456 18234 31512
rect 18290 31456 18295 31512
rect 15377 31454 18295 31456
rect 15377 31451 15443 31454
rect 18229 31451 18295 31454
rect 30005 31378 30071 31381
rect 31200 31378 32000 31408
rect 30005 31376 32000 31378
rect 30005 31320 30010 31376
rect 30066 31320 32000 31376
rect 30005 31318 32000 31320
rect 30005 31315 30071 31318
rect 31200 31288 32000 31318
rect 5909 31040 6229 31041
rect 0 30970 800 31000
rect 5909 30976 5917 31040
rect 5981 30976 5997 31040
rect 6061 30976 6077 31040
rect 6141 30976 6157 31040
rect 6221 30976 6229 31040
rect 5909 30975 6229 30976
rect 15840 31040 16160 31041
rect 15840 30976 15848 31040
rect 15912 30976 15928 31040
rect 15992 30976 16008 31040
rect 16072 30976 16088 31040
rect 16152 30976 16160 31040
rect 15840 30975 16160 30976
rect 25770 31040 26090 31041
rect 25770 30976 25778 31040
rect 25842 30976 25858 31040
rect 25922 30976 25938 31040
rect 26002 30976 26018 31040
rect 26082 30976 26090 31040
rect 25770 30975 26090 30976
rect 1393 30970 1459 30973
rect 0 30968 1459 30970
rect 0 30912 1398 30968
rect 1454 30912 1459 30968
rect 0 30910 1459 30912
rect 0 30880 800 30910
rect 1393 30907 1459 30910
rect 16573 30970 16639 30973
rect 16982 30970 16988 30972
rect 16573 30968 16988 30970
rect 16573 30912 16578 30968
rect 16634 30912 16988 30968
rect 16573 30910 16988 30912
rect 16573 30907 16639 30910
rect 16982 30908 16988 30910
rect 17052 30908 17058 30972
rect 16573 30836 16639 30837
rect 16573 30834 16620 30836
rect 16528 30832 16620 30834
rect 16528 30776 16578 30832
rect 16528 30774 16620 30776
rect 16573 30772 16620 30774
rect 16684 30772 16690 30836
rect 16573 30771 16639 30772
rect 19190 30636 19196 30700
rect 19260 30698 19266 30700
rect 19333 30698 19399 30701
rect 19260 30696 19399 30698
rect 19260 30640 19338 30696
rect 19394 30640 19399 30696
rect 19260 30638 19399 30640
rect 19260 30636 19266 30638
rect 19333 30635 19399 30638
rect 18638 30500 18644 30564
rect 18708 30562 18714 30564
rect 18873 30562 18939 30565
rect 18708 30560 18939 30562
rect 18708 30504 18878 30560
rect 18934 30504 18939 30560
rect 18708 30502 18939 30504
rect 18708 30500 18714 30502
rect 18873 30499 18939 30502
rect 30097 30562 30163 30565
rect 31200 30562 32000 30592
rect 30097 30560 32000 30562
rect 30097 30504 30102 30560
rect 30158 30504 32000 30560
rect 30097 30502 32000 30504
rect 30097 30499 30163 30502
rect 10874 30496 11194 30497
rect 10874 30432 10882 30496
rect 10946 30432 10962 30496
rect 11026 30432 11042 30496
rect 11106 30432 11122 30496
rect 11186 30432 11194 30496
rect 10874 30431 11194 30432
rect 20805 30496 21125 30497
rect 20805 30432 20813 30496
rect 20877 30432 20893 30496
rect 20957 30432 20973 30496
rect 21037 30432 21053 30496
rect 21117 30432 21125 30496
rect 31200 30472 32000 30502
rect 20805 30431 21125 30432
rect 16849 30426 16915 30429
rect 18137 30426 18203 30429
rect 16849 30424 18203 30426
rect 16849 30368 16854 30424
rect 16910 30368 18142 30424
rect 18198 30368 18203 30424
rect 16849 30366 18203 30368
rect 16849 30363 16915 30366
rect 18137 30363 18203 30366
rect 9949 30154 10015 30157
rect 17585 30156 17651 30157
rect 9949 30152 10242 30154
rect 9949 30096 9954 30152
rect 10010 30096 10242 30152
rect 9949 30094 10242 30096
rect 9949 30091 10015 30094
rect 5909 29952 6229 29953
rect 5909 29888 5917 29952
rect 5981 29888 5997 29952
rect 6061 29888 6077 29952
rect 6141 29888 6157 29952
rect 6221 29888 6229 29952
rect 5909 29887 6229 29888
rect 10182 29613 10242 30094
rect 17534 30092 17540 30156
rect 17604 30154 17651 30156
rect 18505 30154 18571 30157
rect 18689 30154 18755 30157
rect 17604 30152 17696 30154
rect 17646 30096 17696 30152
rect 17604 30094 17696 30096
rect 18505 30152 18755 30154
rect 18505 30096 18510 30152
rect 18566 30096 18694 30152
rect 18750 30096 18755 30152
rect 18505 30094 18755 30096
rect 17604 30092 17651 30094
rect 17585 30091 17651 30092
rect 18505 30091 18571 30094
rect 18689 30091 18755 30094
rect 15840 29952 16160 29953
rect 15840 29888 15848 29952
rect 15912 29888 15928 29952
rect 15992 29888 16008 29952
rect 16072 29888 16088 29952
rect 16152 29888 16160 29952
rect 15840 29887 16160 29888
rect 25770 29952 26090 29953
rect 25770 29888 25778 29952
rect 25842 29888 25858 29952
rect 25922 29888 25938 29952
rect 26002 29888 26018 29952
rect 26082 29888 26090 29952
rect 25770 29887 26090 29888
rect 30005 29882 30071 29885
rect 31200 29882 32000 29912
rect 30005 29880 32000 29882
rect 30005 29824 30010 29880
rect 30066 29824 32000 29880
rect 30005 29822 32000 29824
rect 30005 29819 30071 29822
rect 31200 29792 32000 29822
rect 17493 29746 17559 29749
rect 18137 29746 18203 29749
rect 17493 29744 18203 29746
rect 17493 29688 17498 29744
rect 17554 29688 18142 29744
rect 18198 29688 18203 29744
rect 17493 29686 18203 29688
rect 17493 29683 17559 29686
rect 18137 29683 18203 29686
rect 10182 29608 10291 29613
rect 10182 29552 10230 29608
rect 10286 29552 10291 29608
rect 10182 29550 10291 29552
rect 10225 29547 10291 29550
rect 13261 29474 13327 29477
rect 17217 29474 17283 29477
rect 13261 29472 17283 29474
rect 13261 29416 13266 29472
rect 13322 29416 17222 29472
rect 17278 29416 17283 29472
rect 13261 29414 17283 29416
rect 13261 29411 13327 29414
rect 17217 29411 17283 29414
rect 10874 29408 11194 29409
rect 10874 29344 10882 29408
rect 10946 29344 10962 29408
rect 11026 29344 11042 29408
rect 11106 29344 11122 29408
rect 11186 29344 11194 29408
rect 10874 29343 11194 29344
rect 20805 29408 21125 29409
rect 20805 29344 20813 29408
rect 20877 29344 20893 29408
rect 20957 29344 20973 29408
rect 21037 29344 21053 29408
rect 21117 29344 21125 29408
rect 20805 29343 21125 29344
rect 12801 29338 12867 29341
rect 19149 29338 19215 29341
rect 12801 29336 19215 29338
rect 12801 29280 12806 29336
rect 12862 29280 19154 29336
rect 19210 29280 19215 29336
rect 12801 29278 19215 29280
rect 12801 29275 12867 29278
rect 19149 29275 19215 29278
rect 11145 29202 11211 29205
rect 12893 29202 12959 29205
rect 16021 29202 16087 29205
rect 11145 29200 16087 29202
rect 11145 29144 11150 29200
rect 11206 29144 12898 29200
rect 12954 29144 16026 29200
rect 16082 29144 16087 29200
rect 11145 29142 16087 29144
rect 11145 29139 11211 29142
rect 12893 29139 12959 29142
rect 16021 29139 16087 29142
rect 30005 29066 30071 29069
rect 31200 29066 32000 29096
rect 30005 29064 32000 29066
rect 30005 29008 30010 29064
rect 30066 29008 32000 29064
rect 30005 29006 32000 29008
rect 30005 29003 30071 29006
rect 31200 28976 32000 29006
rect 0 28930 800 28960
rect 1577 28930 1643 28933
rect 0 28928 1643 28930
rect 0 28872 1582 28928
rect 1638 28872 1643 28928
rect 0 28870 1643 28872
rect 0 28840 800 28870
rect 1577 28867 1643 28870
rect 5909 28864 6229 28865
rect 5909 28800 5917 28864
rect 5981 28800 5997 28864
rect 6061 28800 6077 28864
rect 6141 28800 6157 28864
rect 6221 28800 6229 28864
rect 5909 28799 6229 28800
rect 15840 28864 16160 28865
rect 15840 28800 15848 28864
rect 15912 28800 15928 28864
rect 15992 28800 16008 28864
rect 16072 28800 16088 28864
rect 16152 28800 16160 28864
rect 15840 28799 16160 28800
rect 25770 28864 26090 28865
rect 25770 28800 25778 28864
rect 25842 28800 25858 28864
rect 25922 28800 25938 28864
rect 26002 28800 26018 28864
rect 26082 28800 26090 28864
rect 25770 28799 26090 28800
rect 19006 28596 19012 28660
rect 19076 28658 19082 28660
rect 19149 28658 19215 28661
rect 19076 28656 19215 28658
rect 19076 28600 19154 28656
rect 19210 28600 19215 28656
rect 19076 28598 19215 28600
rect 19076 28596 19082 28598
rect 19149 28595 19215 28598
rect 19333 28658 19399 28661
rect 21633 28658 21699 28661
rect 24853 28658 24919 28661
rect 19333 28656 21466 28658
rect 19333 28600 19338 28656
rect 19394 28600 21466 28656
rect 19333 28598 21466 28600
rect 19333 28595 19399 28598
rect 21406 28522 21466 28598
rect 21633 28656 24919 28658
rect 21633 28600 21638 28656
rect 21694 28600 24858 28656
rect 24914 28600 24919 28656
rect 21633 28598 24919 28600
rect 21633 28595 21699 28598
rect 24853 28595 24919 28598
rect 22369 28522 22435 28525
rect 21406 28520 22435 28522
rect 21406 28464 22374 28520
rect 22430 28464 22435 28520
rect 21406 28462 22435 28464
rect 22369 28459 22435 28462
rect 18965 28386 19031 28389
rect 19333 28386 19399 28389
rect 20161 28386 20227 28389
rect 18965 28384 19258 28386
rect 18965 28328 18970 28384
rect 19026 28328 19258 28384
rect 18965 28326 19258 28328
rect 18965 28323 19031 28326
rect 10874 28320 11194 28321
rect 10874 28256 10882 28320
rect 10946 28256 10962 28320
rect 11026 28256 11042 28320
rect 11106 28256 11122 28320
rect 11186 28256 11194 28320
rect 10874 28255 11194 28256
rect 17309 28250 17375 28253
rect 19057 28250 19123 28253
rect 17309 28248 19123 28250
rect 17309 28192 17314 28248
rect 17370 28192 19062 28248
rect 19118 28192 19123 28248
rect 17309 28190 19123 28192
rect 17309 28187 17375 28190
rect 19057 28187 19123 28190
rect 18505 28114 18571 28117
rect 18638 28114 18644 28116
rect 18505 28112 18644 28114
rect 18505 28056 18510 28112
rect 18566 28056 18644 28112
rect 18505 28054 18644 28056
rect 18505 28051 18571 28054
rect 18638 28052 18644 28054
rect 18708 28052 18714 28116
rect 19057 28114 19123 28117
rect 19014 28112 19123 28114
rect 19014 28056 19062 28112
rect 19118 28056 19123 28112
rect 19014 28051 19123 28056
rect 17861 27978 17927 27981
rect 19014 27978 19074 28051
rect 17861 27976 19074 27978
rect 17861 27920 17866 27976
rect 17922 27920 19074 27976
rect 17861 27918 19074 27920
rect 17861 27915 17927 27918
rect 18965 27842 19031 27845
rect 19198 27842 19258 28326
rect 19333 28384 20227 28386
rect 19333 28328 19338 28384
rect 19394 28328 20166 28384
rect 20222 28328 20227 28384
rect 19333 28326 20227 28328
rect 19333 28323 19399 28326
rect 20161 28323 20227 28326
rect 30005 28386 30071 28389
rect 31200 28386 32000 28416
rect 30005 28384 32000 28386
rect 30005 28328 30010 28384
rect 30066 28328 32000 28384
rect 30005 28326 32000 28328
rect 30005 28323 30071 28326
rect 20805 28320 21125 28321
rect 20805 28256 20813 28320
rect 20877 28256 20893 28320
rect 20957 28256 20973 28320
rect 21037 28256 21053 28320
rect 21117 28256 21125 28320
rect 31200 28296 32000 28326
rect 20805 28255 21125 28256
rect 19333 28114 19399 28117
rect 19977 28114 20043 28117
rect 19333 28112 20043 28114
rect 19333 28056 19338 28112
rect 19394 28056 19982 28112
rect 20038 28056 20043 28112
rect 19333 28054 20043 28056
rect 19333 28051 19399 28054
rect 19977 28051 20043 28054
rect 18965 27840 19258 27842
rect 18965 27784 18970 27840
rect 19026 27784 19258 27840
rect 18965 27782 19258 27784
rect 18965 27779 19031 27782
rect 5909 27776 6229 27777
rect 5909 27712 5917 27776
rect 5981 27712 5997 27776
rect 6061 27712 6077 27776
rect 6141 27712 6157 27776
rect 6221 27712 6229 27776
rect 5909 27711 6229 27712
rect 15840 27776 16160 27777
rect 15840 27712 15848 27776
rect 15912 27712 15928 27776
rect 15992 27712 16008 27776
rect 16072 27712 16088 27776
rect 16152 27712 16160 27776
rect 15840 27711 16160 27712
rect 25770 27776 26090 27777
rect 25770 27712 25778 27776
rect 25842 27712 25858 27776
rect 25922 27712 25938 27776
rect 26002 27712 26018 27776
rect 26082 27712 26090 27776
rect 25770 27711 26090 27712
rect 18638 27644 18644 27708
rect 18708 27706 18714 27708
rect 19241 27706 19307 27709
rect 18708 27704 19307 27706
rect 18708 27648 19246 27704
rect 19302 27648 19307 27704
rect 18708 27646 19307 27648
rect 18708 27644 18714 27646
rect 19241 27643 19307 27646
rect 30005 27570 30071 27573
rect 31200 27570 32000 27600
rect 30005 27568 32000 27570
rect 30005 27512 30010 27568
rect 30066 27512 32000 27568
rect 30005 27510 32000 27512
rect 30005 27507 30071 27510
rect 31200 27480 32000 27510
rect 10874 27232 11194 27233
rect 10874 27168 10882 27232
rect 10946 27168 10962 27232
rect 11026 27168 11042 27232
rect 11106 27168 11122 27232
rect 11186 27168 11194 27232
rect 10874 27167 11194 27168
rect 20805 27232 21125 27233
rect 20805 27168 20813 27232
rect 20877 27168 20893 27232
rect 20957 27168 20973 27232
rect 21037 27168 21053 27232
rect 21117 27168 21125 27232
rect 20805 27167 21125 27168
rect 19006 27100 19012 27164
rect 19076 27162 19082 27164
rect 19149 27162 19215 27165
rect 19076 27160 19215 27162
rect 19076 27104 19154 27160
rect 19210 27104 19215 27160
rect 19076 27102 19215 27104
rect 19076 27100 19082 27102
rect 19149 27099 19215 27102
rect 0 27026 800 27056
rect 1577 27026 1643 27029
rect 0 27024 1643 27026
rect 0 26968 1582 27024
rect 1638 26968 1643 27024
rect 0 26966 1643 26968
rect 0 26936 800 26966
rect 1577 26963 1643 26966
rect 30005 26890 30071 26893
rect 31200 26890 32000 26920
rect 30005 26888 32000 26890
rect 30005 26832 30010 26888
rect 30066 26832 32000 26888
rect 30005 26830 32000 26832
rect 30005 26827 30071 26830
rect 31200 26800 32000 26830
rect 5909 26688 6229 26689
rect 5909 26624 5917 26688
rect 5981 26624 5997 26688
rect 6061 26624 6077 26688
rect 6141 26624 6157 26688
rect 6221 26624 6229 26688
rect 5909 26623 6229 26624
rect 15840 26688 16160 26689
rect 15840 26624 15848 26688
rect 15912 26624 15928 26688
rect 15992 26624 16008 26688
rect 16072 26624 16088 26688
rect 16152 26624 16160 26688
rect 15840 26623 16160 26624
rect 25770 26688 26090 26689
rect 25770 26624 25778 26688
rect 25842 26624 25858 26688
rect 25922 26624 25938 26688
rect 26002 26624 26018 26688
rect 26082 26624 26090 26688
rect 25770 26623 26090 26624
rect 30005 26210 30071 26213
rect 31200 26210 32000 26240
rect 30005 26208 32000 26210
rect 30005 26152 30010 26208
rect 30066 26152 32000 26208
rect 30005 26150 32000 26152
rect 30005 26147 30071 26150
rect 10874 26144 11194 26145
rect 10874 26080 10882 26144
rect 10946 26080 10962 26144
rect 11026 26080 11042 26144
rect 11106 26080 11122 26144
rect 11186 26080 11194 26144
rect 10874 26079 11194 26080
rect 20805 26144 21125 26145
rect 20805 26080 20813 26144
rect 20877 26080 20893 26144
rect 20957 26080 20973 26144
rect 21037 26080 21053 26144
rect 21117 26080 21125 26144
rect 31200 26120 32000 26150
rect 20805 26079 21125 26080
rect 16205 25938 16271 25941
rect 18045 25938 18111 25941
rect 16205 25936 18111 25938
rect 16205 25880 16210 25936
rect 16266 25880 18050 25936
rect 18106 25880 18111 25936
rect 16205 25878 18111 25880
rect 16205 25875 16271 25878
rect 18045 25875 18111 25878
rect 13353 25802 13419 25805
rect 13997 25802 14063 25805
rect 13353 25800 14063 25802
rect 13353 25744 13358 25800
rect 13414 25744 14002 25800
rect 14058 25744 14063 25800
rect 13353 25742 14063 25744
rect 13353 25739 13419 25742
rect 13997 25739 14063 25742
rect 5909 25600 6229 25601
rect 5909 25536 5917 25600
rect 5981 25536 5997 25600
rect 6061 25536 6077 25600
rect 6141 25536 6157 25600
rect 6221 25536 6229 25600
rect 5909 25535 6229 25536
rect 15840 25600 16160 25601
rect 15840 25536 15848 25600
rect 15912 25536 15928 25600
rect 15992 25536 16008 25600
rect 16072 25536 16088 25600
rect 16152 25536 16160 25600
rect 15840 25535 16160 25536
rect 25770 25600 26090 25601
rect 25770 25536 25778 25600
rect 25842 25536 25858 25600
rect 25922 25536 25938 25600
rect 26002 25536 26018 25600
rect 26082 25536 26090 25600
rect 25770 25535 26090 25536
rect 30005 25394 30071 25397
rect 31200 25394 32000 25424
rect 30005 25392 32000 25394
rect 30005 25336 30010 25392
rect 30066 25336 32000 25392
rect 30005 25334 32000 25336
rect 30005 25331 30071 25334
rect 31200 25304 32000 25334
rect 13353 25122 13419 25125
rect 16297 25122 16363 25125
rect 13353 25120 16363 25122
rect 13353 25064 13358 25120
rect 13414 25064 16302 25120
rect 16358 25064 16363 25120
rect 13353 25062 16363 25064
rect 13353 25059 13419 25062
rect 16297 25059 16363 25062
rect 10874 25056 11194 25057
rect 0 24986 800 25016
rect 10874 24992 10882 25056
rect 10946 24992 10962 25056
rect 11026 24992 11042 25056
rect 11106 24992 11122 25056
rect 11186 24992 11194 25056
rect 10874 24991 11194 24992
rect 20805 25056 21125 25057
rect 20805 24992 20813 25056
rect 20877 24992 20893 25056
rect 20957 24992 20973 25056
rect 21037 24992 21053 25056
rect 21117 24992 21125 25056
rect 20805 24991 21125 24992
rect 1577 24986 1643 24989
rect 0 24984 1643 24986
rect 0 24928 1582 24984
rect 1638 24928 1643 24984
rect 0 24926 1643 24928
rect 0 24896 800 24926
rect 1577 24923 1643 24926
rect 10133 24714 10199 24717
rect 10593 24714 10659 24717
rect 10133 24712 10659 24714
rect 10133 24656 10138 24712
rect 10194 24656 10598 24712
rect 10654 24656 10659 24712
rect 10133 24654 10659 24656
rect 10133 24651 10199 24654
rect 10593 24651 10659 24654
rect 30005 24714 30071 24717
rect 31200 24714 32000 24744
rect 30005 24712 32000 24714
rect 30005 24656 30010 24712
rect 30066 24656 32000 24712
rect 30005 24654 32000 24656
rect 30005 24651 30071 24654
rect 31200 24624 32000 24654
rect 5909 24512 6229 24513
rect 5909 24448 5917 24512
rect 5981 24448 5997 24512
rect 6061 24448 6077 24512
rect 6141 24448 6157 24512
rect 6221 24448 6229 24512
rect 5909 24447 6229 24448
rect 15840 24512 16160 24513
rect 15840 24448 15848 24512
rect 15912 24448 15928 24512
rect 15992 24448 16008 24512
rect 16072 24448 16088 24512
rect 16152 24448 16160 24512
rect 15840 24447 16160 24448
rect 25770 24512 26090 24513
rect 25770 24448 25778 24512
rect 25842 24448 25858 24512
rect 25922 24448 25938 24512
rect 26002 24448 26018 24512
rect 26082 24448 26090 24512
rect 25770 24447 26090 24448
rect 11329 24306 11395 24309
rect 16297 24306 16363 24309
rect 11329 24304 16363 24306
rect 11329 24248 11334 24304
rect 11390 24248 16302 24304
rect 16358 24248 16363 24304
rect 11329 24246 16363 24248
rect 11329 24243 11395 24246
rect 16297 24243 16363 24246
rect 19977 24306 20043 24309
rect 25313 24306 25379 24309
rect 26877 24306 26943 24309
rect 19977 24304 26943 24306
rect 19977 24248 19982 24304
rect 20038 24248 25318 24304
rect 25374 24248 26882 24304
rect 26938 24248 26943 24304
rect 19977 24246 26943 24248
rect 19977 24243 20043 24246
rect 25313 24243 25379 24246
rect 26877 24243 26943 24246
rect 10874 23968 11194 23969
rect 10874 23904 10882 23968
rect 10946 23904 10962 23968
rect 11026 23904 11042 23968
rect 11106 23904 11122 23968
rect 11186 23904 11194 23968
rect 10874 23903 11194 23904
rect 20805 23968 21125 23969
rect 20805 23904 20813 23968
rect 20877 23904 20893 23968
rect 20957 23904 20973 23968
rect 21037 23904 21053 23968
rect 21117 23904 21125 23968
rect 20805 23903 21125 23904
rect 30005 23898 30071 23901
rect 31200 23898 32000 23928
rect 30005 23896 32000 23898
rect 30005 23840 30010 23896
rect 30066 23840 32000 23896
rect 30005 23838 32000 23840
rect 30005 23835 30071 23838
rect 31200 23808 32000 23838
rect 11237 23762 11303 23765
rect 14457 23762 14523 23765
rect 11237 23760 14523 23762
rect 11237 23704 11242 23760
rect 11298 23704 14462 23760
rect 14518 23704 14523 23760
rect 11237 23702 14523 23704
rect 11237 23699 11303 23702
rect 14457 23699 14523 23702
rect 16982 23564 16988 23628
rect 17052 23626 17058 23628
rect 25681 23626 25747 23629
rect 17052 23624 25747 23626
rect 17052 23568 25686 23624
rect 25742 23568 25747 23624
rect 17052 23566 25747 23568
rect 17052 23564 17058 23566
rect 25681 23563 25747 23566
rect 5909 23424 6229 23425
rect 5909 23360 5917 23424
rect 5981 23360 5997 23424
rect 6061 23360 6077 23424
rect 6141 23360 6157 23424
rect 6221 23360 6229 23424
rect 5909 23359 6229 23360
rect 15840 23424 16160 23425
rect 15840 23360 15848 23424
rect 15912 23360 15928 23424
rect 15992 23360 16008 23424
rect 16072 23360 16088 23424
rect 16152 23360 16160 23424
rect 15840 23359 16160 23360
rect 25770 23424 26090 23425
rect 25770 23360 25778 23424
rect 25842 23360 25858 23424
rect 25922 23360 25938 23424
rect 26002 23360 26018 23424
rect 26082 23360 26090 23424
rect 25770 23359 26090 23360
rect 9673 23218 9739 23221
rect 10041 23218 10107 23221
rect 9673 23216 10107 23218
rect 9673 23160 9678 23216
rect 9734 23160 10046 23216
rect 10102 23160 10107 23216
rect 9673 23158 10107 23160
rect 9673 23155 9739 23158
rect 10041 23155 10107 23158
rect 14089 23218 14155 23221
rect 15929 23218 15995 23221
rect 14089 23216 15995 23218
rect 14089 23160 14094 23216
rect 14150 23160 15934 23216
rect 15990 23160 15995 23216
rect 14089 23158 15995 23160
rect 14089 23155 14155 23158
rect 15929 23155 15995 23158
rect 28349 23218 28415 23221
rect 31200 23218 32000 23248
rect 28349 23216 32000 23218
rect 28349 23160 28354 23216
rect 28410 23160 32000 23216
rect 28349 23158 32000 23160
rect 28349 23155 28415 23158
rect 31200 23128 32000 23158
rect 0 22946 800 22976
rect 1577 22946 1643 22949
rect 0 22944 1643 22946
rect 0 22888 1582 22944
rect 1638 22888 1643 22944
rect 0 22886 1643 22888
rect 0 22856 800 22886
rect 1577 22883 1643 22886
rect 10874 22880 11194 22881
rect 10874 22816 10882 22880
rect 10946 22816 10962 22880
rect 11026 22816 11042 22880
rect 11106 22816 11122 22880
rect 11186 22816 11194 22880
rect 10874 22815 11194 22816
rect 20805 22880 21125 22881
rect 20805 22816 20813 22880
rect 20877 22816 20893 22880
rect 20957 22816 20973 22880
rect 21037 22816 21053 22880
rect 21117 22816 21125 22880
rect 20805 22815 21125 22816
rect 16757 22538 16823 22541
rect 18781 22538 18847 22541
rect 21909 22538 21975 22541
rect 16757 22536 17418 22538
rect 16757 22480 16762 22536
rect 16818 22480 17418 22536
rect 16757 22478 17418 22480
rect 16757 22475 16823 22478
rect 11329 22402 11395 22405
rect 12341 22402 12407 22405
rect 11329 22400 12407 22402
rect 11329 22344 11334 22400
rect 11390 22344 12346 22400
rect 12402 22344 12407 22400
rect 11329 22342 12407 22344
rect 11329 22339 11395 22342
rect 12341 22339 12407 22342
rect 16982 22340 16988 22404
rect 17052 22402 17058 22404
rect 17125 22402 17191 22405
rect 17052 22400 17191 22402
rect 17052 22344 17130 22400
rect 17186 22344 17191 22400
rect 17052 22342 17191 22344
rect 17052 22340 17058 22342
rect 17125 22339 17191 22342
rect 5909 22336 6229 22337
rect 5909 22272 5917 22336
rect 5981 22272 5997 22336
rect 6061 22272 6077 22336
rect 6141 22272 6157 22336
rect 6221 22272 6229 22336
rect 5909 22271 6229 22272
rect 15840 22336 16160 22337
rect 15840 22272 15848 22336
rect 15912 22272 15928 22336
rect 15992 22272 16008 22336
rect 16072 22272 16088 22336
rect 16152 22272 16160 22336
rect 15840 22271 16160 22272
rect 17358 22269 17418 22478
rect 18781 22536 21975 22538
rect 18781 22480 18786 22536
rect 18842 22480 21914 22536
rect 21970 22480 21975 22536
rect 18781 22478 21975 22480
rect 18781 22475 18847 22478
rect 21909 22475 21975 22478
rect 28901 22402 28967 22405
rect 31200 22402 32000 22432
rect 28901 22400 32000 22402
rect 28901 22344 28906 22400
rect 28962 22344 32000 22400
rect 28901 22342 32000 22344
rect 28901 22339 28967 22342
rect 25770 22336 26090 22337
rect 25770 22272 25778 22336
rect 25842 22272 25858 22336
rect 25922 22272 25938 22336
rect 26002 22272 26018 22336
rect 26082 22272 26090 22336
rect 31200 22312 32000 22342
rect 25770 22271 26090 22272
rect 17358 22264 17467 22269
rect 17358 22208 17406 22264
rect 17462 22208 17467 22264
rect 17358 22206 17467 22208
rect 17401 22203 17467 22206
rect 12433 22130 12499 22133
rect 19057 22130 19123 22133
rect 12433 22128 19123 22130
rect 12433 22072 12438 22128
rect 12494 22072 19062 22128
rect 19118 22072 19123 22128
rect 12433 22070 19123 22072
rect 12433 22067 12499 22070
rect 19057 22067 19123 22070
rect 27889 22130 27955 22133
rect 28073 22130 28139 22133
rect 28625 22130 28691 22133
rect 27889 22128 28691 22130
rect 27889 22072 27894 22128
rect 27950 22072 28078 22128
rect 28134 22072 28630 22128
rect 28686 22072 28691 22128
rect 27889 22070 28691 22072
rect 27889 22067 27955 22070
rect 28073 22067 28139 22070
rect 28625 22067 28691 22070
rect 10874 21792 11194 21793
rect 10874 21728 10882 21792
rect 10946 21728 10962 21792
rect 11026 21728 11042 21792
rect 11106 21728 11122 21792
rect 11186 21728 11194 21792
rect 10874 21727 11194 21728
rect 20805 21792 21125 21793
rect 20805 21728 20813 21792
rect 20877 21728 20893 21792
rect 20957 21728 20973 21792
rect 21037 21728 21053 21792
rect 21117 21728 21125 21792
rect 20805 21727 21125 21728
rect 17861 21722 17927 21725
rect 18689 21722 18755 21725
rect 17861 21720 18755 21722
rect 17861 21664 17866 21720
rect 17922 21664 18694 21720
rect 18750 21664 18755 21720
rect 17861 21662 18755 21664
rect 17861 21659 17927 21662
rect 18689 21659 18755 21662
rect 28901 21722 28967 21725
rect 31200 21722 32000 21752
rect 28901 21720 32000 21722
rect 28901 21664 28906 21720
rect 28962 21664 32000 21720
rect 28901 21662 32000 21664
rect 28901 21659 28967 21662
rect 31200 21632 32000 21662
rect 11053 21586 11119 21589
rect 11053 21584 12450 21586
rect 11053 21528 11058 21584
rect 11114 21528 12450 21584
rect 11053 21526 12450 21528
rect 11053 21523 11119 21526
rect 10041 21450 10107 21453
rect 12249 21450 12315 21453
rect 10041 21448 12315 21450
rect 10041 21392 10046 21448
rect 10102 21392 12254 21448
rect 12310 21392 12315 21448
rect 10041 21390 12315 21392
rect 12390 21450 12450 21526
rect 17350 21524 17356 21588
rect 17420 21586 17426 21588
rect 18965 21586 19031 21589
rect 17420 21584 19031 21586
rect 17420 21528 18970 21584
rect 19026 21528 19031 21584
rect 17420 21526 19031 21528
rect 17420 21524 17426 21526
rect 18965 21523 19031 21526
rect 20805 21450 20871 21453
rect 21541 21450 21607 21453
rect 12390 21448 21607 21450
rect 12390 21392 20810 21448
rect 20866 21392 21546 21448
rect 21602 21392 21607 21448
rect 12390 21390 21607 21392
rect 10041 21387 10107 21390
rect 12249 21387 12315 21390
rect 20805 21387 20871 21390
rect 21541 21387 21607 21390
rect 11421 21314 11487 21317
rect 12985 21314 13051 21317
rect 11421 21312 13051 21314
rect 11421 21256 11426 21312
rect 11482 21256 12990 21312
rect 13046 21256 13051 21312
rect 11421 21254 13051 21256
rect 11421 21251 11487 21254
rect 12985 21251 13051 21254
rect 20161 21314 20227 21317
rect 24761 21314 24827 21317
rect 20161 21312 24827 21314
rect 20161 21256 20166 21312
rect 20222 21256 24766 21312
rect 24822 21256 24827 21312
rect 20161 21254 24827 21256
rect 20161 21251 20227 21254
rect 24761 21251 24827 21254
rect 5909 21248 6229 21249
rect 5909 21184 5917 21248
rect 5981 21184 5997 21248
rect 6061 21184 6077 21248
rect 6141 21184 6157 21248
rect 6221 21184 6229 21248
rect 5909 21183 6229 21184
rect 15840 21248 16160 21249
rect 15840 21184 15848 21248
rect 15912 21184 15928 21248
rect 15992 21184 16008 21248
rect 16072 21184 16088 21248
rect 16152 21184 16160 21248
rect 15840 21183 16160 21184
rect 25770 21248 26090 21249
rect 25770 21184 25778 21248
rect 25842 21184 25858 21248
rect 25922 21184 25938 21248
rect 26002 21184 26018 21248
rect 26082 21184 26090 21248
rect 25770 21183 26090 21184
rect 11513 21178 11579 21181
rect 12525 21178 12591 21181
rect 11513 21176 12591 21178
rect 11513 21120 11518 21176
rect 11574 21120 12530 21176
rect 12586 21120 12591 21176
rect 11513 21118 12591 21120
rect 11513 21115 11579 21118
rect 12525 21115 12591 21118
rect 0 21042 800 21072
rect 1577 21042 1643 21045
rect 0 21040 1643 21042
rect 0 20984 1582 21040
rect 1638 20984 1643 21040
rect 0 20982 1643 20984
rect 0 20952 800 20982
rect 1577 20979 1643 20982
rect 19609 21042 19675 21045
rect 26233 21042 26299 21045
rect 19609 21040 26299 21042
rect 19609 20984 19614 21040
rect 19670 20984 26238 21040
rect 26294 20984 26299 21040
rect 19609 20982 26299 20984
rect 19609 20979 19675 20982
rect 26233 20979 26299 20982
rect 28533 21042 28599 21045
rect 31200 21042 32000 21072
rect 28533 21040 32000 21042
rect 28533 20984 28538 21040
rect 28594 20984 32000 21040
rect 28533 20982 32000 20984
rect 28533 20979 28599 20982
rect 31200 20952 32000 20982
rect 20621 20906 20687 20909
rect 21541 20906 21607 20909
rect 20621 20904 21607 20906
rect 20621 20848 20626 20904
rect 20682 20848 21546 20904
rect 21602 20848 21607 20904
rect 20621 20846 21607 20848
rect 20621 20843 20687 20846
rect 21541 20843 21607 20846
rect 10874 20704 11194 20705
rect 10874 20640 10882 20704
rect 10946 20640 10962 20704
rect 11026 20640 11042 20704
rect 11106 20640 11122 20704
rect 11186 20640 11194 20704
rect 10874 20639 11194 20640
rect 20805 20704 21125 20705
rect 20805 20640 20813 20704
rect 20877 20640 20893 20704
rect 20957 20640 20973 20704
rect 21037 20640 21053 20704
rect 21117 20640 21125 20704
rect 20805 20639 21125 20640
rect 15009 20634 15075 20637
rect 19190 20634 19196 20636
rect 15009 20632 19196 20634
rect 15009 20576 15014 20632
rect 15070 20576 19196 20632
rect 15009 20574 19196 20576
rect 15009 20571 15075 20574
rect 19190 20572 19196 20574
rect 19260 20572 19266 20636
rect 20069 20498 20135 20501
rect 21725 20498 21791 20501
rect 20069 20496 21791 20498
rect 20069 20440 20074 20496
rect 20130 20440 21730 20496
rect 21786 20440 21791 20496
rect 20069 20438 21791 20440
rect 20069 20435 20135 20438
rect 21725 20435 21791 20438
rect 28257 20226 28323 20229
rect 31200 20226 32000 20256
rect 28257 20224 32000 20226
rect 28257 20168 28262 20224
rect 28318 20168 32000 20224
rect 28257 20166 32000 20168
rect 28257 20163 28323 20166
rect 5909 20160 6229 20161
rect 5909 20096 5917 20160
rect 5981 20096 5997 20160
rect 6061 20096 6077 20160
rect 6141 20096 6157 20160
rect 6221 20096 6229 20160
rect 5909 20095 6229 20096
rect 15840 20160 16160 20161
rect 15840 20096 15848 20160
rect 15912 20096 15928 20160
rect 15992 20096 16008 20160
rect 16072 20096 16088 20160
rect 16152 20096 16160 20160
rect 15840 20095 16160 20096
rect 25770 20160 26090 20161
rect 25770 20096 25778 20160
rect 25842 20096 25858 20160
rect 25922 20096 25938 20160
rect 26002 20096 26018 20160
rect 26082 20096 26090 20160
rect 31200 20136 32000 20166
rect 25770 20095 26090 20096
rect 19425 19818 19491 19821
rect 24761 19818 24827 19821
rect 19425 19816 24827 19818
rect 19425 19760 19430 19816
rect 19486 19760 24766 19816
rect 24822 19760 24827 19816
rect 19425 19758 24827 19760
rect 19425 19755 19491 19758
rect 24761 19755 24827 19758
rect 10874 19616 11194 19617
rect 10874 19552 10882 19616
rect 10946 19552 10962 19616
rect 11026 19552 11042 19616
rect 11106 19552 11122 19616
rect 11186 19552 11194 19616
rect 10874 19551 11194 19552
rect 20805 19616 21125 19617
rect 20805 19552 20813 19616
rect 20877 19552 20893 19616
rect 20957 19552 20973 19616
rect 21037 19552 21053 19616
rect 21117 19552 21125 19616
rect 20805 19551 21125 19552
rect 28809 19546 28875 19549
rect 31200 19546 32000 19576
rect 28809 19544 32000 19546
rect 28809 19488 28814 19544
rect 28870 19488 32000 19544
rect 28809 19486 32000 19488
rect 28809 19483 28875 19486
rect 31200 19456 32000 19486
rect 22001 19410 22067 19413
rect 24669 19410 24735 19413
rect 22001 19408 24735 19410
rect 22001 19352 22006 19408
rect 22062 19352 24674 19408
rect 24730 19352 24735 19408
rect 22001 19350 24735 19352
rect 22001 19347 22067 19350
rect 24669 19347 24735 19350
rect 13813 19138 13879 19141
rect 15009 19138 15075 19141
rect 13813 19136 15075 19138
rect 13813 19080 13818 19136
rect 13874 19080 15014 19136
rect 15070 19080 15075 19136
rect 13813 19078 15075 19080
rect 13813 19075 13879 19078
rect 15009 19075 15075 19078
rect 5909 19072 6229 19073
rect 0 19002 800 19032
rect 5909 19008 5917 19072
rect 5981 19008 5997 19072
rect 6061 19008 6077 19072
rect 6141 19008 6157 19072
rect 6221 19008 6229 19072
rect 5909 19007 6229 19008
rect 15840 19072 16160 19073
rect 15840 19008 15848 19072
rect 15912 19008 15928 19072
rect 15992 19008 16008 19072
rect 16072 19008 16088 19072
rect 16152 19008 16160 19072
rect 15840 19007 16160 19008
rect 25770 19072 26090 19073
rect 25770 19008 25778 19072
rect 25842 19008 25858 19072
rect 25922 19008 25938 19072
rect 26002 19008 26018 19072
rect 26082 19008 26090 19072
rect 25770 19007 26090 19008
rect 1577 19002 1643 19005
rect 0 19000 1643 19002
rect 0 18944 1582 19000
rect 1638 18944 1643 19000
rect 0 18942 1643 18944
rect 0 18912 800 18942
rect 1577 18939 1643 18942
rect 9949 18866 10015 18869
rect 12249 18866 12315 18869
rect 9949 18864 12315 18866
rect 9949 18808 9954 18864
rect 10010 18808 12254 18864
rect 12310 18808 12315 18864
rect 9949 18806 12315 18808
rect 9949 18803 10015 18806
rect 12249 18803 12315 18806
rect 14365 18866 14431 18869
rect 14733 18866 14799 18869
rect 14365 18864 14799 18866
rect 14365 18808 14370 18864
rect 14426 18808 14738 18864
rect 14794 18808 14799 18864
rect 14365 18806 14799 18808
rect 14365 18803 14431 18806
rect 14733 18803 14799 18806
rect 24853 18730 24919 18733
rect 31200 18730 32000 18760
rect 24853 18728 32000 18730
rect 24853 18672 24858 18728
rect 24914 18672 32000 18728
rect 24853 18670 32000 18672
rect 24853 18667 24919 18670
rect 31200 18640 32000 18670
rect 10874 18528 11194 18529
rect 10874 18464 10882 18528
rect 10946 18464 10962 18528
rect 11026 18464 11042 18528
rect 11106 18464 11122 18528
rect 11186 18464 11194 18528
rect 10874 18463 11194 18464
rect 20805 18528 21125 18529
rect 20805 18464 20813 18528
rect 20877 18464 20893 18528
rect 20957 18464 20973 18528
rect 21037 18464 21053 18528
rect 21117 18464 21125 18528
rect 20805 18463 21125 18464
rect 13077 18322 13143 18325
rect 16665 18322 16731 18325
rect 13077 18320 16731 18322
rect 13077 18264 13082 18320
rect 13138 18264 16670 18320
rect 16726 18264 16731 18320
rect 13077 18262 16731 18264
rect 13077 18259 13143 18262
rect 16665 18259 16731 18262
rect 19977 18322 20043 18325
rect 24761 18322 24827 18325
rect 19977 18320 24827 18322
rect 19977 18264 19982 18320
rect 20038 18264 24766 18320
rect 24822 18264 24827 18320
rect 19977 18262 24827 18264
rect 19977 18259 20043 18262
rect 24761 18259 24827 18262
rect 19517 18186 19583 18189
rect 27705 18186 27771 18189
rect 19517 18184 27771 18186
rect 19517 18128 19522 18184
rect 19578 18128 27710 18184
rect 27766 18128 27771 18184
rect 19517 18126 27771 18128
rect 19517 18123 19583 18126
rect 27705 18123 27771 18126
rect 19425 18050 19491 18053
rect 25589 18050 25655 18053
rect 19425 18048 25655 18050
rect 19425 17992 19430 18048
rect 19486 17992 25594 18048
rect 25650 17992 25655 18048
rect 19425 17990 25655 17992
rect 19425 17987 19491 17990
rect 25589 17987 25655 17990
rect 30097 18050 30163 18053
rect 31200 18050 32000 18080
rect 30097 18048 32000 18050
rect 30097 17992 30102 18048
rect 30158 17992 32000 18048
rect 30097 17990 32000 17992
rect 30097 17987 30163 17990
rect 5909 17984 6229 17985
rect 5909 17920 5917 17984
rect 5981 17920 5997 17984
rect 6061 17920 6077 17984
rect 6141 17920 6157 17984
rect 6221 17920 6229 17984
rect 5909 17919 6229 17920
rect 15840 17984 16160 17985
rect 15840 17920 15848 17984
rect 15912 17920 15928 17984
rect 15992 17920 16008 17984
rect 16072 17920 16088 17984
rect 16152 17920 16160 17984
rect 15840 17919 16160 17920
rect 25770 17984 26090 17985
rect 25770 17920 25778 17984
rect 25842 17920 25858 17984
rect 25922 17920 25938 17984
rect 26002 17920 26018 17984
rect 26082 17920 26090 17984
rect 31200 17960 32000 17990
rect 25770 17919 26090 17920
rect 21081 17914 21147 17917
rect 23933 17914 23999 17917
rect 21081 17912 23999 17914
rect 21081 17856 21086 17912
rect 21142 17856 23938 17912
rect 23994 17856 23999 17912
rect 21081 17854 23999 17856
rect 21081 17851 21147 17854
rect 23933 17851 23999 17854
rect 13353 17778 13419 17781
rect 16297 17778 16363 17781
rect 13353 17776 16363 17778
rect 13353 17720 13358 17776
rect 13414 17720 16302 17776
rect 16358 17720 16363 17776
rect 13353 17718 16363 17720
rect 13353 17715 13419 17718
rect 16297 17715 16363 17718
rect 20345 17778 20411 17781
rect 21265 17778 21331 17781
rect 20345 17776 21331 17778
rect 20345 17720 20350 17776
rect 20406 17720 21270 17776
rect 21326 17720 21331 17776
rect 20345 17718 21331 17720
rect 20345 17715 20411 17718
rect 21265 17715 21331 17718
rect 21633 17778 21699 17781
rect 23933 17778 23999 17781
rect 21633 17776 23999 17778
rect 21633 17720 21638 17776
rect 21694 17720 23938 17776
rect 23994 17720 23999 17776
rect 21633 17718 23999 17720
rect 21633 17715 21699 17718
rect 23933 17715 23999 17718
rect 26049 17778 26115 17781
rect 27613 17778 27679 17781
rect 26049 17776 27679 17778
rect 26049 17720 26054 17776
rect 26110 17720 27618 17776
rect 27674 17720 27679 17776
rect 26049 17718 27679 17720
rect 26049 17715 26115 17718
rect 27613 17715 27679 17718
rect 20529 17642 20595 17645
rect 20805 17642 20871 17645
rect 20529 17640 20871 17642
rect 20529 17584 20534 17640
rect 20590 17584 20810 17640
rect 20866 17584 20871 17640
rect 20529 17582 20871 17584
rect 20529 17579 20595 17582
rect 20805 17579 20871 17582
rect 26417 17642 26483 17645
rect 26969 17642 27035 17645
rect 26417 17640 27035 17642
rect 26417 17584 26422 17640
rect 26478 17584 26974 17640
rect 27030 17584 27035 17640
rect 26417 17582 27035 17584
rect 26417 17579 26483 17582
rect 26969 17579 27035 17582
rect 10874 17440 11194 17441
rect 10874 17376 10882 17440
rect 10946 17376 10962 17440
rect 11026 17376 11042 17440
rect 11106 17376 11122 17440
rect 11186 17376 11194 17440
rect 10874 17375 11194 17376
rect 20805 17440 21125 17441
rect 20805 17376 20813 17440
rect 20877 17376 20893 17440
rect 20957 17376 20973 17440
rect 21037 17376 21053 17440
rect 21117 17376 21125 17440
rect 20805 17375 21125 17376
rect 19793 17370 19859 17373
rect 19793 17368 20730 17370
rect 19793 17312 19798 17368
rect 19854 17312 20730 17368
rect 19793 17310 20730 17312
rect 19793 17307 19859 17310
rect 20670 17234 20730 17310
rect 31200 17234 32000 17264
rect 20670 17174 32000 17234
rect 31200 17144 32000 17174
rect 15745 17098 15811 17101
rect 15929 17098 15995 17101
rect 15745 17096 15995 17098
rect 15745 17040 15750 17096
rect 15806 17040 15934 17096
rect 15990 17040 15995 17096
rect 15745 17038 15995 17040
rect 15745 17035 15811 17038
rect 15929 17035 15995 17038
rect 0 16962 800 16992
rect 1577 16962 1643 16965
rect 0 16960 1643 16962
rect 0 16904 1582 16960
rect 1638 16904 1643 16960
rect 0 16902 1643 16904
rect 0 16872 800 16902
rect 1577 16899 1643 16902
rect 5909 16896 6229 16897
rect 5909 16832 5917 16896
rect 5981 16832 5997 16896
rect 6061 16832 6077 16896
rect 6141 16832 6157 16896
rect 6221 16832 6229 16896
rect 5909 16831 6229 16832
rect 15840 16896 16160 16897
rect 15840 16832 15848 16896
rect 15912 16832 15928 16896
rect 15992 16832 16008 16896
rect 16072 16832 16088 16896
rect 16152 16832 16160 16896
rect 15840 16831 16160 16832
rect 25770 16896 26090 16897
rect 25770 16832 25778 16896
rect 25842 16832 25858 16896
rect 25922 16832 25938 16896
rect 26002 16832 26018 16896
rect 26082 16832 26090 16896
rect 25770 16831 26090 16832
rect 21265 16826 21331 16829
rect 21265 16824 24410 16826
rect 21265 16768 21270 16824
rect 21326 16768 24410 16824
rect 21265 16766 24410 16768
rect 21265 16763 21331 16766
rect 21173 16690 21239 16693
rect 21449 16690 21515 16693
rect 21173 16688 21515 16690
rect 21173 16632 21178 16688
rect 21234 16632 21454 16688
rect 21510 16632 21515 16688
rect 21173 16630 21515 16632
rect 21173 16627 21239 16630
rect 21449 16627 21515 16630
rect 24350 16554 24410 16766
rect 31200 16554 32000 16584
rect 24350 16494 32000 16554
rect 31200 16464 32000 16494
rect 10874 16352 11194 16353
rect 10874 16288 10882 16352
rect 10946 16288 10962 16352
rect 11026 16288 11042 16352
rect 11106 16288 11122 16352
rect 11186 16288 11194 16352
rect 10874 16287 11194 16288
rect 20805 16352 21125 16353
rect 20805 16288 20813 16352
rect 20877 16288 20893 16352
rect 20957 16288 20973 16352
rect 21037 16288 21053 16352
rect 21117 16288 21125 16352
rect 20805 16287 21125 16288
rect 28901 15874 28967 15877
rect 31200 15874 32000 15904
rect 28901 15872 32000 15874
rect 28901 15816 28906 15872
rect 28962 15816 32000 15872
rect 28901 15814 32000 15816
rect 28901 15811 28967 15814
rect 5909 15808 6229 15809
rect 5909 15744 5917 15808
rect 5981 15744 5997 15808
rect 6061 15744 6077 15808
rect 6141 15744 6157 15808
rect 6221 15744 6229 15808
rect 5909 15743 6229 15744
rect 15840 15808 16160 15809
rect 15840 15744 15848 15808
rect 15912 15744 15928 15808
rect 15992 15744 16008 15808
rect 16072 15744 16088 15808
rect 16152 15744 16160 15808
rect 15840 15743 16160 15744
rect 25770 15808 26090 15809
rect 25770 15744 25778 15808
rect 25842 15744 25858 15808
rect 25922 15744 25938 15808
rect 26002 15744 26018 15808
rect 26082 15744 26090 15808
rect 31200 15784 32000 15814
rect 25770 15743 26090 15744
rect 10874 15264 11194 15265
rect 10874 15200 10882 15264
rect 10946 15200 10962 15264
rect 11026 15200 11042 15264
rect 11106 15200 11122 15264
rect 11186 15200 11194 15264
rect 10874 15199 11194 15200
rect 20805 15264 21125 15265
rect 20805 15200 20813 15264
rect 20877 15200 20893 15264
rect 20957 15200 20973 15264
rect 21037 15200 21053 15264
rect 21117 15200 21125 15264
rect 20805 15199 21125 15200
rect 28533 15058 28599 15061
rect 31200 15058 32000 15088
rect 28533 15056 32000 15058
rect 28533 15000 28538 15056
rect 28594 15000 32000 15056
rect 28533 14998 32000 15000
rect 28533 14995 28599 14998
rect 31200 14968 32000 14998
rect 0 14922 800 14952
rect 1577 14922 1643 14925
rect 0 14920 1643 14922
rect 0 14864 1582 14920
rect 1638 14864 1643 14920
rect 0 14862 1643 14864
rect 0 14832 800 14862
rect 1577 14859 1643 14862
rect 20621 14922 20687 14925
rect 22185 14922 22251 14925
rect 20621 14920 22251 14922
rect 20621 14864 20626 14920
rect 20682 14864 22190 14920
rect 22246 14864 22251 14920
rect 20621 14862 22251 14864
rect 20621 14859 20687 14862
rect 22185 14859 22251 14862
rect 5909 14720 6229 14721
rect 5909 14656 5917 14720
rect 5981 14656 5997 14720
rect 6061 14656 6077 14720
rect 6141 14656 6157 14720
rect 6221 14656 6229 14720
rect 5909 14655 6229 14656
rect 15840 14720 16160 14721
rect 15840 14656 15848 14720
rect 15912 14656 15928 14720
rect 15992 14656 16008 14720
rect 16072 14656 16088 14720
rect 16152 14656 16160 14720
rect 15840 14655 16160 14656
rect 25770 14720 26090 14721
rect 25770 14656 25778 14720
rect 25842 14656 25858 14720
rect 25922 14656 25938 14720
rect 26002 14656 26018 14720
rect 26082 14656 26090 14720
rect 25770 14655 26090 14656
rect 21265 14378 21331 14381
rect 21398 14378 21404 14380
rect 21265 14376 21404 14378
rect 21265 14320 21270 14376
rect 21326 14320 21404 14376
rect 21265 14318 21404 14320
rect 21265 14315 21331 14318
rect 21398 14316 21404 14318
rect 21468 14378 21474 14380
rect 23197 14378 23263 14381
rect 21468 14376 23263 14378
rect 21468 14320 23202 14376
rect 23258 14320 23263 14376
rect 21468 14318 23263 14320
rect 21468 14316 21474 14318
rect 23197 14315 23263 14318
rect 28625 14378 28691 14381
rect 31200 14378 32000 14408
rect 28625 14376 32000 14378
rect 28625 14320 28630 14376
rect 28686 14320 32000 14376
rect 28625 14318 32000 14320
rect 28625 14315 28691 14318
rect 31200 14288 32000 14318
rect 10874 14176 11194 14177
rect 10874 14112 10882 14176
rect 10946 14112 10962 14176
rect 11026 14112 11042 14176
rect 11106 14112 11122 14176
rect 11186 14112 11194 14176
rect 10874 14111 11194 14112
rect 20805 14176 21125 14177
rect 20805 14112 20813 14176
rect 20877 14112 20893 14176
rect 20957 14112 20973 14176
rect 21037 14112 21053 14176
rect 21117 14112 21125 14176
rect 20805 14111 21125 14112
rect 5909 13632 6229 13633
rect 5909 13568 5917 13632
rect 5981 13568 5997 13632
rect 6061 13568 6077 13632
rect 6141 13568 6157 13632
rect 6221 13568 6229 13632
rect 5909 13567 6229 13568
rect 15840 13632 16160 13633
rect 15840 13568 15848 13632
rect 15912 13568 15928 13632
rect 15992 13568 16008 13632
rect 16072 13568 16088 13632
rect 16152 13568 16160 13632
rect 15840 13567 16160 13568
rect 25770 13632 26090 13633
rect 25770 13568 25778 13632
rect 25842 13568 25858 13632
rect 25922 13568 25938 13632
rect 26002 13568 26018 13632
rect 26082 13568 26090 13632
rect 25770 13567 26090 13568
rect 28809 13562 28875 13565
rect 31200 13562 32000 13592
rect 28809 13560 32000 13562
rect 28809 13504 28814 13560
rect 28870 13504 32000 13560
rect 28809 13502 32000 13504
rect 28809 13499 28875 13502
rect 31200 13472 32000 13502
rect 10874 13088 11194 13089
rect 0 13018 800 13048
rect 10874 13024 10882 13088
rect 10946 13024 10962 13088
rect 11026 13024 11042 13088
rect 11106 13024 11122 13088
rect 11186 13024 11194 13088
rect 10874 13023 11194 13024
rect 20805 13088 21125 13089
rect 20805 13024 20813 13088
rect 20877 13024 20893 13088
rect 20957 13024 20973 13088
rect 21037 13024 21053 13088
rect 21117 13024 21125 13088
rect 20805 13023 21125 13024
rect 1577 13018 1643 13021
rect 0 13016 1643 13018
rect 0 12960 1582 13016
rect 1638 12960 1643 13016
rect 0 12958 1643 12960
rect 0 12928 800 12958
rect 1577 12955 1643 12958
rect 28901 12882 28967 12885
rect 31200 12882 32000 12912
rect 28901 12880 32000 12882
rect 28901 12824 28906 12880
rect 28962 12824 32000 12880
rect 28901 12822 32000 12824
rect 28901 12819 28967 12822
rect 31200 12792 32000 12822
rect 20478 12548 20484 12612
rect 20548 12610 20554 12612
rect 20713 12610 20779 12613
rect 20548 12608 20779 12610
rect 20548 12552 20718 12608
rect 20774 12552 20779 12608
rect 20548 12550 20779 12552
rect 20548 12548 20554 12550
rect 20713 12547 20779 12550
rect 5909 12544 6229 12545
rect 5909 12480 5917 12544
rect 5981 12480 5997 12544
rect 6061 12480 6077 12544
rect 6141 12480 6157 12544
rect 6221 12480 6229 12544
rect 5909 12479 6229 12480
rect 15840 12544 16160 12545
rect 15840 12480 15848 12544
rect 15912 12480 15928 12544
rect 15992 12480 16008 12544
rect 16072 12480 16088 12544
rect 16152 12480 16160 12544
rect 15840 12479 16160 12480
rect 25770 12544 26090 12545
rect 25770 12480 25778 12544
rect 25842 12480 25858 12544
rect 25922 12480 25938 12544
rect 26002 12480 26018 12544
rect 26082 12480 26090 12544
rect 25770 12479 26090 12480
rect 28809 12066 28875 12069
rect 31200 12066 32000 12096
rect 28809 12064 32000 12066
rect 28809 12008 28814 12064
rect 28870 12008 32000 12064
rect 28809 12006 32000 12008
rect 28809 12003 28875 12006
rect 10874 12000 11194 12001
rect 10874 11936 10882 12000
rect 10946 11936 10962 12000
rect 11026 11936 11042 12000
rect 11106 11936 11122 12000
rect 11186 11936 11194 12000
rect 10874 11935 11194 11936
rect 20805 12000 21125 12001
rect 20805 11936 20813 12000
rect 20877 11936 20893 12000
rect 20957 11936 20973 12000
rect 21037 11936 21053 12000
rect 21117 11936 21125 12000
rect 31200 11976 32000 12006
rect 20805 11935 21125 11936
rect 21817 11930 21883 11933
rect 23013 11930 23079 11933
rect 21817 11928 23079 11930
rect 21817 11872 21822 11928
rect 21878 11872 23018 11928
rect 23074 11872 23079 11928
rect 21817 11870 23079 11872
rect 21817 11867 21883 11870
rect 22050 11661 22110 11870
rect 23013 11867 23079 11870
rect 22050 11656 22159 11661
rect 22050 11600 22098 11656
rect 22154 11600 22159 11656
rect 22050 11598 22159 11600
rect 22093 11595 22159 11598
rect 5909 11456 6229 11457
rect 5909 11392 5917 11456
rect 5981 11392 5997 11456
rect 6061 11392 6077 11456
rect 6141 11392 6157 11456
rect 6221 11392 6229 11456
rect 5909 11391 6229 11392
rect 15840 11456 16160 11457
rect 15840 11392 15848 11456
rect 15912 11392 15928 11456
rect 15992 11392 16008 11456
rect 16072 11392 16088 11456
rect 16152 11392 16160 11456
rect 15840 11391 16160 11392
rect 25770 11456 26090 11457
rect 25770 11392 25778 11456
rect 25842 11392 25858 11456
rect 25922 11392 25938 11456
rect 26002 11392 26018 11456
rect 26082 11392 26090 11456
rect 25770 11391 26090 11392
rect 27797 11386 27863 11389
rect 31200 11386 32000 11416
rect 27797 11384 32000 11386
rect 27797 11328 27802 11384
rect 27858 11328 32000 11384
rect 27797 11326 32000 11328
rect 27797 11323 27863 11326
rect 31200 11296 32000 11326
rect 21449 11116 21515 11117
rect 21398 11114 21404 11116
rect 21358 11054 21404 11114
rect 21468 11112 21515 11116
rect 21510 11056 21515 11112
rect 21398 11052 21404 11054
rect 21468 11052 21515 11056
rect 21449 11051 21515 11052
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 10874 10912 11194 10913
rect 10874 10848 10882 10912
rect 10946 10848 10962 10912
rect 11026 10848 11042 10912
rect 11106 10848 11122 10912
rect 11186 10848 11194 10912
rect 10874 10847 11194 10848
rect 20805 10912 21125 10913
rect 20805 10848 20813 10912
rect 20877 10848 20893 10912
rect 20957 10848 20973 10912
rect 21037 10848 21053 10912
rect 21117 10848 21125 10912
rect 20805 10847 21125 10848
rect 20437 10708 20503 10709
rect 20437 10706 20484 10708
rect 20392 10704 20484 10706
rect 20392 10648 20442 10704
rect 20392 10646 20484 10648
rect 20437 10644 20484 10646
rect 20548 10644 20554 10708
rect 29177 10706 29243 10709
rect 31200 10706 32000 10736
rect 29177 10704 32000 10706
rect 29177 10648 29182 10704
rect 29238 10648 32000 10704
rect 29177 10646 32000 10648
rect 20437 10643 20503 10644
rect 29177 10643 29243 10646
rect 31200 10616 32000 10646
rect 5909 10368 6229 10369
rect 5909 10304 5917 10368
rect 5981 10304 5997 10368
rect 6061 10304 6077 10368
rect 6141 10304 6157 10368
rect 6221 10304 6229 10368
rect 5909 10303 6229 10304
rect 15840 10368 16160 10369
rect 15840 10304 15848 10368
rect 15912 10304 15928 10368
rect 15992 10304 16008 10368
rect 16072 10304 16088 10368
rect 16152 10304 16160 10368
rect 15840 10303 16160 10304
rect 25770 10368 26090 10369
rect 25770 10304 25778 10368
rect 25842 10304 25858 10368
rect 25922 10304 25938 10368
rect 26002 10304 26018 10368
rect 26082 10304 26090 10368
rect 25770 10303 26090 10304
rect 30189 9890 30255 9893
rect 31200 9890 32000 9920
rect 30189 9888 32000 9890
rect 30189 9832 30194 9888
rect 30250 9832 32000 9888
rect 30189 9830 32000 9832
rect 30189 9827 30255 9830
rect 10874 9824 11194 9825
rect 10874 9760 10882 9824
rect 10946 9760 10962 9824
rect 11026 9760 11042 9824
rect 11106 9760 11122 9824
rect 11186 9760 11194 9824
rect 10874 9759 11194 9760
rect 20805 9824 21125 9825
rect 20805 9760 20813 9824
rect 20877 9760 20893 9824
rect 20957 9760 20973 9824
rect 21037 9760 21053 9824
rect 21117 9760 21125 9824
rect 31200 9800 32000 9830
rect 20805 9759 21125 9760
rect 5909 9280 6229 9281
rect 5909 9216 5917 9280
rect 5981 9216 5997 9280
rect 6061 9216 6077 9280
rect 6141 9216 6157 9280
rect 6221 9216 6229 9280
rect 5909 9215 6229 9216
rect 15840 9280 16160 9281
rect 15840 9216 15848 9280
rect 15912 9216 15928 9280
rect 15992 9216 16008 9280
rect 16072 9216 16088 9280
rect 16152 9216 16160 9280
rect 15840 9215 16160 9216
rect 25770 9280 26090 9281
rect 25770 9216 25778 9280
rect 25842 9216 25858 9280
rect 25922 9216 25938 9280
rect 26002 9216 26018 9280
rect 26082 9216 26090 9280
rect 25770 9215 26090 9216
rect 20529 9210 20595 9213
rect 22185 9210 22251 9213
rect 20529 9208 22251 9210
rect 20529 9152 20534 9208
rect 20590 9152 22190 9208
rect 22246 9152 22251 9208
rect 20529 9150 22251 9152
rect 20529 9147 20595 9150
rect 22185 9147 22251 9150
rect 30097 9210 30163 9213
rect 31200 9210 32000 9240
rect 30097 9208 32000 9210
rect 30097 9152 30102 9208
rect 30158 9152 32000 9208
rect 30097 9150 32000 9152
rect 30097 9147 30163 9150
rect 31200 9120 32000 9150
rect 20897 9074 20963 9077
rect 21173 9074 21239 9077
rect 22185 9074 22251 9077
rect 20897 9072 22251 9074
rect 20897 9016 20902 9072
rect 20958 9016 21178 9072
rect 21234 9016 22190 9072
rect 22246 9016 22251 9072
rect 20897 9014 22251 9016
rect 20897 9011 20963 9014
rect 21173 9011 21239 9014
rect 22185 9011 22251 9014
rect 0 8938 800 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 800 8878
rect 1577 8875 1643 8878
rect 10874 8736 11194 8737
rect 10874 8672 10882 8736
rect 10946 8672 10962 8736
rect 11026 8672 11042 8736
rect 11106 8672 11122 8736
rect 11186 8672 11194 8736
rect 10874 8671 11194 8672
rect 20805 8736 21125 8737
rect 20805 8672 20813 8736
rect 20877 8672 20893 8736
rect 20957 8672 20973 8736
rect 21037 8672 21053 8736
rect 21117 8672 21125 8736
rect 20805 8671 21125 8672
rect 23105 8530 23171 8533
rect 25221 8530 25287 8533
rect 23105 8528 25287 8530
rect 23105 8472 23110 8528
rect 23166 8472 25226 8528
rect 25282 8472 25287 8528
rect 23105 8470 25287 8472
rect 23105 8467 23171 8470
rect 25221 8467 25287 8470
rect 30097 8394 30163 8397
rect 31200 8394 32000 8424
rect 30097 8392 32000 8394
rect 30097 8336 30102 8392
rect 30158 8336 32000 8392
rect 30097 8334 32000 8336
rect 30097 8331 30163 8334
rect 31200 8304 32000 8334
rect 5909 8192 6229 8193
rect 5909 8128 5917 8192
rect 5981 8128 5997 8192
rect 6061 8128 6077 8192
rect 6141 8128 6157 8192
rect 6221 8128 6229 8192
rect 5909 8127 6229 8128
rect 15840 8192 16160 8193
rect 15840 8128 15848 8192
rect 15912 8128 15928 8192
rect 15992 8128 16008 8192
rect 16072 8128 16088 8192
rect 16152 8128 16160 8192
rect 15840 8127 16160 8128
rect 25770 8192 26090 8193
rect 25770 8128 25778 8192
rect 25842 8128 25858 8192
rect 25922 8128 25938 8192
rect 26002 8128 26018 8192
rect 26082 8128 26090 8192
rect 25770 8127 26090 8128
rect 30097 7714 30163 7717
rect 31200 7714 32000 7744
rect 30097 7712 32000 7714
rect 30097 7656 30102 7712
rect 30158 7656 32000 7712
rect 30097 7654 32000 7656
rect 30097 7651 30163 7654
rect 10874 7648 11194 7649
rect 10874 7584 10882 7648
rect 10946 7584 10962 7648
rect 11026 7584 11042 7648
rect 11106 7584 11122 7648
rect 11186 7584 11194 7648
rect 10874 7583 11194 7584
rect 20805 7648 21125 7649
rect 20805 7584 20813 7648
rect 20877 7584 20893 7648
rect 20957 7584 20973 7648
rect 21037 7584 21053 7648
rect 21117 7584 21125 7648
rect 31200 7624 32000 7654
rect 20805 7583 21125 7584
rect 5909 7104 6229 7105
rect 0 7034 800 7064
rect 5909 7040 5917 7104
rect 5981 7040 5997 7104
rect 6061 7040 6077 7104
rect 6141 7040 6157 7104
rect 6221 7040 6229 7104
rect 5909 7039 6229 7040
rect 15840 7104 16160 7105
rect 15840 7040 15848 7104
rect 15912 7040 15928 7104
rect 15992 7040 16008 7104
rect 16072 7040 16088 7104
rect 16152 7040 16160 7104
rect 15840 7039 16160 7040
rect 25770 7104 26090 7105
rect 25770 7040 25778 7104
rect 25842 7040 25858 7104
rect 25922 7040 25938 7104
rect 26002 7040 26018 7104
rect 26082 7040 26090 7104
rect 25770 7039 26090 7040
rect 1577 7034 1643 7037
rect 0 7032 1643 7034
rect 0 6976 1582 7032
rect 1638 6976 1643 7032
rect 0 6974 1643 6976
rect 0 6944 800 6974
rect 1577 6971 1643 6974
rect 30097 6898 30163 6901
rect 31200 6898 32000 6928
rect 30097 6896 32000 6898
rect 30097 6840 30102 6896
rect 30158 6840 32000 6896
rect 30097 6838 32000 6840
rect 30097 6835 30163 6838
rect 31200 6808 32000 6838
rect 10874 6560 11194 6561
rect 10874 6496 10882 6560
rect 10946 6496 10962 6560
rect 11026 6496 11042 6560
rect 11106 6496 11122 6560
rect 11186 6496 11194 6560
rect 10874 6495 11194 6496
rect 20805 6560 21125 6561
rect 20805 6496 20813 6560
rect 20877 6496 20893 6560
rect 20957 6496 20973 6560
rect 21037 6496 21053 6560
rect 21117 6496 21125 6560
rect 20805 6495 21125 6496
rect 30097 6218 30163 6221
rect 31200 6218 32000 6248
rect 30097 6216 32000 6218
rect 30097 6160 30102 6216
rect 30158 6160 32000 6216
rect 30097 6158 32000 6160
rect 30097 6155 30163 6158
rect 31200 6128 32000 6158
rect 5909 6016 6229 6017
rect 5909 5952 5917 6016
rect 5981 5952 5997 6016
rect 6061 5952 6077 6016
rect 6141 5952 6157 6016
rect 6221 5952 6229 6016
rect 5909 5951 6229 5952
rect 15840 6016 16160 6017
rect 15840 5952 15848 6016
rect 15912 5952 15928 6016
rect 15992 5952 16008 6016
rect 16072 5952 16088 6016
rect 16152 5952 16160 6016
rect 15840 5951 16160 5952
rect 25770 6016 26090 6017
rect 25770 5952 25778 6016
rect 25842 5952 25858 6016
rect 25922 5952 25938 6016
rect 26002 5952 26018 6016
rect 26082 5952 26090 6016
rect 25770 5951 26090 5952
rect 21357 5810 21423 5813
rect 22277 5810 22343 5813
rect 21357 5808 22343 5810
rect 21357 5752 21362 5808
rect 21418 5752 22282 5808
rect 22338 5752 22343 5808
rect 21357 5750 22343 5752
rect 21357 5747 21423 5750
rect 22277 5747 22343 5750
rect 20989 5674 21055 5677
rect 21449 5674 21515 5677
rect 20989 5672 21515 5674
rect 20989 5616 20994 5672
rect 21050 5616 21454 5672
rect 21510 5616 21515 5672
rect 20989 5614 21515 5616
rect 20989 5611 21055 5614
rect 21449 5611 21515 5614
rect 29913 5538 29979 5541
rect 31200 5538 32000 5568
rect 29913 5536 32000 5538
rect 29913 5480 29918 5536
rect 29974 5480 32000 5536
rect 29913 5478 32000 5480
rect 29913 5475 29979 5478
rect 10874 5472 11194 5473
rect 10874 5408 10882 5472
rect 10946 5408 10962 5472
rect 11026 5408 11042 5472
rect 11106 5408 11122 5472
rect 11186 5408 11194 5472
rect 10874 5407 11194 5408
rect 20805 5472 21125 5473
rect 20805 5408 20813 5472
rect 20877 5408 20893 5472
rect 20957 5408 20973 5472
rect 21037 5408 21053 5472
rect 21117 5408 21125 5472
rect 31200 5448 32000 5478
rect 20805 5407 21125 5408
rect 0 4994 800 5024
rect 1577 4994 1643 4997
rect 0 4992 1643 4994
rect 0 4936 1582 4992
rect 1638 4936 1643 4992
rect 0 4934 1643 4936
rect 0 4904 800 4934
rect 1577 4931 1643 4934
rect 5909 4928 6229 4929
rect 5909 4864 5917 4928
rect 5981 4864 5997 4928
rect 6061 4864 6077 4928
rect 6141 4864 6157 4928
rect 6221 4864 6229 4928
rect 5909 4863 6229 4864
rect 15840 4928 16160 4929
rect 15840 4864 15848 4928
rect 15912 4864 15928 4928
rect 15992 4864 16008 4928
rect 16072 4864 16088 4928
rect 16152 4864 16160 4928
rect 15840 4863 16160 4864
rect 25770 4928 26090 4929
rect 25770 4864 25778 4928
rect 25842 4864 25858 4928
rect 25922 4864 25938 4928
rect 26002 4864 26018 4928
rect 26082 4864 26090 4928
rect 25770 4863 26090 4864
rect 29913 4722 29979 4725
rect 31200 4722 32000 4752
rect 29913 4720 32000 4722
rect 29913 4664 29918 4720
rect 29974 4664 32000 4720
rect 29913 4662 32000 4664
rect 29913 4659 29979 4662
rect 31200 4632 32000 4662
rect 10874 4384 11194 4385
rect 10874 4320 10882 4384
rect 10946 4320 10962 4384
rect 11026 4320 11042 4384
rect 11106 4320 11122 4384
rect 11186 4320 11194 4384
rect 10874 4319 11194 4320
rect 20805 4384 21125 4385
rect 20805 4320 20813 4384
rect 20877 4320 20893 4384
rect 20957 4320 20973 4384
rect 21037 4320 21053 4384
rect 21117 4320 21125 4384
rect 20805 4319 21125 4320
rect 29913 4042 29979 4045
rect 31200 4042 32000 4072
rect 29913 4040 32000 4042
rect 29913 3984 29918 4040
rect 29974 3984 32000 4040
rect 29913 3982 32000 3984
rect 29913 3979 29979 3982
rect 31200 3952 32000 3982
rect 5909 3840 6229 3841
rect 5909 3776 5917 3840
rect 5981 3776 5997 3840
rect 6061 3776 6077 3840
rect 6141 3776 6157 3840
rect 6221 3776 6229 3840
rect 5909 3775 6229 3776
rect 15840 3840 16160 3841
rect 15840 3776 15848 3840
rect 15912 3776 15928 3840
rect 15992 3776 16008 3840
rect 16072 3776 16088 3840
rect 16152 3776 16160 3840
rect 15840 3775 16160 3776
rect 25770 3840 26090 3841
rect 25770 3776 25778 3840
rect 25842 3776 25858 3840
rect 25922 3776 25938 3840
rect 26002 3776 26018 3840
rect 26082 3776 26090 3840
rect 25770 3775 26090 3776
rect 10874 3296 11194 3297
rect 10874 3232 10882 3296
rect 10946 3232 10962 3296
rect 11026 3232 11042 3296
rect 11106 3232 11122 3296
rect 11186 3232 11194 3296
rect 10874 3231 11194 3232
rect 20805 3296 21125 3297
rect 20805 3232 20813 3296
rect 20877 3232 20893 3296
rect 20957 3232 20973 3296
rect 21037 3232 21053 3296
rect 21117 3232 21125 3296
rect 20805 3231 21125 3232
rect 30005 3226 30071 3229
rect 31200 3226 32000 3256
rect 30005 3224 32000 3226
rect 30005 3168 30010 3224
rect 30066 3168 32000 3224
rect 30005 3166 32000 3168
rect 30005 3163 30071 3166
rect 31200 3136 32000 3166
rect 0 2954 800 2984
rect 1577 2954 1643 2957
rect 0 2952 1643 2954
rect 0 2896 1582 2952
rect 1638 2896 1643 2952
rect 0 2894 1643 2896
rect 0 2864 800 2894
rect 1577 2891 1643 2894
rect 5909 2752 6229 2753
rect 5909 2688 5917 2752
rect 5981 2688 5997 2752
rect 6061 2688 6077 2752
rect 6141 2688 6157 2752
rect 6221 2688 6229 2752
rect 5909 2687 6229 2688
rect 15840 2752 16160 2753
rect 15840 2688 15848 2752
rect 15912 2688 15928 2752
rect 15992 2688 16008 2752
rect 16072 2688 16088 2752
rect 16152 2688 16160 2752
rect 15840 2687 16160 2688
rect 25770 2752 26090 2753
rect 25770 2688 25778 2752
rect 25842 2688 25858 2752
rect 25922 2688 25938 2752
rect 26002 2688 26018 2752
rect 26082 2688 26090 2752
rect 25770 2687 26090 2688
rect 29821 2546 29887 2549
rect 31200 2546 32000 2576
rect 29821 2544 32000 2546
rect 29821 2488 29826 2544
rect 29882 2488 32000 2544
rect 29821 2486 32000 2488
rect 29821 2483 29887 2486
rect 31200 2456 32000 2486
rect 10874 2208 11194 2209
rect 10874 2144 10882 2208
rect 10946 2144 10962 2208
rect 11026 2144 11042 2208
rect 11106 2144 11122 2208
rect 11186 2144 11194 2208
rect 10874 2143 11194 2144
rect 20805 2208 21125 2209
rect 20805 2144 20813 2208
rect 20877 2144 20893 2208
rect 20957 2144 20973 2208
rect 21037 2144 21053 2208
rect 21117 2144 21125 2208
rect 20805 2143 21125 2144
rect 29913 1730 29979 1733
rect 31200 1730 32000 1760
rect 29913 1728 32000 1730
rect 29913 1672 29918 1728
rect 29974 1672 32000 1728
rect 29913 1670 32000 1672
rect 29913 1667 29979 1670
rect 31200 1640 32000 1670
rect 0 1050 800 1080
rect 1577 1050 1643 1053
rect 0 1048 1643 1050
rect 0 992 1582 1048
rect 1638 992 1643 1048
rect 0 990 1643 992
rect 0 960 800 990
rect 1577 987 1643 990
rect 28717 1050 28783 1053
rect 31200 1050 32000 1080
rect 28717 1048 32000 1050
rect 28717 992 28722 1048
rect 28778 992 32000 1048
rect 28717 990 32000 992
rect 28717 987 28783 990
rect 31200 960 32000 990
rect 29729 370 29795 373
rect 31200 370 32000 400
rect 29729 368 32000 370
rect 29729 312 29734 368
rect 29790 312 32000 368
rect 29729 310 32000 312
rect 29729 307 29795 310
rect 31200 280 32000 310
<< via3 >>
rect 10882 45724 10946 45728
rect 10882 45668 10886 45724
rect 10886 45668 10942 45724
rect 10942 45668 10946 45724
rect 10882 45664 10946 45668
rect 10962 45724 11026 45728
rect 10962 45668 10966 45724
rect 10966 45668 11022 45724
rect 11022 45668 11026 45724
rect 10962 45664 11026 45668
rect 11042 45724 11106 45728
rect 11042 45668 11046 45724
rect 11046 45668 11102 45724
rect 11102 45668 11106 45724
rect 11042 45664 11106 45668
rect 11122 45724 11186 45728
rect 11122 45668 11126 45724
rect 11126 45668 11182 45724
rect 11182 45668 11186 45724
rect 11122 45664 11186 45668
rect 20813 45724 20877 45728
rect 20813 45668 20817 45724
rect 20817 45668 20873 45724
rect 20873 45668 20877 45724
rect 20813 45664 20877 45668
rect 20893 45724 20957 45728
rect 20893 45668 20897 45724
rect 20897 45668 20953 45724
rect 20953 45668 20957 45724
rect 20893 45664 20957 45668
rect 20973 45724 21037 45728
rect 20973 45668 20977 45724
rect 20977 45668 21033 45724
rect 21033 45668 21037 45724
rect 20973 45664 21037 45668
rect 21053 45724 21117 45728
rect 21053 45668 21057 45724
rect 21057 45668 21113 45724
rect 21113 45668 21117 45724
rect 21053 45664 21117 45668
rect 5917 45180 5981 45184
rect 5917 45124 5921 45180
rect 5921 45124 5977 45180
rect 5977 45124 5981 45180
rect 5917 45120 5981 45124
rect 5997 45180 6061 45184
rect 5997 45124 6001 45180
rect 6001 45124 6057 45180
rect 6057 45124 6061 45180
rect 5997 45120 6061 45124
rect 6077 45180 6141 45184
rect 6077 45124 6081 45180
rect 6081 45124 6137 45180
rect 6137 45124 6141 45180
rect 6077 45120 6141 45124
rect 6157 45180 6221 45184
rect 6157 45124 6161 45180
rect 6161 45124 6217 45180
rect 6217 45124 6221 45180
rect 6157 45120 6221 45124
rect 15848 45180 15912 45184
rect 15848 45124 15852 45180
rect 15852 45124 15908 45180
rect 15908 45124 15912 45180
rect 15848 45120 15912 45124
rect 15928 45180 15992 45184
rect 15928 45124 15932 45180
rect 15932 45124 15988 45180
rect 15988 45124 15992 45180
rect 15928 45120 15992 45124
rect 16008 45180 16072 45184
rect 16008 45124 16012 45180
rect 16012 45124 16068 45180
rect 16068 45124 16072 45180
rect 16008 45120 16072 45124
rect 16088 45180 16152 45184
rect 16088 45124 16092 45180
rect 16092 45124 16148 45180
rect 16148 45124 16152 45180
rect 16088 45120 16152 45124
rect 25778 45180 25842 45184
rect 25778 45124 25782 45180
rect 25782 45124 25838 45180
rect 25838 45124 25842 45180
rect 25778 45120 25842 45124
rect 25858 45180 25922 45184
rect 25858 45124 25862 45180
rect 25862 45124 25918 45180
rect 25918 45124 25922 45180
rect 25858 45120 25922 45124
rect 25938 45180 26002 45184
rect 25938 45124 25942 45180
rect 25942 45124 25998 45180
rect 25998 45124 26002 45180
rect 25938 45120 26002 45124
rect 26018 45180 26082 45184
rect 26018 45124 26022 45180
rect 26022 45124 26078 45180
rect 26078 45124 26082 45180
rect 26018 45120 26082 45124
rect 21220 44780 21284 44844
rect 10882 44636 10946 44640
rect 10882 44580 10886 44636
rect 10886 44580 10942 44636
rect 10942 44580 10946 44636
rect 10882 44576 10946 44580
rect 10962 44636 11026 44640
rect 10962 44580 10966 44636
rect 10966 44580 11022 44636
rect 11022 44580 11026 44636
rect 10962 44576 11026 44580
rect 11042 44636 11106 44640
rect 11042 44580 11046 44636
rect 11046 44580 11102 44636
rect 11102 44580 11106 44636
rect 11042 44576 11106 44580
rect 11122 44636 11186 44640
rect 11122 44580 11126 44636
rect 11126 44580 11182 44636
rect 11182 44580 11186 44636
rect 11122 44576 11186 44580
rect 20813 44636 20877 44640
rect 20813 44580 20817 44636
rect 20817 44580 20873 44636
rect 20873 44580 20877 44636
rect 20813 44576 20877 44580
rect 20893 44636 20957 44640
rect 20893 44580 20897 44636
rect 20897 44580 20953 44636
rect 20953 44580 20957 44636
rect 20893 44576 20957 44580
rect 20973 44636 21037 44640
rect 20973 44580 20977 44636
rect 20977 44580 21033 44636
rect 21033 44580 21037 44636
rect 20973 44576 21037 44580
rect 21053 44636 21117 44640
rect 21053 44580 21057 44636
rect 21057 44580 21113 44636
rect 21113 44580 21117 44636
rect 21053 44576 21117 44580
rect 5917 44092 5981 44096
rect 5917 44036 5921 44092
rect 5921 44036 5977 44092
rect 5977 44036 5981 44092
rect 5917 44032 5981 44036
rect 5997 44092 6061 44096
rect 5997 44036 6001 44092
rect 6001 44036 6057 44092
rect 6057 44036 6061 44092
rect 5997 44032 6061 44036
rect 6077 44092 6141 44096
rect 6077 44036 6081 44092
rect 6081 44036 6137 44092
rect 6137 44036 6141 44092
rect 6077 44032 6141 44036
rect 6157 44092 6221 44096
rect 6157 44036 6161 44092
rect 6161 44036 6217 44092
rect 6217 44036 6221 44092
rect 6157 44032 6221 44036
rect 15848 44092 15912 44096
rect 15848 44036 15852 44092
rect 15852 44036 15908 44092
rect 15908 44036 15912 44092
rect 15848 44032 15912 44036
rect 15928 44092 15992 44096
rect 15928 44036 15932 44092
rect 15932 44036 15988 44092
rect 15988 44036 15992 44092
rect 15928 44032 15992 44036
rect 16008 44092 16072 44096
rect 16008 44036 16012 44092
rect 16012 44036 16068 44092
rect 16068 44036 16072 44092
rect 16008 44032 16072 44036
rect 16088 44092 16152 44096
rect 16088 44036 16092 44092
rect 16092 44036 16148 44092
rect 16148 44036 16152 44092
rect 16088 44032 16152 44036
rect 25778 44092 25842 44096
rect 25778 44036 25782 44092
rect 25782 44036 25838 44092
rect 25838 44036 25842 44092
rect 25778 44032 25842 44036
rect 25858 44092 25922 44096
rect 25858 44036 25862 44092
rect 25862 44036 25918 44092
rect 25918 44036 25922 44092
rect 25858 44032 25922 44036
rect 25938 44092 26002 44096
rect 25938 44036 25942 44092
rect 25942 44036 25998 44092
rect 25998 44036 26002 44092
rect 25938 44032 26002 44036
rect 26018 44092 26082 44096
rect 26018 44036 26022 44092
rect 26022 44036 26078 44092
rect 26078 44036 26082 44092
rect 26018 44032 26082 44036
rect 10882 43548 10946 43552
rect 10882 43492 10886 43548
rect 10886 43492 10942 43548
rect 10942 43492 10946 43548
rect 10882 43488 10946 43492
rect 10962 43548 11026 43552
rect 10962 43492 10966 43548
rect 10966 43492 11022 43548
rect 11022 43492 11026 43548
rect 10962 43488 11026 43492
rect 11042 43548 11106 43552
rect 11042 43492 11046 43548
rect 11046 43492 11102 43548
rect 11102 43492 11106 43548
rect 11042 43488 11106 43492
rect 11122 43548 11186 43552
rect 11122 43492 11126 43548
rect 11126 43492 11182 43548
rect 11182 43492 11186 43548
rect 11122 43488 11186 43492
rect 20813 43548 20877 43552
rect 20813 43492 20817 43548
rect 20817 43492 20873 43548
rect 20873 43492 20877 43548
rect 20813 43488 20877 43492
rect 20893 43548 20957 43552
rect 20893 43492 20897 43548
rect 20897 43492 20953 43548
rect 20953 43492 20957 43548
rect 20893 43488 20957 43492
rect 20973 43548 21037 43552
rect 20973 43492 20977 43548
rect 20977 43492 21033 43548
rect 21033 43492 21037 43548
rect 20973 43488 21037 43492
rect 21053 43548 21117 43552
rect 21053 43492 21057 43548
rect 21057 43492 21113 43548
rect 21113 43492 21117 43548
rect 21053 43488 21117 43492
rect 5917 43004 5981 43008
rect 5917 42948 5921 43004
rect 5921 42948 5977 43004
rect 5977 42948 5981 43004
rect 5917 42944 5981 42948
rect 5997 43004 6061 43008
rect 5997 42948 6001 43004
rect 6001 42948 6057 43004
rect 6057 42948 6061 43004
rect 5997 42944 6061 42948
rect 6077 43004 6141 43008
rect 6077 42948 6081 43004
rect 6081 42948 6137 43004
rect 6137 42948 6141 43004
rect 6077 42944 6141 42948
rect 6157 43004 6221 43008
rect 6157 42948 6161 43004
rect 6161 42948 6217 43004
rect 6217 42948 6221 43004
rect 6157 42944 6221 42948
rect 15848 43004 15912 43008
rect 15848 42948 15852 43004
rect 15852 42948 15908 43004
rect 15908 42948 15912 43004
rect 15848 42944 15912 42948
rect 15928 43004 15992 43008
rect 15928 42948 15932 43004
rect 15932 42948 15988 43004
rect 15988 42948 15992 43004
rect 15928 42944 15992 42948
rect 16008 43004 16072 43008
rect 16008 42948 16012 43004
rect 16012 42948 16068 43004
rect 16068 42948 16072 43004
rect 16008 42944 16072 42948
rect 16088 43004 16152 43008
rect 16088 42948 16092 43004
rect 16092 42948 16148 43004
rect 16148 42948 16152 43004
rect 16088 42944 16152 42948
rect 25778 43004 25842 43008
rect 25778 42948 25782 43004
rect 25782 42948 25838 43004
rect 25838 42948 25842 43004
rect 25778 42944 25842 42948
rect 25858 43004 25922 43008
rect 25858 42948 25862 43004
rect 25862 42948 25918 43004
rect 25918 42948 25922 43004
rect 25858 42944 25922 42948
rect 25938 43004 26002 43008
rect 25938 42948 25942 43004
rect 25942 42948 25998 43004
rect 25998 42948 26002 43004
rect 25938 42944 26002 42948
rect 26018 43004 26082 43008
rect 26018 42948 26022 43004
rect 26022 42948 26078 43004
rect 26078 42948 26082 43004
rect 26018 42944 26082 42948
rect 10882 42460 10946 42464
rect 10882 42404 10886 42460
rect 10886 42404 10942 42460
rect 10942 42404 10946 42460
rect 10882 42400 10946 42404
rect 10962 42460 11026 42464
rect 10962 42404 10966 42460
rect 10966 42404 11022 42460
rect 11022 42404 11026 42460
rect 10962 42400 11026 42404
rect 11042 42460 11106 42464
rect 11042 42404 11046 42460
rect 11046 42404 11102 42460
rect 11102 42404 11106 42460
rect 11042 42400 11106 42404
rect 11122 42460 11186 42464
rect 11122 42404 11126 42460
rect 11126 42404 11182 42460
rect 11182 42404 11186 42460
rect 11122 42400 11186 42404
rect 20813 42460 20877 42464
rect 20813 42404 20817 42460
rect 20817 42404 20873 42460
rect 20873 42404 20877 42460
rect 20813 42400 20877 42404
rect 20893 42460 20957 42464
rect 20893 42404 20897 42460
rect 20897 42404 20953 42460
rect 20953 42404 20957 42460
rect 20893 42400 20957 42404
rect 20973 42460 21037 42464
rect 20973 42404 20977 42460
rect 20977 42404 21033 42460
rect 21033 42404 21037 42460
rect 20973 42400 21037 42404
rect 21053 42460 21117 42464
rect 21053 42404 21057 42460
rect 21057 42404 21113 42460
rect 21113 42404 21117 42460
rect 21053 42400 21117 42404
rect 5917 41916 5981 41920
rect 5917 41860 5921 41916
rect 5921 41860 5977 41916
rect 5977 41860 5981 41916
rect 5917 41856 5981 41860
rect 5997 41916 6061 41920
rect 5997 41860 6001 41916
rect 6001 41860 6057 41916
rect 6057 41860 6061 41916
rect 5997 41856 6061 41860
rect 6077 41916 6141 41920
rect 6077 41860 6081 41916
rect 6081 41860 6137 41916
rect 6137 41860 6141 41916
rect 6077 41856 6141 41860
rect 6157 41916 6221 41920
rect 6157 41860 6161 41916
rect 6161 41860 6217 41916
rect 6217 41860 6221 41916
rect 6157 41856 6221 41860
rect 15848 41916 15912 41920
rect 15848 41860 15852 41916
rect 15852 41860 15908 41916
rect 15908 41860 15912 41916
rect 15848 41856 15912 41860
rect 15928 41916 15992 41920
rect 15928 41860 15932 41916
rect 15932 41860 15988 41916
rect 15988 41860 15992 41916
rect 15928 41856 15992 41860
rect 16008 41916 16072 41920
rect 16008 41860 16012 41916
rect 16012 41860 16068 41916
rect 16068 41860 16072 41916
rect 16008 41856 16072 41860
rect 16088 41916 16152 41920
rect 16088 41860 16092 41916
rect 16092 41860 16148 41916
rect 16148 41860 16152 41916
rect 16088 41856 16152 41860
rect 25778 41916 25842 41920
rect 25778 41860 25782 41916
rect 25782 41860 25838 41916
rect 25838 41860 25842 41916
rect 25778 41856 25842 41860
rect 25858 41916 25922 41920
rect 25858 41860 25862 41916
rect 25862 41860 25918 41916
rect 25918 41860 25922 41916
rect 25858 41856 25922 41860
rect 25938 41916 26002 41920
rect 25938 41860 25942 41916
rect 25942 41860 25998 41916
rect 25998 41860 26002 41916
rect 25938 41856 26002 41860
rect 26018 41916 26082 41920
rect 26018 41860 26022 41916
rect 26022 41860 26078 41916
rect 26078 41860 26082 41916
rect 26018 41856 26082 41860
rect 10882 41372 10946 41376
rect 10882 41316 10886 41372
rect 10886 41316 10942 41372
rect 10942 41316 10946 41372
rect 10882 41312 10946 41316
rect 10962 41372 11026 41376
rect 10962 41316 10966 41372
rect 10966 41316 11022 41372
rect 11022 41316 11026 41372
rect 10962 41312 11026 41316
rect 11042 41372 11106 41376
rect 11042 41316 11046 41372
rect 11046 41316 11102 41372
rect 11102 41316 11106 41372
rect 11042 41312 11106 41316
rect 11122 41372 11186 41376
rect 11122 41316 11126 41372
rect 11126 41316 11182 41372
rect 11182 41316 11186 41372
rect 11122 41312 11186 41316
rect 20813 41372 20877 41376
rect 20813 41316 20817 41372
rect 20817 41316 20873 41372
rect 20873 41316 20877 41372
rect 20813 41312 20877 41316
rect 20893 41372 20957 41376
rect 20893 41316 20897 41372
rect 20897 41316 20953 41372
rect 20953 41316 20957 41372
rect 20893 41312 20957 41316
rect 20973 41372 21037 41376
rect 20973 41316 20977 41372
rect 20977 41316 21033 41372
rect 21033 41316 21037 41372
rect 20973 41312 21037 41316
rect 21053 41372 21117 41376
rect 21053 41316 21057 41372
rect 21057 41316 21113 41372
rect 21113 41316 21117 41372
rect 21053 41312 21117 41316
rect 5917 40828 5981 40832
rect 5917 40772 5921 40828
rect 5921 40772 5977 40828
rect 5977 40772 5981 40828
rect 5917 40768 5981 40772
rect 5997 40828 6061 40832
rect 5997 40772 6001 40828
rect 6001 40772 6057 40828
rect 6057 40772 6061 40828
rect 5997 40768 6061 40772
rect 6077 40828 6141 40832
rect 6077 40772 6081 40828
rect 6081 40772 6137 40828
rect 6137 40772 6141 40828
rect 6077 40768 6141 40772
rect 6157 40828 6221 40832
rect 6157 40772 6161 40828
rect 6161 40772 6217 40828
rect 6217 40772 6221 40828
rect 6157 40768 6221 40772
rect 15848 40828 15912 40832
rect 15848 40772 15852 40828
rect 15852 40772 15908 40828
rect 15908 40772 15912 40828
rect 15848 40768 15912 40772
rect 15928 40828 15992 40832
rect 15928 40772 15932 40828
rect 15932 40772 15988 40828
rect 15988 40772 15992 40828
rect 15928 40768 15992 40772
rect 16008 40828 16072 40832
rect 16008 40772 16012 40828
rect 16012 40772 16068 40828
rect 16068 40772 16072 40828
rect 16008 40768 16072 40772
rect 16088 40828 16152 40832
rect 16088 40772 16092 40828
rect 16092 40772 16148 40828
rect 16148 40772 16152 40828
rect 16088 40768 16152 40772
rect 25778 40828 25842 40832
rect 25778 40772 25782 40828
rect 25782 40772 25838 40828
rect 25838 40772 25842 40828
rect 25778 40768 25842 40772
rect 25858 40828 25922 40832
rect 25858 40772 25862 40828
rect 25862 40772 25918 40828
rect 25918 40772 25922 40828
rect 25858 40768 25922 40772
rect 25938 40828 26002 40832
rect 25938 40772 25942 40828
rect 25942 40772 25998 40828
rect 25998 40772 26002 40828
rect 25938 40768 26002 40772
rect 26018 40828 26082 40832
rect 26018 40772 26022 40828
rect 26022 40772 26078 40828
rect 26078 40772 26082 40828
rect 26018 40768 26082 40772
rect 21220 40564 21284 40628
rect 10882 40284 10946 40288
rect 10882 40228 10886 40284
rect 10886 40228 10942 40284
rect 10942 40228 10946 40284
rect 10882 40224 10946 40228
rect 10962 40284 11026 40288
rect 10962 40228 10966 40284
rect 10966 40228 11022 40284
rect 11022 40228 11026 40284
rect 10962 40224 11026 40228
rect 11042 40284 11106 40288
rect 11042 40228 11046 40284
rect 11046 40228 11102 40284
rect 11102 40228 11106 40284
rect 11042 40224 11106 40228
rect 11122 40284 11186 40288
rect 11122 40228 11126 40284
rect 11126 40228 11182 40284
rect 11182 40228 11186 40284
rect 11122 40224 11186 40228
rect 20813 40284 20877 40288
rect 20813 40228 20817 40284
rect 20817 40228 20873 40284
rect 20873 40228 20877 40284
rect 20813 40224 20877 40228
rect 20893 40284 20957 40288
rect 20893 40228 20897 40284
rect 20897 40228 20953 40284
rect 20953 40228 20957 40284
rect 20893 40224 20957 40228
rect 20973 40284 21037 40288
rect 20973 40228 20977 40284
rect 20977 40228 21033 40284
rect 21033 40228 21037 40284
rect 20973 40224 21037 40228
rect 21053 40284 21117 40288
rect 21053 40228 21057 40284
rect 21057 40228 21113 40284
rect 21113 40228 21117 40284
rect 21053 40224 21117 40228
rect 5917 39740 5981 39744
rect 5917 39684 5921 39740
rect 5921 39684 5977 39740
rect 5977 39684 5981 39740
rect 5917 39680 5981 39684
rect 5997 39740 6061 39744
rect 5997 39684 6001 39740
rect 6001 39684 6057 39740
rect 6057 39684 6061 39740
rect 5997 39680 6061 39684
rect 6077 39740 6141 39744
rect 6077 39684 6081 39740
rect 6081 39684 6137 39740
rect 6137 39684 6141 39740
rect 6077 39680 6141 39684
rect 6157 39740 6221 39744
rect 6157 39684 6161 39740
rect 6161 39684 6217 39740
rect 6217 39684 6221 39740
rect 6157 39680 6221 39684
rect 15848 39740 15912 39744
rect 15848 39684 15852 39740
rect 15852 39684 15908 39740
rect 15908 39684 15912 39740
rect 15848 39680 15912 39684
rect 15928 39740 15992 39744
rect 15928 39684 15932 39740
rect 15932 39684 15988 39740
rect 15988 39684 15992 39740
rect 15928 39680 15992 39684
rect 16008 39740 16072 39744
rect 16008 39684 16012 39740
rect 16012 39684 16068 39740
rect 16068 39684 16072 39740
rect 16008 39680 16072 39684
rect 16088 39740 16152 39744
rect 16088 39684 16092 39740
rect 16092 39684 16148 39740
rect 16148 39684 16152 39740
rect 16088 39680 16152 39684
rect 25778 39740 25842 39744
rect 25778 39684 25782 39740
rect 25782 39684 25838 39740
rect 25838 39684 25842 39740
rect 25778 39680 25842 39684
rect 25858 39740 25922 39744
rect 25858 39684 25862 39740
rect 25862 39684 25918 39740
rect 25918 39684 25922 39740
rect 25858 39680 25922 39684
rect 25938 39740 26002 39744
rect 25938 39684 25942 39740
rect 25942 39684 25998 39740
rect 25998 39684 26002 39740
rect 25938 39680 26002 39684
rect 26018 39740 26082 39744
rect 26018 39684 26022 39740
rect 26022 39684 26078 39740
rect 26078 39684 26082 39740
rect 26018 39680 26082 39684
rect 10882 39196 10946 39200
rect 10882 39140 10886 39196
rect 10886 39140 10942 39196
rect 10942 39140 10946 39196
rect 10882 39136 10946 39140
rect 10962 39196 11026 39200
rect 10962 39140 10966 39196
rect 10966 39140 11022 39196
rect 11022 39140 11026 39196
rect 10962 39136 11026 39140
rect 11042 39196 11106 39200
rect 11042 39140 11046 39196
rect 11046 39140 11102 39196
rect 11102 39140 11106 39196
rect 11042 39136 11106 39140
rect 11122 39196 11186 39200
rect 11122 39140 11126 39196
rect 11126 39140 11182 39196
rect 11182 39140 11186 39196
rect 11122 39136 11186 39140
rect 20813 39196 20877 39200
rect 20813 39140 20817 39196
rect 20817 39140 20873 39196
rect 20873 39140 20877 39196
rect 20813 39136 20877 39140
rect 20893 39196 20957 39200
rect 20893 39140 20897 39196
rect 20897 39140 20953 39196
rect 20953 39140 20957 39196
rect 20893 39136 20957 39140
rect 20973 39196 21037 39200
rect 20973 39140 20977 39196
rect 20977 39140 21033 39196
rect 21033 39140 21037 39196
rect 20973 39136 21037 39140
rect 21053 39196 21117 39200
rect 21053 39140 21057 39196
rect 21057 39140 21113 39196
rect 21113 39140 21117 39196
rect 21053 39136 21117 39140
rect 5917 38652 5981 38656
rect 5917 38596 5921 38652
rect 5921 38596 5977 38652
rect 5977 38596 5981 38652
rect 5917 38592 5981 38596
rect 5997 38652 6061 38656
rect 5997 38596 6001 38652
rect 6001 38596 6057 38652
rect 6057 38596 6061 38652
rect 5997 38592 6061 38596
rect 6077 38652 6141 38656
rect 6077 38596 6081 38652
rect 6081 38596 6137 38652
rect 6137 38596 6141 38652
rect 6077 38592 6141 38596
rect 6157 38652 6221 38656
rect 6157 38596 6161 38652
rect 6161 38596 6217 38652
rect 6217 38596 6221 38652
rect 6157 38592 6221 38596
rect 15848 38652 15912 38656
rect 15848 38596 15852 38652
rect 15852 38596 15908 38652
rect 15908 38596 15912 38652
rect 15848 38592 15912 38596
rect 15928 38652 15992 38656
rect 15928 38596 15932 38652
rect 15932 38596 15988 38652
rect 15988 38596 15992 38652
rect 15928 38592 15992 38596
rect 16008 38652 16072 38656
rect 16008 38596 16012 38652
rect 16012 38596 16068 38652
rect 16068 38596 16072 38652
rect 16008 38592 16072 38596
rect 16088 38652 16152 38656
rect 16088 38596 16092 38652
rect 16092 38596 16148 38652
rect 16148 38596 16152 38652
rect 16088 38592 16152 38596
rect 25778 38652 25842 38656
rect 25778 38596 25782 38652
rect 25782 38596 25838 38652
rect 25838 38596 25842 38652
rect 25778 38592 25842 38596
rect 25858 38652 25922 38656
rect 25858 38596 25862 38652
rect 25862 38596 25918 38652
rect 25918 38596 25922 38652
rect 25858 38592 25922 38596
rect 25938 38652 26002 38656
rect 25938 38596 25942 38652
rect 25942 38596 25998 38652
rect 25998 38596 26002 38652
rect 25938 38592 26002 38596
rect 26018 38652 26082 38656
rect 26018 38596 26022 38652
rect 26022 38596 26078 38652
rect 26078 38596 26082 38652
rect 26018 38592 26082 38596
rect 10882 38108 10946 38112
rect 10882 38052 10886 38108
rect 10886 38052 10942 38108
rect 10942 38052 10946 38108
rect 10882 38048 10946 38052
rect 10962 38108 11026 38112
rect 10962 38052 10966 38108
rect 10966 38052 11022 38108
rect 11022 38052 11026 38108
rect 10962 38048 11026 38052
rect 11042 38108 11106 38112
rect 11042 38052 11046 38108
rect 11046 38052 11102 38108
rect 11102 38052 11106 38108
rect 11042 38048 11106 38052
rect 11122 38108 11186 38112
rect 11122 38052 11126 38108
rect 11126 38052 11182 38108
rect 11182 38052 11186 38108
rect 11122 38048 11186 38052
rect 20813 38108 20877 38112
rect 20813 38052 20817 38108
rect 20817 38052 20873 38108
rect 20873 38052 20877 38108
rect 20813 38048 20877 38052
rect 20893 38108 20957 38112
rect 20893 38052 20897 38108
rect 20897 38052 20953 38108
rect 20953 38052 20957 38108
rect 20893 38048 20957 38052
rect 20973 38108 21037 38112
rect 20973 38052 20977 38108
rect 20977 38052 21033 38108
rect 21033 38052 21037 38108
rect 20973 38048 21037 38052
rect 21053 38108 21117 38112
rect 21053 38052 21057 38108
rect 21057 38052 21113 38108
rect 21113 38052 21117 38108
rect 21053 38048 21117 38052
rect 5917 37564 5981 37568
rect 5917 37508 5921 37564
rect 5921 37508 5977 37564
rect 5977 37508 5981 37564
rect 5917 37504 5981 37508
rect 5997 37564 6061 37568
rect 5997 37508 6001 37564
rect 6001 37508 6057 37564
rect 6057 37508 6061 37564
rect 5997 37504 6061 37508
rect 6077 37564 6141 37568
rect 6077 37508 6081 37564
rect 6081 37508 6137 37564
rect 6137 37508 6141 37564
rect 6077 37504 6141 37508
rect 6157 37564 6221 37568
rect 6157 37508 6161 37564
rect 6161 37508 6217 37564
rect 6217 37508 6221 37564
rect 6157 37504 6221 37508
rect 15848 37564 15912 37568
rect 15848 37508 15852 37564
rect 15852 37508 15908 37564
rect 15908 37508 15912 37564
rect 15848 37504 15912 37508
rect 15928 37564 15992 37568
rect 15928 37508 15932 37564
rect 15932 37508 15988 37564
rect 15988 37508 15992 37564
rect 15928 37504 15992 37508
rect 16008 37564 16072 37568
rect 16008 37508 16012 37564
rect 16012 37508 16068 37564
rect 16068 37508 16072 37564
rect 16008 37504 16072 37508
rect 16088 37564 16152 37568
rect 16088 37508 16092 37564
rect 16092 37508 16148 37564
rect 16148 37508 16152 37564
rect 16088 37504 16152 37508
rect 25778 37564 25842 37568
rect 25778 37508 25782 37564
rect 25782 37508 25838 37564
rect 25838 37508 25842 37564
rect 25778 37504 25842 37508
rect 25858 37564 25922 37568
rect 25858 37508 25862 37564
rect 25862 37508 25918 37564
rect 25918 37508 25922 37564
rect 25858 37504 25922 37508
rect 25938 37564 26002 37568
rect 25938 37508 25942 37564
rect 25942 37508 25998 37564
rect 25998 37508 26002 37564
rect 25938 37504 26002 37508
rect 26018 37564 26082 37568
rect 26018 37508 26022 37564
rect 26022 37508 26078 37564
rect 26078 37508 26082 37564
rect 26018 37504 26082 37508
rect 10882 37020 10946 37024
rect 10882 36964 10886 37020
rect 10886 36964 10942 37020
rect 10942 36964 10946 37020
rect 10882 36960 10946 36964
rect 10962 37020 11026 37024
rect 10962 36964 10966 37020
rect 10966 36964 11022 37020
rect 11022 36964 11026 37020
rect 10962 36960 11026 36964
rect 11042 37020 11106 37024
rect 11042 36964 11046 37020
rect 11046 36964 11102 37020
rect 11102 36964 11106 37020
rect 11042 36960 11106 36964
rect 11122 37020 11186 37024
rect 11122 36964 11126 37020
rect 11126 36964 11182 37020
rect 11182 36964 11186 37020
rect 11122 36960 11186 36964
rect 20813 37020 20877 37024
rect 20813 36964 20817 37020
rect 20817 36964 20873 37020
rect 20873 36964 20877 37020
rect 20813 36960 20877 36964
rect 20893 37020 20957 37024
rect 20893 36964 20897 37020
rect 20897 36964 20953 37020
rect 20953 36964 20957 37020
rect 20893 36960 20957 36964
rect 20973 37020 21037 37024
rect 20973 36964 20977 37020
rect 20977 36964 21033 37020
rect 21033 36964 21037 37020
rect 20973 36960 21037 36964
rect 21053 37020 21117 37024
rect 21053 36964 21057 37020
rect 21057 36964 21113 37020
rect 21113 36964 21117 37020
rect 21053 36960 21117 36964
rect 5917 36476 5981 36480
rect 5917 36420 5921 36476
rect 5921 36420 5977 36476
rect 5977 36420 5981 36476
rect 5917 36416 5981 36420
rect 5997 36476 6061 36480
rect 5997 36420 6001 36476
rect 6001 36420 6057 36476
rect 6057 36420 6061 36476
rect 5997 36416 6061 36420
rect 6077 36476 6141 36480
rect 6077 36420 6081 36476
rect 6081 36420 6137 36476
rect 6137 36420 6141 36476
rect 6077 36416 6141 36420
rect 6157 36476 6221 36480
rect 6157 36420 6161 36476
rect 6161 36420 6217 36476
rect 6217 36420 6221 36476
rect 6157 36416 6221 36420
rect 15848 36476 15912 36480
rect 15848 36420 15852 36476
rect 15852 36420 15908 36476
rect 15908 36420 15912 36476
rect 15848 36416 15912 36420
rect 15928 36476 15992 36480
rect 15928 36420 15932 36476
rect 15932 36420 15988 36476
rect 15988 36420 15992 36476
rect 15928 36416 15992 36420
rect 16008 36476 16072 36480
rect 16008 36420 16012 36476
rect 16012 36420 16068 36476
rect 16068 36420 16072 36476
rect 16008 36416 16072 36420
rect 16088 36476 16152 36480
rect 16088 36420 16092 36476
rect 16092 36420 16148 36476
rect 16148 36420 16152 36476
rect 16088 36416 16152 36420
rect 25778 36476 25842 36480
rect 25778 36420 25782 36476
rect 25782 36420 25838 36476
rect 25838 36420 25842 36476
rect 25778 36416 25842 36420
rect 25858 36476 25922 36480
rect 25858 36420 25862 36476
rect 25862 36420 25918 36476
rect 25918 36420 25922 36476
rect 25858 36416 25922 36420
rect 25938 36476 26002 36480
rect 25938 36420 25942 36476
rect 25942 36420 25998 36476
rect 25998 36420 26002 36476
rect 25938 36416 26002 36420
rect 26018 36476 26082 36480
rect 26018 36420 26022 36476
rect 26022 36420 26078 36476
rect 26078 36420 26082 36476
rect 26018 36416 26082 36420
rect 18644 36272 18708 36276
rect 18644 36216 18658 36272
rect 18658 36216 18708 36272
rect 18644 36212 18708 36216
rect 10882 35932 10946 35936
rect 10882 35876 10886 35932
rect 10886 35876 10942 35932
rect 10942 35876 10946 35932
rect 10882 35872 10946 35876
rect 10962 35932 11026 35936
rect 10962 35876 10966 35932
rect 10966 35876 11022 35932
rect 11022 35876 11026 35932
rect 10962 35872 11026 35876
rect 11042 35932 11106 35936
rect 11042 35876 11046 35932
rect 11046 35876 11102 35932
rect 11102 35876 11106 35932
rect 11042 35872 11106 35876
rect 11122 35932 11186 35936
rect 11122 35876 11126 35932
rect 11126 35876 11182 35932
rect 11182 35876 11186 35932
rect 11122 35872 11186 35876
rect 20813 35932 20877 35936
rect 20813 35876 20817 35932
rect 20817 35876 20873 35932
rect 20873 35876 20877 35932
rect 20813 35872 20877 35876
rect 20893 35932 20957 35936
rect 20893 35876 20897 35932
rect 20897 35876 20953 35932
rect 20953 35876 20957 35932
rect 20893 35872 20957 35876
rect 20973 35932 21037 35936
rect 20973 35876 20977 35932
rect 20977 35876 21033 35932
rect 21033 35876 21037 35932
rect 20973 35872 21037 35876
rect 21053 35932 21117 35936
rect 21053 35876 21057 35932
rect 21057 35876 21113 35932
rect 21113 35876 21117 35932
rect 21053 35872 21117 35876
rect 5917 35388 5981 35392
rect 5917 35332 5921 35388
rect 5921 35332 5977 35388
rect 5977 35332 5981 35388
rect 5917 35328 5981 35332
rect 5997 35388 6061 35392
rect 5997 35332 6001 35388
rect 6001 35332 6057 35388
rect 6057 35332 6061 35388
rect 5997 35328 6061 35332
rect 6077 35388 6141 35392
rect 6077 35332 6081 35388
rect 6081 35332 6137 35388
rect 6137 35332 6141 35388
rect 6077 35328 6141 35332
rect 6157 35388 6221 35392
rect 6157 35332 6161 35388
rect 6161 35332 6217 35388
rect 6217 35332 6221 35388
rect 6157 35328 6221 35332
rect 15848 35388 15912 35392
rect 15848 35332 15852 35388
rect 15852 35332 15908 35388
rect 15908 35332 15912 35388
rect 15848 35328 15912 35332
rect 15928 35388 15992 35392
rect 15928 35332 15932 35388
rect 15932 35332 15988 35388
rect 15988 35332 15992 35388
rect 15928 35328 15992 35332
rect 16008 35388 16072 35392
rect 16008 35332 16012 35388
rect 16012 35332 16068 35388
rect 16068 35332 16072 35388
rect 16008 35328 16072 35332
rect 16088 35388 16152 35392
rect 16088 35332 16092 35388
rect 16092 35332 16148 35388
rect 16148 35332 16152 35388
rect 16088 35328 16152 35332
rect 25778 35388 25842 35392
rect 25778 35332 25782 35388
rect 25782 35332 25838 35388
rect 25838 35332 25842 35388
rect 25778 35328 25842 35332
rect 25858 35388 25922 35392
rect 25858 35332 25862 35388
rect 25862 35332 25918 35388
rect 25918 35332 25922 35388
rect 25858 35328 25922 35332
rect 25938 35388 26002 35392
rect 25938 35332 25942 35388
rect 25942 35332 25998 35388
rect 25998 35332 26002 35388
rect 25938 35328 26002 35332
rect 26018 35388 26082 35392
rect 26018 35332 26022 35388
rect 26022 35332 26078 35388
rect 26078 35332 26082 35388
rect 26018 35328 26082 35332
rect 19012 35048 19076 35052
rect 19012 34992 19062 35048
rect 19062 34992 19076 35048
rect 19012 34988 19076 34992
rect 10882 34844 10946 34848
rect 10882 34788 10886 34844
rect 10886 34788 10942 34844
rect 10942 34788 10946 34844
rect 10882 34784 10946 34788
rect 10962 34844 11026 34848
rect 10962 34788 10966 34844
rect 10966 34788 11022 34844
rect 11022 34788 11026 34844
rect 10962 34784 11026 34788
rect 11042 34844 11106 34848
rect 11042 34788 11046 34844
rect 11046 34788 11102 34844
rect 11102 34788 11106 34844
rect 11042 34784 11106 34788
rect 11122 34844 11186 34848
rect 11122 34788 11126 34844
rect 11126 34788 11182 34844
rect 11182 34788 11186 34844
rect 11122 34784 11186 34788
rect 17356 34580 17420 34644
rect 20813 34844 20877 34848
rect 20813 34788 20817 34844
rect 20817 34788 20873 34844
rect 20873 34788 20877 34844
rect 20813 34784 20877 34788
rect 20893 34844 20957 34848
rect 20893 34788 20897 34844
rect 20897 34788 20953 34844
rect 20953 34788 20957 34844
rect 20893 34784 20957 34788
rect 20973 34844 21037 34848
rect 20973 34788 20977 34844
rect 20977 34788 21033 34844
rect 21033 34788 21037 34844
rect 20973 34784 21037 34788
rect 21053 34844 21117 34848
rect 21053 34788 21057 34844
rect 21057 34788 21113 34844
rect 21113 34788 21117 34844
rect 21053 34784 21117 34788
rect 5917 34300 5981 34304
rect 5917 34244 5921 34300
rect 5921 34244 5977 34300
rect 5977 34244 5981 34300
rect 5917 34240 5981 34244
rect 5997 34300 6061 34304
rect 5997 34244 6001 34300
rect 6001 34244 6057 34300
rect 6057 34244 6061 34300
rect 5997 34240 6061 34244
rect 6077 34300 6141 34304
rect 6077 34244 6081 34300
rect 6081 34244 6137 34300
rect 6137 34244 6141 34300
rect 6077 34240 6141 34244
rect 6157 34300 6221 34304
rect 6157 34244 6161 34300
rect 6161 34244 6217 34300
rect 6217 34244 6221 34300
rect 6157 34240 6221 34244
rect 15848 34300 15912 34304
rect 15848 34244 15852 34300
rect 15852 34244 15908 34300
rect 15908 34244 15912 34300
rect 15848 34240 15912 34244
rect 15928 34300 15992 34304
rect 15928 34244 15932 34300
rect 15932 34244 15988 34300
rect 15988 34244 15992 34300
rect 15928 34240 15992 34244
rect 16008 34300 16072 34304
rect 16008 34244 16012 34300
rect 16012 34244 16068 34300
rect 16068 34244 16072 34300
rect 16008 34240 16072 34244
rect 16088 34300 16152 34304
rect 16088 34244 16092 34300
rect 16092 34244 16148 34300
rect 16148 34244 16152 34300
rect 16088 34240 16152 34244
rect 25778 34300 25842 34304
rect 25778 34244 25782 34300
rect 25782 34244 25838 34300
rect 25838 34244 25842 34300
rect 25778 34240 25842 34244
rect 25858 34300 25922 34304
rect 25858 34244 25862 34300
rect 25862 34244 25918 34300
rect 25918 34244 25922 34300
rect 25858 34240 25922 34244
rect 25938 34300 26002 34304
rect 25938 34244 25942 34300
rect 25942 34244 25998 34300
rect 25998 34244 26002 34300
rect 25938 34240 26002 34244
rect 26018 34300 26082 34304
rect 26018 34244 26022 34300
rect 26022 34244 26078 34300
rect 26078 34244 26082 34300
rect 26018 34240 26082 34244
rect 16620 33900 16684 33964
rect 19012 33764 19076 33828
rect 10882 33756 10946 33760
rect 10882 33700 10886 33756
rect 10886 33700 10942 33756
rect 10942 33700 10946 33756
rect 10882 33696 10946 33700
rect 10962 33756 11026 33760
rect 10962 33700 10966 33756
rect 10966 33700 11022 33756
rect 11022 33700 11026 33756
rect 10962 33696 11026 33700
rect 11042 33756 11106 33760
rect 11042 33700 11046 33756
rect 11046 33700 11102 33756
rect 11102 33700 11106 33756
rect 11042 33696 11106 33700
rect 11122 33756 11186 33760
rect 11122 33700 11126 33756
rect 11126 33700 11182 33756
rect 11182 33700 11186 33756
rect 11122 33696 11186 33700
rect 20813 33756 20877 33760
rect 20813 33700 20817 33756
rect 20817 33700 20873 33756
rect 20873 33700 20877 33756
rect 20813 33696 20877 33700
rect 20893 33756 20957 33760
rect 20893 33700 20897 33756
rect 20897 33700 20953 33756
rect 20953 33700 20957 33756
rect 20893 33696 20957 33700
rect 20973 33756 21037 33760
rect 20973 33700 20977 33756
rect 20977 33700 21033 33756
rect 21033 33700 21037 33756
rect 20973 33696 21037 33700
rect 21053 33756 21117 33760
rect 21053 33700 21057 33756
rect 21057 33700 21113 33756
rect 21113 33700 21117 33756
rect 21053 33696 21117 33700
rect 5917 33212 5981 33216
rect 5917 33156 5921 33212
rect 5921 33156 5977 33212
rect 5977 33156 5981 33212
rect 5917 33152 5981 33156
rect 5997 33212 6061 33216
rect 5997 33156 6001 33212
rect 6001 33156 6057 33212
rect 6057 33156 6061 33212
rect 5997 33152 6061 33156
rect 6077 33212 6141 33216
rect 6077 33156 6081 33212
rect 6081 33156 6137 33212
rect 6137 33156 6141 33212
rect 6077 33152 6141 33156
rect 6157 33212 6221 33216
rect 6157 33156 6161 33212
rect 6161 33156 6217 33212
rect 6217 33156 6221 33212
rect 6157 33152 6221 33156
rect 15848 33212 15912 33216
rect 15848 33156 15852 33212
rect 15852 33156 15908 33212
rect 15908 33156 15912 33212
rect 15848 33152 15912 33156
rect 15928 33212 15992 33216
rect 15928 33156 15932 33212
rect 15932 33156 15988 33212
rect 15988 33156 15992 33212
rect 15928 33152 15992 33156
rect 16008 33212 16072 33216
rect 16008 33156 16012 33212
rect 16012 33156 16068 33212
rect 16068 33156 16072 33212
rect 16008 33152 16072 33156
rect 16088 33212 16152 33216
rect 16088 33156 16092 33212
rect 16092 33156 16148 33212
rect 16148 33156 16152 33212
rect 16088 33152 16152 33156
rect 25778 33212 25842 33216
rect 25778 33156 25782 33212
rect 25782 33156 25838 33212
rect 25838 33156 25842 33212
rect 25778 33152 25842 33156
rect 25858 33212 25922 33216
rect 25858 33156 25862 33212
rect 25862 33156 25918 33212
rect 25918 33156 25922 33212
rect 25858 33152 25922 33156
rect 25938 33212 26002 33216
rect 25938 33156 25942 33212
rect 25942 33156 25998 33212
rect 25998 33156 26002 33212
rect 25938 33152 26002 33156
rect 26018 33212 26082 33216
rect 26018 33156 26022 33212
rect 26022 33156 26078 33212
rect 26078 33156 26082 33212
rect 26018 33152 26082 33156
rect 10882 32668 10946 32672
rect 10882 32612 10886 32668
rect 10886 32612 10942 32668
rect 10942 32612 10946 32668
rect 10882 32608 10946 32612
rect 10962 32668 11026 32672
rect 10962 32612 10966 32668
rect 10966 32612 11022 32668
rect 11022 32612 11026 32668
rect 10962 32608 11026 32612
rect 11042 32668 11106 32672
rect 11042 32612 11046 32668
rect 11046 32612 11102 32668
rect 11102 32612 11106 32668
rect 11042 32608 11106 32612
rect 11122 32668 11186 32672
rect 11122 32612 11126 32668
rect 11126 32612 11182 32668
rect 11182 32612 11186 32668
rect 11122 32608 11186 32612
rect 20813 32668 20877 32672
rect 20813 32612 20817 32668
rect 20817 32612 20873 32668
rect 20873 32612 20877 32668
rect 20813 32608 20877 32612
rect 20893 32668 20957 32672
rect 20893 32612 20897 32668
rect 20897 32612 20953 32668
rect 20953 32612 20957 32668
rect 20893 32608 20957 32612
rect 20973 32668 21037 32672
rect 20973 32612 20977 32668
rect 20977 32612 21033 32668
rect 21033 32612 21037 32668
rect 20973 32608 21037 32612
rect 21053 32668 21117 32672
rect 21053 32612 21057 32668
rect 21057 32612 21113 32668
rect 21113 32612 21117 32668
rect 21053 32608 21117 32612
rect 5917 32124 5981 32128
rect 5917 32068 5921 32124
rect 5921 32068 5977 32124
rect 5977 32068 5981 32124
rect 5917 32064 5981 32068
rect 5997 32124 6061 32128
rect 5997 32068 6001 32124
rect 6001 32068 6057 32124
rect 6057 32068 6061 32124
rect 5997 32064 6061 32068
rect 6077 32124 6141 32128
rect 6077 32068 6081 32124
rect 6081 32068 6137 32124
rect 6137 32068 6141 32124
rect 6077 32064 6141 32068
rect 6157 32124 6221 32128
rect 6157 32068 6161 32124
rect 6161 32068 6217 32124
rect 6217 32068 6221 32124
rect 6157 32064 6221 32068
rect 15848 32124 15912 32128
rect 15848 32068 15852 32124
rect 15852 32068 15908 32124
rect 15908 32068 15912 32124
rect 15848 32064 15912 32068
rect 15928 32124 15992 32128
rect 15928 32068 15932 32124
rect 15932 32068 15988 32124
rect 15988 32068 15992 32124
rect 15928 32064 15992 32068
rect 16008 32124 16072 32128
rect 16008 32068 16012 32124
rect 16012 32068 16068 32124
rect 16068 32068 16072 32124
rect 16008 32064 16072 32068
rect 16088 32124 16152 32128
rect 16088 32068 16092 32124
rect 16092 32068 16148 32124
rect 16148 32068 16152 32124
rect 16088 32064 16152 32068
rect 25778 32124 25842 32128
rect 25778 32068 25782 32124
rect 25782 32068 25838 32124
rect 25838 32068 25842 32124
rect 25778 32064 25842 32068
rect 25858 32124 25922 32128
rect 25858 32068 25862 32124
rect 25862 32068 25918 32124
rect 25918 32068 25922 32124
rect 25858 32064 25922 32068
rect 25938 32124 26002 32128
rect 25938 32068 25942 32124
rect 25942 32068 25998 32124
rect 25998 32068 26002 32124
rect 25938 32064 26002 32068
rect 26018 32124 26082 32128
rect 26018 32068 26022 32124
rect 26022 32068 26078 32124
rect 26078 32068 26082 32124
rect 26018 32064 26082 32068
rect 17540 31860 17604 31924
rect 10882 31580 10946 31584
rect 10882 31524 10886 31580
rect 10886 31524 10942 31580
rect 10942 31524 10946 31580
rect 10882 31520 10946 31524
rect 10962 31580 11026 31584
rect 10962 31524 10966 31580
rect 10966 31524 11022 31580
rect 11022 31524 11026 31580
rect 10962 31520 11026 31524
rect 11042 31580 11106 31584
rect 11042 31524 11046 31580
rect 11046 31524 11102 31580
rect 11102 31524 11106 31580
rect 11042 31520 11106 31524
rect 11122 31580 11186 31584
rect 11122 31524 11126 31580
rect 11126 31524 11182 31580
rect 11182 31524 11186 31580
rect 11122 31520 11186 31524
rect 20813 31580 20877 31584
rect 20813 31524 20817 31580
rect 20817 31524 20873 31580
rect 20873 31524 20877 31580
rect 20813 31520 20877 31524
rect 20893 31580 20957 31584
rect 20893 31524 20897 31580
rect 20897 31524 20953 31580
rect 20953 31524 20957 31580
rect 20893 31520 20957 31524
rect 20973 31580 21037 31584
rect 20973 31524 20977 31580
rect 20977 31524 21033 31580
rect 21033 31524 21037 31580
rect 20973 31520 21037 31524
rect 21053 31580 21117 31584
rect 21053 31524 21057 31580
rect 21057 31524 21113 31580
rect 21113 31524 21117 31580
rect 21053 31520 21117 31524
rect 5917 31036 5981 31040
rect 5917 30980 5921 31036
rect 5921 30980 5977 31036
rect 5977 30980 5981 31036
rect 5917 30976 5981 30980
rect 5997 31036 6061 31040
rect 5997 30980 6001 31036
rect 6001 30980 6057 31036
rect 6057 30980 6061 31036
rect 5997 30976 6061 30980
rect 6077 31036 6141 31040
rect 6077 30980 6081 31036
rect 6081 30980 6137 31036
rect 6137 30980 6141 31036
rect 6077 30976 6141 30980
rect 6157 31036 6221 31040
rect 6157 30980 6161 31036
rect 6161 30980 6217 31036
rect 6217 30980 6221 31036
rect 6157 30976 6221 30980
rect 15848 31036 15912 31040
rect 15848 30980 15852 31036
rect 15852 30980 15908 31036
rect 15908 30980 15912 31036
rect 15848 30976 15912 30980
rect 15928 31036 15992 31040
rect 15928 30980 15932 31036
rect 15932 30980 15988 31036
rect 15988 30980 15992 31036
rect 15928 30976 15992 30980
rect 16008 31036 16072 31040
rect 16008 30980 16012 31036
rect 16012 30980 16068 31036
rect 16068 30980 16072 31036
rect 16008 30976 16072 30980
rect 16088 31036 16152 31040
rect 16088 30980 16092 31036
rect 16092 30980 16148 31036
rect 16148 30980 16152 31036
rect 16088 30976 16152 30980
rect 25778 31036 25842 31040
rect 25778 30980 25782 31036
rect 25782 30980 25838 31036
rect 25838 30980 25842 31036
rect 25778 30976 25842 30980
rect 25858 31036 25922 31040
rect 25858 30980 25862 31036
rect 25862 30980 25918 31036
rect 25918 30980 25922 31036
rect 25858 30976 25922 30980
rect 25938 31036 26002 31040
rect 25938 30980 25942 31036
rect 25942 30980 25998 31036
rect 25998 30980 26002 31036
rect 25938 30976 26002 30980
rect 26018 31036 26082 31040
rect 26018 30980 26022 31036
rect 26022 30980 26078 31036
rect 26078 30980 26082 31036
rect 26018 30976 26082 30980
rect 16988 30908 17052 30972
rect 16620 30832 16684 30836
rect 16620 30776 16634 30832
rect 16634 30776 16684 30832
rect 16620 30772 16684 30776
rect 19196 30636 19260 30700
rect 18644 30500 18708 30564
rect 10882 30492 10946 30496
rect 10882 30436 10886 30492
rect 10886 30436 10942 30492
rect 10942 30436 10946 30492
rect 10882 30432 10946 30436
rect 10962 30492 11026 30496
rect 10962 30436 10966 30492
rect 10966 30436 11022 30492
rect 11022 30436 11026 30492
rect 10962 30432 11026 30436
rect 11042 30492 11106 30496
rect 11042 30436 11046 30492
rect 11046 30436 11102 30492
rect 11102 30436 11106 30492
rect 11042 30432 11106 30436
rect 11122 30492 11186 30496
rect 11122 30436 11126 30492
rect 11126 30436 11182 30492
rect 11182 30436 11186 30492
rect 11122 30432 11186 30436
rect 20813 30492 20877 30496
rect 20813 30436 20817 30492
rect 20817 30436 20873 30492
rect 20873 30436 20877 30492
rect 20813 30432 20877 30436
rect 20893 30492 20957 30496
rect 20893 30436 20897 30492
rect 20897 30436 20953 30492
rect 20953 30436 20957 30492
rect 20893 30432 20957 30436
rect 20973 30492 21037 30496
rect 20973 30436 20977 30492
rect 20977 30436 21033 30492
rect 21033 30436 21037 30492
rect 20973 30432 21037 30436
rect 21053 30492 21117 30496
rect 21053 30436 21057 30492
rect 21057 30436 21113 30492
rect 21113 30436 21117 30492
rect 21053 30432 21117 30436
rect 5917 29948 5981 29952
rect 5917 29892 5921 29948
rect 5921 29892 5977 29948
rect 5977 29892 5981 29948
rect 5917 29888 5981 29892
rect 5997 29948 6061 29952
rect 5997 29892 6001 29948
rect 6001 29892 6057 29948
rect 6057 29892 6061 29948
rect 5997 29888 6061 29892
rect 6077 29948 6141 29952
rect 6077 29892 6081 29948
rect 6081 29892 6137 29948
rect 6137 29892 6141 29948
rect 6077 29888 6141 29892
rect 6157 29948 6221 29952
rect 6157 29892 6161 29948
rect 6161 29892 6217 29948
rect 6217 29892 6221 29948
rect 6157 29888 6221 29892
rect 17540 30152 17604 30156
rect 17540 30096 17590 30152
rect 17590 30096 17604 30152
rect 17540 30092 17604 30096
rect 15848 29948 15912 29952
rect 15848 29892 15852 29948
rect 15852 29892 15908 29948
rect 15908 29892 15912 29948
rect 15848 29888 15912 29892
rect 15928 29948 15992 29952
rect 15928 29892 15932 29948
rect 15932 29892 15988 29948
rect 15988 29892 15992 29948
rect 15928 29888 15992 29892
rect 16008 29948 16072 29952
rect 16008 29892 16012 29948
rect 16012 29892 16068 29948
rect 16068 29892 16072 29948
rect 16008 29888 16072 29892
rect 16088 29948 16152 29952
rect 16088 29892 16092 29948
rect 16092 29892 16148 29948
rect 16148 29892 16152 29948
rect 16088 29888 16152 29892
rect 25778 29948 25842 29952
rect 25778 29892 25782 29948
rect 25782 29892 25838 29948
rect 25838 29892 25842 29948
rect 25778 29888 25842 29892
rect 25858 29948 25922 29952
rect 25858 29892 25862 29948
rect 25862 29892 25918 29948
rect 25918 29892 25922 29948
rect 25858 29888 25922 29892
rect 25938 29948 26002 29952
rect 25938 29892 25942 29948
rect 25942 29892 25998 29948
rect 25998 29892 26002 29948
rect 25938 29888 26002 29892
rect 26018 29948 26082 29952
rect 26018 29892 26022 29948
rect 26022 29892 26078 29948
rect 26078 29892 26082 29948
rect 26018 29888 26082 29892
rect 10882 29404 10946 29408
rect 10882 29348 10886 29404
rect 10886 29348 10942 29404
rect 10942 29348 10946 29404
rect 10882 29344 10946 29348
rect 10962 29404 11026 29408
rect 10962 29348 10966 29404
rect 10966 29348 11022 29404
rect 11022 29348 11026 29404
rect 10962 29344 11026 29348
rect 11042 29404 11106 29408
rect 11042 29348 11046 29404
rect 11046 29348 11102 29404
rect 11102 29348 11106 29404
rect 11042 29344 11106 29348
rect 11122 29404 11186 29408
rect 11122 29348 11126 29404
rect 11126 29348 11182 29404
rect 11182 29348 11186 29404
rect 11122 29344 11186 29348
rect 20813 29404 20877 29408
rect 20813 29348 20817 29404
rect 20817 29348 20873 29404
rect 20873 29348 20877 29404
rect 20813 29344 20877 29348
rect 20893 29404 20957 29408
rect 20893 29348 20897 29404
rect 20897 29348 20953 29404
rect 20953 29348 20957 29404
rect 20893 29344 20957 29348
rect 20973 29404 21037 29408
rect 20973 29348 20977 29404
rect 20977 29348 21033 29404
rect 21033 29348 21037 29404
rect 20973 29344 21037 29348
rect 21053 29404 21117 29408
rect 21053 29348 21057 29404
rect 21057 29348 21113 29404
rect 21113 29348 21117 29404
rect 21053 29344 21117 29348
rect 5917 28860 5981 28864
rect 5917 28804 5921 28860
rect 5921 28804 5977 28860
rect 5977 28804 5981 28860
rect 5917 28800 5981 28804
rect 5997 28860 6061 28864
rect 5997 28804 6001 28860
rect 6001 28804 6057 28860
rect 6057 28804 6061 28860
rect 5997 28800 6061 28804
rect 6077 28860 6141 28864
rect 6077 28804 6081 28860
rect 6081 28804 6137 28860
rect 6137 28804 6141 28860
rect 6077 28800 6141 28804
rect 6157 28860 6221 28864
rect 6157 28804 6161 28860
rect 6161 28804 6217 28860
rect 6217 28804 6221 28860
rect 6157 28800 6221 28804
rect 15848 28860 15912 28864
rect 15848 28804 15852 28860
rect 15852 28804 15908 28860
rect 15908 28804 15912 28860
rect 15848 28800 15912 28804
rect 15928 28860 15992 28864
rect 15928 28804 15932 28860
rect 15932 28804 15988 28860
rect 15988 28804 15992 28860
rect 15928 28800 15992 28804
rect 16008 28860 16072 28864
rect 16008 28804 16012 28860
rect 16012 28804 16068 28860
rect 16068 28804 16072 28860
rect 16008 28800 16072 28804
rect 16088 28860 16152 28864
rect 16088 28804 16092 28860
rect 16092 28804 16148 28860
rect 16148 28804 16152 28860
rect 16088 28800 16152 28804
rect 25778 28860 25842 28864
rect 25778 28804 25782 28860
rect 25782 28804 25838 28860
rect 25838 28804 25842 28860
rect 25778 28800 25842 28804
rect 25858 28860 25922 28864
rect 25858 28804 25862 28860
rect 25862 28804 25918 28860
rect 25918 28804 25922 28860
rect 25858 28800 25922 28804
rect 25938 28860 26002 28864
rect 25938 28804 25942 28860
rect 25942 28804 25998 28860
rect 25998 28804 26002 28860
rect 25938 28800 26002 28804
rect 26018 28860 26082 28864
rect 26018 28804 26022 28860
rect 26022 28804 26078 28860
rect 26078 28804 26082 28860
rect 26018 28800 26082 28804
rect 19012 28596 19076 28660
rect 10882 28316 10946 28320
rect 10882 28260 10886 28316
rect 10886 28260 10942 28316
rect 10942 28260 10946 28316
rect 10882 28256 10946 28260
rect 10962 28316 11026 28320
rect 10962 28260 10966 28316
rect 10966 28260 11022 28316
rect 11022 28260 11026 28316
rect 10962 28256 11026 28260
rect 11042 28316 11106 28320
rect 11042 28260 11046 28316
rect 11046 28260 11102 28316
rect 11102 28260 11106 28316
rect 11042 28256 11106 28260
rect 11122 28316 11186 28320
rect 11122 28260 11126 28316
rect 11126 28260 11182 28316
rect 11182 28260 11186 28316
rect 11122 28256 11186 28260
rect 18644 28052 18708 28116
rect 20813 28316 20877 28320
rect 20813 28260 20817 28316
rect 20817 28260 20873 28316
rect 20873 28260 20877 28316
rect 20813 28256 20877 28260
rect 20893 28316 20957 28320
rect 20893 28260 20897 28316
rect 20897 28260 20953 28316
rect 20953 28260 20957 28316
rect 20893 28256 20957 28260
rect 20973 28316 21037 28320
rect 20973 28260 20977 28316
rect 20977 28260 21033 28316
rect 21033 28260 21037 28316
rect 20973 28256 21037 28260
rect 21053 28316 21117 28320
rect 21053 28260 21057 28316
rect 21057 28260 21113 28316
rect 21113 28260 21117 28316
rect 21053 28256 21117 28260
rect 5917 27772 5981 27776
rect 5917 27716 5921 27772
rect 5921 27716 5977 27772
rect 5977 27716 5981 27772
rect 5917 27712 5981 27716
rect 5997 27772 6061 27776
rect 5997 27716 6001 27772
rect 6001 27716 6057 27772
rect 6057 27716 6061 27772
rect 5997 27712 6061 27716
rect 6077 27772 6141 27776
rect 6077 27716 6081 27772
rect 6081 27716 6137 27772
rect 6137 27716 6141 27772
rect 6077 27712 6141 27716
rect 6157 27772 6221 27776
rect 6157 27716 6161 27772
rect 6161 27716 6217 27772
rect 6217 27716 6221 27772
rect 6157 27712 6221 27716
rect 15848 27772 15912 27776
rect 15848 27716 15852 27772
rect 15852 27716 15908 27772
rect 15908 27716 15912 27772
rect 15848 27712 15912 27716
rect 15928 27772 15992 27776
rect 15928 27716 15932 27772
rect 15932 27716 15988 27772
rect 15988 27716 15992 27772
rect 15928 27712 15992 27716
rect 16008 27772 16072 27776
rect 16008 27716 16012 27772
rect 16012 27716 16068 27772
rect 16068 27716 16072 27772
rect 16008 27712 16072 27716
rect 16088 27772 16152 27776
rect 16088 27716 16092 27772
rect 16092 27716 16148 27772
rect 16148 27716 16152 27772
rect 16088 27712 16152 27716
rect 25778 27772 25842 27776
rect 25778 27716 25782 27772
rect 25782 27716 25838 27772
rect 25838 27716 25842 27772
rect 25778 27712 25842 27716
rect 25858 27772 25922 27776
rect 25858 27716 25862 27772
rect 25862 27716 25918 27772
rect 25918 27716 25922 27772
rect 25858 27712 25922 27716
rect 25938 27772 26002 27776
rect 25938 27716 25942 27772
rect 25942 27716 25998 27772
rect 25998 27716 26002 27772
rect 25938 27712 26002 27716
rect 26018 27772 26082 27776
rect 26018 27716 26022 27772
rect 26022 27716 26078 27772
rect 26078 27716 26082 27772
rect 26018 27712 26082 27716
rect 18644 27644 18708 27708
rect 10882 27228 10946 27232
rect 10882 27172 10886 27228
rect 10886 27172 10942 27228
rect 10942 27172 10946 27228
rect 10882 27168 10946 27172
rect 10962 27228 11026 27232
rect 10962 27172 10966 27228
rect 10966 27172 11022 27228
rect 11022 27172 11026 27228
rect 10962 27168 11026 27172
rect 11042 27228 11106 27232
rect 11042 27172 11046 27228
rect 11046 27172 11102 27228
rect 11102 27172 11106 27228
rect 11042 27168 11106 27172
rect 11122 27228 11186 27232
rect 11122 27172 11126 27228
rect 11126 27172 11182 27228
rect 11182 27172 11186 27228
rect 11122 27168 11186 27172
rect 20813 27228 20877 27232
rect 20813 27172 20817 27228
rect 20817 27172 20873 27228
rect 20873 27172 20877 27228
rect 20813 27168 20877 27172
rect 20893 27228 20957 27232
rect 20893 27172 20897 27228
rect 20897 27172 20953 27228
rect 20953 27172 20957 27228
rect 20893 27168 20957 27172
rect 20973 27228 21037 27232
rect 20973 27172 20977 27228
rect 20977 27172 21033 27228
rect 21033 27172 21037 27228
rect 20973 27168 21037 27172
rect 21053 27228 21117 27232
rect 21053 27172 21057 27228
rect 21057 27172 21113 27228
rect 21113 27172 21117 27228
rect 21053 27168 21117 27172
rect 19012 27100 19076 27164
rect 5917 26684 5981 26688
rect 5917 26628 5921 26684
rect 5921 26628 5977 26684
rect 5977 26628 5981 26684
rect 5917 26624 5981 26628
rect 5997 26684 6061 26688
rect 5997 26628 6001 26684
rect 6001 26628 6057 26684
rect 6057 26628 6061 26684
rect 5997 26624 6061 26628
rect 6077 26684 6141 26688
rect 6077 26628 6081 26684
rect 6081 26628 6137 26684
rect 6137 26628 6141 26684
rect 6077 26624 6141 26628
rect 6157 26684 6221 26688
rect 6157 26628 6161 26684
rect 6161 26628 6217 26684
rect 6217 26628 6221 26684
rect 6157 26624 6221 26628
rect 15848 26684 15912 26688
rect 15848 26628 15852 26684
rect 15852 26628 15908 26684
rect 15908 26628 15912 26684
rect 15848 26624 15912 26628
rect 15928 26684 15992 26688
rect 15928 26628 15932 26684
rect 15932 26628 15988 26684
rect 15988 26628 15992 26684
rect 15928 26624 15992 26628
rect 16008 26684 16072 26688
rect 16008 26628 16012 26684
rect 16012 26628 16068 26684
rect 16068 26628 16072 26684
rect 16008 26624 16072 26628
rect 16088 26684 16152 26688
rect 16088 26628 16092 26684
rect 16092 26628 16148 26684
rect 16148 26628 16152 26684
rect 16088 26624 16152 26628
rect 25778 26684 25842 26688
rect 25778 26628 25782 26684
rect 25782 26628 25838 26684
rect 25838 26628 25842 26684
rect 25778 26624 25842 26628
rect 25858 26684 25922 26688
rect 25858 26628 25862 26684
rect 25862 26628 25918 26684
rect 25918 26628 25922 26684
rect 25858 26624 25922 26628
rect 25938 26684 26002 26688
rect 25938 26628 25942 26684
rect 25942 26628 25998 26684
rect 25998 26628 26002 26684
rect 25938 26624 26002 26628
rect 26018 26684 26082 26688
rect 26018 26628 26022 26684
rect 26022 26628 26078 26684
rect 26078 26628 26082 26684
rect 26018 26624 26082 26628
rect 10882 26140 10946 26144
rect 10882 26084 10886 26140
rect 10886 26084 10942 26140
rect 10942 26084 10946 26140
rect 10882 26080 10946 26084
rect 10962 26140 11026 26144
rect 10962 26084 10966 26140
rect 10966 26084 11022 26140
rect 11022 26084 11026 26140
rect 10962 26080 11026 26084
rect 11042 26140 11106 26144
rect 11042 26084 11046 26140
rect 11046 26084 11102 26140
rect 11102 26084 11106 26140
rect 11042 26080 11106 26084
rect 11122 26140 11186 26144
rect 11122 26084 11126 26140
rect 11126 26084 11182 26140
rect 11182 26084 11186 26140
rect 11122 26080 11186 26084
rect 20813 26140 20877 26144
rect 20813 26084 20817 26140
rect 20817 26084 20873 26140
rect 20873 26084 20877 26140
rect 20813 26080 20877 26084
rect 20893 26140 20957 26144
rect 20893 26084 20897 26140
rect 20897 26084 20953 26140
rect 20953 26084 20957 26140
rect 20893 26080 20957 26084
rect 20973 26140 21037 26144
rect 20973 26084 20977 26140
rect 20977 26084 21033 26140
rect 21033 26084 21037 26140
rect 20973 26080 21037 26084
rect 21053 26140 21117 26144
rect 21053 26084 21057 26140
rect 21057 26084 21113 26140
rect 21113 26084 21117 26140
rect 21053 26080 21117 26084
rect 5917 25596 5981 25600
rect 5917 25540 5921 25596
rect 5921 25540 5977 25596
rect 5977 25540 5981 25596
rect 5917 25536 5981 25540
rect 5997 25596 6061 25600
rect 5997 25540 6001 25596
rect 6001 25540 6057 25596
rect 6057 25540 6061 25596
rect 5997 25536 6061 25540
rect 6077 25596 6141 25600
rect 6077 25540 6081 25596
rect 6081 25540 6137 25596
rect 6137 25540 6141 25596
rect 6077 25536 6141 25540
rect 6157 25596 6221 25600
rect 6157 25540 6161 25596
rect 6161 25540 6217 25596
rect 6217 25540 6221 25596
rect 6157 25536 6221 25540
rect 15848 25596 15912 25600
rect 15848 25540 15852 25596
rect 15852 25540 15908 25596
rect 15908 25540 15912 25596
rect 15848 25536 15912 25540
rect 15928 25596 15992 25600
rect 15928 25540 15932 25596
rect 15932 25540 15988 25596
rect 15988 25540 15992 25596
rect 15928 25536 15992 25540
rect 16008 25596 16072 25600
rect 16008 25540 16012 25596
rect 16012 25540 16068 25596
rect 16068 25540 16072 25596
rect 16008 25536 16072 25540
rect 16088 25596 16152 25600
rect 16088 25540 16092 25596
rect 16092 25540 16148 25596
rect 16148 25540 16152 25596
rect 16088 25536 16152 25540
rect 25778 25596 25842 25600
rect 25778 25540 25782 25596
rect 25782 25540 25838 25596
rect 25838 25540 25842 25596
rect 25778 25536 25842 25540
rect 25858 25596 25922 25600
rect 25858 25540 25862 25596
rect 25862 25540 25918 25596
rect 25918 25540 25922 25596
rect 25858 25536 25922 25540
rect 25938 25596 26002 25600
rect 25938 25540 25942 25596
rect 25942 25540 25998 25596
rect 25998 25540 26002 25596
rect 25938 25536 26002 25540
rect 26018 25596 26082 25600
rect 26018 25540 26022 25596
rect 26022 25540 26078 25596
rect 26078 25540 26082 25596
rect 26018 25536 26082 25540
rect 10882 25052 10946 25056
rect 10882 24996 10886 25052
rect 10886 24996 10942 25052
rect 10942 24996 10946 25052
rect 10882 24992 10946 24996
rect 10962 25052 11026 25056
rect 10962 24996 10966 25052
rect 10966 24996 11022 25052
rect 11022 24996 11026 25052
rect 10962 24992 11026 24996
rect 11042 25052 11106 25056
rect 11042 24996 11046 25052
rect 11046 24996 11102 25052
rect 11102 24996 11106 25052
rect 11042 24992 11106 24996
rect 11122 25052 11186 25056
rect 11122 24996 11126 25052
rect 11126 24996 11182 25052
rect 11182 24996 11186 25052
rect 11122 24992 11186 24996
rect 20813 25052 20877 25056
rect 20813 24996 20817 25052
rect 20817 24996 20873 25052
rect 20873 24996 20877 25052
rect 20813 24992 20877 24996
rect 20893 25052 20957 25056
rect 20893 24996 20897 25052
rect 20897 24996 20953 25052
rect 20953 24996 20957 25052
rect 20893 24992 20957 24996
rect 20973 25052 21037 25056
rect 20973 24996 20977 25052
rect 20977 24996 21033 25052
rect 21033 24996 21037 25052
rect 20973 24992 21037 24996
rect 21053 25052 21117 25056
rect 21053 24996 21057 25052
rect 21057 24996 21113 25052
rect 21113 24996 21117 25052
rect 21053 24992 21117 24996
rect 5917 24508 5981 24512
rect 5917 24452 5921 24508
rect 5921 24452 5977 24508
rect 5977 24452 5981 24508
rect 5917 24448 5981 24452
rect 5997 24508 6061 24512
rect 5997 24452 6001 24508
rect 6001 24452 6057 24508
rect 6057 24452 6061 24508
rect 5997 24448 6061 24452
rect 6077 24508 6141 24512
rect 6077 24452 6081 24508
rect 6081 24452 6137 24508
rect 6137 24452 6141 24508
rect 6077 24448 6141 24452
rect 6157 24508 6221 24512
rect 6157 24452 6161 24508
rect 6161 24452 6217 24508
rect 6217 24452 6221 24508
rect 6157 24448 6221 24452
rect 15848 24508 15912 24512
rect 15848 24452 15852 24508
rect 15852 24452 15908 24508
rect 15908 24452 15912 24508
rect 15848 24448 15912 24452
rect 15928 24508 15992 24512
rect 15928 24452 15932 24508
rect 15932 24452 15988 24508
rect 15988 24452 15992 24508
rect 15928 24448 15992 24452
rect 16008 24508 16072 24512
rect 16008 24452 16012 24508
rect 16012 24452 16068 24508
rect 16068 24452 16072 24508
rect 16008 24448 16072 24452
rect 16088 24508 16152 24512
rect 16088 24452 16092 24508
rect 16092 24452 16148 24508
rect 16148 24452 16152 24508
rect 16088 24448 16152 24452
rect 25778 24508 25842 24512
rect 25778 24452 25782 24508
rect 25782 24452 25838 24508
rect 25838 24452 25842 24508
rect 25778 24448 25842 24452
rect 25858 24508 25922 24512
rect 25858 24452 25862 24508
rect 25862 24452 25918 24508
rect 25918 24452 25922 24508
rect 25858 24448 25922 24452
rect 25938 24508 26002 24512
rect 25938 24452 25942 24508
rect 25942 24452 25998 24508
rect 25998 24452 26002 24508
rect 25938 24448 26002 24452
rect 26018 24508 26082 24512
rect 26018 24452 26022 24508
rect 26022 24452 26078 24508
rect 26078 24452 26082 24508
rect 26018 24448 26082 24452
rect 10882 23964 10946 23968
rect 10882 23908 10886 23964
rect 10886 23908 10942 23964
rect 10942 23908 10946 23964
rect 10882 23904 10946 23908
rect 10962 23964 11026 23968
rect 10962 23908 10966 23964
rect 10966 23908 11022 23964
rect 11022 23908 11026 23964
rect 10962 23904 11026 23908
rect 11042 23964 11106 23968
rect 11042 23908 11046 23964
rect 11046 23908 11102 23964
rect 11102 23908 11106 23964
rect 11042 23904 11106 23908
rect 11122 23964 11186 23968
rect 11122 23908 11126 23964
rect 11126 23908 11182 23964
rect 11182 23908 11186 23964
rect 11122 23904 11186 23908
rect 20813 23964 20877 23968
rect 20813 23908 20817 23964
rect 20817 23908 20873 23964
rect 20873 23908 20877 23964
rect 20813 23904 20877 23908
rect 20893 23964 20957 23968
rect 20893 23908 20897 23964
rect 20897 23908 20953 23964
rect 20953 23908 20957 23964
rect 20893 23904 20957 23908
rect 20973 23964 21037 23968
rect 20973 23908 20977 23964
rect 20977 23908 21033 23964
rect 21033 23908 21037 23964
rect 20973 23904 21037 23908
rect 21053 23964 21117 23968
rect 21053 23908 21057 23964
rect 21057 23908 21113 23964
rect 21113 23908 21117 23964
rect 21053 23904 21117 23908
rect 16988 23564 17052 23628
rect 5917 23420 5981 23424
rect 5917 23364 5921 23420
rect 5921 23364 5977 23420
rect 5977 23364 5981 23420
rect 5917 23360 5981 23364
rect 5997 23420 6061 23424
rect 5997 23364 6001 23420
rect 6001 23364 6057 23420
rect 6057 23364 6061 23420
rect 5997 23360 6061 23364
rect 6077 23420 6141 23424
rect 6077 23364 6081 23420
rect 6081 23364 6137 23420
rect 6137 23364 6141 23420
rect 6077 23360 6141 23364
rect 6157 23420 6221 23424
rect 6157 23364 6161 23420
rect 6161 23364 6217 23420
rect 6217 23364 6221 23420
rect 6157 23360 6221 23364
rect 15848 23420 15912 23424
rect 15848 23364 15852 23420
rect 15852 23364 15908 23420
rect 15908 23364 15912 23420
rect 15848 23360 15912 23364
rect 15928 23420 15992 23424
rect 15928 23364 15932 23420
rect 15932 23364 15988 23420
rect 15988 23364 15992 23420
rect 15928 23360 15992 23364
rect 16008 23420 16072 23424
rect 16008 23364 16012 23420
rect 16012 23364 16068 23420
rect 16068 23364 16072 23420
rect 16008 23360 16072 23364
rect 16088 23420 16152 23424
rect 16088 23364 16092 23420
rect 16092 23364 16148 23420
rect 16148 23364 16152 23420
rect 16088 23360 16152 23364
rect 25778 23420 25842 23424
rect 25778 23364 25782 23420
rect 25782 23364 25838 23420
rect 25838 23364 25842 23420
rect 25778 23360 25842 23364
rect 25858 23420 25922 23424
rect 25858 23364 25862 23420
rect 25862 23364 25918 23420
rect 25918 23364 25922 23420
rect 25858 23360 25922 23364
rect 25938 23420 26002 23424
rect 25938 23364 25942 23420
rect 25942 23364 25998 23420
rect 25998 23364 26002 23420
rect 25938 23360 26002 23364
rect 26018 23420 26082 23424
rect 26018 23364 26022 23420
rect 26022 23364 26078 23420
rect 26078 23364 26082 23420
rect 26018 23360 26082 23364
rect 10882 22876 10946 22880
rect 10882 22820 10886 22876
rect 10886 22820 10942 22876
rect 10942 22820 10946 22876
rect 10882 22816 10946 22820
rect 10962 22876 11026 22880
rect 10962 22820 10966 22876
rect 10966 22820 11022 22876
rect 11022 22820 11026 22876
rect 10962 22816 11026 22820
rect 11042 22876 11106 22880
rect 11042 22820 11046 22876
rect 11046 22820 11102 22876
rect 11102 22820 11106 22876
rect 11042 22816 11106 22820
rect 11122 22876 11186 22880
rect 11122 22820 11126 22876
rect 11126 22820 11182 22876
rect 11182 22820 11186 22876
rect 11122 22816 11186 22820
rect 20813 22876 20877 22880
rect 20813 22820 20817 22876
rect 20817 22820 20873 22876
rect 20873 22820 20877 22876
rect 20813 22816 20877 22820
rect 20893 22876 20957 22880
rect 20893 22820 20897 22876
rect 20897 22820 20953 22876
rect 20953 22820 20957 22876
rect 20893 22816 20957 22820
rect 20973 22876 21037 22880
rect 20973 22820 20977 22876
rect 20977 22820 21033 22876
rect 21033 22820 21037 22876
rect 20973 22816 21037 22820
rect 21053 22876 21117 22880
rect 21053 22820 21057 22876
rect 21057 22820 21113 22876
rect 21113 22820 21117 22876
rect 21053 22816 21117 22820
rect 16988 22340 17052 22404
rect 5917 22332 5981 22336
rect 5917 22276 5921 22332
rect 5921 22276 5977 22332
rect 5977 22276 5981 22332
rect 5917 22272 5981 22276
rect 5997 22332 6061 22336
rect 5997 22276 6001 22332
rect 6001 22276 6057 22332
rect 6057 22276 6061 22332
rect 5997 22272 6061 22276
rect 6077 22332 6141 22336
rect 6077 22276 6081 22332
rect 6081 22276 6137 22332
rect 6137 22276 6141 22332
rect 6077 22272 6141 22276
rect 6157 22332 6221 22336
rect 6157 22276 6161 22332
rect 6161 22276 6217 22332
rect 6217 22276 6221 22332
rect 6157 22272 6221 22276
rect 15848 22332 15912 22336
rect 15848 22276 15852 22332
rect 15852 22276 15908 22332
rect 15908 22276 15912 22332
rect 15848 22272 15912 22276
rect 15928 22332 15992 22336
rect 15928 22276 15932 22332
rect 15932 22276 15988 22332
rect 15988 22276 15992 22332
rect 15928 22272 15992 22276
rect 16008 22332 16072 22336
rect 16008 22276 16012 22332
rect 16012 22276 16068 22332
rect 16068 22276 16072 22332
rect 16008 22272 16072 22276
rect 16088 22332 16152 22336
rect 16088 22276 16092 22332
rect 16092 22276 16148 22332
rect 16148 22276 16152 22332
rect 16088 22272 16152 22276
rect 25778 22332 25842 22336
rect 25778 22276 25782 22332
rect 25782 22276 25838 22332
rect 25838 22276 25842 22332
rect 25778 22272 25842 22276
rect 25858 22332 25922 22336
rect 25858 22276 25862 22332
rect 25862 22276 25918 22332
rect 25918 22276 25922 22332
rect 25858 22272 25922 22276
rect 25938 22332 26002 22336
rect 25938 22276 25942 22332
rect 25942 22276 25998 22332
rect 25998 22276 26002 22332
rect 25938 22272 26002 22276
rect 26018 22332 26082 22336
rect 26018 22276 26022 22332
rect 26022 22276 26078 22332
rect 26078 22276 26082 22332
rect 26018 22272 26082 22276
rect 10882 21788 10946 21792
rect 10882 21732 10886 21788
rect 10886 21732 10942 21788
rect 10942 21732 10946 21788
rect 10882 21728 10946 21732
rect 10962 21788 11026 21792
rect 10962 21732 10966 21788
rect 10966 21732 11022 21788
rect 11022 21732 11026 21788
rect 10962 21728 11026 21732
rect 11042 21788 11106 21792
rect 11042 21732 11046 21788
rect 11046 21732 11102 21788
rect 11102 21732 11106 21788
rect 11042 21728 11106 21732
rect 11122 21788 11186 21792
rect 11122 21732 11126 21788
rect 11126 21732 11182 21788
rect 11182 21732 11186 21788
rect 11122 21728 11186 21732
rect 20813 21788 20877 21792
rect 20813 21732 20817 21788
rect 20817 21732 20873 21788
rect 20873 21732 20877 21788
rect 20813 21728 20877 21732
rect 20893 21788 20957 21792
rect 20893 21732 20897 21788
rect 20897 21732 20953 21788
rect 20953 21732 20957 21788
rect 20893 21728 20957 21732
rect 20973 21788 21037 21792
rect 20973 21732 20977 21788
rect 20977 21732 21033 21788
rect 21033 21732 21037 21788
rect 20973 21728 21037 21732
rect 21053 21788 21117 21792
rect 21053 21732 21057 21788
rect 21057 21732 21113 21788
rect 21113 21732 21117 21788
rect 21053 21728 21117 21732
rect 17356 21524 17420 21588
rect 5917 21244 5981 21248
rect 5917 21188 5921 21244
rect 5921 21188 5977 21244
rect 5977 21188 5981 21244
rect 5917 21184 5981 21188
rect 5997 21244 6061 21248
rect 5997 21188 6001 21244
rect 6001 21188 6057 21244
rect 6057 21188 6061 21244
rect 5997 21184 6061 21188
rect 6077 21244 6141 21248
rect 6077 21188 6081 21244
rect 6081 21188 6137 21244
rect 6137 21188 6141 21244
rect 6077 21184 6141 21188
rect 6157 21244 6221 21248
rect 6157 21188 6161 21244
rect 6161 21188 6217 21244
rect 6217 21188 6221 21244
rect 6157 21184 6221 21188
rect 15848 21244 15912 21248
rect 15848 21188 15852 21244
rect 15852 21188 15908 21244
rect 15908 21188 15912 21244
rect 15848 21184 15912 21188
rect 15928 21244 15992 21248
rect 15928 21188 15932 21244
rect 15932 21188 15988 21244
rect 15988 21188 15992 21244
rect 15928 21184 15992 21188
rect 16008 21244 16072 21248
rect 16008 21188 16012 21244
rect 16012 21188 16068 21244
rect 16068 21188 16072 21244
rect 16008 21184 16072 21188
rect 16088 21244 16152 21248
rect 16088 21188 16092 21244
rect 16092 21188 16148 21244
rect 16148 21188 16152 21244
rect 16088 21184 16152 21188
rect 25778 21244 25842 21248
rect 25778 21188 25782 21244
rect 25782 21188 25838 21244
rect 25838 21188 25842 21244
rect 25778 21184 25842 21188
rect 25858 21244 25922 21248
rect 25858 21188 25862 21244
rect 25862 21188 25918 21244
rect 25918 21188 25922 21244
rect 25858 21184 25922 21188
rect 25938 21244 26002 21248
rect 25938 21188 25942 21244
rect 25942 21188 25998 21244
rect 25998 21188 26002 21244
rect 25938 21184 26002 21188
rect 26018 21244 26082 21248
rect 26018 21188 26022 21244
rect 26022 21188 26078 21244
rect 26078 21188 26082 21244
rect 26018 21184 26082 21188
rect 10882 20700 10946 20704
rect 10882 20644 10886 20700
rect 10886 20644 10942 20700
rect 10942 20644 10946 20700
rect 10882 20640 10946 20644
rect 10962 20700 11026 20704
rect 10962 20644 10966 20700
rect 10966 20644 11022 20700
rect 11022 20644 11026 20700
rect 10962 20640 11026 20644
rect 11042 20700 11106 20704
rect 11042 20644 11046 20700
rect 11046 20644 11102 20700
rect 11102 20644 11106 20700
rect 11042 20640 11106 20644
rect 11122 20700 11186 20704
rect 11122 20644 11126 20700
rect 11126 20644 11182 20700
rect 11182 20644 11186 20700
rect 11122 20640 11186 20644
rect 20813 20700 20877 20704
rect 20813 20644 20817 20700
rect 20817 20644 20873 20700
rect 20873 20644 20877 20700
rect 20813 20640 20877 20644
rect 20893 20700 20957 20704
rect 20893 20644 20897 20700
rect 20897 20644 20953 20700
rect 20953 20644 20957 20700
rect 20893 20640 20957 20644
rect 20973 20700 21037 20704
rect 20973 20644 20977 20700
rect 20977 20644 21033 20700
rect 21033 20644 21037 20700
rect 20973 20640 21037 20644
rect 21053 20700 21117 20704
rect 21053 20644 21057 20700
rect 21057 20644 21113 20700
rect 21113 20644 21117 20700
rect 21053 20640 21117 20644
rect 19196 20572 19260 20636
rect 5917 20156 5981 20160
rect 5917 20100 5921 20156
rect 5921 20100 5977 20156
rect 5977 20100 5981 20156
rect 5917 20096 5981 20100
rect 5997 20156 6061 20160
rect 5997 20100 6001 20156
rect 6001 20100 6057 20156
rect 6057 20100 6061 20156
rect 5997 20096 6061 20100
rect 6077 20156 6141 20160
rect 6077 20100 6081 20156
rect 6081 20100 6137 20156
rect 6137 20100 6141 20156
rect 6077 20096 6141 20100
rect 6157 20156 6221 20160
rect 6157 20100 6161 20156
rect 6161 20100 6217 20156
rect 6217 20100 6221 20156
rect 6157 20096 6221 20100
rect 15848 20156 15912 20160
rect 15848 20100 15852 20156
rect 15852 20100 15908 20156
rect 15908 20100 15912 20156
rect 15848 20096 15912 20100
rect 15928 20156 15992 20160
rect 15928 20100 15932 20156
rect 15932 20100 15988 20156
rect 15988 20100 15992 20156
rect 15928 20096 15992 20100
rect 16008 20156 16072 20160
rect 16008 20100 16012 20156
rect 16012 20100 16068 20156
rect 16068 20100 16072 20156
rect 16008 20096 16072 20100
rect 16088 20156 16152 20160
rect 16088 20100 16092 20156
rect 16092 20100 16148 20156
rect 16148 20100 16152 20156
rect 16088 20096 16152 20100
rect 25778 20156 25842 20160
rect 25778 20100 25782 20156
rect 25782 20100 25838 20156
rect 25838 20100 25842 20156
rect 25778 20096 25842 20100
rect 25858 20156 25922 20160
rect 25858 20100 25862 20156
rect 25862 20100 25918 20156
rect 25918 20100 25922 20156
rect 25858 20096 25922 20100
rect 25938 20156 26002 20160
rect 25938 20100 25942 20156
rect 25942 20100 25998 20156
rect 25998 20100 26002 20156
rect 25938 20096 26002 20100
rect 26018 20156 26082 20160
rect 26018 20100 26022 20156
rect 26022 20100 26078 20156
rect 26078 20100 26082 20156
rect 26018 20096 26082 20100
rect 10882 19612 10946 19616
rect 10882 19556 10886 19612
rect 10886 19556 10942 19612
rect 10942 19556 10946 19612
rect 10882 19552 10946 19556
rect 10962 19612 11026 19616
rect 10962 19556 10966 19612
rect 10966 19556 11022 19612
rect 11022 19556 11026 19612
rect 10962 19552 11026 19556
rect 11042 19612 11106 19616
rect 11042 19556 11046 19612
rect 11046 19556 11102 19612
rect 11102 19556 11106 19612
rect 11042 19552 11106 19556
rect 11122 19612 11186 19616
rect 11122 19556 11126 19612
rect 11126 19556 11182 19612
rect 11182 19556 11186 19612
rect 11122 19552 11186 19556
rect 20813 19612 20877 19616
rect 20813 19556 20817 19612
rect 20817 19556 20873 19612
rect 20873 19556 20877 19612
rect 20813 19552 20877 19556
rect 20893 19612 20957 19616
rect 20893 19556 20897 19612
rect 20897 19556 20953 19612
rect 20953 19556 20957 19612
rect 20893 19552 20957 19556
rect 20973 19612 21037 19616
rect 20973 19556 20977 19612
rect 20977 19556 21033 19612
rect 21033 19556 21037 19612
rect 20973 19552 21037 19556
rect 21053 19612 21117 19616
rect 21053 19556 21057 19612
rect 21057 19556 21113 19612
rect 21113 19556 21117 19612
rect 21053 19552 21117 19556
rect 5917 19068 5981 19072
rect 5917 19012 5921 19068
rect 5921 19012 5977 19068
rect 5977 19012 5981 19068
rect 5917 19008 5981 19012
rect 5997 19068 6061 19072
rect 5997 19012 6001 19068
rect 6001 19012 6057 19068
rect 6057 19012 6061 19068
rect 5997 19008 6061 19012
rect 6077 19068 6141 19072
rect 6077 19012 6081 19068
rect 6081 19012 6137 19068
rect 6137 19012 6141 19068
rect 6077 19008 6141 19012
rect 6157 19068 6221 19072
rect 6157 19012 6161 19068
rect 6161 19012 6217 19068
rect 6217 19012 6221 19068
rect 6157 19008 6221 19012
rect 15848 19068 15912 19072
rect 15848 19012 15852 19068
rect 15852 19012 15908 19068
rect 15908 19012 15912 19068
rect 15848 19008 15912 19012
rect 15928 19068 15992 19072
rect 15928 19012 15932 19068
rect 15932 19012 15988 19068
rect 15988 19012 15992 19068
rect 15928 19008 15992 19012
rect 16008 19068 16072 19072
rect 16008 19012 16012 19068
rect 16012 19012 16068 19068
rect 16068 19012 16072 19068
rect 16008 19008 16072 19012
rect 16088 19068 16152 19072
rect 16088 19012 16092 19068
rect 16092 19012 16148 19068
rect 16148 19012 16152 19068
rect 16088 19008 16152 19012
rect 25778 19068 25842 19072
rect 25778 19012 25782 19068
rect 25782 19012 25838 19068
rect 25838 19012 25842 19068
rect 25778 19008 25842 19012
rect 25858 19068 25922 19072
rect 25858 19012 25862 19068
rect 25862 19012 25918 19068
rect 25918 19012 25922 19068
rect 25858 19008 25922 19012
rect 25938 19068 26002 19072
rect 25938 19012 25942 19068
rect 25942 19012 25998 19068
rect 25998 19012 26002 19068
rect 25938 19008 26002 19012
rect 26018 19068 26082 19072
rect 26018 19012 26022 19068
rect 26022 19012 26078 19068
rect 26078 19012 26082 19068
rect 26018 19008 26082 19012
rect 10882 18524 10946 18528
rect 10882 18468 10886 18524
rect 10886 18468 10942 18524
rect 10942 18468 10946 18524
rect 10882 18464 10946 18468
rect 10962 18524 11026 18528
rect 10962 18468 10966 18524
rect 10966 18468 11022 18524
rect 11022 18468 11026 18524
rect 10962 18464 11026 18468
rect 11042 18524 11106 18528
rect 11042 18468 11046 18524
rect 11046 18468 11102 18524
rect 11102 18468 11106 18524
rect 11042 18464 11106 18468
rect 11122 18524 11186 18528
rect 11122 18468 11126 18524
rect 11126 18468 11182 18524
rect 11182 18468 11186 18524
rect 11122 18464 11186 18468
rect 20813 18524 20877 18528
rect 20813 18468 20817 18524
rect 20817 18468 20873 18524
rect 20873 18468 20877 18524
rect 20813 18464 20877 18468
rect 20893 18524 20957 18528
rect 20893 18468 20897 18524
rect 20897 18468 20953 18524
rect 20953 18468 20957 18524
rect 20893 18464 20957 18468
rect 20973 18524 21037 18528
rect 20973 18468 20977 18524
rect 20977 18468 21033 18524
rect 21033 18468 21037 18524
rect 20973 18464 21037 18468
rect 21053 18524 21117 18528
rect 21053 18468 21057 18524
rect 21057 18468 21113 18524
rect 21113 18468 21117 18524
rect 21053 18464 21117 18468
rect 5917 17980 5981 17984
rect 5917 17924 5921 17980
rect 5921 17924 5977 17980
rect 5977 17924 5981 17980
rect 5917 17920 5981 17924
rect 5997 17980 6061 17984
rect 5997 17924 6001 17980
rect 6001 17924 6057 17980
rect 6057 17924 6061 17980
rect 5997 17920 6061 17924
rect 6077 17980 6141 17984
rect 6077 17924 6081 17980
rect 6081 17924 6137 17980
rect 6137 17924 6141 17980
rect 6077 17920 6141 17924
rect 6157 17980 6221 17984
rect 6157 17924 6161 17980
rect 6161 17924 6217 17980
rect 6217 17924 6221 17980
rect 6157 17920 6221 17924
rect 15848 17980 15912 17984
rect 15848 17924 15852 17980
rect 15852 17924 15908 17980
rect 15908 17924 15912 17980
rect 15848 17920 15912 17924
rect 15928 17980 15992 17984
rect 15928 17924 15932 17980
rect 15932 17924 15988 17980
rect 15988 17924 15992 17980
rect 15928 17920 15992 17924
rect 16008 17980 16072 17984
rect 16008 17924 16012 17980
rect 16012 17924 16068 17980
rect 16068 17924 16072 17980
rect 16008 17920 16072 17924
rect 16088 17980 16152 17984
rect 16088 17924 16092 17980
rect 16092 17924 16148 17980
rect 16148 17924 16152 17980
rect 16088 17920 16152 17924
rect 25778 17980 25842 17984
rect 25778 17924 25782 17980
rect 25782 17924 25838 17980
rect 25838 17924 25842 17980
rect 25778 17920 25842 17924
rect 25858 17980 25922 17984
rect 25858 17924 25862 17980
rect 25862 17924 25918 17980
rect 25918 17924 25922 17980
rect 25858 17920 25922 17924
rect 25938 17980 26002 17984
rect 25938 17924 25942 17980
rect 25942 17924 25998 17980
rect 25998 17924 26002 17980
rect 25938 17920 26002 17924
rect 26018 17980 26082 17984
rect 26018 17924 26022 17980
rect 26022 17924 26078 17980
rect 26078 17924 26082 17980
rect 26018 17920 26082 17924
rect 10882 17436 10946 17440
rect 10882 17380 10886 17436
rect 10886 17380 10942 17436
rect 10942 17380 10946 17436
rect 10882 17376 10946 17380
rect 10962 17436 11026 17440
rect 10962 17380 10966 17436
rect 10966 17380 11022 17436
rect 11022 17380 11026 17436
rect 10962 17376 11026 17380
rect 11042 17436 11106 17440
rect 11042 17380 11046 17436
rect 11046 17380 11102 17436
rect 11102 17380 11106 17436
rect 11042 17376 11106 17380
rect 11122 17436 11186 17440
rect 11122 17380 11126 17436
rect 11126 17380 11182 17436
rect 11182 17380 11186 17436
rect 11122 17376 11186 17380
rect 20813 17436 20877 17440
rect 20813 17380 20817 17436
rect 20817 17380 20873 17436
rect 20873 17380 20877 17436
rect 20813 17376 20877 17380
rect 20893 17436 20957 17440
rect 20893 17380 20897 17436
rect 20897 17380 20953 17436
rect 20953 17380 20957 17436
rect 20893 17376 20957 17380
rect 20973 17436 21037 17440
rect 20973 17380 20977 17436
rect 20977 17380 21033 17436
rect 21033 17380 21037 17436
rect 20973 17376 21037 17380
rect 21053 17436 21117 17440
rect 21053 17380 21057 17436
rect 21057 17380 21113 17436
rect 21113 17380 21117 17436
rect 21053 17376 21117 17380
rect 5917 16892 5981 16896
rect 5917 16836 5921 16892
rect 5921 16836 5977 16892
rect 5977 16836 5981 16892
rect 5917 16832 5981 16836
rect 5997 16892 6061 16896
rect 5997 16836 6001 16892
rect 6001 16836 6057 16892
rect 6057 16836 6061 16892
rect 5997 16832 6061 16836
rect 6077 16892 6141 16896
rect 6077 16836 6081 16892
rect 6081 16836 6137 16892
rect 6137 16836 6141 16892
rect 6077 16832 6141 16836
rect 6157 16892 6221 16896
rect 6157 16836 6161 16892
rect 6161 16836 6217 16892
rect 6217 16836 6221 16892
rect 6157 16832 6221 16836
rect 15848 16892 15912 16896
rect 15848 16836 15852 16892
rect 15852 16836 15908 16892
rect 15908 16836 15912 16892
rect 15848 16832 15912 16836
rect 15928 16892 15992 16896
rect 15928 16836 15932 16892
rect 15932 16836 15988 16892
rect 15988 16836 15992 16892
rect 15928 16832 15992 16836
rect 16008 16892 16072 16896
rect 16008 16836 16012 16892
rect 16012 16836 16068 16892
rect 16068 16836 16072 16892
rect 16008 16832 16072 16836
rect 16088 16892 16152 16896
rect 16088 16836 16092 16892
rect 16092 16836 16148 16892
rect 16148 16836 16152 16892
rect 16088 16832 16152 16836
rect 25778 16892 25842 16896
rect 25778 16836 25782 16892
rect 25782 16836 25838 16892
rect 25838 16836 25842 16892
rect 25778 16832 25842 16836
rect 25858 16892 25922 16896
rect 25858 16836 25862 16892
rect 25862 16836 25918 16892
rect 25918 16836 25922 16892
rect 25858 16832 25922 16836
rect 25938 16892 26002 16896
rect 25938 16836 25942 16892
rect 25942 16836 25998 16892
rect 25998 16836 26002 16892
rect 25938 16832 26002 16836
rect 26018 16892 26082 16896
rect 26018 16836 26022 16892
rect 26022 16836 26078 16892
rect 26078 16836 26082 16892
rect 26018 16832 26082 16836
rect 10882 16348 10946 16352
rect 10882 16292 10886 16348
rect 10886 16292 10942 16348
rect 10942 16292 10946 16348
rect 10882 16288 10946 16292
rect 10962 16348 11026 16352
rect 10962 16292 10966 16348
rect 10966 16292 11022 16348
rect 11022 16292 11026 16348
rect 10962 16288 11026 16292
rect 11042 16348 11106 16352
rect 11042 16292 11046 16348
rect 11046 16292 11102 16348
rect 11102 16292 11106 16348
rect 11042 16288 11106 16292
rect 11122 16348 11186 16352
rect 11122 16292 11126 16348
rect 11126 16292 11182 16348
rect 11182 16292 11186 16348
rect 11122 16288 11186 16292
rect 20813 16348 20877 16352
rect 20813 16292 20817 16348
rect 20817 16292 20873 16348
rect 20873 16292 20877 16348
rect 20813 16288 20877 16292
rect 20893 16348 20957 16352
rect 20893 16292 20897 16348
rect 20897 16292 20953 16348
rect 20953 16292 20957 16348
rect 20893 16288 20957 16292
rect 20973 16348 21037 16352
rect 20973 16292 20977 16348
rect 20977 16292 21033 16348
rect 21033 16292 21037 16348
rect 20973 16288 21037 16292
rect 21053 16348 21117 16352
rect 21053 16292 21057 16348
rect 21057 16292 21113 16348
rect 21113 16292 21117 16348
rect 21053 16288 21117 16292
rect 5917 15804 5981 15808
rect 5917 15748 5921 15804
rect 5921 15748 5977 15804
rect 5977 15748 5981 15804
rect 5917 15744 5981 15748
rect 5997 15804 6061 15808
rect 5997 15748 6001 15804
rect 6001 15748 6057 15804
rect 6057 15748 6061 15804
rect 5997 15744 6061 15748
rect 6077 15804 6141 15808
rect 6077 15748 6081 15804
rect 6081 15748 6137 15804
rect 6137 15748 6141 15804
rect 6077 15744 6141 15748
rect 6157 15804 6221 15808
rect 6157 15748 6161 15804
rect 6161 15748 6217 15804
rect 6217 15748 6221 15804
rect 6157 15744 6221 15748
rect 15848 15804 15912 15808
rect 15848 15748 15852 15804
rect 15852 15748 15908 15804
rect 15908 15748 15912 15804
rect 15848 15744 15912 15748
rect 15928 15804 15992 15808
rect 15928 15748 15932 15804
rect 15932 15748 15988 15804
rect 15988 15748 15992 15804
rect 15928 15744 15992 15748
rect 16008 15804 16072 15808
rect 16008 15748 16012 15804
rect 16012 15748 16068 15804
rect 16068 15748 16072 15804
rect 16008 15744 16072 15748
rect 16088 15804 16152 15808
rect 16088 15748 16092 15804
rect 16092 15748 16148 15804
rect 16148 15748 16152 15804
rect 16088 15744 16152 15748
rect 25778 15804 25842 15808
rect 25778 15748 25782 15804
rect 25782 15748 25838 15804
rect 25838 15748 25842 15804
rect 25778 15744 25842 15748
rect 25858 15804 25922 15808
rect 25858 15748 25862 15804
rect 25862 15748 25918 15804
rect 25918 15748 25922 15804
rect 25858 15744 25922 15748
rect 25938 15804 26002 15808
rect 25938 15748 25942 15804
rect 25942 15748 25998 15804
rect 25998 15748 26002 15804
rect 25938 15744 26002 15748
rect 26018 15804 26082 15808
rect 26018 15748 26022 15804
rect 26022 15748 26078 15804
rect 26078 15748 26082 15804
rect 26018 15744 26082 15748
rect 10882 15260 10946 15264
rect 10882 15204 10886 15260
rect 10886 15204 10942 15260
rect 10942 15204 10946 15260
rect 10882 15200 10946 15204
rect 10962 15260 11026 15264
rect 10962 15204 10966 15260
rect 10966 15204 11022 15260
rect 11022 15204 11026 15260
rect 10962 15200 11026 15204
rect 11042 15260 11106 15264
rect 11042 15204 11046 15260
rect 11046 15204 11102 15260
rect 11102 15204 11106 15260
rect 11042 15200 11106 15204
rect 11122 15260 11186 15264
rect 11122 15204 11126 15260
rect 11126 15204 11182 15260
rect 11182 15204 11186 15260
rect 11122 15200 11186 15204
rect 20813 15260 20877 15264
rect 20813 15204 20817 15260
rect 20817 15204 20873 15260
rect 20873 15204 20877 15260
rect 20813 15200 20877 15204
rect 20893 15260 20957 15264
rect 20893 15204 20897 15260
rect 20897 15204 20953 15260
rect 20953 15204 20957 15260
rect 20893 15200 20957 15204
rect 20973 15260 21037 15264
rect 20973 15204 20977 15260
rect 20977 15204 21033 15260
rect 21033 15204 21037 15260
rect 20973 15200 21037 15204
rect 21053 15260 21117 15264
rect 21053 15204 21057 15260
rect 21057 15204 21113 15260
rect 21113 15204 21117 15260
rect 21053 15200 21117 15204
rect 5917 14716 5981 14720
rect 5917 14660 5921 14716
rect 5921 14660 5977 14716
rect 5977 14660 5981 14716
rect 5917 14656 5981 14660
rect 5997 14716 6061 14720
rect 5997 14660 6001 14716
rect 6001 14660 6057 14716
rect 6057 14660 6061 14716
rect 5997 14656 6061 14660
rect 6077 14716 6141 14720
rect 6077 14660 6081 14716
rect 6081 14660 6137 14716
rect 6137 14660 6141 14716
rect 6077 14656 6141 14660
rect 6157 14716 6221 14720
rect 6157 14660 6161 14716
rect 6161 14660 6217 14716
rect 6217 14660 6221 14716
rect 6157 14656 6221 14660
rect 15848 14716 15912 14720
rect 15848 14660 15852 14716
rect 15852 14660 15908 14716
rect 15908 14660 15912 14716
rect 15848 14656 15912 14660
rect 15928 14716 15992 14720
rect 15928 14660 15932 14716
rect 15932 14660 15988 14716
rect 15988 14660 15992 14716
rect 15928 14656 15992 14660
rect 16008 14716 16072 14720
rect 16008 14660 16012 14716
rect 16012 14660 16068 14716
rect 16068 14660 16072 14716
rect 16008 14656 16072 14660
rect 16088 14716 16152 14720
rect 16088 14660 16092 14716
rect 16092 14660 16148 14716
rect 16148 14660 16152 14716
rect 16088 14656 16152 14660
rect 25778 14716 25842 14720
rect 25778 14660 25782 14716
rect 25782 14660 25838 14716
rect 25838 14660 25842 14716
rect 25778 14656 25842 14660
rect 25858 14716 25922 14720
rect 25858 14660 25862 14716
rect 25862 14660 25918 14716
rect 25918 14660 25922 14716
rect 25858 14656 25922 14660
rect 25938 14716 26002 14720
rect 25938 14660 25942 14716
rect 25942 14660 25998 14716
rect 25998 14660 26002 14716
rect 25938 14656 26002 14660
rect 26018 14716 26082 14720
rect 26018 14660 26022 14716
rect 26022 14660 26078 14716
rect 26078 14660 26082 14716
rect 26018 14656 26082 14660
rect 21404 14316 21468 14380
rect 10882 14172 10946 14176
rect 10882 14116 10886 14172
rect 10886 14116 10942 14172
rect 10942 14116 10946 14172
rect 10882 14112 10946 14116
rect 10962 14172 11026 14176
rect 10962 14116 10966 14172
rect 10966 14116 11022 14172
rect 11022 14116 11026 14172
rect 10962 14112 11026 14116
rect 11042 14172 11106 14176
rect 11042 14116 11046 14172
rect 11046 14116 11102 14172
rect 11102 14116 11106 14172
rect 11042 14112 11106 14116
rect 11122 14172 11186 14176
rect 11122 14116 11126 14172
rect 11126 14116 11182 14172
rect 11182 14116 11186 14172
rect 11122 14112 11186 14116
rect 20813 14172 20877 14176
rect 20813 14116 20817 14172
rect 20817 14116 20873 14172
rect 20873 14116 20877 14172
rect 20813 14112 20877 14116
rect 20893 14172 20957 14176
rect 20893 14116 20897 14172
rect 20897 14116 20953 14172
rect 20953 14116 20957 14172
rect 20893 14112 20957 14116
rect 20973 14172 21037 14176
rect 20973 14116 20977 14172
rect 20977 14116 21033 14172
rect 21033 14116 21037 14172
rect 20973 14112 21037 14116
rect 21053 14172 21117 14176
rect 21053 14116 21057 14172
rect 21057 14116 21113 14172
rect 21113 14116 21117 14172
rect 21053 14112 21117 14116
rect 5917 13628 5981 13632
rect 5917 13572 5921 13628
rect 5921 13572 5977 13628
rect 5977 13572 5981 13628
rect 5917 13568 5981 13572
rect 5997 13628 6061 13632
rect 5997 13572 6001 13628
rect 6001 13572 6057 13628
rect 6057 13572 6061 13628
rect 5997 13568 6061 13572
rect 6077 13628 6141 13632
rect 6077 13572 6081 13628
rect 6081 13572 6137 13628
rect 6137 13572 6141 13628
rect 6077 13568 6141 13572
rect 6157 13628 6221 13632
rect 6157 13572 6161 13628
rect 6161 13572 6217 13628
rect 6217 13572 6221 13628
rect 6157 13568 6221 13572
rect 15848 13628 15912 13632
rect 15848 13572 15852 13628
rect 15852 13572 15908 13628
rect 15908 13572 15912 13628
rect 15848 13568 15912 13572
rect 15928 13628 15992 13632
rect 15928 13572 15932 13628
rect 15932 13572 15988 13628
rect 15988 13572 15992 13628
rect 15928 13568 15992 13572
rect 16008 13628 16072 13632
rect 16008 13572 16012 13628
rect 16012 13572 16068 13628
rect 16068 13572 16072 13628
rect 16008 13568 16072 13572
rect 16088 13628 16152 13632
rect 16088 13572 16092 13628
rect 16092 13572 16148 13628
rect 16148 13572 16152 13628
rect 16088 13568 16152 13572
rect 25778 13628 25842 13632
rect 25778 13572 25782 13628
rect 25782 13572 25838 13628
rect 25838 13572 25842 13628
rect 25778 13568 25842 13572
rect 25858 13628 25922 13632
rect 25858 13572 25862 13628
rect 25862 13572 25918 13628
rect 25918 13572 25922 13628
rect 25858 13568 25922 13572
rect 25938 13628 26002 13632
rect 25938 13572 25942 13628
rect 25942 13572 25998 13628
rect 25998 13572 26002 13628
rect 25938 13568 26002 13572
rect 26018 13628 26082 13632
rect 26018 13572 26022 13628
rect 26022 13572 26078 13628
rect 26078 13572 26082 13628
rect 26018 13568 26082 13572
rect 10882 13084 10946 13088
rect 10882 13028 10886 13084
rect 10886 13028 10942 13084
rect 10942 13028 10946 13084
rect 10882 13024 10946 13028
rect 10962 13084 11026 13088
rect 10962 13028 10966 13084
rect 10966 13028 11022 13084
rect 11022 13028 11026 13084
rect 10962 13024 11026 13028
rect 11042 13084 11106 13088
rect 11042 13028 11046 13084
rect 11046 13028 11102 13084
rect 11102 13028 11106 13084
rect 11042 13024 11106 13028
rect 11122 13084 11186 13088
rect 11122 13028 11126 13084
rect 11126 13028 11182 13084
rect 11182 13028 11186 13084
rect 11122 13024 11186 13028
rect 20813 13084 20877 13088
rect 20813 13028 20817 13084
rect 20817 13028 20873 13084
rect 20873 13028 20877 13084
rect 20813 13024 20877 13028
rect 20893 13084 20957 13088
rect 20893 13028 20897 13084
rect 20897 13028 20953 13084
rect 20953 13028 20957 13084
rect 20893 13024 20957 13028
rect 20973 13084 21037 13088
rect 20973 13028 20977 13084
rect 20977 13028 21033 13084
rect 21033 13028 21037 13084
rect 20973 13024 21037 13028
rect 21053 13084 21117 13088
rect 21053 13028 21057 13084
rect 21057 13028 21113 13084
rect 21113 13028 21117 13084
rect 21053 13024 21117 13028
rect 20484 12548 20548 12612
rect 5917 12540 5981 12544
rect 5917 12484 5921 12540
rect 5921 12484 5977 12540
rect 5977 12484 5981 12540
rect 5917 12480 5981 12484
rect 5997 12540 6061 12544
rect 5997 12484 6001 12540
rect 6001 12484 6057 12540
rect 6057 12484 6061 12540
rect 5997 12480 6061 12484
rect 6077 12540 6141 12544
rect 6077 12484 6081 12540
rect 6081 12484 6137 12540
rect 6137 12484 6141 12540
rect 6077 12480 6141 12484
rect 6157 12540 6221 12544
rect 6157 12484 6161 12540
rect 6161 12484 6217 12540
rect 6217 12484 6221 12540
rect 6157 12480 6221 12484
rect 15848 12540 15912 12544
rect 15848 12484 15852 12540
rect 15852 12484 15908 12540
rect 15908 12484 15912 12540
rect 15848 12480 15912 12484
rect 15928 12540 15992 12544
rect 15928 12484 15932 12540
rect 15932 12484 15988 12540
rect 15988 12484 15992 12540
rect 15928 12480 15992 12484
rect 16008 12540 16072 12544
rect 16008 12484 16012 12540
rect 16012 12484 16068 12540
rect 16068 12484 16072 12540
rect 16008 12480 16072 12484
rect 16088 12540 16152 12544
rect 16088 12484 16092 12540
rect 16092 12484 16148 12540
rect 16148 12484 16152 12540
rect 16088 12480 16152 12484
rect 25778 12540 25842 12544
rect 25778 12484 25782 12540
rect 25782 12484 25838 12540
rect 25838 12484 25842 12540
rect 25778 12480 25842 12484
rect 25858 12540 25922 12544
rect 25858 12484 25862 12540
rect 25862 12484 25918 12540
rect 25918 12484 25922 12540
rect 25858 12480 25922 12484
rect 25938 12540 26002 12544
rect 25938 12484 25942 12540
rect 25942 12484 25998 12540
rect 25998 12484 26002 12540
rect 25938 12480 26002 12484
rect 26018 12540 26082 12544
rect 26018 12484 26022 12540
rect 26022 12484 26078 12540
rect 26078 12484 26082 12540
rect 26018 12480 26082 12484
rect 10882 11996 10946 12000
rect 10882 11940 10886 11996
rect 10886 11940 10942 11996
rect 10942 11940 10946 11996
rect 10882 11936 10946 11940
rect 10962 11996 11026 12000
rect 10962 11940 10966 11996
rect 10966 11940 11022 11996
rect 11022 11940 11026 11996
rect 10962 11936 11026 11940
rect 11042 11996 11106 12000
rect 11042 11940 11046 11996
rect 11046 11940 11102 11996
rect 11102 11940 11106 11996
rect 11042 11936 11106 11940
rect 11122 11996 11186 12000
rect 11122 11940 11126 11996
rect 11126 11940 11182 11996
rect 11182 11940 11186 11996
rect 11122 11936 11186 11940
rect 20813 11996 20877 12000
rect 20813 11940 20817 11996
rect 20817 11940 20873 11996
rect 20873 11940 20877 11996
rect 20813 11936 20877 11940
rect 20893 11996 20957 12000
rect 20893 11940 20897 11996
rect 20897 11940 20953 11996
rect 20953 11940 20957 11996
rect 20893 11936 20957 11940
rect 20973 11996 21037 12000
rect 20973 11940 20977 11996
rect 20977 11940 21033 11996
rect 21033 11940 21037 11996
rect 20973 11936 21037 11940
rect 21053 11996 21117 12000
rect 21053 11940 21057 11996
rect 21057 11940 21113 11996
rect 21113 11940 21117 11996
rect 21053 11936 21117 11940
rect 5917 11452 5981 11456
rect 5917 11396 5921 11452
rect 5921 11396 5977 11452
rect 5977 11396 5981 11452
rect 5917 11392 5981 11396
rect 5997 11452 6061 11456
rect 5997 11396 6001 11452
rect 6001 11396 6057 11452
rect 6057 11396 6061 11452
rect 5997 11392 6061 11396
rect 6077 11452 6141 11456
rect 6077 11396 6081 11452
rect 6081 11396 6137 11452
rect 6137 11396 6141 11452
rect 6077 11392 6141 11396
rect 6157 11452 6221 11456
rect 6157 11396 6161 11452
rect 6161 11396 6217 11452
rect 6217 11396 6221 11452
rect 6157 11392 6221 11396
rect 15848 11452 15912 11456
rect 15848 11396 15852 11452
rect 15852 11396 15908 11452
rect 15908 11396 15912 11452
rect 15848 11392 15912 11396
rect 15928 11452 15992 11456
rect 15928 11396 15932 11452
rect 15932 11396 15988 11452
rect 15988 11396 15992 11452
rect 15928 11392 15992 11396
rect 16008 11452 16072 11456
rect 16008 11396 16012 11452
rect 16012 11396 16068 11452
rect 16068 11396 16072 11452
rect 16008 11392 16072 11396
rect 16088 11452 16152 11456
rect 16088 11396 16092 11452
rect 16092 11396 16148 11452
rect 16148 11396 16152 11452
rect 16088 11392 16152 11396
rect 25778 11452 25842 11456
rect 25778 11396 25782 11452
rect 25782 11396 25838 11452
rect 25838 11396 25842 11452
rect 25778 11392 25842 11396
rect 25858 11452 25922 11456
rect 25858 11396 25862 11452
rect 25862 11396 25918 11452
rect 25918 11396 25922 11452
rect 25858 11392 25922 11396
rect 25938 11452 26002 11456
rect 25938 11396 25942 11452
rect 25942 11396 25998 11452
rect 25998 11396 26002 11452
rect 25938 11392 26002 11396
rect 26018 11452 26082 11456
rect 26018 11396 26022 11452
rect 26022 11396 26078 11452
rect 26078 11396 26082 11452
rect 26018 11392 26082 11396
rect 21404 11112 21468 11116
rect 21404 11056 21454 11112
rect 21454 11056 21468 11112
rect 21404 11052 21468 11056
rect 10882 10908 10946 10912
rect 10882 10852 10886 10908
rect 10886 10852 10942 10908
rect 10942 10852 10946 10908
rect 10882 10848 10946 10852
rect 10962 10908 11026 10912
rect 10962 10852 10966 10908
rect 10966 10852 11022 10908
rect 11022 10852 11026 10908
rect 10962 10848 11026 10852
rect 11042 10908 11106 10912
rect 11042 10852 11046 10908
rect 11046 10852 11102 10908
rect 11102 10852 11106 10908
rect 11042 10848 11106 10852
rect 11122 10908 11186 10912
rect 11122 10852 11126 10908
rect 11126 10852 11182 10908
rect 11182 10852 11186 10908
rect 11122 10848 11186 10852
rect 20813 10908 20877 10912
rect 20813 10852 20817 10908
rect 20817 10852 20873 10908
rect 20873 10852 20877 10908
rect 20813 10848 20877 10852
rect 20893 10908 20957 10912
rect 20893 10852 20897 10908
rect 20897 10852 20953 10908
rect 20953 10852 20957 10908
rect 20893 10848 20957 10852
rect 20973 10908 21037 10912
rect 20973 10852 20977 10908
rect 20977 10852 21033 10908
rect 21033 10852 21037 10908
rect 20973 10848 21037 10852
rect 21053 10908 21117 10912
rect 21053 10852 21057 10908
rect 21057 10852 21113 10908
rect 21113 10852 21117 10908
rect 21053 10848 21117 10852
rect 20484 10704 20548 10708
rect 20484 10648 20498 10704
rect 20498 10648 20548 10704
rect 20484 10644 20548 10648
rect 5917 10364 5981 10368
rect 5917 10308 5921 10364
rect 5921 10308 5977 10364
rect 5977 10308 5981 10364
rect 5917 10304 5981 10308
rect 5997 10364 6061 10368
rect 5997 10308 6001 10364
rect 6001 10308 6057 10364
rect 6057 10308 6061 10364
rect 5997 10304 6061 10308
rect 6077 10364 6141 10368
rect 6077 10308 6081 10364
rect 6081 10308 6137 10364
rect 6137 10308 6141 10364
rect 6077 10304 6141 10308
rect 6157 10364 6221 10368
rect 6157 10308 6161 10364
rect 6161 10308 6217 10364
rect 6217 10308 6221 10364
rect 6157 10304 6221 10308
rect 15848 10364 15912 10368
rect 15848 10308 15852 10364
rect 15852 10308 15908 10364
rect 15908 10308 15912 10364
rect 15848 10304 15912 10308
rect 15928 10364 15992 10368
rect 15928 10308 15932 10364
rect 15932 10308 15988 10364
rect 15988 10308 15992 10364
rect 15928 10304 15992 10308
rect 16008 10364 16072 10368
rect 16008 10308 16012 10364
rect 16012 10308 16068 10364
rect 16068 10308 16072 10364
rect 16008 10304 16072 10308
rect 16088 10364 16152 10368
rect 16088 10308 16092 10364
rect 16092 10308 16148 10364
rect 16148 10308 16152 10364
rect 16088 10304 16152 10308
rect 25778 10364 25842 10368
rect 25778 10308 25782 10364
rect 25782 10308 25838 10364
rect 25838 10308 25842 10364
rect 25778 10304 25842 10308
rect 25858 10364 25922 10368
rect 25858 10308 25862 10364
rect 25862 10308 25918 10364
rect 25918 10308 25922 10364
rect 25858 10304 25922 10308
rect 25938 10364 26002 10368
rect 25938 10308 25942 10364
rect 25942 10308 25998 10364
rect 25998 10308 26002 10364
rect 25938 10304 26002 10308
rect 26018 10364 26082 10368
rect 26018 10308 26022 10364
rect 26022 10308 26078 10364
rect 26078 10308 26082 10364
rect 26018 10304 26082 10308
rect 10882 9820 10946 9824
rect 10882 9764 10886 9820
rect 10886 9764 10942 9820
rect 10942 9764 10946 9820
rect 10882 9760 10946 9764
rect 10962 9820 11026 9824
rect 10962 9764 10966 9820
rect 10966 9764 11022 9820
rect 11022 9764 11026 9820
rect 10962 9760 11026 9764
rect 11042 9820 11106 9824
rect 11042 9764 11046 9820
rect 11046 9764 11102 9820
rect 11102 9764 11106 9820
rect 11042 9760 11106 9764
rect 11122 9820 11186 9824
rect 11122 9764 11126 9820
rect 11126 9764 11182 9820
rect 11182 9764 11186 9820
rect 11122 9760 11186 9764
rect 20813 9820 20877 9824
rect 20813 9764 20817 9820
rect 20817 9764 20873 9820
rect 20873 9764 20877 9820
rect 20813 9760 20877 9764
rect 20893 9820 20957 9824
rect 20893 9764 20897 9820
rect 20897 9764 20953 9820
rect 20953 9764 20957 9820
rect 20893 9760 20957 9764
rect 20973 9820 21037 9824
rect 20973 9764 20977 9820
rect 20977 9764 21033 9820
rect 21033 9764 21037 9820
rect 20973 9760 21037 9764
rect 21053 9820 21117 9824
rect 21053 9764 21057 9820
rect 21057 9764 21113 9820
rect 21113 9764 21117 9820
rect 21053 9760 21117 9764
rect 5917 9276 5981 9280
rect 5917 9220 5921 9276
rect 5921 9220 5977 9276
rect 5977 9220 5981 9276
rect 5917 9216 5981 9220
rect 5997 9276 6061 9280
rect 5997 9220 6001 9276
rect 6001 9220 6057 9276
rect 6057 9220 6061 9276
rect 5997 9216 6061 9220
rect 6077 9276 6141 9280
rect 6077 9220 6081 9276
rect 6081 9220 6137 9276
rect 6137 9220 6141 9276
rect 6077 9216 6141 9220
rect 6157 9276 6221 9280
rect 6157 9220 6161 9276
rect 6161 9220 6217 9276
rect 6217 9220 6221 9276
rect 6157 9216 6221 9220
rect 15848 9276 15912 9280
rect 15848 9220 15852 9276
rect 15852 9220 15908 9276
rect 15908 9220 15912 9276
rect 15848 9216 15912 9220
rect 15928 9276 15992 9280
rect 15928 9220 15932 9276
rect 15932 9220 15988 9276
rect 15988 9220 15992 9276
rect 15928 9216 15992 9220
rect 16008 9276 16072 9280
rect 16008 9220 16012 9276
rect 16012 9220 16068 9276
rect 16068 9220 16072 9276
rect 16008 9216 16072 9220
rect 16088 9276 16152 9280
rect 16088 9220 16092 9276
rect 16092 9220 16148 9276
rect 16148 9220 16152 9276
rect 16088 9216 16152 9220
rect 25778 9276 25842 9280
rect 25778 9220 25782 9276
rect 25782 9220 25838 9276
rect 25838 9220 25842 9276
rect 25778 9216 25842 9220
rect 25858 9276 25922 9280
rect 25858 9220 25862 9276
rect 25862 9220 25918 9276
rect 25918 9220 25922 9276
rect 25858 9216 25922 9220
rect 25938 9276 26002 9280
rect 25938 9220 25942 9276
rect 25942 9220 25998 9276
rect 25998 9220 26002 9276
rect 25938 9216 26002 9220
rect 26018 9276 26082 9280
rect 26018 9220 26022 9276
rect 26022 9220 26078 9276
rect 26078 9220 26082 9276
rect 26018 9216 26082 9220
rect 10882 8732 10946 8736
rect 10882 8676 10886 8732
rect 10886 8676 10942 8732
rect 10942 8676 10946 8732
rect 10882 8672 10946 8676
rect 10962 8732 11026 8736
rect 10962 8676 10966 8732
rect 10966 8676 11022 8732
rect 11022 8676 11026 8732
rect 10962 8672 11026 8676
rect 11042 8732 11106 8736
rect 11042 8676 11046 8732
rect 11046 8676 11102 8732
rect 11102 8676 11106 8732
rect 11042 8672 11106 8676
rect 11122 8732 11186 8736
rect 11122 8676 11126 8732
rect 11126 8676 11182 8732
rect 11182 8676 11186 8732
rect 11122 8672 11186 8676
rect 20813 8732 20877 8736
rect 20813 8676 20817 8732
rect 20817 8676 20873 8732
rect 20873 8676 20877 8732
rect 20813 8672 20877 8676
rect 20893 8732 20957 8736
rect 20893 8676 20897 8732
rect 20897 8676 20953 8732
rect 20953 8676 20957 8732
rect 20893 8672 20957 8676
rect 20973 8732 21037 8736
rect 20973 8676 20977 8732
rect 20977 8676 21033 8732
rect 21033 8676 21037 8732
rect 20973 8672 21037 8676
rect 21053 8732 21117 8736
rect 21053 8676 21057 8732
rect 21057 8676 21113 8732
rect 21113 8676 21117 8732
rect 21053 8672 21117 8676
rect 5917 8188 5981 8192
rect 5917 8132 5921 8188
rect 5921 8132 5977 8188
rect 5977 8132 5981 8188
rect 5917 8128 5981 8132
rect 5997 8188 6061 8192
rect 5997 8132 6001 8188
rect 6001 8132 6057 8188
rect 6057 8132 6061 8188
rect 5997 8128 6061 8132
rect 6077 8188 6141 8192
rect 6077 8132 6081 8188
rect 6081 8132 6137 8188
rect 6137 8132 6141 8188
rect 6077 8128 6141 8132
rect 6157 8188 6221 8192
rect 6157 8132 6161 8188
rect 6161 8132 6217 8188
rect 6217 8132 6221 8188
rect 6157 8128 6221 8132
rect 15848 8188 15912 8192
rect 15848 8132 15852 8188
rect 15852 8132 15908 8188
rect 15908 8132 15912 8188
rect 15848 8128 15912 8132
rect 15928 8188 15992 8192
rect 15928 8132 15932 8188
rect 15932 8132 15988 8188
rect 15988 8132 15992 8188
rect 15928 8128 15992 8132
rect 16008 8188 16072 8192
rect 16008 8132 16012 8188
rect 16012 8132 16068 8188
rect 16068 8132 16072 8188
rect 16008 8128 16072 8132
rect 16088 8188 16152 8192
rect 16088 8132 16092 8188
rect 16092 8132 16148 8188
rect 16148 8132 16152 8188
rect 16088 8128 16152 8132
rect 25778 8188 25842 8192
rect 25778 8132 25782 8188
rect 25782 8132 25838 8188
rect 25838 8132 25842 8188
rect 25778 8128 25842 8132
rect 25858 8188 25922 8192
rect 25858 8132 25862 8188
rect 25862 8132 25918 8188
rect 25918 8132 25922 8188
rect 25858 8128 25922 8132
rect 25938 8188 26002 8192
rect 25938 8132 25942 8188
rect 25942 8132 25998 8188
rect 25998 8132 26002 8188
rect 25938 8128 26002 8132
rect 26018 8188 26082 8192
rect 26018 8132 26022 8188
rect 26022 8132 26078 8188
rect 26078 8132 26082 8188
rect 26018 8128 26082 8132
rect 10882 7644 10946 7648
rect 10882 7588 10886 7644
rect 10886 7588 10942 7644
rect 10942 7588 10946 7644
rect 10882 7584 10946 7588
rect 10962 7644 11026 7648
rect 10962 7588 10966 7644
rect 10966 7588 11022 7644
rect 11022 7588 11026 7644
rect 10962 7584 11026 7588
rect 11042 7644 11106 7648
rect 11042 7588 11046 7644
rect 11046 7588 11102 7644
rect 11102 7588 11106 7644
rect 11042 7584 11106 7588
rect 11122 7644 11186 7648
rect 11122 7588 11126 7644
rect 11126 7588 11182 7644
rect 11182 7588 11186 7644
rect 11122 7584 11186 7588
rect 20813 7644 20877 7648
rect 20813 7588 20817 7644
rect 20817 7588 20873 7644
rect 20873 7588 20877 7644
rect 20813 7584 20877 7588
rect 20893 7644 20957 7648
rect 20893 7588 20897 7644
rect 20897 7588 20953 7644
rect 20953 7588 20957 7644
rect 20893 7584 20957 7588
rect 20973 7644 21037 7648
rect 20973 7588 20977 7644
rect 20977 7588 21033 7644
rect 21033 7588 21037 7644
rect 20973 7584 21037 7588
rect 21053 7644 21117 7648
rect 21053 7588 21057 7644
rect 21057 7588 21113 7644
rect 21113 7588 21117 7644
rect 21053 7584 21117 7588
rect 5917 7100 5981 7104
rect 5917 7044 5921 7100
rect 5921 7044 5977 7100
rect 5977 7044 5981 7100
rect 5917 7040 5981 7044
rect 5997 7100 6061 7104
rect 5997 7044 6001 7100
rect 6001 7044 6057 7100
rect 6057 7044 6061 7100
rect 5997 7040 6061 7044
rect 6077 7100 6141 7104
rect 6077 7044 6081 7100
rect 6081 7044 6137 7100
rect 6137 7044 6141 7100
rect 6077 7040 6141 7044
rect 6157 7100 6221 7104
rect 6157 7044 6161 7100
rect 6161 7044 6217 7100
rect 6217 7044 6221 7100
rect 6157 7040 6221 7044
rect 15848 7100 15912 7104
rect 15848 7044 15852 7100
rect 15852 7044 15908 7100
rect 15908 7044 15912 7100
rect 15848 7040 15912 7044
rect 15928 7100 15992 7104
rect 15928 7044 15932 7100
rect 15932 7044 15988 7100
rect 15988 7044 15992 7100
rect 15928 7040 15992 7044
rect 16008 7100 16072 7104
rect 16008 7044 16012 7100
rect 16012 7044 16068 7100
rect 16068 7044 16072 7100
rect 16008 7040 16072 7044
rect 16088 7100 16152 7104
rect 16088 7044 16092 7100
rect 16092 7044 16148 7100
rect 16148 7044 16152 7100
rect 16088 7040 16152 7044
rect 25778 7100 25842 7104
rect 25778 7044 25782 7100
rect 25782 7044 25838 7100
rect 25838 7044 25842 7100
rect 25778 7040 25842 7044
rect 25858 7100 25922 7104
rect 25858 7044 25862 7100
rect 25862 7044 25918 7100
rect 25918 7044 25922 7100
rect 25858 7040 25922 7044
rect 25938 7100 26002 7104
rect 25938 7044 25942 7100
rect 25942 7044 25998 7100
rect 25998 7044 26002 7100
rect 25938 7040 26002 7044
rect 26018 7100 26082 7104
rect 26018 7044 26022 7100
rect 26022 7044 26078 7100
rect 26078 7044 26082 7100
rect 26018 7040 26082 7044
rect 10882 6556 10946 6560
rect 10882 6500 10886 6556
rect 10886 6500 10942 6556
rect 10942 6500 10946 6556
rect 10882 6496 10946 6500
rect 10962 6556 11026 6560
rect 10962 6500 10966 6556
rect 10966 6500 11022 6556
rect 11022 6500 11026 6556
rect 10962 6496 11026 6500
rect 11042 6556 11106 6560
rect 11042 6500 11046 6556
rect 11046 6500 11102 6556
rect 11102 6500 11106 6556
rect 11042 6496 11106 6500
rect 11122 6556 11186 6560
rect 11122 6500 11126 6556
rect 11126 6500 11182 6556
rect 11182 6500 11186 6556
rect 11122 6496 11186 6500
rect 20813 6556 20877 6560
rect 20813 6500 20817 6556
rect 20817 6500 20873 6556
rect 20873 6500 20877 6556
rect 20813 6496 20877 6500
rect 20893 6556 20957 6560
rect 20893 6500 20897 6556
rect 20897 6500 20953 6556
rect 20953 6500 20957 6556
rect 20893 6496 20957 6500
rect 20973 6556 21037 6560
rect 20973 6500 20977 6556
rect 20977 6500 21033 6556
rect 21033 6500 21037 6556
rect 20973 6496 21037 6500
rect 21053 6556 21117 6560
rect 21053 6500 21057 6556
rect 21057 6500 21113 6556
rect 21113 6500 21117 6556
rect 21053 6496 21117 6500
rect 5917 6012 5981 6016
rect 5917 5956 5921 6012
rect 5921 5956 5977 6012
rect 5977 5956 5981 6012
rect 5917 5952 5981 5956
rect 5997 6012 6061 6016
rect 5997 5956 6001 6012
rect 6001 5956 6057 6012
rect 6057 5956 6061 6012
rect 5997 5952 6061 5956
rect 6077 6012 6141 6016
rect 6077 5956 6081 6012
rect 6081 5956 6137 6012
rect 6137 5956 6141 6012
rect 6077 5952 6141 5956
rect 6157 6012 6221 6016
rect 6157 5956 6161 6012
rect 6161 5956 6217 6012
rect 6217 5956 6221 6012
rect 6157 5952 6221 5956
rect 15848 6012 15912 6016
rect 15848 5956 15852 6012
rect 15852 5956 15908 6012
rect 15908 5956 15912 6012
rect 15848 5952 15912 5956
rect 15928 6012 15992 6016
rect 15928 5956 15932 6012
rect 15932 5956 15988 6012
rect 15988 5956 15992 6012
rect 15928 5952 15992 5956
rect 16008 6012 16072 6016
rect 16008 5956 16012 6012
rect 16012 5956 16068 6012
rect 16068 5956 16072 6012
rect 16008 5952 16072 5956
rect 16088 6012 16152 6016
rect 16088 5956 16092 6012
rect 16092 5956 16148 6012
rect 16148 5956 16152 6012
rect 16088 5952 16152 5956
rect 25778 6012 25842 6016
rect 25778 5956 25782 6012
rect 25782 5956 25838 6012
rect 25838 5956 25842 6012
rect 25778 5952 25842 5956
rect 25858 6012 25922 6016
rect 25858 5956 25862 6012
rect 25862 5956 25918 6012
rect 25918 5956 25922 6012
rect 25858 5952 25922 5956
rect 25938 6012 26002 6016
rect 25938 5956 25942 6012
rect 25942 5956 25998 6012
rect 25998 5956 26002 6012
rect 25938 5952 26002 5956
rect 26018 6012 26082 6016
rect 26018 5956 26022 6012
rect 26022 5956 26078 6012
rect 26078 5956 26082 6012
rect 26018 5952 26082 5956
rect 10882 5468 10946 5472
rect 10882 5412 10886 5468
rect 10886 5412 10942 5468
rect 10942 5412 10946 5468
rect 10882 5408 10946 5412
rect 10962 5468 11026 5472
rect 10962 5412 10966 5468
rect 10966 5412 11022 5468
rect 11022 5412 11026 5468
rect 10962 5408 11026 5412
rect 11042 5468 11106 5472
rect 11042 5412 11046 5468
rect 11046 5412 11102 5468
rect 11102 5412 11106 5468
rect 11042 5408 11106 5412
rect 11122 5468 11186 5472
rect 11122 5412 11126 5468
rect 11126 5412 11182 5468
rect 11182 5412 11186 5468
rect 11122 5408 11186 5412
rect 20813 5468 20877 5472
rect 20813 5412 20817 5468
rect 20817 5412 20873 5468
rect 20873 5412 20877 5468
rect 20813 5408 20877 5412
rect 20893 5468 20957 5472
rect 20893 5412 20897 5468
rect 20897 5412 20953 5468
rect 20953 5412 20957 5468
rect 20893 5408 20957 5412
rect 20973 5468 21037 5472
rect 20973 5412 20977 5468
rect 20977 5412 21033 5468
rect 21033 5412 21037 5468
rect 20973 5408 21037 5412
rect 21053 5468 21117 5472
rect 21053 5412 21057 5468
rect 21057 5412 21113 5468
rect 21113 5412 21117 5468
rect 21053 5408 21117 5412
rect 5917 4924 5981 4928
rect 5917 4868 5921 4924
rect 5921 4868 5977 4924
rect 5977 4868 5981 4924
rect 5917 4864 5981 4868
rect 5997 4924 6061 4928
rect 5997 4868 6001 4924
rect 6001 4868 6057 4924
rect 6057 4868 6061 4924
rect 5997 4864 6061 4868
rect 6077 4924 6141 4928
rect 6077 4868 6081 4924
rect 6081 4868 6137 4924
rect 6137 4868 6141 4924
rect 6077 4864 6141 4868
rect 6157 4924 6221 4928
rect 6157 4868 6161 4924
rect 6161 4868 6217 4924
rect 6217 4868 6221 4924
rect 6157 4864 6221 4868
rect 15848 4924 15912 4928
rect 15848 4868 15852 4924
rect 15852 4868 15908 4924
rect 15908 4868 15912 4924
rect 15848 4864 15912 4868
rect 15928 4924 15992 4928
rect 15928 4868 15932 4924
rect 15932 4868 15988 4924
rect 15988 4868 15992 4924
rect 15928 4864 15992 4868
rect 16008 4924 16072 4928
rect 16008 4868 16012 4924
rect 16012 4868 16068 4924
rect 16068 4868 16072 4924
rect 16008 4864 16072 4868
rect 16088 4924 16152 4928
rect 16088 4868 16092 4924
rect 16092 4868 16148 4924
rect 16148 4868 16152 4924
rect 16088 4864 16152 4868
rect 25778 4924 25842 4928
rect 25778 4868 25782 4924
rect 25782 4868 25838 4924
rect 25838 4868 25842 4924
rect 25778 4864 25842 4868
rect 25858 4924 25922 4928
rect 25858 4868 25862 4924
rect 25862 4868 25918 4924
rect 25918 4868 25922 4924
rect 25858 4864 25922 4868
rect 25938 4924 26002 4928
rect 25938 4868 25942 4924
rect 25942 4868 25998 4924
rect 25998 4868 26002 4924
rect 25938 4864 26002 4868
rect 26018 4924 26082 4928
rect 26018 4868 26022 4924
rect 26022 4868 26078 4924
rect 26078 4868 26082 4924
rect 26018 4864 26082 4868
rect 10882 4380 10946 4384
rect 10882 4324 10886 4380
rect 10886 4324 10942 4380
rect 10942 4324 10946 4380
rect 10882 4320 10946 4324
rect 10962 4380 11026 4384
rect 10962 4324 10966 4380
rect 10966 4324 11022 4380
rect 11022 4324 11026 4380
rect 10962 4320 11026 4324
rect 11042 4380 11106 4384
rect 11042 4324 11046 4380
rect 11046 4324 11102 4380
rect 11102 4324 11106 4380
rect 11042 4320 11106 4324
rect 11122 4380 11186 4384
rect 11122 4324 11126 4380
rect 11126 4324 11182 4380
rect 11182 4324 11186 4380
rect 11122 4320 11186 4324
rect 20813 4380 20877 4384
rect 20813 4324 20817 4380
rect 20817 4324 20873 4380
rect 20873 4324 20877 4380
rect 20813 4320 20877 4324
rect 20893 4380 20957 4384
rect 20893 4324 20897 4380
rect 20897 4324 20953 4380
rect 20953 4324 20957 4380
rect 20893 4320 20957 4324
rect 20973 4380 21037 4384
rect 20973 4324 20977 4380
rect 20977 4324 21033 4380
rect 21033 4324 21037 4380
rect 20973 4320 21037 4324
rect 21053 4380 21117 4384
rect 21053 4324 21057 4380
rect 21057 4324 21113 4380
rect 21113 4324 21117 4380
rect 21053 4320 21117 4324
rect 5917 3836 5981 3840
rect 5917 3780 5921 3836
rect 5921 3780 5977 3836
rect 5977 3780 5981 3836
rect 5917 3776 5981 3780
rect 5997 3836 6061 3840
rect 5997 3780 6001 3836
rect 6001 3780 6057 3836
rect 6057 3780 6061 3836
rect 5997 3776 6061 3780
rect 6077 3836 6141 3840
rect 6077 3780 6081 3836
rect 6081 3780 6137 3836
rect 6137 3780 6141 3836
rect 6077 3776 6141 3780
rect 6157 3836 6221 3840
rect 6157 3780 6161 3836
rect 6161 3780 6217 3836
rect 6217 3780 6221 3836
rect 6157 3776 6221 3780
rect 15848 3836 15912 3840
rect 15848 3780 15852 3836
rect 15852 3780 15908 3836
rect 15908 3780 15912 3836
rect 15848 3776 15912 3780
rect 15928 3836 15992 3840
rect 15928 3780 15932 3836
rect 15932 3780 15988 3836
rect 15988 3780 15992 3836
rect 15928 3776 15992 3780
rect 16008 3836 16072 3840
rect 16008 3780 16012 3836
rect 16012 3780 16068 3836
rect 16068 3780 16072 3836
rect 16008 3776 16072 3780
rect 16088 3836 16152 3840
rect 16088 3780 16092 3836
rect 16092 3780 16148 3836
rect 16148 3780 16152 3836
rect 16088 3776 16152 3780
rect 25778 3836 25842 3840
rect 25778 3780 25782 3836
rect 25782 3780 25838 3836
rect 25838 3780 25842 3836
rect 25778 3776 25842 3780
rect 25858 3836 25922 3840
rect 25858 3780 25862 3836
rect 25862 3780 25918 3836
rect 25918 3780 25922 3836
rect 25858 3776 25922 3780
rect 25938 3836 26002 3840
rect 25938 3780 25942 3836
rect 25942 3780 25998 3836
rect 25998 3780 26002 3836
rect 25938 3776 26002 3780
rect 26018 3836 26082 3840
rect 26018 3780 26022 3836
rect 26022 3780 26078 3836
rect 26078 3780 26082 3836
rect 26018 3776 26082 3780
rect 10882 3292 10946 3296
rect 10882 3236 10886 3292
rect 10886 3236 10942 3292
rect 10942 3236 10946 3292
rect 10882 3232 10946 3236
rect 10962 3292 11026 3296
rect 10962 3236 10966 3292
rect 10966 3236 11022 3292
rect 11022 3236 11026 3292
rect 10962 3232 11026 3236
rect 11042 3292 11106 3296
rect 11042 3236 11046 3292
rect 11046 3236 11102 3292
rect 11102 3236 11106 3292
rect 11042 3232 11106 3236
rect 11122 3292 11186 3296
rect 11122 3236 11126 3292
rect 11126 3236 11182 3292
rect 11182 3236 11186 3292
rect 11122 3232 11186 3236
rect 20813 3292 20877 3296
rect 20813 3236 20817 3292
rect 20817 3236 20873 3292
rect 20873 3236 20877 3292
rect 20813 3232 20877 3236
rect 20893 3292 20957 3296
rect 20893 3236 20897 3292
rect 20897 3236 20953 3292
rect 20953 3236 20957 3292
rect 20893 3232 20957 3236
rect 20973 3292 21037 3296
rect 20973 3236 20977 3292
rect 20977 3236 21033 3292
rect 21033 3236 21037 3292
rect 20973 3232 21037 3236
rect 21053 3292 21117 3296
rect 21053 3236 21057 3292
rect 21057 3236 21113 3292
rect 21113 3236 21117 3292
rect 21053 3232 21117 3236
rect 5917 2748 5981 2752
rect 5917 2692 5921 2748
rect 5921 2692 5977 2748
rect 5977 2692 5981 2748
rect 5917 2688 5981 2692
rect 5997 2748 6061 2752
rect 5997 2692 6001 2748
rect 6001 2692 6057 2748
rect 6057 2692 6061 2748
rect 5997 2688 6061 2692
rect 6077 2748 6141 2752
rect 6077 2692 6081 2748
rect 6081 2692 6137 2748
rect 6137 2692 6141 2748
rect 6077 2688 6141 2692
rect 6157 2748 6221 2752
rect 6157 2692 6161 2748
rect 6161 2692 6217 2748
rect 6217 2692 6221 2748
rect 6157 2688 6221 2692
rect 15848 2748 15912 2752
rect 15848 2692 15852 2748
rect 15852 2692 15908 2748
rect 15908 2692 15912 2748
rect 15848 2688 15912 2692
rect 15928 2748 15992 2752
rect 15928 2692 15932 2748
rect 15932 2692 15988 2748
rect 15988 2692 15992 2748
rect 15928 2688 15992 2692
rect 16008 2748 16072 2752
rect 16008 2692 16012 2748
rect 16012 2692 16068 2748
rect 16068 2692 16072 2748
rect 16008 2688 16072 2692
rect 16088 2748 16152 2752
rect 16088 2692 16092 2748
rect 16092 2692 16148 2748
rect 16148 2692 16152 2748
rect 16088 2688 16152 2692
rect 25778 2748 25842 2752
rect 25778 2692 25782 2748
rect 25782 2692 25838 2748
rect 25838 2692 25842 2748
rect 25778 2688 25842 2692
rect 25858 2748 25922 2752
rect 25858 2692 25862 2748
rect 25862 2692 25918 2748
rect 25918 2692 25922 2748
rect 25858 2688 25922 2692
rect 25938 2748 26002 2752
rect 25938 2692 25942 2748
rect 25942 2692 25998 2748
rect 25998 2692 26002 2748
rect 25938 2688 26002 2692
rect 26018 2748 26082 2752
rect 26018 2692 26022 2748
rect 26022 2692 26078 2748
rect 26078 2692 26082 2748
rect 26018 2688 26082 2692
rect 10882 2204 10946 2208
rect 10882 2148 10886 2204
rect 10886 2148 10942 2204
rect 10942 2148 10946 2204
rect 10882 2144 10946 2148
rect 10962 2204 11026 2208
rect 10962 2148 10966 2204
rect 10966 2148 11022 2204
rect 11022 2148 11026 2204
rect 10962 2144 11026 2148
rect 11042 2204 11106 2208
rect 11042 2148 11046 2204
rect 11046 2148 11102 2204
rect 11102 2148 11106 2204
rect 11042 2144 11106 2148
rect 11122 2204 11186 2208
rect 11122 2148 11126 2204
rect 11126 2148 11182 2204
rect 11182 2148 11186 2204
rect 11122 2144 11186 2148
rect 20813 2204 20877 2208
rect 20813 2148 20817 2204
rect 20817 2148 20873 2204
rect 20873 2148 20877 2204
rect 20813 2144 20877 2148
rect 20893 2204 20957 2208
rect 20893 2148 20897 2204
rect 20897 2148 20953 2204
rect 20953 2148 20957 2204
rect 20893 2144 20957 2148
rect 20973 2204 21037 2208
rect 20973 2148 20977 2204
rect 20977 2148 21033 2204
rect 21033 2148 21037 2204
rect 20973 2144 21037 2148
rect 21053 2204 21117 2208
rect 21053 2148 21057 2204
rect 21057 2148 21113 2204
rect 21113 2148 21117 2204
rect 21053 2144 21117 2148
<< metal4 >>
rect 5909 45184 6229 45744
rect 5909 45120 5917 45184
rect 5981 45120 5997 45184
rect 6061 45120 6077 45184
rect 6141 45120 6157 45184
rect 6221 45120 6229 45184
rect 5909 44096 6229 45120
rect 5909 44032 5917 44096
rect 5981 44032 5997 44096
rect 6061 44032 6077 44096
rect 6141 44032 6157 44096
rect 6221 44032 6229 44096
rect 5909 43008 6229 44032
rect 5909 42944 5917 43008
rect 5981 42944 5997 43008
rect 6061 42944 6077 43008
rect 6141 42944 6157 43008
rect 6221 42944 6229 43008
rect 5909 41920 6229 42944
rect 5909 41856 5917 41920
rect 5981 41856 5997 41920
rect 6061 41856 6077 41920
rect 6141 41856 6157 41920
rect 6221 41856 6229 41920
rect 5909 40832 6229 41856
rect 5909 40768 5917 40832
rect 5981 40768 5997 40832
rect 6061 40768 6077 40832
rect 6141 40768 6157 40832
rect 6221 40768 6229 40832
rect 5909 39744 6229 40768
rect 5909 39680 5917 39744
rect 5981 39680 5997 39744
rect 6061 39680 6077 39744
rect 6141 39680 6157 39744
rect 6221 39680 6229 39744
rect 5909 38656 6229 39680
rect 5909 38592 5917 38656
rect 5981 38592 5997 38656
rect 6061 38592 6077 38656
rect 6141 38592 6157 38656
rect 6221 38592 6229 38656
rect 5909 37568 6229 38592
rect 5909 37504 5917 37568
rect 5981 37504 5997 37568
rect 6061 37504 6077 37568
rect 6141 37504 6157 37568
rect 6221 37504 6229 37568
rect 5909 36480 6229 37504
rect 5909 36416 5917 36480
rect 5981 36416 5997 36480
rect 6061 36416 6077 36480
rect 6141 36416 6157 36480
rect 6221 36416 6229 36480
rect 5909 35392 6229 36416
rect 5909 35328 5917 35392
rect 5981 35328 5997 35392
rect 6061 35328 6077 35392
rect 6141 35328 6157 35392
rect 6221 35328 6229 35392
rect 5909 34304 6229 35328
rect 5909 34240 5917 34304
rect 5981 34240 5997 34304
rect 6061 34240 6077 34304
rect 6141 34240 6157 34304
rect 6221 34240 6229 34304
rect 5909 33216 6229 34240
rect 5909 33152 5917 33216
rect 5981 33152 5997 33216
rect 6061 33152 6077 33216
rect 6141 33152 6157 33216
rect 6221 33152 6229 33216
rect 5909 32128 6229 33152
rect 5909 32064 5917 32128
rect 5981 32064 5997 32128
rect 6061 32064 6077 32128
rect 6141 32064 6157 32128
rect 6221 32064 6229 32128
rect 5909 31040 6229 32064
rect 5909 30976 5917 31040
rect 5981 30976 5997 31040
rect 6061 30976 6077 31040
rect 6141 30976 6157 31040
rect 6221 30976 6229 31040
rect 5909 29952 6229 30976
rect 5909 29888 5917 29952
rect 5981 29888 5997 29952
rect 6061 29888 6077 29952
rect 6141 29888 6157 29952
rect 6221 29888 6229 29952
rect 5909 28864 6229 29888
rect 5909 28800 5917 28864
rect 5981 28800 5997 28864
rect 6061 28800 6077 28864
rect 6141 28800 6157 28864
rect 6221 28800 6229 28864
rect 5909 27776 6229 28800
rect 5909 27712 5917 27776
rect 5981 27712 5997 27776
rect 6061 27712 6077 27776
rect 6141 27712 6157 27776
rect 6221 27712 6229 27776
rect 5909 26688 6229 27712
rect 5909 26624 5917 26688
rect 5981 26624 5997 26688
rect 6061 26624 6077 26688
rect 6141 26624 6157 26688
rect 6221 26624 6229 26688
rect 5909 25600 6229 26624
rect 5909 25536 5917 25600
rect 5981 25536 5997 25600
rect 6061 25536 6077 25600
rect 6141 25536 6157 25600
rect 6221 25536 6229 25600
rect 5909 24512 6229 25536
rect 5909 24448 5917 24512
rect 5981 24448 5997 24512
rect 6061 24448 6077 24512
rect 6141 24448 6157 24512
rect 6221 24448 6229 24512
rect 5909 23424 6229 24448
rect 5909 23360 5917 23424
rect 5981 23360 5997 23424
rect 6061 23360 6077 23424
rect 6141 23360 6157 23424
rect 6221 23360 6229 23424
rect 5909 22336 6229 23360
rect 5909 22272 5917 22336
rect 5981 22272 5997 22336
rect 6061 22272 6077 22336
rect 6141 22272 6157 22336
rect 6221 22272 6229 22336
rect 5909 21248 6229 22272
rect 5909 21184 5917 21248
rect 5981 21184 5997 21248
rect 6061 21184 6077 21248
rect 6141 21184 6157 21248
rect 6221 21184 6229 21248
rect 5909 20160 6229 21184
rect 5909 20096 5917 20160
rect 5981 20096 5997 20160
rect 6061 20096 6077 20160
rect 6141 20096 6157 20160
rect 6221 20096 6229 20160
rect 5909 19072 6229 20096
rect 5909 19008 5917 19072
rect 5981 19008 5997 19072
rect 6061 19008 6077 19072
rect 6141 19008 6157 19072
rect 6221 19008 6229 19072
rect 5909 17984 6229 19008
rect 5909 17920 5917 17984
rect 5981 17920 5997 17984
rect 6061 17920 6077 17984
rect 6141 17920 6157 17984
rect 6221 17920 6229 17984
rect 5909 16896 6229 17920
rect 5909 16832 5917 16896
rect 5981 16832 5997 16896
rect 6061 16832 6077 16896
rect 6141 16832 6157 16896
rect 6221 16832 6229 16896
rect 5909 15808 6229 16832
rect 5909 15744 5917 15808
rect 5981 15744 5997 15808
rect 6061 15744 6077 15808
rect 6141 15744 6157 15808
rect 6221 15744 6229 15808
rect 5909 14720 6229 15744
rect 5909 14656 5917 14720
rect 5981 14656 5997 14720
rect 6061 14656 6077 14720
rect 6141 14656 6157 14720
rect 6221 14656 6229 14720
rect 5909 13632 6229 14656
rect 5909 13568 5917 13632
rect 5981 13568 5997 13632
rect 6061 13568 6077 13632
rect 6141 13568 6157 13632
rect 6221 13568 6229 13632
rect 5909 12544 6229 13568
rect 5909 12480 5917 12544
rect 5981 12480 5997 12544
rect 6061 12480 6077 12544
rect 6141 12480 6157 12544
rect 6221 12480 6229 12544
rect 5909 11456 6229 12480
rect 5909 11392 5917 11456
rect 5981 11392 5997 11456
rect 6061 11392 6077 11456
rect 6141 11392 6157 11456
rect 6221 11392 6229 11456
rect 5909 10368 6229 11392
rect 5909 10304 5917 10368
rect 5981 10304 5997 10368
rect 6061 10304 6077 10368
rect 6141 10304 6157 10368
rect 6221 10304 6229 10368
rect 5909 9280 6229 10304
rect 5909 9216 5917 9280
rect 5981 9216 5997 9280
rect 6061 9216 6077 9280
rect 6141 9216 6157 9280
rect 6221 9216 6229 9280
rect 5909 8192 6229 9216
rect 5909 8128 5917 8192
rect 5981 8128 5997 8192
rect 6061 8128 6077 8192
rect 6141 8128 6157 8192
rect 6221 8128 6229 8192
rect 5909 7104 6229 8128
rect 5909 7040 5917 7104
rect 5981 7040 5997 7104
rect 6061 7040 6077 7104
rect 6141 7040 6157 7104
rect 6221 7040 6229 7104
rect 5909 6016 6229 7040
rect 5909 5952 5917 6016
rect 5981 5952 5997 6016
rect 6061 5952 6077 6016
rect 6141 5952 6157 6016
rect 6221 5952 6229 6016
rect 5909 4928 6229 5952
rect 5909 4864 5917 4928
rect 5981 4864 5997 4928
rect 6061 4864 6077 4928
rect 6141 4864 6157 4928
rect 6221 4864 6229 4928
rect 5909 3840 6229 4864
rect 5909 3776 5917 3840
rect 5981 3776 5997 3840
rect 6061 3776 6077 3840
rect 6141 3776 6157 3840
rect 6221 3776 6229 3840
rect 5909 2752 6229 3776
rect 5909 2688 5917 2752
rect 5981 2688 5997 2752
rect 6061 2688 6077 2752
rect 6141 2688 6157 2752
rect 6221 2688 6229 2752
rect 5909 2128 6229 2688
rect 10874 45728 11194 45744
rect 10874 45664 10882 45728
rect 10946 45664 10962 45728
rect 11026 45664 11042 45728
rect 11106 45664 11122 45728
rect 11186 45664 11194 45728
rect 10874 44640 11194 45664
rect 10874 44576 10882 44640
rect 10946 44576 10962 44640
rect 11026 44576 11042 44640
rect 11106 44576 11122 44640
rect 11186 44576 11194 44640
rect 10874 43552 11194 44576
rect 10874 43488 10882 43552
rect 10946 43488 10962 43552
rect 11026 43488 11042 43552
rect 11106 43488 11122 43552
rect 11186 43488 11194 43552
rect 10874 42464 11194 43488
rect 10874 42400 10882 42464
rect 10946 42400 10962 42464
rect 11026 42400 11042 42464
rect 11106 42400 11122 42464
rect 11186 42400 11194 42464
rect 10874 41376 11194 42400
rect 10874 41312 10882 41376
rect 10946 41312 10962 41376
rect 11026 41312 11042 41376
rect 11106 41312 11122 41376
rect 11186 41312 11194 41376
rect 10874 40288 11194 41312
rect 10874 40224 10882 40288
rect 10946 40224 10962 40288
rect 11026 40224 11042 40288
rect 11106 40224 11122 40288
rect 11186 40224 11194 40288
rect 10874 39200 11194 40224
rect 10874 39136 10882 39200
rect 10946 39136 10962 39200
rect 11026 39136 11042 39200
rect 11106 39136 11122 39200
rect 11186 39136 11194 39200
rect 10874 38112 11194 39136
rect 10874 38048 10882 38112
rect 10946 38048 10962 38112
rect 11026 38048 11042 38112
rect 11106 38048 11122 38112
rect 11186 38048 11194 38112
rect 10874 37024 11194 38048
rect 10874 36960 10882 37024
rect 10946 36960 10962 37024
rect 11026 36960 11042 37024
rect 11106 36960 11122 37024
rect 11186 36960 11194 37024
rect 10874 35936 11194 36960
rect 10874 35872 10882 35936
rect 10946 35872 10962 35936
rect 11026 35872 11042 35936
rect 11106 35872 11122 35936
rect 11186 35872 11194 35936
rect 10874 34848 11194 35872
rect 10874 34784 10882 34848
rect 10946 34784 10962 34848
rect 11026 34784 11042 34848
rect 11106 34784 11122 34848
rect 11186 34784 11194 34848
rect 10874 33760 11194 34784
rect 10874 33696 10882 33760
rect 10946 33696 10962 33760
rect 11026 33696 11042 33760
rect 11106 33696 11122 33760
rect 11186 33696 11194 33760
rect 10874 32672 11194 33696
rect 10874 32608 10882 32672
rect 10946 32608 10962 32672
rect 11026 32608 11042 32672
rect 11106 32608 11122 32672
rect 11186 32608 11194 32672
rect 10874 31584 11194 32608
rect 10874 31520 10882 31584
rect 10946 31520 10962 31584
rect 11026 31520 11042 31584
rect 11106 31520 11122 31584
rect 11186 31520 11194 31584
rect 10874 30496 11194 31520
rect 10874 30432 10882 30496
rect 10946 30432 10962 30496
rect 11026 30432 11042 30496
rect 11106 30432 11122 30496
rect 11186 30432 11194 30496
rect 10874 29408 11194 30432
rect 10874 29344 10882 29408
rect 10946 29344 10962 29408
rect 11026 29344 11042 29408
rect 11106 29344 11122 29408
rect 11186 29344 11194 29408
rect 10874 28320 11194 29344
rect 10874 28256 10882 28320
rect 10946 28256 10962 28320
rect 11026 28256 11042 28320
rect 11106 28256 11122 28320
rect 11186 28256 11194 28320
rect 10874 27232 11194 28256
rect 10874 27168 10882 27232
rect 10946 27168 10962 27232
rect 11026 27168 11042 27232
rect 11106 27168 11122 27232
rect 11186 27168 11194 27232
rect 10874 26144 11194 27168
rect 10874 26080 10882 26144
rect 10946 26080 10962 26144
rect 11026 26080 11042 26144
rect 11106 26080 11122 26144
rect 11186 26080 11194 26144
rect 10874 25056 11194 26080
rect 10874 24992 10882 25056
rect 10946 24992 10962 25056
rect 11026 24992 11042 25056
rect 11106 24992 11122 25056
rect 11186 24992 11194 25056
rect 10874 23968 11194 24992
rect 10874 23904 10882 23968
rect 10946 23904 10962 23968
rect 11026 23904 11042 23968
rect 11106 23904 11122 23968
rect 11186 23904 11194 23968
rect 10874 22880 11194 23904
rect 10874 22816 10882 22880
rect 10946 22816 10962 22880
rect 11026 22816 11042 22880
rect 11106 22816 11122 22880
rect 11186 22816 11194 22880
rect 10874 21792 11194 22816
rect 10874 21728 10882 21792
rect 10946 21728 10962 21792
rect 11026 21728 11042 21792
rect 11106 21728 11122 21792
rect 11186 21728 11194 21792
rect 10874 20704 11194 21728
rect 10874 20640 10882 20704
rect 10946 20640 10962 20704
rect 11026 20640 11042 20704
rect 11106 20640 11122 20704
rect 11186 20640 11194 20704
rect 10874 19616 11194 20640
rect 10874 19552 10882 19616
rect 10946 19552 10962 19616
rect 11026 19552 11042 19616
rect 11106 19552 11122 19616
rect 11186 19552 11194 19616
rect 10874 18528 11194 19552
rect 10874 18464 10882 18528
rect 10946 18464 10962 18528
rect 11026 18464 11042 18528
rect 11106 18464 11122 18528
rect 11186 18464 11194 18528
rect 10874 17440 11194 18464
rect 10874 17376 10882 17440
rect 10946 17376 10962 17440
rect 11026 17376 11042 17440
rect 11106 17376 11122 17440
rect 11186 17376 11194 17440
rect 10874 16352 11194 17376
rect 10874 16288 10882 16352
rect 10946 16288 10962 16352
rect 11026 16288 11042 16352
rect 11106 16288 11122 16352
rect 11186 16288 11194 16352
rect 10874 15264 11194 16288
rect 10874 15200 10882 15264
rect 10946 15200 10962 15264
rect 11026 15200 11042 15264
rect 11106 15200 11122 15264
rect 11186 15200 11194 15264
rect 10874 14176 11194 15200
rect 10874 14112 10882 14176
rect 10946 14112 10962 14176
rect 11026 14112 11042 14176
rect 11106 14112 11122 14176
rect 11186 14112 11194 14176
rect 10874 13088 11194 14112
rect 10874 13024 10882 13088
rect 10946 13024 10962 13088
rect 11026 13024 11042 13088
rect 11106 13024 11122 13088
rect 11186 13024 11194 13088
rect 10874 12000 11194 13024
rect 10874 11936 10882 12000
rect 10946 11936 10962 12000
rect 11026 11936 11042 12000
rect 11106 11936 11122 12000
rect 11186 11936 11194 12000
rect 10874 10912 11194 11936
rect 10874 10848 10882 10912
rect 10946 10848 10962 10912
rect 11026 10848 11042 10912
rect 11106 10848 11122 10912
rect 11186 10848 11194 10912
rect 10874 9824 11194 10848
rect 10874 9760 10882 9824
rect 10946 9760 10962 9824
rect 11026 9760 11042 9824
rect 11106 9760 11122 9824
rect 11186 9760 11194 9824
rect 10874 8736 11194 9760
rect 10874 8672 10882 8736
rect 10946 8672 10962 8736
rect 11026 8672 11042 8736
rect 11106 8672 11122 8736
rect 11186 8672 11194 8736
rect 10874 7648 11194 8672
rect 10874 7584 10882 7648
rect 10946 7584 10962 7648
rect 11026 7584 11042 7648
rect 11106 7584 11122 7648
rect 11186 7584 11194 7648
rect 10874 6560 11194 7584
rect 10874 6496 10882 6560
rect 10946 6496 10962 6560
rect 11026 6496 11042 6560
rect 11106 6496 11122 6560
rect 11186 6496 11194 6560
rect 10874 5472 11194 6496
rect 10874 5408 10882 5472
rect 10946 5408 10962 5472
rect 11026 5408 11042 5472
rect 11106 5408 11122 5472
rect 11186 5408 11194 5472
rect 10874 4384 11194 5408
rect 10874 4320 10882 4384
rect 10946 4320 10962 4384
rect 11026 4320 11042 4384
rect 11106 4320 11122 4384
rect 11186 4320 11194 4384
rect 10874 3296 11194 4320
rect 10874 3232 10882 3296
rect 10946 3232 10962 3296
rect 11026 3232 11042 3296
rect 11106 3232 11122 3296
rect 11186 3232 11194 3296
rect 10874 2208 11194 3232
rect 10874 2144 10882 2208
rect 10946 2144 10962 2208
rect 11026 2144 11042 2208
rect 11106 2144 11122 2208
rect 11186 2144 11194 2208
rect 10874 2128 11194 2144
rect 15839 45184 16160 45744
rect 15839 45120 15848 45184
rect 15912 45120 15928 45184
rect 15992 45120 16008 45184
rect 16072 45120 16088 45184
rect 16152 45120 16160 45184
rect 15839 44096 16160 45120
rect 15839 44032 15848 44096
rect 15912 44032 15928 44096
rect 15992 44032 16008 44096
rect 16072 44032 16088 44096
rect 16152 44032 16160 44096
rect 15839 43008 16160 44032
rect 15839 42944 15848 43008
rect 15912 42944 15928 43008
rect 15992 42944 16008 43008
rect 16072 42944 16088 43008
rect 16152 42944 16160 43008
rect 15839 41920 16160 42944
rect 15839 41856 15848 41920
rect 15912 41856 15928 41920
rect 15992 41856 16008 41920
rect 16072 41856 16088 41920
rect 16152 41856 16160 41920
rect 15839 40832 16160 41856
rect 15839 40768 15848 40832
rect 15912 40768 15928 40832
rect 15992 40768 16008 40832
rect 16072 40768 16088 40832
rect 16152 40768 16160 40832
rect 15839 39744 16160 40768
rect 15839 39680 15848 39744
rect 15912 39680 15928 39744
rect 15992 39680 16008 39744
rect 16072 39680 16088 39744
rect 16152 39680 16160 39744
rect 15839 38656 16160 39680
rect 15839 38592 15848 38656
rect 15912 38592 15928 38656
rect 15992 38592 16008 38656
rect 16072 38592 16088 38656
rect 16152 38592 16160 38656
rect 15839 37568 16160 38592
rect 15839 37504 15848 37568
rect 15912 37504 15928 37568
rect 15992 37504 16008 37568
rect 16072 37504 16088 37568
rect 16152 37504 16160 37568
rect 15839 36480 16160 37504
rect 15839 36416 15848 36480
rect 15912 36416 15928 36480
rect 15992 36416 16008 36480
rect 16072 36416 16088 36480
rect 16152 36416 16160 36480
rect 15839 35392 16160 36416
rect 20805 45728 21125 45744
rect 20805 45664 20813 45728
rect 20877 45664 20893 45728
rect 20957 45664 20973 45728
rect 21037 45664 21053 45728
rect 21117 45664 21125 45728
rect 20805 44640 21125 45664
rect 25770 45184 26090 45744
rect 25770 45120 25778 45184
rect 25842 45120 25858 45184
rect 25922 45120 25938 45184
rect 26002 45120 26018 45184
rect 26082 45120 26090 45184
rect 21219 44844 21285 44845
rect 21219 44780 21220 44844
rect 21284 44780 21285 44844
rect 21219 44779 21285 44780
rect 20805 44576 20813 44640
rect 20877 44576 20893 44640
rect 20957 44576 20973 44640
rect 21037 44576 21053 44640
rect 21117 44576 21125 44640
rect 20805 43552 21125 44576
rect 20805 43488 20813 43552
rect 20877 43488 20893 43552
rect 20957 43488 20973 43552
rect 21037 43488 21053 43552
rect 21117 43488 21125 43552
rect 20805 42464 21125 43488
rect 20805 42400 20813 42464
rect 20877 42400 20893 42464
rect 20957 42400 20973 42464
rect 21037 42400 21053 42464
rect 21117 42400 21125 42464
rect 20805 41376 21125 42400
rect 20805 41312 20813 41376
rect 20877 41312 20893 41376
rect 20957 41312 20973 41376
rect 21037 41312 21053 41376
rect 21117 41312 21125 41376
rect 20805 40288 21125 41312
rect 21222 40629 21282 44779
rect 25770 44096 26090 45120
rect 25770 44032 25778 44096
rect 25842 44032 25858 44096
rect 25922 44032 25938 44096
rect 26002 44032 26018 44096
rect 26082 44032 26090 44096
rect 25770 43008 26090 44032
rect 25770 42944 25778 43008
rect 25842 42944 25858 43008
rect 25922 42944 25938 43008
rect 26002 42944 26018 43008
rect 26082 42944 26090 43008
rect 25770 41920 26090 42944
rect 25770 41856 25778 41920
rect 25842 41856 25858 41920
rect 25922 41856 25938 41920
rect 26002 41856 26018 41920
rect 26082 41856 26090 41920
rect 25770 40832 26090 41856
rect 25770 40768 25778 40832
rect 25842 40768 25858 40832
rect 25922 40768 25938 40832
rect 26002 40768 26018 40832
rect 26082 40768 26090 40832
rect 21219 40628 21285 40629
rect 21219 40564 21220 40628
rect 21284 40564 21285 40628
rect 21219 40563 21285 40564
rect 20805 40224 20813 40288
rect 20877 40224 20893 40288
rect 20957 40224 20973 40288
rect 21037 40224 21053 40288
rect 21117 40224 21125 40288
rect 20805 39200 21125 40224
rect 20805 39136 20813 39200
rect 20877 39136 20893 39200
rect 20957 39136 20973 39200
rect 21037 39136 21053 39200
rect 21117 39136 21125 39200
rect 20805 38112 21125 39136
rect 20805 38048 20813 38112
rect 20877 38048 20893 38112
rect 20957 38048 20973 38112
rect 21037 38048 21053 38112
rect 21117 38048 21125 38112
rect 20805 37024 21125 38048
rect 20805 36960 20813 37024
rect 20877 36960 20893 37024
rect 20957 36960 20973 37024
rect 21037 36960 21053 37024
rect 21117 36960 21125 37024
rect 18643 36276 18709 36277
rect 18643 36212 18644 36276
rect 18708 36212 18709 36276
rect 18643 36211 18709 36212
rect 15839 35328 15848 35392
rect 15912 35328 15928 35392
rect 15992 35328 16008 35392
rect 16072 35328 16088 35392
rect 16152 35328 16160 35392
rect 15839 34304 16160 35328
rect 17355 34644 17421 34645
rect 17355 34580 17356 34644
rect 17420 34580 17421 34644
rect 17355 34579 17421 34580
rect 15839 34240 15848 34304
rect 15912 34240 15928 34304
rect 15992 34240 16008 34304
rect 16072 34240 16088 34304
rect 16152 34240 16160 34304
rect 15839 33216 16160 34240
rect 16619 33964 16685 33965
rect 16619 33900 16620 33964
rect 16684 33900 16685 33964
rect 16619 33899 16685 33900
rect 15839 33152 15848 33216
rect 15912 33152 15928 33216
rect 15992 33152 16008 33216
rect 16072 33152 16088 33216
rect 16152 33152 16160 33216
rect 15839 32128 16160 33152
rect 15839 32064 15848 32128
rect 15912 32064 15928 32128
rect 15992 32064 16008 32128
rect 16072 32064 16088 32128
rect 16152 32064 16160 32128
rect 15839 31040 16160 32064
rect 15839 30976 15848 31040
rect 15912 30976 15928 31040
rect 15992 30976 16008 31040
rect 16072 30976 16088 31040
rect 16152 30976 16160 31040
rect 15839 29952 16160 30976
rect 16622 30837 16682 33899
rect 16987 30972 17053 30973
rect 16987 30908 16988 30972
rect 17052 30908 17053 30972
rect 16987 30907 17053 30908
rect 16619 30836 16685 30837
rect 16619 30772 16620 30836
rect 16684 30772 16685 30836
rect 16619 30771 16685 30772
rect 15839 29888 15848 29952
rect 15912 29888 15928 29952
rect 15992 29888 16008 29952
rect 16072 29888 16088 29952
rect 16152 29888 16160 29952
rect 15839 28864 16160 29888
rect 15839 28800 15848 28864
rect 15912 28800 15928 28864
rect 15992 28800 16008 28864
rect 16072 28800 16088 28864
rect 16152 28800 16160 28864
rect 15839 27776 16160 28800
rect 15839 27712 15848 27776
rect 15912 27712 15928 27776
rect 15992 27712 16008 27776
rect 16072 27712 16088 27776
rect 16152 27712 16160 27776
rect 15839 26688 16160 27712
rect 15839 26624 15848 26688
rect 15912 26624 15928 26688
rect 15992 26624 16008 26688
rect 16072 26624 16088 26688
rect 16152 26624 16160 26688
rect 15839 25600 16160 26624
rect 15839 25536 15848 25600
rect 15912 25536 15928 25600
rect 15992 25536 16008 25600
rect 16072 25536 16088 25600
rect 16152 25536 16160 25600
rect 15839 24512 16160 25536
rect 15839 24448 15848 24512
rect 15912 24448 15928 24512
rect 15992 24448 16008 24512
rect 16072 24448 16088 24512
rect 16152 24448 16160 24512
rect 15839 23424 16160 24448
rect 16990 23629 17050 30907
rect 16987 23628 17053 23629
rect 16987 23564 16988 23628
rect 17052 23564 17053 23628
rect 16987 23563 17053 23564
rect 15839 23360 15848 23424
rect 15912 23360 15928 23424
rect 15992 23360 16008 23424
rect 16072 23360 16088 23424
rect 16152 23360 16160 23424
rect 15839 22336 16160 23360
rect 16990 22405 17050 23563
rect 16987 22404 17053 22405
rect 16987 22340 16988 22404
rect 17052 22340 17053 22404
rect 16987 22339 17053 22340
rect 15839 22272 15848 22336
rect 15912 22272 15928 22336
rect 15992 22272 16008 22336
rect 16072 22272 16088 22336
rect 16152 22272 16160 22336
rect 15839 21248 16160 22272
rect 17358 21589 17418 34579
rect 17539 31924 17605 31925
rect 17539 31860 17540 31924
rect 17604 31860 17605 31924
rect 17539 31859 17605 31860
rect 17542 30157 17602 31859
rect 18646 30565 18706 36211
rect 20805 35936 21125 36960
rect 20805 35872 20813 35936
rect 20877 35872 20893 35936
rect 20957 35872 20973 35936
rect 21037 35872 21053 35936
rect 21117 35872 21125 35936
rect 19011 35052 19077 35053
rect 19011 34988 19012 35052
rect 19076 34988 19077 35052
rect 19011 34987 19077 34988
rect 19014 33829 19074 34987
rect 20805 34848 21125 35872
rect 20805 34784 20813 34848
rect 20877 34784 20893 34848
rect 20957 34784 20973 34848
rect 21037 34784 21053 34848
rect 21117 34784 21125 34848
rect 19011 33828 19077 33829
rect 19011 33764 19012 33828
rect 19076 33764 19077 33828
rect 19011 33763 19077 33764
rect 20805 33760 21125 34784
rect 20805 33696 20813 33760
rect 20877 33696 20893 33760
rect 20957 33696 20973 33760
rect 21037 33696 21053 33760
rect 21117 33696 21125 33760
rect 20805 32672 21125 33696
rect 20805 32608 20813 32672
rect 20877 32608 20893 32672
rect 20957 32608 20973 32672
rect 21037 32608 21053 32672
rect 21117 32608 21125 32672
rect 20805 31584 21125 32608
rect 20805 31520 20813 31584
rect 20877 31520 20893 31584
rect 20957 31520 20973 31584
rect 21037 31520 21053 31584
rect 21117 31520 21125 31584
rect 19195 30700 19261 30701
rect 19195 30636 19196 30700
rect 19260 30636 19261 30700
rect 19195 30635 19261 30636
rect 18643 30564 18709 30565
rect 18643 30500 18644 30564
rect 18708 30500 18709 30564
rect 18643 30499 18709 30500
rect 17539 30156 17605 30157
rect 17539 30092 17540 30156
rect 17604 30092 17605 30156
rect 17539 30091 17605 30092
rect 19011 28660 19077 28661
rect 19011 28596 19012 28660
rect 19076 28596 19077 28660
rect 19011 28595 19077 28596
rect 18643 28116 18709 28117
rect 18643 28052 18644 28116
rect 18708 28052 18709 28116
rect 18643 28051 18709 28052
rect 18646 27709 18706 28051
rect 18643 27708 18709 27709
rect 18643 27644 18644 27708
rect 18708 27644 18709 27708
rect 18643 27643 18709 27644
rect 19014 27165 19074 28595
rect 19011 27164 19077 27165
rect 19011 27100 19012 27164
rect 19076 27100 19077 27164
rect 19011 27099 19077 27100
rect 17355 21588 17421 21589
rect 17355 21524 17356 21588
rect 17420 21524 17421 21588
rect 17355 21523 17421 21524
rect 15839 21184 15848 21248
rect 15912 21184 15928 21248
rect 15992 21184 16008 21248
rect 16072 21184 16088 21248
rect 16152 21184 16160 21248
rect 15839 20160 16160 21184
rect 19198 20637 19258 30635
rect 20805 30496 21125 31520
rect 20805 30432 20813 30496
rect 20877 30432 20893 30496
rect 20957 30432 20973 30496
rect 21037 30432 21053 30496
rect 21117 30432 21125 30496
rect 20805 29408 21125 30432
rect 20805 29344 20813 29408
rect 20877 29344 20893 29408
rect 20957 29344 20973 29408
rect 21037 29344 21053 29408
rect 21117 29344 21125 29408
rect 20805 28320 21125 29344
rect 20805 28256 20813 28320
rect 20877 28256 20893 28320
rect 20957 28256 20973 28320
rect 21037 28256 21053 28320
rect 21117 28256 21125 28320
rect 20805 27232 21125 28256
rect 20805 27168 20813 27232
rect 20877 27168 20893 27232
rect 20957 27168 20973 27232
rect 21037 27168 21053 27232
rect 21117 27168 21125 27232
rect 20805 26144 21125 27168
rect 20805 26080 20813 26144
rect 20877 26080 20893 26144
rect 20957 26080 20973 26144
rect 21037 26080 21053 26144
rect 21117 26080 21125 26144
rect 20805 25056 21125 26080
rect 20805 24992 20813 25056
rect 20877 24992 20893 25056
rect 20957 24992 20973 25056
rect 21037 24992 21053 25056
rect 21117 24992 21125 25056
rect 20805 23968 21125 24992
rect 20805 23904 20813 23968
rect 20877 23904 20893 23968
rect 20957 23904 20973 23968
rect 21037 23904 21053 23968
rect 21117 23904 21125 23968
rect 20805 22880 21125 23904
rect 20805 22816 20813 22880
rect 20877 22816 20893 22880
rect 20957 22816 20973 22880
rect 21037 22816 21053 22880
rect 21117 22816 21125 22880
rect 20805 21792 21125 22816
rect 20805 21728 20813 21792
rect 20877 21728 20893 21792
rect 20957 21728 20973 21792
rect 21037 21728 21053 21792
rect 21117 21728 21125 21792
rect 20805 20704 21125 21728
rect 20805 20640 20813 20704
rect 20877 20640 20893 20704
rect 20957 20640 20973 20704
rect 21037 20640 21053 20704
rect 21117 20640 21125 20704
rect 19195 20636 19261 20637
rect 19195 20572 19196 20636
rect 19260 20572 19261 20636
rect 19195 20571 19261 20572
rect 15839 20096 15848 20160
rect 15912 20096 15928 20160
rect 15992 20096 16008 20160
rect 16072 20096 16088 20160
rect 16152 20096 16160 20160
rect 15839 19072 16160 20096
rect 15839 19008 15848 19072
rect 15912 19008 15928 19072
rect 15992 19008 16008 19072
rect 16072 19008 16088 19072
rect 16152 19008 16160 19072
rect 15839 17984 16160 19008
rect 15839 17920 15848 17984
rect 15912 17920 15928 17984
rect 15992 17920 16008 17984
rect 16072 17920 16088 17984
rect 16152 17920 16160 17984
rect 15839 16896 16160 17920
rect 15839 16832 15848 16896
rect 15912 16832 15928 16896
rect 15992 16832 16008 16896
rect 16072 16832 16088 16896
rect 16152 16832 16160 16896
rect 15839 15808 16160 16832
rect 15839 15744 15848 15808
rect 15912 15744 15928 15808
rect 15992 15744 16008 15808
rect 16072 15744 16088 15808
rect 16152 15744 16160 15808
rect 15839 14720 16160 15744
rect 15839 14656 15848 14720
rect 15912 14656 15928 14720
rect 15992 14656 16008 14720
rect 16072 14656 16088 14720
rect 16152 14656 16160 14720
rect 15839 13632 16160 14656
rect 15839 13568 15848 13632
rect 15912 13568 15928 13632
rect 15992 13568 16008 13632
rect 16072 13568 16088 13632
rect 16152 13568 16160 13632
rect 15839 12544 16160 13568
rect 20805 19616 21125 20640
rect 20805 19552 20813 19616
rect 20877 19552 20893 19616
rect 20957 19552 20973 19616
rect 21037 19552 21053 19616
rect 21117 19552 21125 19616
rect 20805 18528 21125 19552
rect 20805 18464 20813 18528
rect 20877 18464 20893 18528
rect 20957 18464 20973 18528
rect 21037 18464 21053 18528
rect 21117 18464 21125 18528
rect 20805 17440 21125 18464
rect 20805 17376 20813 17440
rect 20877 17376 20893 17440
rect 20957 17376 20973 17440
rect 21037 17376 21053 17440
rect 21117 17376 21125 17440
rect 20805 16352 21125 17376
rect 20805 16288 20813 16352
rect 20877 16288 20893 16352
rect 20957 16288 20973 16352
rect 21037 16288 21053 16352
rect 21117 16288 21125 16352
rect 20805 15264 21125 16288
rect 20805 15200 20813 15264
rect 20877 15200 20893 15264
rect 20957 15200 20973 15264
rect 21037 15200 21053 15264
rect 21117 15200 21125 15264
rect 20805 14176 21125 15200
rect 25770 39744 26090 40768
rect 25770 39680 25778 39744
rect 25842 39680 25858 39744
rect 25922 39680 25938 39744
rect 26002 39680 26018 39744
rect 26082 39680 26090 39744
rect 25770 38656 26090 39680
rect 25770 38592 25778 38656
rect 25842 38592 25858 38656
rect 25922 38592 25938 38656
rect 26002 38592 26018 38656
rect 26082 38592 26090 38656
rect 25770 37568 26090 38592
rect 25770 37504 25778 37568
rect 25842 37504 25858 37568
rect 25922 37504 25938 37568
rect 26002 37504 26018 37568
rect 26082 37504 26090 37568
rect 25770 36480 26090 37504
rect 25770 36416 25778 36480
rect 25842 36416 25858 36480
rect 25922 36416 25938 36480
rect 26002 36416 26018 36480
rect 26082 36416 26090 36480
rect 25770 35392 26090 36416
rect 25770 35328 25778 35392
rect 25842 35328 25858 35392
rect 25922 35328 25938 35392
rect 26002 35328 26018 35392
rect 26082 35328 26090 35392
rect 25770 34304 26090 35328
rect 25770 34240 25778 34304
rect 25842 34240 25858 34304
rect 25922 34240 25938 34304
rect 26002 34240 26018 34304
rect 26082 34240 26090 34304
rect 25770 33216 26090 34240
rect 25770 33152 25778 33216
rect 25842 33152 25858 33216
rect 25922 33152 25938 33216
rect 26002 33152 26018 33216
rect 26082 33152 26090 33216
rect 25770 32128 26090 33152
rect 25770 32064 25778 32128
rect 25842 32064 25858 32128
rect 25922 32064 25938 32128
rect 26002 32064 26018 32128
rect 26082 32064 26090 32128
rect 25770 31040 26090 32064
rect 25770 30976 25778 31040
rect 25842 30976 25858 31040
rect 25922 30976 25938 31040
rect 26002 30976 26018 31040
rect 26082 30976 26090 31040
rect 25770 29952 26090 30976
rect 25770 29888 25778 29952
rect 25842 29888 25858 29952
rect 25922 29888 25938 29952
rect 26002 29888 26018 29952
rect 26082 29888 26090 29952
rect 25770 28864 26090 29888
rect 25770 28800 25778 28864
rect 25842 28800 25858 28864
rect 25922 28800 25938 28864
rect 26002 28800 26018 28864
rect 26082 28800 26090 28864
rect 25770 27776 26090 28800
rect 25770 27712 25778 27776
rect 25842 27712 25858 27776
rect 25922 27712 25938 27776
rect 26002 27712 26018 27776
rect 26082 27712 26090 27776
rect 25770 26688 26090 27712
rect 25770 26624 25778 26688
rect 25842 26624 25858 26688
rect 25922 26624 25938 26688
rect 26002 26624 26018 26688
rect 26082 26624 26090 26688
rect 25770 25600 26090 26624
rect 25770 25536 25778 25600
rect 25842 25536 25858 25600
rect 25922 25536 25938 25600
rect 26002 25536 26018 25600
rect 26082 25536 26090 25600
rect 25770 24512 26090 25536
rect 25770 24448 25778 24512
rect 25842 24448 25858 24512
rect 25922 24448 25938 24512
rect 26002 24448 26018 24512
rect 26082 24448 26090 24512
rect 25770 23424 26090 24448
rect 25770 23360 25778 23424
rect 25842 23360 25858 23424
rect 25922 23360 25938 23424
rect 26002 23360 26018 23424
rect 26082 23360 26090 23424
rect 25770 22336 26090 23360
rect 25770 22272 25778 22336
rect 25842 22272 25858 22336
rect 25922 22272 25938 22336
rect 26002 22272 26018 22336
rect 26082 22272 26090 22336
rect 25770 21248 26090 22272
rect 25770 21184 25778 21248
rect 25842 21184 25858 21248
rect 25922 21184 25938 21248
rect 26002 21184 26018 21248
rect 26082 21184 26090 21248
rect 25770 20160 26090 21184
rect 25770 20096 25778 20160
rect 25842 20096 25858 20160
rect 25922 20096 25938 20160
rect 26002 20096 26018 20160
rect 26082 20096 26090 20160
rect 25770 19072 26090 20096
rect 25770 19008 25778 19072
rect 25842 19008 25858 19072
rect 25922 19008 25938 19072
rect 26002 19008 26018 19072
rect 26082 19008 26090 19072
rect 25770 17984 26090 19008
rect 25770 17920 25778 17984
rect 25842 17920 25858 17984
rect 25922 17920 25938 17984
rect 26002 17920 26018 17984
rect 26082 17920 26090 17984
rect 25770 16896 26090 17920
rect 25770 16832 25778 16896
rect 25842 16832 25858 16896
rect 25922 16832 25938 16896
rect 26002 16832 26018 16896
rect 26082 16832 26090 16896
rect 25770 15808 26090 16832
rect 25770 15744 25778 15808
rect 25842 15744 25858 15808
rect 25922 15744 25938 15808
rect 26002 15744 26018 15808
rect 26082 15744 26090 15808
rect 25770 14720 26090 15744
rect 25770 14656 25778 14720
rect 25842 14656 25858 14720
rect 25922 14656 25938 14720
rect 26002 14656 26018 14720
rect 26082 14656 26090 14720
rect 21403 14380 21469 14381
rect 21403 14316 21404 14380
rect 21468 14316 21469 14380
rect 21403 14315 21469 14316
rect 20805 14112 20813 14176
rect 20877 14112 20893 14176
rect 20957 14112 20973 14176
rect 21037 14112 21053 14176
rect 21117 14112 21125 14176
rect 20805 13088 21125 14112
rect 20805 13024 20813 13088
rect 20877 13024 20893 13088
rect 20957 13024 20973 13088
rect 21037 13024 21053 13088
rect 21117 13024 21125 13088
rect 20483 12612 20549 12613
rect 20483 12548 20484 12612
rect 20548 12548 20549 12612
rect 20483 12547 20549 12548
rect 15839 12480 15848 12544
rect 15912 12480 15928 12544
rect 15992 12480 16008 12544
rect 16072 12480 16088 12544
rect 16152 12480 16160 12544
rect 15839 11456 16160 12480
rect 15839 11392 15848 11456
rect 15912 11392 15928 11456
rect 15992 11392 16008 11456
rect 16072 11392 16088 11456
rect 16152 11392 16160 11456
rect 15839 10368 16160 11392
rect 20486 10709 20546 12547
rect 20805 12000 21125 13024
rect 20805 11936 20813 12000
rect 20877 11936 20893 12000
rect 20957 11936 20973 12000
rect 21037 11936 21053 12000
rect 21117 11936 21125 12000
rect 20805 10912 21125 11936
rect 21406 11117 21466 14315
rect 25770 13632 26090 14656
rect 25770 13568 25778 13632
rect 25842 13568 25858 13632
rect 25922 13568 25938 13632
rect 26002 13568 26018 13632
rect 26082 13568 26090 13632
rect 25770 12544 26090 13568
rect 25770 12480 25778 12544
rect 25842 12480 25858 12544
rect 25922 12480 25938 12544
rect 26002 12480 26018 12544
rect 26082 12480 26090 12544
rect 25770 11456 26090 12480
rect 25770 11392 25778 11456
rect 25842 11392 25858 11456
rect 25922 11392 25938 11456
rect 26002 11392 26018 11456
rect 26082 11392 26090 11456
rect 21403 11116 21469 11117
rect 21403 11052 21404 11116
rect 21468 11052 21469 11116
rect 21403 11051 21469 11052
rect 20805 10848 20813 10912
rect 20877 10848 20893 10912
rect 20957 10848 20973 10912
rect 21037 10848 21053 10912
rect 21117 10848 21125 10912
rect 20483 10708 20549 10709
rect 20483 10644 20484 10708
rect 20548 10644 20549 10708
rect 20483 10643 20549 10644
rect 15839 10304 15848 10368
rect 15912 10304 15928 10368
rect 15992 10304 16008 10368
rect 16072 10304 16088 10368
rect 16152 10304 16160 10368
rect 15839 9280 16160 10304
rect 15839 9216 15848 9280
rect 15912 9216 15928 9280
rect 15992 9216 16008 9280
rect 16072 9216 16088 9280
rect 16152 9216 16160 9280
rect 15839 8192 16160 9216
rect 15839 8128 15848 8192
rect 15912 8128 15928 8192
rect 15992 8128 16008 8192
rect 16072 8128 16088 8192
rect 16152 8128 16160 8192
rect 15839 7104 16160 8128
rect 15839 7040 15848 7104
rect 15912 7040 15928 7104
rect 15992 7040 16008 7104
rect 16072 7040 16088 7104
rect 16152 7040 16160 7104
rect 15839 6016 16160 7040
rect 15839 5952 15848 6016
rect 15912 5952 15928 6016
rect 15992 5952 16008 6016
rect 16072 5952 16088 6016
rect 16152 5952 16160 6016
rect 15839 4928 16160 5952
rect 15839 4864 15848 4928
rect 15912 4864 15928 4928
rect 15992 4864 16008 4928
rect 16072 4864 16088 4928
rect 16152 4864 16160 4928
rect 15839 3840 16160 4864
rect 15839 3776 15848 3840
rect 15912 3776 15928 3840
rect 15992 3776 16008 3840
rect 16072 3776 16088 3840
rect 16152 3776 16160 3840
rect 15839 2752 16160 3776
rect 15839 2688 15848 2752
rect 15912 2688 15928 2752
rect 15992 2688 16008 2752
rect 16072 2688 16088 2752
rect 16152 2688 16160 2752
rect 15839 2128 16160 2688
rect 20805 9824 21125 10848
rect 20805 9760 20813 9824
rect 20877 9760 20893 9824
rect 20957 9760 20973 9824
rect 21037 9760 21053 9824
rect 21117 9760 21125 9824
rect 20805 8736 21125 9760
rect 20805 8672 20813 8736
rect 20877 8672 20893 8736
rect 20957 8672 20973 8736
rect 21037 8672 21053 8736
rect 21117 8672 21125 8736
rect 20805 7648 21125 8672
rect 20805 7584 20813 7648
rect 20877 7584 20893 7648
rect 20957 7584 20973 7648
rect 21037 7584 21053 7648
rect 21117 7584 21125 7648
rect 20805 6560 21125 7584
rect 20805 6496 20813 6560
rect 20877 6496 20893 6560
rect 20957 6496 20973 6560
rect 21037 6496 21053 6560
rect 21117 6496 21125 6560
rect 20805 5472 21125 6496
rect 20805 5408 20813 5472
rect 20877 5408 20893 5472
rect 20957 5408 20973 5472
rect 21037 5408 21053 5472
rect 21117 5408 21125 5472
rect 20805 4384 21125 5408
rect 20805 4320 20813 4384
rect 20877 4320 20893 4384
rect 20957 4320 20973 4384
rect 21037 4320 21053 4384
rect 21117 4320 21125 4384
rect 20805 3296 21125 4320
rect 20805 3232 20813 3296
rect 20877 3232 20893 3296
rect 20957 3232 20973 3296
rect 21037 3232 21053 3296
rect 21117 3232 21125 3296
rect 20805 2208 21125 3232
rect 20805 2144 20813 2208
rect 20877 2144 20893 2208
rect 20957 2144 20973 2208
rect 21037 2144 21053 2208
rect 21117 2144 21125 2208
rect 20805 2128 21125 2144
rect 25770 10368 26090 11392
rect 25770 10304 25778 10368
rect 25842 10304 25858 10368
rect 25922 10304 25938 10368
rect 26002 10304 26018 10368
rect 26082 10304 26090 10368
rect 25770 9280 26090 10304
rect 25770 9216 25778 9280
rect 25842 9216 25858 9280
rect 25922 9216 25938 9280
rect 26002 9216 26018 9280
rect 26082 9216 26090 9280
rect 25770 8192 26090 9216
rect 25770 8128 25778 8192
rect 25842 8128 25858 8192
rect 25922 8128 25938 8192
rect 26002 8128 26018 8192
rect 26082 8128 26090 8192
rect 25770 7104 26090 8128
rect 25770 7040 25778 7104
rect 25842 7040 25858 7104
rect 25922 7040 25938 7104
rect 26002 7040 26018 7104
rect 26082 7040 26090 7104
rect 25770 6016 26090 7040
rect 25770 5952 25778 6016
rect 25842 5952 25858 6016
rect 25922 5952 25938 6016
rect 26002 5952 26018 6016
rect 26082 5952 26090 6016
rect 25770 4928 26090 5952
rect 25770 4864 25778 4928
rect 25842 4864 25858 4928
rect 25922 4864 25938 4928
rect 26002 4864 26018 4928
rect 26082 4864 26090 4928
rect 25770 3840 26090 4864
rect 25770 3776 25778 3840
rect 25842 3776 25858 3840
rect 25922 3776 25938 3840
rect 26002 3776 26018 3840
rect 26082 3776 26090 3840
rect 25770 2752 26090 3776
rect 25770 2688 25778 2752
rect 25842 2688 25858 2752
rect 25922 2688 25938 2752
rect 26002 2688 26018 2752
rect 26082 2688 26090 2752
rect 25770 2128 26090 2688
use sky130_fd_sc_hd__decap_8  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_19
timestamp 1635444444
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_7
timestamp 1635444444
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635444444
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1635444444
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1635444444
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1635444444
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_31
timestamp 1635444444
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_43
timestamp 1635444444
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1635444444
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1635444444
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1635444444
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1635444444
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1635444444
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1635444444
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1635444444
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1635444444
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1635444444
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1635444444
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1635444444
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1635444444
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1635444444
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1635444444
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1635444444
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1635444444
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp 1635444444
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1635444444
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1635444444
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1635444444
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1615_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 12880 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _1815_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1635444444
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1635444444
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_144
timestamp 1635444444
transform 1 0 14352 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_134
timestamp 1635444444
transform 1 0 13432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_142
timestamp 1635444444
transform 1 0 14168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1635444444
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1571_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1823_
timestamp 1635444444
transform 1 0 14260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1635444444
transform 1 0 15456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1635444444
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1635444444
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1635444444
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1635444444
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1635444444
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1635444444
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1635444444
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1635444444
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1635444444
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1635444444
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1635444444
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1635444444
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1635444444
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1635444444
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1635444444
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1635444444
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1635444444
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1635444444
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1635444444
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1635444444
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1635444444
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1635444444
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1635444444
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1635444444
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1635444444
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1635444444
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1635444444
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1635444444
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1635444444
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1635444444
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1635444444
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1635444444
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1635444444
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1635444444
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293
timestamp 1635444444
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_299
timestamp 1635444444
transform 1 0 28612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1635444444
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1635444444
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_305
timestamp 1635444444
transform 1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1635444444
transform 1 0 28704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_309
timestamp 1635444444
transform 1 0 29532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_316
timestamp 1635444444
transform 1 0 30176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_309
timestamp 1635444444
transform 1 0 29532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_316
timestamp 1635444444
transform 1 0 30176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635444444
transform -1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635444444
transform -1 0 30820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1635444444
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 29624 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input67
timestamp 1635444444
transform 1 0 29624 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1635444444
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1635444444
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635444444
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1635444444
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1635444444
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1635444444
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1635444444
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1635444444
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1635444444
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1635444444
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1635444444
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1635444444
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1635444444
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1635444444
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_105
timestamp 1635444444
transform 1 0 10764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1635444444
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 10488 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1814_
timestamp 1635444444
transform 1 0 11132 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp 1635444444
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1635444444
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1635444444
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1822_
timestamp 1635444444
transform 1 0 14352 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1635444444
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1635444444
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1635444444
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1635444444
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1635444444
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1635444444
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1635444444
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1635444444
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1635444444
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1635444444
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1635444444
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1635444444
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1635444444
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1635444444
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1635444444
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1635444444
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1635444444
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1635444444
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_309
timestamp 1635444444
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_316
timestamp 1635444444
transform 1 0 30176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635444444
transform -1 0 30820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1635444444
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1635444444
transform 1 0 29808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1635444444
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1635444444
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635444444
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1635444444
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1635444444
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1635444444
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1635444444
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1635444444
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1635444444
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1635444444
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1635444444
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1635444444
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1635444444
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1635444444
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_116
timestamp 1635444444
transform 1 0 11776 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1635444444
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1635444444
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1616_
timestamp 1635444444
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _1617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 12972 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1632_
timestamp 1635444444
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_138
timestamp 1635444444
transform 1 0 13800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_149
timestamp 1635444444
transform 1 0 14812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _1572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14168 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_3_156
timestamp 1635444444
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1635444444
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 15180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1810_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_178
timestamp 1635444444
transform 1 0 17480 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1874_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 18216 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_3_203
timestamp 1635444444
transform 1 0 19780 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1635444444
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1635444444
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1635444444
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1635444444
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1635444444
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1635444444
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1635444444
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1635444444
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1635444444
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1635444444
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1635444444
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1635444444
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_305
timestamp 1635444444
transform 1 0 29164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_311
timestamp 1635444444
transform 1 0 29716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_316
timestamp 1635444444
transform 1 0 30176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635444444
transform -1 0 30820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1635444444
transform 1 0 29808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1635444444
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1635444444
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635444444
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1635444444
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1635444444
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1635444444
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1635444444
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1635444444
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1635444444
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1635444444
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1635444444
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1635444444
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1635444444
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1635444444
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1635444444
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_121
timestamp 1635444444
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_125
timestamp 1635444444
transform 1 0 12604 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1736_
timestamp 1635444444
transform 1 0 12696 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1635444444
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1635444444
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_147
timestamp 1635444444
transform 1 0 14628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1635444444
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1593_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_154
timestamp 1635444444
transform 1 0 15272 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_162
timestamp 1635444444
transform 1 0 16008 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1875_
timestamp 1635444444
transform 1 0 16100 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_4_180
timestamp 1635444444
transform 1 0 17664 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1635444444
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1635444444
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_197
timestamp 1635444444
transform 1 0 19228 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 19964 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_221
timestamp 1635444444
transform 1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1635444444
transform 1 0 21804 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1635444444
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1635444444
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1635444444
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_261
timestamp 1635444444
transform 1 0 25116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1635444444
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_273
timestamp 1635444444
transform 1 0 26220 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _1170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 25392 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_285
timestamp 1635444444
transform 1 0 27324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_297
timestamp 1635444444
transform 1 0 28428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1635444444
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_309
timestamp 1635444444
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_316
timestamp 1635444444
transform 1 0 30176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635444444
transform -1 0 30820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1635444444
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 29808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_19
timestamp 1635444444
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_7
timestamp 1635444444
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635444444
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1635444444
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_31
timestamp 1635444444
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_43
timestamp 1635444444
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1635444444
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1635444444
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1635444444
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1635444444
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1635444444
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1635444444
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1635444444
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1635444444
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_118
timestamp 1635444444
transform 1 0 11960 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_126
timestamp 1635444444
transform 1 0 12696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1635444444
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1611_
timestamp 1635444444
transform 1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 11500 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1635444444
transform 1 0 13248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_141
timestamp 1635444444
transform 1 0 14076 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1594_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14812 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1610_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 13616 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_5_156
timestamp 1635444444
transform 1 0 15456 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1635444444
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1635444444
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1888_
timestamp 1635444444
transform 1 0 17020 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_5_190
timestamp 1635444444
transform 1 0 18584 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1635444444
transform 1 0 18952 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_5_210
timestamp 1635444444
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1635444444
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_234
timestamp 1635444444
transform 1 0 22632 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1635444444
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1309_
timestamp 1635444444
transform 1 0 21804 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_246
timestamp 1635444444
transform 1 0 23736 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_258
timestamp 1635444444
transform 1 0 24840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1169_
timestamp 1635444444
transform 1 0 25024 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1635444444
transform 1 0 25852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 1635444444
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1635444444
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1635444444
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1635444444
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_305
timestamp 1635444444
transform 1 0 29164 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_311
timestamp 1635444444
transform 1 0 29716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_316
timestamp 1635444444
transform 1 0 30176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635444444
transform -1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1635444444
transform 1 0 29808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1635444444
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1635444444
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1635444444
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1635444444
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635444444
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635444444
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1635444444
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1635444444
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1635444444
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1635444444
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1635444444
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1635444444
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1635444444
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1635444444
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1635444444
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1635444444
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1635444444
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1635444444
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1635444444
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1635444444
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1635444444
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1635444444
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1635444444
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1635444444
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1635444444
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1635444444
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1635444444
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1635444444
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1614_
timestamp 1635444444
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1819_
timestamp 1635444444
transform 1 0 10580 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_6_124
timestamp 1635444444
transform 1 0 12512 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1635444444
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1635444444
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp 1635444444
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_127
timestamp 1635444444
transform 1 0 12788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1635444444
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1547_
timestamp 1635444444
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1778_
timestamp 1635444444
transform 1 0 11960 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1635444444
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_134
timestamp 1635444444
transform 1 0 13432 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_140
timestamp 1635444444
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1635444444
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1612_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 13248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1816_
timestamp 1635444444
transform 1 0 14076 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1817_
timestamp 1635444444
transform 1 0 14076 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_6_162
timestamp 1635444444
transform 1 0 16008 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_169
timestamp 1635444444
transform 1 0 16652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1635444444
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp 1635444444
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1635444444
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1210_
timestamp 1635444444
transform 1 0 16376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_181
timestamp 1635444444
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1635444444
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_185
timestamp 1635444444
transform 1 0 18124 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1635444444
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 17388 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1206_
timestamp 1635444444
transform 1 0 18676 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1635444444
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_206
timestamp 1635444444
transform 1 0 20056 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_200
timestamp 1635444444
transform 1 0 19504 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_208
timestamp 1635444444
transform 1 0 20240 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__o31a_1  _1212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 19412 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 20424 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1306_
timestamp 1635444444
transform 1 0 20792 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1635444444
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_235
timestamp 1635444444
transform 1 0 22724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1635444444
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_228
timestamp 1635444444
transform 1 0 22080 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1635444444
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1305_
timestamp 1635444444
transform 1 0 21988 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1417_
timestamp 1635444444
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1635444444
transform 1 0 22448 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1635444444
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1635444444
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_253
timestamp 1635444444
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_261
timestamp 1635444444
transform 1 0 25116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_248
timestamp 1635444444
transform 1 0 23920 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1635444444
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1635444444
transform 1 0 24288 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_279
timestamp 1635444444
transform 1 0 26772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_268
timestamp 1635444444
transform 1 0 25760 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1635444444
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1635444444
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1164_
timestamp 1635444444
transform 1 0 27140 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1635444444
transform 1 0 25300 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1635444444
transform 1 0 27140 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_6_299
timestamp 1635444444
transform 1 0 28612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_292
timestamp 1635444444
transform 1 0 27968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_305
timestamp 1635444444
transform 1 0 29164 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1162_
timestamp 1635444444
transform 1 0 28336 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1635444444
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp 1635444444
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_316
timestamp 1635444444
transform 1 0 30176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_316
timestamp 1635444444
transform 1 0 30176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635444444
transform -1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635444444
transform -1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1635444444
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1635444444
transform 1 0 29808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1635444444
transform 1 0 29900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1635444444
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1635444444
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635444444
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1635444444
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1635444444
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1635444444
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1635444444
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1635444444
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1635444444
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1635444444
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1635444444
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1635444444
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1635444444
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1635444444
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _1820_
timestamp 1635444444
transform 1 0 10580 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_8_124
timestamp 1635444444
transform 1 0 12512 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1551_
timestamp 1635444444
transform 1 0 12880 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1635444444
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1635444444
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1635444444
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1635444444
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_153
timestamp 1635444444
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_165
timestamp 1635444444
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _1211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 16652 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1761_
timestamp 1635444444
transform 1 0 15456 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_176
timestamp 1635444444
transform 1 0 17296 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_182
timestamp 1635444444
transform 1 0 17848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1635444444
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1635444444
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1213_
timestamp 1635444444
transform 1 0 17940 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_197
timestamp 1635444444
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_211
timestamp 1635444444
transform 1 0 20516 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1308_
timestamp 1635444444
transform 1 0 19780 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1635444444
transform 1 0 20884 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_231
timestamp 1635444444
transform 1 0 22356 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1304_
timestamp 1635444444
transform 1 0 22724 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_243
timestamp 1635444444
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1635444444
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_253
timestamp 1635444444
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_261
timestamp 1635444444
transform 1 0 25116 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1635444444
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1168_
timestamp 1635444444
transform 1 0 25208 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_271
timestamp 1635444444
transform 1 0 26036 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1166_
timestamp 1635444444
transform 1 0 26404 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_284
timestamp 1635444444
transform 1 0 27232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1635444444
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1635444444
transform 1 0 27600 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 1635444444
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_316
timestamp 1635444444
transform 1 0 30176 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635444444
transform -1 0 30820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1635444444
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1635444444
transform 1 0 29900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_19
timestamp 1635444444
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_7
timestamp 1635444444
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635444444
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1635444444
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_31
timestamp 1635444444
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1635444444
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1635444444
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1635444444
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1635444444
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1635444444
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1635444444
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1635444444
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1635444444
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1635444444
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1635444444
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1635444444
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1635444444
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1818_
timestamp 1635444444
transform 1 0 12328 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_9_143
timestamp 1635444444
transform 1 0 14260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_150
timestamp 1635444444
transform 1 0 14904 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1552_
timestamp 1635444444
transform 1 0 14628 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1635444444
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp 1635444444
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1635444444
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1887_
timestamp 1635444444
transform 1 0 16744 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_9_187
timestamp 1635444444
transform 1 0 18308 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_195
timestamp 1635444444
transform 1 0 19044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_214
timestamp 1635444444
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1635444444
transform 1 0 19320 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1635444444
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_228
timestamp 1635444444
transform 1 0 22080 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_234
timestamp 1635444444
transform 1 0 22632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1635444444
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1301_
timestamp 1635444444
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1635444444
transform 1 0 22724 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_9_251
timestamp 1635444444
transform 1 0 24196 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_259
timestamp 1635444444
transform 1 0 24932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1171_
timestamp 1635444444
transform 1 0 25024 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_9_270
timestamp 1635444444
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1635444444
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1635444444
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1635444444
transform 1 0 26956 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_297
timestamp 1635444444
transform 1 0 28428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1161_
timestamp 1635444444
transform 1 0 28796 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_310
timestamp 1635444444
transform 1 0 29624 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_318
timestamp 1635444444
transform 1 0 30360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635444444
transform -1 0 30820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1635444444
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1635444444
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635444444
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1635444444
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1635444444
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1635444444
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1635444444
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1635444444
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1635444444
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1635444444
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1635444444
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1635444444
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1635444444
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1635444444
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1635444444
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_126
timestamp 1635444444
transform 1 0 12696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1548_
timestamp 1635444444
transform 1 0 12236 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1550_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1635444444
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_145
timestamp 1635444444
transform 1 0 14444 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1635444444
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1553_
timestamp 1635444444
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_157
timestamp 1635444444
transform 1 0 15548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_161
timestamp 1635444444
transform 1 0 15916 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_165
timestamp 1635444444
transform 1 0 16284 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_173
timestamp 1635444444
transform 1 0 17020 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1577_
timestamp 1635444444
transform 1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_184
timestamp 1635444444
transform 1 0 18032 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1635444444
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1635444444
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1184_
timestamp 1635444444
transform 1 0 17296 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_wb_clk_i
timestamp 1635444444
transform 1 0 18400 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_203
timestamp 1635444444
transform 1 0 19780 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1635444444
transform 1 0 20424 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1208_
timestamp 1635444444
transform 1 0 20148 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1209_
timestamp 1635444444
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1303_
timestamp 1635444444
transform 1 0 20792 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_10_224
timestamp 1635444444
transform 1 0 21712 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_236
timestamp 1635444444
transform 1 0 22816 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1307_
timestamp 1635444444
transform 1 0 22080 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1635444444
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1635444444
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_256
timestamp 1635444444
transform 1 0 24656 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_262
timestamp 1635444444
transform 1 0 25208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1635444444
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1424_
timestamp 1635444444
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1431_
timestamp 1635444444
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_279
timestamp 1635444444
transform 1 0 26772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1635444444
transform 1 0 25300 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_287
timestamp 1635444444
transform 1 0 27508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_297
timestamp 1635444444
transform 1 0 28428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp 1635444444
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1160_
timestamp 1635444444
transform 1 0 27600 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_309
timestamp 1635444444
transform 1 0 29532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_316
timestamp 1635444444
transform 1 0 30176 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635444444
transform -1 0 30820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1635444444
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1635444444
transform 1 0 29900 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1635444444
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1635444444
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635444444
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1635444444
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1635444444
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1635444444
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1635444444
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1635444444
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1635444444
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1635444444
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1635444444
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1635444444
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1635444444
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1619_
timestamp 1635444444
transform 1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1635444444
transform 1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1635444444
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1635444444
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1549_
timestamp 1635444444
transform 1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1618_
timestamp 1635444444
transform 1 0 11500 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_11_137
timestamp 1635444444
transform 1 0 13708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1635444444
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_150
timestamp 1635444444
transform 1 0 14904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1597_
timestamp 1635444444
transform 1 0 14444 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1598_
timestamp 1635444444
transform 1 0 13800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_154
timestamp 1635444444
transform 1 0 15272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1635444444
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_174
timestamp 1635444444
transform 1 0 17112 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1635444444
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1576_
timestamp 1635444444
transform 1 0 16652 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1804_
timestamp 1635444444
transform 1 0 15364 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_182
timestamp 1635444444
transform 1 0 17848 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1635444444
transform 1 0 18032 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_200
timestamp 1635444444
transform 1 0 19504 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_208
timestamp 1635444444
transform 1 0 20240 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_213
timestamp 1635444444
transform 1 0 20700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1203_
timestamp 1635444444
transform 1 0 20332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1635444444
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_229
timestamp 1635444444
transform 1 0 22172 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_235
timestamp 1635444444
transform 1 0 22724 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1635444444
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1172_
timestamp 1635444444
transform 1 0 22816 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_wb_clk_i
timestamp 1635444444
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_245
timestamp 1635444444
transform 1 0 23644 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1635444444
transform 1 0 24012 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_265
timestamp 1635444444
transform 1 0 25484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1635444444
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1635444444
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1163_
timestamp 1635444444
transform 1 0 26956 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_11_291
timestamp 1635444444
transform 1 0 27876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_299
timestamp 1635444444
transform 1 0 28612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1635444444
transform 1 0 28704 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_316
timestamp 1635444444
transform 1 0 30176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635444444
transform -1 0 30820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_19
timestamp 1635444444
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_7
timestamp 1635444444
transform 1 0 1748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635444444
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1635444444
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1635444444
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1635444444
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1635444444
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1635444444
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1635444444
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1635444444
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1635444444
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1635444444
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1635444444
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1635444444
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_105
timestamp 1635444444
transform 1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_97
timestamp 1635444444
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1776_
timestamp 1635444444
transform 1 0 10948 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_116
timestamp 1635444444
transform 1 0 11776 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_124
timestamp 1635444444
transform 1 0 12512 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1633_
timestamp 1635444444
transform 1 0 12788 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp 1635444444
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1635444444
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_151
timestamp 1635444444
transform 1 0 14996 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1635444444
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1759_
timestamp 1635444444
transform 1 0 14168 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_160
timestamp 1635444444
transform 1 0 15824 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_168
timestamp 1635444444
transform 1 0 16560 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_173
timestamp 1635444444
transform 1 0 17020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1635444444
transform 1 0 16744 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1608_
timestamp 1635444444
transform 1 0 15548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1635444444
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1635444444
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1635444444
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1182_
timestamp 1635444444
transform 1 0 17388 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1635444444
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_205
timestamp 1635444444
transform 1 0 19964 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1185_
timestamp 1635444444
transform 1 0 19596 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1274_
timestamp 1635444444
transform 1 0 20700 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_221
timestamp 1635444444
transform 1 0 21436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_225
timestamp 1635444444
transform 1 0 21804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_234
timestamp 1635444444
transform 1 0 22632 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_238
timestamp 1635444444
transform 1 0 23000 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1174_
timestamp 1635444444
transform 1 0 23092 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1269_
timestamp 1635444444
transform 1 0 21896 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1635444444
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_253
timestamp 1635444444
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_261
timestamp 1635444444
transform 1 0 25116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1635444444
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_274
timestamp 1635444444
transform 1 0 26312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_281
timestamp 1635444444
transform 1 0 26956 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1635444444
transform 1 0 26680 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1165_
timestamp 1635444444
transform 1 0 25392 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_12_295
timestamp 1635444444
transform 1 0 28244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_302
timestamp 1635444444
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1155_
timestamp 1635444444
transform 1 0 27324 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1635444444
transform 1 0 28612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_309
timestamp 1635444444
transform 1 0 29532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_316
timestamp 1635444444
transform 1 0 30176 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635444444
transform -1 0 30820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1635444444
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1635444444
transform 1 0 29900 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1635444444
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1635444444
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1635444444
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1635444444
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635444444
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635444444
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1635444444
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1635444444
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1635444444
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1635444444
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1635444444
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1635444444
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1635444444
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1635444444
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1635444444
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1635444444
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1635444444
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1635444444
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1635444444
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1635444444
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1635444444
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1635444444
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1635444444
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1635444444
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1635444444
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_93
timestamp 1635444444
transform 1 0 9660 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1635444444
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1777_
timestamp 1635444444
transform 1 0 10580 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1781_
timestamp 1635444444
transform 1 0 10212 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1635444444
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 1635444444
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_121
timestamp 1635444444
transform 1 0 12236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_112
timestamp 1635444444
transform 1 0 11408 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_120
timestamp 1635444444
transform 1 0 12144 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1635444444
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1635444444
transform 1 0 11960 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1738_
timestamp 1635444444
transform 1 0 12604 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1762_
timestamp 1635444444
transform 1 0 12420 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_13_134
timestamp 1635444444
transform 1 0 13432 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1635444444
transform 1 0 14444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_149
timestamp 1635444444
transform 1 0 14812 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1635444444
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_150
timestamp 1635444444
transform 1 0 14904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1635444444
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1554_
timestamp 1635444444
transform 1 0 13984 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14904 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1779_
timestamp 1635444444
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1630_
timestamp 1635444444
transform 1 0 15272 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1635444444
transform 1 0 15824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_162
timestamp 1635444444
transform 1 0 16008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1635444444
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1635444444
transform 1 0 15456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1207_
timestamp 1635444444
transform 1 0 17112 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1193_
timestamp 1635444444
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1635444444
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_170
timestamp 1635444444
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1635444444
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1635444444
transform 1 0 16652 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_185
timestamp 1635444444
transform 1 0 18124 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_182
timestamp 1635444444
transform 1 0 17848 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1635444444
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1635444444
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1181_
timestamp 1635444444
transform 1 0 18216 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1186_
timestamp 1635444444
transform 1 0 18492 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_197
timestamp 1635444444
transform 1 0 19228 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_203
timestamp 1635444444
transform 1 0 19780 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_213
timestamp 1635444444
transform 1 0 20700 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1635444444
transform 1 0 19872 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1635444444
transform 1 0 19228 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1635444444
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1635444444
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1635444444
transform 1 0 21252 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_229
timestamp 1635444444
transform 1 0 22172 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1635444444
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1273_
timestamp 1635444444
transform 1 0 21344 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1860_
timestamp 1635444444
transform 1 0 21988 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1635444444
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_241
timestamp 1635444444
transform 1 0 23276 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1635444444
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1635444444
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1635444444
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1167_
timestamp 1635444444
transform 1 0 24932 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_2  _1861_
timestamp 1635444444
transform 1 0 23920 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  _1159_
timestamp 1635444444
transform 1 0 26128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_269
timestamp 1635444444
transform 1 0 25852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_271
timestamp 1635444444
transform 1 0 26036 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_265
timestamp 1635444444
transform 1 0 25484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_wb_clk_i
timestamp 1635444444
transform 1 0 26220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1635444444
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_277
timestamp 1635444444
transform 1 0 26588 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1635444444
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1635444444
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1635444444
transform 1 0 27140 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_13_285
timestamp 1635444444
transform 1 0 27324 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_296
timestamp 1635444444
transform 1 0 28336 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_299
timestamp 1635444444
transform 1 0 28612 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1157_
timestamp 1635444444
transform 1 0 27416 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1635444444
transform 1 0 28704 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_316
timestamp 1635444444
transform 1 0 30176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1635444444
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_309
timestamp 1635444444
transform 1 0 29532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_316
timestamp 1635444444
transform 1 0 30176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635444444
transform -1 0 30820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635444444
transform -1 0 30820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1635444444
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1635444444
transform 1 0 29900 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1635444444
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1635444444
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635444444
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1635444444
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1635444444
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1635444444
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1635444444
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1635444444
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1635444444
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1635444444
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1635444444
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1635444444
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_93
timestamp 1635444444
transform 1 0 9660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1621_
timestamp 1635444444
transform 1 0 10396 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1635444444
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_131
timestamp 1635444444
transform 1 0 13156 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1635444444
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1636_
timestamp 1635444444
transform 1 0 11500 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1739_
timestamp 1635444444
transform 1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_143
timestamp 1635444444
transform 1 0 14260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_149
timestamp 1635444444
transform 1 0 14812 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1628_
timestamp 1635444444
transform 1 0 14904 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1635444444
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1635444444
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_172
timestamp 1635444444
transform 1 0 16928 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1635444444
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1607_
timestamp 1635444444
transform 1 0 15548 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1629_
timestamp 1635444444
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_182
timestamp 1635444444
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1635444444
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1187_
timestamp 1635444444
transform 1 0 18216 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1188_
timestamp 1635444444
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_210
timestamp 1635444444
transform 1 0 20424 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1635444444
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1189_
timestamp 1635444444
transform 1 0 19504 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1635444444
transform 1 0 20792 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_228
timestamp 1635444444
transform 1 0 22080 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_240
timestamp 1635444444
transform 1 0 23184 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1635444444
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1408_
timestamp 1635444444
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_248
timestamp 1635444444
transform 1 0 23920 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_259
timestamp 1635444444
transform 1 0 24932 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1173_
timestamp 1635444444
transform 1 0 24012 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_15_265
timestamp 1635444444
transform 1 0 25484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1635444444
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1635444444
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_2  _1700_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 26956 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a22oi_2  _1721_
timestamp 1635444444
transform 1 0 25576 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_15_291
timestamp 1635444444
transform 1 0 27876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_299
timestamp 1635444444
transform 1 0 28612 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1635444444
transform 1 0 28704 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_316
timestamp 1635444444
transform 1 0 30176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635444444
transform -1 0 30820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_14
timestamp 1635444444
transform 1 0 2392 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_7
timestamp 1635444444
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635444444
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1729_
timestamp 1635444444
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1635444444
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1635444444
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1635444444
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1635444444
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1635444444
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1635444444
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1635444444
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1635444444
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1635444444
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1635444444
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1635444444
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_105
timestamp 1635444444
transform 1 0 10764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp 1635444444
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1635444444
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_97
timestamp 1635444444
transform 1 0 10028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1375_
timestamp 1635444444
transform 1 0 9384 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_1  _1622_
timestamp 1635444444
transform 1 0 10120 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_16_120
timestamp 1635444444
transform 1 0 12144 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__o221ai_1  _1637_
timestamp 1635444444
transform 1 0 11500 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_16_132
timestamp 1635444444
transform 1 0 13248 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1635444444
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1635444444
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_156
timestamp 1635444444
transform 1 0 15456 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_160
timestamp 1635444444
transform 1 0 15824 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1635444444
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_173
timestamp 1635444444
transform 1 0 17020 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1567_
timestamp 1635444444
transform 1 0 16744 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1589_
timestamp 1635444444
transform 1 0 15916 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1590_
timestamp 1635444444
transform 1 0 15180 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_185
timestamp 1635444444
transform 1 0 18124 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp 1635444444
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1635444444
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_206
timestamp 1635444444
transform 1 0 20056 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_212
timestamp 1635444444
transform 1 0 20608 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_216
timestamp 1635444444
transform 1 0 20976 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1190_
timestamp 1635444444
transform 1 0 19228 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1191_
timestamp 1635444444
transform 1 0 20700 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_229
timestamp 1635444444
transform 1 0 22172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _1275_
timestamp 1635444444
transform 1 0 21344 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_241
timestamp 1635444444
transform 1 0 23276 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1635444444
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1635444444
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1423_
timestamp 1635444444
transform 1 0 23644 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1635444444
transform 1 0 24380 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_269
timestamp 1635444444
transform 1 0 25852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_273
timestamp 1635444444
transform 1 0 26220 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_2  _1711_
timestamp 1635444444
transform 1 0 26312 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_16_284
timestamp 1635444444
transform 1 0 27232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_291
timestamp 1635444444
transform 1 0 27876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1635444444
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1156_
timestamp 1635444444
transform 1 0 28244 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1635444444
transform 1 0 27600 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_313
timestamp 1635444444
transform 1 0 29900 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_319
timestamp 1635444444
transform 1 0 30452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635444444
transform -1 0 30820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1635444444
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_wb_clk_i
timestamp 1635444444
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1635444444
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1635444444
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635444444
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1635444444
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1635444444
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1635444444
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1635444444
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1635444444
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1635444444
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1635444444
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1635444444
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_100
timestamp 1635444444
transform 1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1635444444
transform 1 0 9660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _1374_
timestamp 1635444444
transform 1 0 9844 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1635444444
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_117
timestamp 1635444444
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_121
timestamp 1635444444
transform 1 0 12236 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_127
timestamp 1635444444
transform 1 0 12788 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_131
timestamp 1635444444
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1635444444
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1626_
timestamp 1635444444
transform 1 0 12880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1627_
timestamp 1635444444
transform 1 0 11960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1635444444
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_148
timestamp 1635444444
transform 1 0 14720 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1592_
timestamp 1635444444
transform 1 0 14812 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1760_
timestamp 1635444444
transform 1 0 13524 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1635444444
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp 1635444444
transform 1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1635444444
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1635444444
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1591_
timestamp 1635444444
transform 1 0 15548 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1635444444
transform 1 0 16652 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_17_185
timestamp 1635444444
transform 1 0 18124 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_191
timestamp 1635444444
transform 1 0 18676 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1197_
timestamp 1635444444
transform 1 0 18768 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_201
timestamp 1635444444
transform 1 0 19596 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_209
timestamp 1635444444
transform 1 0 20332 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1276_
timestamp 1635444444
transform 1 0 20516 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1635444444
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1635444444
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1635444444
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1635444444
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1635444444
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1635444444
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_264
timestamp 1635444444
transform 1 0 25392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_272
timestamp 1635444444
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_281
timestamp 1635444444
transform 1 0 26956 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1635444444
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1635444444
transform 1 0 25760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_296
timestamp 1635444444
transform 1 0 28336 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1158_
timestamp 1635444444
transform 1 0 27508 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1635444444
transform 1 0 28704 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_316
timestamp 1635444444
transform 1 0 30176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635444444
transform -1 0 30820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1635444444
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1635444444
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635444444
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1635444444
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1635444444
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1635444444
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1635444444
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1635444444
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1635444444
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1635444444
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1635444444
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1635444444
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1635444444
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1635444444
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_97
timestamp 1635444444
transform 1 0 10028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1782_
timestamp 1635444444
transform 1 0 10304 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_122
timestamp 1635444444
transform 1 0 12328 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp 1635444444
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1625_
timestamp 1635444444
transform 1 0 12696 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1774_
timestamp 1635444444
transform 1 0 11500 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1635444444
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_150
timestamp 1635444444
transform 1 0 14904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1635444444
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1811_
timestamp 1635444444
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_160
timestamp 1635444444
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_172
timestamp 1635444444
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1028_
timestamp 1635444444
transform 1 0 15272 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1194_
timestamp 1635444444
transform 1 0 16192 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1635444444
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1635444444
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1635444444
transform 1 0 17296 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 1635444444
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1192_
timestamp 1635444444
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1635444444
transform 1 0 19228 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_221
timestamp 1635444444
transform 1 0 21436 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1635444444
transform 1 0 21988 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1635444444
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1635444444
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_262
timestamp 1635444444
transform 1 0 25208 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1635444444
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1176_
timestamp 1635444444
transform 1 0 24380 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_270
timestamp 1635444444
transform 1 0 25944 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_282
timestamp 1635444444
transform 1 0 27048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_2  _1673_
timestamp 1635444444
transform 1 0 26128 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_18_286
timestamp 1635444444
transform 1 0 27416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_297
timestamp 1635444444
transform 1 0 28428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1635444444
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1149_
timestamp 1635444444
transform 1 0 27508 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1635444444
transform 1 0 28796 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_309
timestamp 1635444444
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_316
timestamp 1635444444
transform 1 0 30176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635444444
transform -1 0 30820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1635444444
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1635444444
transform 1 0 29900 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1635444444
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1635444444
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_19
timestamp 1635444444
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_7
timestamp 1635444444
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635444444
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635444444
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1635444444
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1635444444
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1635444444
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1635444444
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1635444444
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1635444444
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1635444444
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1635444444
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1635444444
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1635444444
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1635444444
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1635444444
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1635444444
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1635444444
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_81
timestamp 1635444444
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1635444444
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1635444444
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1635444444
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1635444444
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1635444444
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_89
timestamp 1635444444
transform 1 0 9292 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1635444444
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_103
timestamp 1635444444
transform 1 0 10580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1635444444
transform 1 0 9660 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1605_
timestamp 1635444444
transform 1 0 10948 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1606_
timestamp 1635444444
transform 1 0 9384 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1620_
timestamp 1635444444
transform 1 0 9936 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1773_
timestamp 1635444444
transform 1 0 10028 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1635444444
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1635444444
transform 1 0 11960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_131
timestamp 1635444444
transform 1 0 13156 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1635444444
transform 1 0 11592 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_125
timestamp 1635444444
transform 1 0 12604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1635444444
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1623_
timestamp 1635444444
transform 1 0 11684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1635_
timestamp 1635444444
transform 1 0 11960 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1732_
timestamp 1635444444
transform 1 0 12328 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_137
timestamp 1635444444
transform 1 0 13708 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_147
timestamp 1635444444
transform 1 0 14628 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1635444444
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1635444444
transform 1 0 14352 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1635444444
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1635444444
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1775_
timestamp 1635444444
transform 1 0 14720 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1780_
timestamp 1635444444
transform 1 0 13800 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1635444444
transform 1 0 15364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1635444444
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1635444444
transform 1 0 16928 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_157
timestamp 1635444444
transform 1 0 15548 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1635444444
transform 1 0 16376 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1635444444
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1545_
timestamp 1635444444
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1568_
timestamp 1635444444
transform 1 0 15548 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1569_
timestamp 1635444444
transform 1 0 15916 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_19_184
timestamp 1635444444
transform 1 0 18032 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1635444444
transform 1 0 18952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_178
timestamp 1635444444
transform 1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_182
timestamp 1635444444
transform 1 0 17848 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1635444444
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1635444444
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1635444444
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1195_
timestamp 1635444444
transform 1 0 17940 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1199_
timestamp 1635444444
transform 1 0 18124 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1635444444
transform 1 0 19688 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1198_
timestamp 1635444444
transform 1 0 19320 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1635444444
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1635444444
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1635444444
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_205
timestamp 1635444444
transform 1 0 19964 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1272_
timestamp 1635444444
transform 1 0 21068 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1267_
timestamp 1635444444
transform 1 0 20424 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1196_
timestamp 1635444444
transform 1 0 20332 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_20_213
timestamp 1635444444
transform 1 0 20700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_216
timestamp 1635444444
transform 1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_235
timestamp 1635444444
transform 1 0 22724 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_227
timestamp 1635444444
transform 1 0 21988 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_238
timestamp 1635444444
transform 1 0 23000 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1635444444
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1268_
timestamp 1635444444
transform 1 0 21804 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1398_
timestamp 1635444444
transform 1 0 22724 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1646_
timestamp 1635444444
transform 1 0 23368 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1415_
timestamp 1635444444
transform 1 0 23368 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1177_
timestamp 1635444444
transform 1 0 24104 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1635444444
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_246
timestamp 1635444444
transform 1 0 23736 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_241
timestamp 1635444444
transform 1 0 23276 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1175_
timestamp 1635444444
transform 1 0 24380 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1635444444
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1635444444
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_259
timestamp 1635444444
transform 1 0 24932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_262
timestamp 1635444444
transform 1 0 25208 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_2  _1694_
timestamp 1635444444
transform 1 0 25576 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22oi_1  _1662_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 25852 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_268
timestamp 1635444444
transform 1 0 25760 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1635444444
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1154_
timestamp 1635444444
transform 1 0 27048 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1635444444
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_281
timestamp 1635444444
transform 1 0 26956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_275
timestamp 1635444444
transform 1 0 26404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1635444444
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1635444444
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1635444444
transform 1 0 27140 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_19_299
timestamp 1635444444
transform 1 0 28612 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_291
timestamp 1635444444
transform 1 0 27876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1635444444
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1152_
timestamp 1635444444
transform 1 0 28244 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1153_
timestamp 1635444444
transform 1 0 28980 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_312
timestamp 1635444444
transform 1 0 29808 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_312
timestamp 1635444444
transform 1 0 29808 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635444444
transform -1 0 30820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635444444
transform -1 0 30820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1635444444
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1638_
timestamp 1635444444
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1635444444
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1635444444
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635444444
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1635444444
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1635444444
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1635444444
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1635444444
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1635444444
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1635444444
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1635444444
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_81
timestamp 1635444444
transform 1 0 8556 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_100
timestamp 1635444444
transform 1 0 10304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1635444444
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1635444444
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _0898_
timestamp 1635444444
transform 1 0 9476 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1604_
timestamp 1635444444
transform 1 0 10672 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1635444444
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1635444444
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_120
timestamp 1635444444
transform 1 0 12144 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1635444444
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1624_
timestamp 1635444444
transform 1 0 11776 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_132
timestamp 1635444444
transform 1 0 13248 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1635444444
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1556_
timestamp 1635444444
transform 1 0 14352 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1635444444
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_172
timestamp 1635444444
transform 1 0 16928 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1635444444
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1544_
timestamp 1635444444
transform 1 0 15548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1546_
timestamp 1635444444
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_179
timestamp 1635444444
transform 1 0 17572 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_189
timestamp 1635444444
transform 1 0 18492 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1570_
timestamp 1635444444
transform 1 0 17296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1635444444
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_201
timestamp 1635444444
transform 1 0 19596 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_213
timestamp 1635444444
transform 1 0 20700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1635444444
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_228
timestamp 1635444444
transform 1 0 22080 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_236
timestamp 1635444444
transform 1 0 22816 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1635444444
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1386_
timestamp 1635444444
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1635444444
transform 1 0 22908 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_253
timestamp 1635444444
transform 1 0 24380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_257
timestamp 1635444444
transform 1 0 24748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_262
timestamp 1635444444
transform 1 0 25208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1645_
timestamp 1635444444
transform 1 0 24840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1635444444
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1635444444
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1635444444
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_2  _1686_
timestamp 1635444444
transform 1 0 25576 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_21_285
timestamp 1635444444
transform 1 0 27324 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_295
timestamp 1635444444
transform 1 0 28244 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_299
timestamp 1635444444
transform 1 0 28612 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1147_
timestamp 1635444444
transform 1 0 27416 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1635444444
transform 1 0 28704 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_316
timestamp 1635444444
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635444444
transform -1 0 30820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1635444444
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1635444444
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635444444
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1635444444
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1635444444
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1635444444
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1635444444
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1635444444
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1635444444
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1635444444
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1635444444
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1635444444
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1977_
timestamp 1635444444
transform 1 0 8924 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_101
timestamp 1635444444
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_109
timestamp 1635444444
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 1635444444
transform 1 0 11684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1635444444
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1020_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 12052 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1584_
timestamp 1635444444
transform 1 0 11408 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1600_
timestamp 1635444444
transform 1 0 12880 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1635444444
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1635444444
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_150
timestamp 1635444444
transform 1 0 14904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1635444444
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1809_
timestamp 1635444444
transform 1 0 14076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1635444444
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_167
timestamp 1635444444
transform 1 0 16468 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_171
timestamp 1635444444
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1543_
timestamp 1635444444
transform 1 0 16560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1813_
timestamp 1635444444
transform 1 0 15272 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_178
timestamp 1635444444
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_182
timestamp 1635444444
transform 1 0 17848 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1635444444
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1635444444
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1202_
timestamp 1635444444
transform 1 0 17940 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1587_
timestamp 1635444444
transform 1 0 17204 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1635444444
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1280_
timestamp 1635444444
transform 1 0 21068 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1635444444
transform 1 0 19228 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_226
timestamp 1635444444
transform 1 0 21896 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1635444444
transform 1 0 22448 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1635444444
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_253
timestamp 1635444444
transform 1 0 24380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1635444444
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1635444444
transform 1 0 24472 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_270
timestamp 1635444444
transform 1 0 25944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1150_
timestamp 1635444444
transform 1 0 26680 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_287
timestamp 1635444444
transform 1 0 27508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1635444444
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1151_
timestamp 1635444444
transform 1 0 27876 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1635444444
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_312
timestamp 1635444444
transform 1 0 29808 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635444444
transform -1 0 30820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1635444444
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1660_
timestamp 1635444444
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_19
timestamp 1635444444
transform 1 0 2852 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_7
timestamp 1635444444
transform 1 0 1748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1635444444
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1635444444
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_31
timestamp 1635444444
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_43
timestamp 1635444444
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1635444444
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1635444444
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1635444444
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1635444444
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1635444444
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_106
timestamp 1635444444
transform 1 0 10856 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1635444444
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1978_
timestamp 1635444444
transform 1 0 9384 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_23_122
timestamp 1635444444
transform 1 0 12328 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1635444444
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1730_
timestamp 1635444444
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1807_
timestamp 1635444444
transform 1 0 12880 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_137
timestamp 1635444444
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_145
timestamp 1635444444
transform 1 0 14444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1557_
timestamp 1635444444
transform 1 0 14628 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_156
timestamp 1635444444
transform 1 0 15456 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1635444444
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp 1635444444
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1635444444
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1635444444
transform 1 0 16744 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_wb_clk_i
timestamp 1635444444
transform 1 0 15824 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_186
timestamp 1635444444
transform 1 0 18216 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1200_
timestamp 1635444444
transform 1 0 18584 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_199
timestamp 1635444444
transform 1 0 19412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_203
timestamp 1635444444
transform 1 0 19780 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1635444444
transform 1 0 19872 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1635444444
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_234
timestamp 1635444444
transform 1 0 22632 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1635444444
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1282_
timestamp 1635444444
transform 1 0 21804 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1294_
timestamp 1635444444
transform 1 0 23000 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_247
timestamp 1635444444
transform 1 0 23828 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_254
timestamp 1635444444
transform 1 0 24472 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1414_
timestamp 1635444444
transform 1 0 24196 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1635444444
transform 1 0 25208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_266
timestamp 1635444444
transform 1 0 25576 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1635444444
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1635444444
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1635444444
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_1  _1647_
timestamp 1635444444
transform 1 0 25944 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_285
timestamp 1635444444
transform 1 0 27324 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_296
timestamp 1635444444
transform 1 0 28336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1142_
timestamp 1635444444
transform 1 0 27416 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1635444444
transform 1 0 28704 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_316
timestamp 1635444444
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1635444444
transform -1 0 30820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1635444444
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1635444444
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_8
timestamp 1635444444
transform 1 0 1840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1635444444
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1658_
timestamp 1635444444
transform 1 0 1564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1635444444
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1635444444
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1635444444
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1635444444
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1635444444
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1635444444
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1635444444
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1635444444
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1635444444
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1635444444
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_106
timestamp 1635444444
transform 1 0 10856 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1635444444
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1046_
timestamp 1635444444
transform 1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_118
timestamp 1635444444
transform 1 0 11960 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_126
timestamp 1635444444
transform 1 0 12696 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1601_
timestamp 1635444444
transform 1 0 12788 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _1602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 11224 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1635444444
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1635444444
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_151
timestamp 1635444444
transform 1 0 14996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1635444444
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1812_
timestamp 1635444444
transform 1 0 14168 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_164
timestamp 1635444444
transform 1 0 16192 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_172
timestamp 1635444444
transform 1 0 16928 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1783_
timestamp 1635444444
transform 1 0 15364 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1635444444
transform 1 0 17112 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1635444444
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1635444444
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_206
timestamp 1635444444
transform 1 0 20056 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_214
timestamp 1635444444
transform 1 0 20792 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1214_
timestamp 1635444444
transform 1 0 19228 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1635444444
transform 1 0 20884 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_231
timestamp 1635444444
transform 1 0 22356 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1296_
timestamp 1635444444
transform 1 0 22724 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_244
timestamp 1635444444
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1635444444
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1635444444
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1178_
timestamp 1635444444
transform 1 0 24564 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_24_264
timestamp 1635444444
transform 1 0 25392 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_270
timestamp 1635444444
transform 1 0 25944 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_274
timestamp 1635444444
transform 1 0 26312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1685_
timestamp 1635444444
transform 1 0 26036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1635444444
transform 1 0 26680 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_294
timestamp 1635444444
transform 1 0 28152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1635444444
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1671_
timestamp 1635444444
transform 1 0 28520 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1635444444
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_309
timestamp 1635444444
transform 1 0 29532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_316
timestamp 1635444444
transform 1 0 30176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1635444444
transform -1 0 30820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1635444444
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1635444444
transform 1 0 29900 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1635444444
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1635444444
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1635444444
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1635444444
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1635444444
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1635444444
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1635444444
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1635444444
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1635444444
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1635444444
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1635444444
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1635444444
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_93
timestamp 1635444444
transform 1 0 9660 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1599_
timestamp 1635444444
transform 1 0 10396 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1635444444
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_128
timestamp 1635444444
transform 1 0 12880 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1635444444
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1806_
timestamp 1635444444
transform 1 0 12052 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_143
timestamp 1635444444
transform 1 0 14260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__o221ai_1  _1558_
timestamp 1635444444
transform 1 0 13616 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1635444444
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1635444444
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1803_
timestamp 1635444444
transform 1 0 15364 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1805_
timestamp 1635444444
transform 1 0 16652 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1635444444
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_185
timestamp 1635444444
transform 1 0 18124 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_191
timestamp 1635444444
transform 1 0 18676 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1216_
timestamp 1635444444
transform 1 0 18768 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1588_
timestamp 1635444444
transform 1 0 17848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_201
timestamp 1635444444
transform 1 0 19596 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_207
timestamp 1635444444
transform 1 0 20148 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_212
timestamp 1635444444
transform 1 0 20608 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1635444444
transform 1 0 20976 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_wb_clk_i
timestamp 1635444444
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1635444444
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_232
timestamp 1635444444
transform 1 0 22448 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1635444444
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1396_
timestamp 1635444444
transform 1 0 23000 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1418_
timestamp 1635444444
transform 1 0 21804 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_25_241
timestamp 1635444444
transform 1 0 23276 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_249
timestamp 1635444444
transform 1 0 24012 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_254
timestamp 1635444444
transform 1 0 24472 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1071_
timestamp 1635444444
transform 1 0 24104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1635444444
transform 1 0 24840 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1635444444
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_281
timestamp 1635444444
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1635444444
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_285
timestamp 1635444444
transform 1 0 27324 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_296
timestamp 1635444444
transform 1 0 28336 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1146_
timestamp 1635444444
transform 1 0 27416 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1635444444
transform 1 0 28704 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1635444444
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1635444444
transform -1 0 30820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1635444444
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1635444444
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_14
timestamp 1635444444
transform 1 0 2392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_7
timestamp 1635444444
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1635444444
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1635444444
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1363_
timestamp 1635444444
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1635444444
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1635444444
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1635444444
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1635444444
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_26
timestamp 1635444444
transform 1 0 3496 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_38
timestamp 1635444444
transform 1 0 4600 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1635444444
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1635444444
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1635444444
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1635444444
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1635444444
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1635444444
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1635444444
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1635444444
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1635444444
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1635444444
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1635444444
transform 1 0 8556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1635444444
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1976_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8740 0 -1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_26_102
timestamp 1635444444
transform 1 0 10488 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_102
timestamp 1635444444
transform 1 0 10488 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0899_
timestamp 1635444444
transform 1 0 9660 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1772_
timestamp 1635444444
transform 1 0 10856 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_115
timestamp 1635444444
transform 1 0 11684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_126
timestamp 1635444444
transform 1 0 12696 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1635444444
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1635444444
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1635444444
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_127
timestamp 1635444444
transform 1 0 12788 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1635444444
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1585_
timestamp 1635444444
transform 1 0 12052 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1808_
timestamp 1635444444
transform 1 0 11960 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1635444444
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_150
timestamp 1635444444
transform 1 0 14904 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_135
timestamp 1635444444
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_146
timestamp 1635444444
transform 1 0 14536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1635444444
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1541_
timestamp 1635444444
transform 1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1542_
timestamp 1635444444
transform 1 0 13248 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1767_
timestamp 1635444444
transform 1 0 13708 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1802_
timestamp 1635444444
transform 1 0 14076 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_159
timestamp 1635444444
transform 1 0 15732 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_171
timestamp 1635444444
transform 1 0 16836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1635444444
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1635444444
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1635444444
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1578_
timestamp 1635444444
transform 1 0 15548 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1580_
timestamp 1635444444
transform 1 0 15272 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1801_
timestamp 1635444444
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_183
timestamp 1635444444
transform 1 0 17940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1635444444
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1635444444
transform 1 0 17480 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_185
timestamp 1635444444
transform 1 0 18124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1635444444
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1566_
timestamp 1635444444
transform 1 0 17848 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_213
timestamp 1635444444
transform 1 0 20700 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_197
timestamp 1635444444
transform 1 0 19228 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_202
timestamp 1635444444
transform 1 0 19688 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_209
timestamp 1635444444
transform 1 0 20332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1399_
timestamp 1635444444
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1401_
timestamp 1635444444
transform 1 0 21068 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1409_
timestamp 1635444444
transform 1 0 20700 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1416_
timestamp 1635444444
transform 1 0 19412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1635444444
transform 1 0 19228 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_26_224
timestamp 1635444444
transform 1 0 21712 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_232
timestamp 1635444444
transform 1 0 22448 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1635444444
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_228
timestamp 1635444444
transform 1 0 22080 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_232
timestamp 1635444444
transform 1 0 22448 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1635444444
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1292_
timestamp 1635444444
transform 1 0 22540 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1402_
timestamp 1635444444
transform 1 0 22540 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1407_
timestamp 1635444444
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_242
timestamp 1635444444
transform 1 0 23368 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1635444444
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_260
timestamp 1635444444
transform 1 0 25024 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_242
timestamp 1635444444
transform 1 0 23368 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_262
timestamp 1635444444
transform 1 0 25208 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1635444444
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1432_
timestamp 1635444444
transform 1 0 24380 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1635444444
transform 1 0 23736 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1640_
timestamp 1635444444
transform 1 0 25668 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_270
timestamp 1635444444
transform 1 0 25944 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_270
timestamp 1635444444
transform 1 0 25944 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_266
timestamp 1635444444
transform 1 0 25576 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1635444444
transform 1 0 26128 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1112_
timestamp 1635444444
transform 1 0 26312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1635444444
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1635444444
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1635444444
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_278
timestamp 1635444444
transform 1 0 26680 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1145_
timestamp 1635444444
transform 1 0 27048 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_291
timestamp 1635444444
transform 1 0 27876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1635444444
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1635444444
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1635444444
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1141_
timestamp 1635444444
transform 1 0 28244 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1143_
timestamp 1635444444
transform 1 0 27324 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1635444444
transform 1 0 28612 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_26_312
timestamp 1635444444
transform 1 0 29808 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_315
timestamp 1635444444
transform 1 0 30084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_319
timestamp 1635444444
transform 1 0 30452 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1635444444
transform -1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1635444444
transform -1 0 30820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1635444444
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1635444444
transform 1 0 29532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_20
timestamp 1635444444
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1635444444
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_8
timestamp 1635444444
transform 1 0 1840 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1635444444
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1670_
timestamp 1635444444
transform 1 0 1564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1635444444
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1635444444
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1635444444
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1635444444
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1635444444
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1635444444
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1635444444
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1635444444
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1368_
timestamp 1635444444
transform 1 0 8188 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_106
timestamp 1635444444
transform 1 0 10856 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_89
timestamp 1635444444
transform 1 0 9292 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1635444444
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1367_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9384 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _1603_
timestamp 1635444444
transform 1 0 10488 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_119
timestamp 1635444444
transform 1 0 12052 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_125
timestamp 1635444444
transform 1 0 12604 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1768_
timestamp 1635444444
transform 1 0 12696 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1771_
timestamp 1635444444
transform 1 0 11224 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_135
timestamp 1635444444
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1635444444
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_148
timestamp 1635444444
transform 1 0 14720 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1635444444
transform 1 0 15088 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1635444444
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _1559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14076 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_28_156
timestamp 1635444444
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_169
timestamp 1635444444
transform 1 0 16652 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1579_
timestamp 1635444444
transform 1 0 15180 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1799_
timestamp 1635444444
transform 1 0 15824 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_175
timestamp 1635444444
transform 1 0 17204 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1635444444
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1635444444
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1635444444
transform 1 0 17296 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1635444444
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_203
timestamp 1635444444
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_215
timestamp 1635444444
transform 1 0 20884 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1281_
timestamp 1635444444
transform 1 0 20148 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1635444444
transform 1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_232
timestamp 1635444444
transform 1 0 22448 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1410_
timestamp 1635444444
transform 1 0 21620 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1419_
timestamp 1635444444
transform 1 0 22816 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1635444444
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1635444444
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_256
timestamp 1635444444
transform 1 0 24656 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1635444444
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1430_
timestamp 1635444444
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_264
timestamp 1635444444
transform 1 0 25392 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_268
timestamp 1635444444
transform 1 0 25760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_281
timestamp 1635444444
transform 1 0 26956 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1648_
timestamp 1635444444
transform 1 0 26128 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1661_
timestamp 1635444444
transform 1 0 25484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_297
timestamp 1635444444
transform 1 0 28428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1635444444
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1138_
timestamp 1635444444
transform 1 0 27508 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1635444444
transform 1 0 28796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1635444444
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_316
timestamp 1635444444
transform 1 0 30176 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1635444444
transform -1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1635444444
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1635444444
transform 1 0 29900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1635444444
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1635444444
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1635444444
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1635444444
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1635444444
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1635444444
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1635444444
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1635444444
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1635444444
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_69
timestamp 1635444444
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1635444444
transform 1 0 7728 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_100
timestamp 1635444444
transform 1 0 10304 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_88
timestamp 1635444444
transform 1 0 9200 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_117
timestamp 1635444444
transform 1 0 11868 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1635444444
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1635444444
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1563_
timestamp 1635444444
transform 1 0 12972 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1583_
timestamp 1635444444
transform 1 0 12236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1586_
timestamp 1635444444
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_132
timestamp 1635444444
transform 1 0 13248 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_144
timestamp 1635444444
transform 1 0 14352 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1581_
timestamp 1635444444
transform 1 0 14720 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_157
timestamp 1635444444
transform 1 0 15548 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1635444444
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1635444444
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1564_
timestamp 1635444444
transform 1 0 15916 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1657_
timestamp 1635444444
transform 1 0 16652 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_29_176
timestamp 1635444444
transform 1 0 17296 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1635444444
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1635444444
transform 1 0 17664 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_216
timestamp 1635444444
transform 1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1635444444
transform 1 0 19504 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1635444444
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_230
timestamp 1635444444
transform 1 0 22264 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_238
timestamp 1635444444
transform 1 0 23000 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1635444444
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1288_
timestamp 1635444444
transform 1 0 22632 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1406_
timestamp 1635444444
transform 1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_251
timestamp 1635444444
transform 1 0 24196 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_259
timestamp 1635444444
transform 1 0 24932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1290_
timestamp 1635444444
transform 1 0 23368 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1635444444
transform 1 0 25024 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1635444444
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1635444444
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1635444444
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1635444444
transform 1 0 27140 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_299
timestamp 1635444444
transform 1 0 28612 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1139_
timestamp 1635444444
transform 1 0 28980 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_312
timestamp 1635444444
transform 1 0 29808 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1635444444
transform -1 0 30820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1635444444
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1635444444
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1635444444
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1635444444
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1635444444
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1635444444
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1635444444
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1635444444
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1635444444
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1635444444
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1635444444
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1635444444
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1635444444
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1635444444
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _1974_
timestamp 1635444444
transform 1 0 9844 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_30_112
timestamp 1635444444
transform 1 0 11408 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_125
timestamp 1635444444
transform 1 0 12604 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0903_
timestamp 1635444444
transform 1 0 11776 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1635444444
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_145
timestamp 1635444444
transform 1 0 14444 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1635444444
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1539_
timestamp 1635444444
transform 1 0 13340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1540_
timestamp 1635444444
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_159
timestamp 1635444444
transform 1 0 15732 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_163
timestamp 1635444444
transform 1 0 16100 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_173
timestamp 1635444444
transform 1 0 17020 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1582_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 15180 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1800_
timestamp 1635444444
transform 1 0 16192 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1635444444
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1635444444
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1635444444
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1201_
timestamp 1635444444
transform 1 0 17572 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_197
timestamp 1635444444
transform 1 0 19228 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_201
timestamp 1635444444
transform 1 0 19596 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 1635444444
transform 1 0 20240 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_216
timestamp 1635444444
transform 1 0 20976 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1283_
timestamp 1635444444
transform 1 0 20608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1635444444
transform 1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1635444444
transform 1 0 19320 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_223
timestamp 1635444444
transform 1 0 21620 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1270_
timestamp 1635444444
transform 1 0 21344 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1289_
timestamp 1635444444
transform 1 0 22356 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_30_241
timestamp 1635444444
transform 1 0 23276 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1635444444
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_257
timestamp 1635444444
transform 1 0 24748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1635444444
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1663_
timestamp 1635444444
transform 1 0 25116 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1719_
timestamp 1635444444
transform 1 0 23644 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_wb_clk_i
timestamp 1635444444
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_270
timestamp 1635444444
transform 1 0 25944 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1140_
timestamp 1635444444
transform 1 0 26312 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1635444444
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1635444444
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1635444444
transform 1 0 27600 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1635444444
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_316
timestamp 1635444444
transform 1 0 30176 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1635444444
transform -1 0 30820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1635444444
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1635444444
transform 1 0 29900 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_19
timestamp 1635444444
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_7
timestamp 1635444444
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1635444444
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1635444444
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_31
timestamp 1635444444
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_43
timestamp 1635444444
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1635444444
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1635444444
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1635444444
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1635444444
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1635444444
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_101
timestamp 1635444444
transform 1 0 10396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1635444444
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0902_
timestamp 1635444444
transform 1 0 9660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1635444444
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1635444444
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_126
timestamp 1635444444
transform 1 0 12696 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1635444444
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1561_
timestamp 1635444444
transform 1 0 13064 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1562_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 11960 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_135
timestamp 1635444444
transform 1 0 13524 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_152
timestamp 1635444444
transform 1 0 15088 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 13892 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1635444444
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1635444444
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_173
timestamp 1635444444
transform 1 0 17020 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1635444444
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1560_
timestamp 1635444444
transform 1 0 15456 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1565_
timestamp 1635444444
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_187
timestamp 1635444444
transform 1 0 18308 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _1215_
timestamp 1635444444
transform 1 0 17572 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1635444444
transform 1 0 19412 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_204
timestamp 1635444444
transform 1 0 19872 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_212
timestamp 1635444444
transform 1 0 20608 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1635444444
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1105_
timestamp 1635444444
transform 1 0 19504 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1271_
timestamp 1635444444
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1635444444
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1635444444
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1635444444
transform 1 0 21804 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_31_241
timestamp 1635444444
transform 1 0 23276 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_247
timestamp 1635444444
transform 1 0 23828 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1635444444
transform 1 0 23920 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_264
timestamp 1635444444
transform 1 0 25392 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1635444444
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1635444444
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1635444444
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1132_
timestamp 1635444444
transform 1 0 27140 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_wb_clk_i
timestamp 1635444444
transform 1 0 26128 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1635444444
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_299
timestamp 1635444444
transform 1 0 28612 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1635444444
transform 1 0 28704 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_316
timestamp 1635444444
transform 1 0 30176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1635444444
transform -1 0 30820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1635444444
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1635444444
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_8
timestamp 1635444444
transform 1 0 1840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1635444444
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1681_
timestamp 1635444444
transform 1 0 1564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1635444444
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1635444444
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1635444444
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1635444444
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1635444444
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1635444444
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1635444444
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1635444444
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1975_
timestamp 1635444444
transform 1 0 8924 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_32_102
timestamp 1635444444
transform 1 0 10488 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_114
timestamp 1635444444
transform 1 0 11592 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_122
timestamp 1635444444
transform 1 0 12328 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_130
timestamp 1635444444
transform 1 0 13064 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1022_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 11776 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1643_
timestamp 1635444444
transform 1 0 13156 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1635444444
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_147
timestamp 1635444444
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1635444444
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _1573_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1770_
timestamp 1635444444
transform 1 0 14996 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_160
timestamp 1635444444
transform 1 0 15824 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_173
timestamp 1635444444
transform 1 0 17020 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1796_
timestamp 1635444444
transform 1 0 16192 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_32_184
timestamp 1635444444
transform 1 0 18032 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1635444444
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1669_
timestamp 1635444444
transform 1 0 17388 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1635444444
transform 1 0 20056 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_214
timestamp 1635444444
transform 1 0 20792 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1148_
timestamp 1635444444
transform 1 0 20424 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1205_
timestamp 1635444444
transform 1 0 19228 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_220
timestamp 1635444444
transform 1 0 21344 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_229
timestamp 1635444444
transform 1 0 22172 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_237
timestamp 1635444444
transform 1 0 22908 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1293_
timestamp 1635444444
transform 1 0 23092 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1295_
timestamp 1635444444
transform 1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1635444444
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1635444444
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1635444444
transform 1 0 24380 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_32_269
timestamp 1635444444
transform 1 0 25852 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1712_
timestamp 1635444444
transform 1 0 26404 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_284
timestamp 1635444444
transform 1 0 27232 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_297
timestamp 1635444444
transform 1 0 28428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1635444444
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1144_
timestamp 1635444444
transform 1 0 27600 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1698_
timestamp 1635444444
transform 1 0 28796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_312
timestamp 1635444444
transform 1 0 29808 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1635444444
transform -1 0 30820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1635444444
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1709_
timestamp 1635444444
transform 1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1635444444
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1635444444
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1635444444
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1635444444
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1635444444
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1635444444
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1635444444
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1635444444
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1635444444
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1635444444
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1635444444
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1635444444
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1635444444
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1635444444
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1635444444
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1635444444
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1635444444
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1635444444
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1635444444
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_81
timestamp 1635444444
transform 1 0 8556 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_86
timestamp 1635444444
transform 1 0 9016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1635444444
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1635444444
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1635444444
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0900_
timestamp 1635444444
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0901_
timestamp 1635444444
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0897_
timestamp 1635444444
transform 1 0 9384 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1635444444
transform 1 0 9936 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_95
timestamp 1635444444
transform 1 0 9844 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_89
timestamp 1635444444
transform 1 0 9292 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_94
timestamp 1635444444
transform 1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1031_
timestamp 1635444444
transform 1 0 10580 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0896_
timestamp 1635444444
transform 1 0 10120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1635444444
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1635444444
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_108
timestamp 1635444444
transform 1 0 11040 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1021_
timestamp 1635444444
transform 1 0 11684 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0905_
timestamp 1635444444
transform 1 0 11408 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1635444444
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1635444444
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1635444444
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_2  _1032_
timestamp 1635444444
transform 1 0 12696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1635444444
transform 1 0 12604 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_34_125
timestamp 1635444444
transform 1 0 12604 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_121
timestamp 1635444444
transform 1 0 12236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_124
timestamp 1635444444
transform 1 0 12512 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_120
timestamp 1635444444
transform 1 0 12144 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_130
timestamp 1635444444
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_130
timestamp 1635444444
transform 1 0 13064 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_134
timestamp 1635444444
transform 1 0 13432 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_152
timestamp 1635444444
transform 1 0 15088 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1635444444
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1635444444
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_150
timestamp 1635444444
transform 1 0 14904 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1635444444
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _1654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 13524 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_2  _1704_
timestamp 1635444444
transform 1 0 14352 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1641_
timestamp 1635444444
transform 1 0 15456 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1574_
timestamp 1635444444
transform 1 0 15272 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_34_159
timestamp 1635444444
transform 1 0 15732 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1635444444
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1769_
timestamp 1635444444
transform 1 0 16652 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1659_
timestamp 1635444444
transform 1 0 17112 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1535_
timestamp 1635444444
transform 1 0 16376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1635444444
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_170
timestamp 1635444444
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_165
timestamp 1635444444
transform 1 0 16284 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1635444444
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_178
timestamp 1635444444
transform 1 0 17480 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_186
timestamp 1635444444
transform 1 0 18216 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_184
timestamp 1635444444
transform 1 0 18032 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1635444444
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1635444444
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1204_
timestamp 1635444444
transform 1 0 18400 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1635444444
transform 1 0 18308 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_33_203
timestamp 1635444444
transform 1 0 19780 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1635444444
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_203
timestamp 1635444444
transform 1 0 19780 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_216
timestamp 1635444444
transform 1 0 20976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0883_
timestamp 1635444444
transform 1 0 19412 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1278_
timestamp 1635444444
transform 1 0 20516 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1284_
timestamp 1635444444
transform 1 0 20516 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1297_
timestamp 1635444444
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1291_
timestamp 1635444444
transform 1 0 21988 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 1635444444
transform 1 0 21344 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1635444444
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1635444444
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1635444444
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1400_
timestamp 1635444444
transform 1 0 23000 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1635444444
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_234
timestamp 1635444444
transform 1 0 22632 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1426_
timestamp 1635444444
transform 1 0 23092 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_242
timestamp 1635444444
transform 1 0 23368 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_249
timestamp 1635444444
transform 1 0 24012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_253
timestamp 1635444444
transform 1 0 24380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1635444444
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_253
timestamp 1635444444
transform 1 0 24380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1635444444
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1635444444
transform 1 0 23736 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1687_
timestamp 1635444444
transform 1 0 24472 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1722_
timestamp 1635444444
transform 1 0 24472 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_263
timestamp 1635444444
transform 1 0 25300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1635444444
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_281
timestamp 1635444444
transform 1 0 26956 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_263
timestamp 1635444444
transform 1 0 25300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_277
timestamp 1635444444
transform 1 0 26588 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1635444444
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1642_
timestamp 1635444444
transform 1 0 25668 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1674_
timestamp 1635444444
transform 1 0 25668 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_296
timestamp 1635444444
transform 1 0 28336 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_288
timestamp 1635444444
transform 1 0 27600 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_302
timestamp 1635444444
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1134_
timestamp 1635444444
transform 1 0 27968 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1137_
timestamp 1635444444
transform 1 0 27508 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1672_
timestamp 1635444444
transform 1 0 27324 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1635444444
transform 1 0 28704 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 1635444444
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_309
timestamp 1635444444
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_316
timestamp 1635444444
transform 1 0 30176 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1635444444
transform -1 0 30820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1635444444
transform -1 0 30820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1635444444
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1635444444
transform 1 0 29900 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_14
timestamp 1635444444
transform 1 0 2392 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_7
timestamp 1635444444
transform 1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1635444444
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1689_
timestamp 1635444444
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1635444444
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_26
timestamp 1635444444
transform 1 0 3496 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_38
timestamp 1635444444
transform 1 0 4600 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_50
timestamp 1635444444
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1635444444
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1635444444
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_69
timestamp 1635444444
transform 1 0 7452 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1954_
timestamp 1635444444
transform 1 0 7728 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_35_101
timestamp 1635444444
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1635444444
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_89
timestamp 1635444444
transform 1 0 9292 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_93
timestamp 1635444444
transform 1 0 9660 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _1042_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9752 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1635444444
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1635444444
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1973_
timestamp 1635444444
transform 1 0 11776 0 -1 21760
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_35_135
timestamp 1635444444
transform 1 0 13524 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_143
timestamp 1635444444
transform 1 0 14260 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_152
timestamp 1635444444
transform 1 0 15088 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1026_
timestamp 1635444444
transform 1 0 13892 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1179_
timestamp 1635444444
transform 1 0 14628 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1635444444
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1635444444
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_173
timestamp 1635444444
transform 1 0 17020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1635444444
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1635444444
transform 1 0 15456 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1526_
timestamp 1635444444
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_177
timestamp 1635444444
transform 1 0 17388 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_185
timestamp 1635444444
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1635444444
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1680_
timestamp 1635444444
transform 1 0 17480 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1688_
timestamp 1635444444
transform 1 0 18492 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_35_204
timestamp 1635444444
transform 1 0 19872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_213
timestamp 1635444444
transform 1 0 20700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1635444444
transform 1 0 21068 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0979_
timestamp 1635444444
transform 1 0 19504 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1635444444
transform 1 0 20240 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1635444444
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_230
timestamp 1635444444
transform 1 0 22264 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1635444444
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1300_
timestamp 1635444444
transform 1 0 21804 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1635444444
transform 1 0 22632 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_35_250
timestamp 1635444444
transform 1 0 24104 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_256
timestamp 1635444444
transform 1 0 24656 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1652_
timestamp 1635444444
transform 1 0 24748 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_35_267
timestamp 1635444444
transform 1 0 25668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1635444444
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1635444444
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1635444444
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1635444444
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1653_
timestamp 1635444444
transform 1 0 26036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_296
timestamp 1635444444
transform 1 0 28336 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1136_
timestamp 1635444444
transform 1 0 27508 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1635444444
transform 1 0 28704 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_316
timestamp 1635444444
transform 1 0 30176 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1635444444
transform -1 0 30820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1635444444
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1635444444
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1635444444
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1635444444
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1635444444
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1635444444
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1635444444
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1635444444
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1635444444
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1635444444
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1635444444
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1635444444
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1635444444
transform 1 0 8188 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1635444444
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1039_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 10580 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1047_
timestamp 1635444444
transform 1 0 9476 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_111
timestamp 1635444444
transform 1 0 11316 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_121
timestamp 1635444444
transform 1 0 12236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_128
timestamp 1635444444
transform 1 0 12880 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1041_
timestamp 1635444444
transform 1 0 11684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1527_
timestamp 1635444444
transform 1 0 12604 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_146
timestamp 1635444444
transform 1 0 14536 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_150
timestamp 1635444444
transform 1 0 14904 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1635444444
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1024_
timestamp 1635444444
transform 1 0 14076 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1766_
timestamp 1635444444
transform 1 0 14996 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_160
timestamp 1635444444
transform 1 0 15824 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_173
timestamp 1635444444
transform 1 0 17020 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1765_
timestamp 1635444444
transform 1 0 16192 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_36_181
timestamp 1635444444
transform 1 0 17756 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1635444444
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1635444444
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1218_
timestamp 1635444444
transform 1 0 17940 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1635444444
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_205
timestamp 1635444444
transform 1 0 19964 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_209
timestamp 1635444444
transform 1 0 20332 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1217_
timestamp 1635444444
transform 1 0 19596 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1635444444
transform 1 0 20424 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_36_226
timestamp 1635444444
transform 1 0 21896 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_234
timestamp 1635444444
transform 1 0 22632 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1425_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 22908 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1635444444
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1635444444
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_259
timestamp 1635444444
transform 1 0 24932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1635444444
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _1437_
timestamp 1635444444
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_263
timestamp 1635444444
transform 1 0 25300 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_273
timestamp 1635444444
transform 1 0 26220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_277
timestamp 1635444444
transform 1 0 26588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1695_
timestamp 1635444444
transform 1 0 25392 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1701_
timestamp 1635444444
transform 1 0 26680 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_36_287
timestamp 1635444444
transform 1 0 27508 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1635444444
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1135_
timestamp 1635444444
transform 1 0 28244 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_36_312
timestamp 1635444444
transform 1 0 29808 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1635444444
transform -1 0 30820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1635444444
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1635444444
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1635444444
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1635444444
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1635444444
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1635444444
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1635444444
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1635444444
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1635444444
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1635444444
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1635444444
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp 1635444444
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_77
timestamp 1635444444
transform 1 0 8188 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_87
timestamp 1635444444
transform 1 0 9108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_1  _1048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8464 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_37_106
timestamp 1635444444
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_91
timestamp 1635444444
transform 1 0 9476 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_95
timestamp 1635444444
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_99
timestamp 1635444444
transform 1 0 10212 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1635444444
transform 1 0 9568 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1045_
timestamp 1635444444
transform 1 0 10304 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_116
timestamp 1635444444
transform 1 0 11776 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_123
timestamp 1635444444
transform 1 0 12420 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_131
timestamp 1635444444
transform 1 0 13156 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1635444444
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1635444444
transform 1 0 11500 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1635444444
transform 1 0 12144 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_136
timestamp 1635444444
transform 1 0 13616 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_149
timestamp 1635444444
transform 1 0 14812 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1055_
timestamp 1635444444
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1763_
timestamp 1635444444
transform 1 0 13984 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_37_160
timestamp 1635444444
transform 1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1635444444
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_1  _1538_
timestamp 1635444444
transform 1 0 15180 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1784_
timestamp 1635444444
transform 1 0 16652 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_37_178
timestamp 1635444444
transform 1 0 17480 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_186
timestamp 1635444444
transform 1 0 18216 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 18400 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_37_208
timestamp 1635444444
transform 1 0 20240 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1635444444
transform 1 0 20792 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 1635444444
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1635444444
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1635444444
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1635444444
transform 1 0 21804 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_37_241
timestamp 1635444444
transform 1 0 23276 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_249
timestamp 1635444444
transform 1 0 24012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_253
timestamp 1635444444
transform 1 0 24380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_258
timestamp 1635444444
transform 1 0 24840 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1397_
timestamp 1635444444
transform 1 0 23644 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1639_
timestamp 1635444444
transform 1 0 24472 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1676_
timestamp 1635444444
transform 1 0 25208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_266
timestamp 1635444444
transform 1 0 25576 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_272
timestamp 1635444444
transform 1 0 26128 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1635444444
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_281
timestamp 1635444444
transform 1 0 26956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1635444444
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1684_
timestamp 1635444444
transform 1 0 26220 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_293
timestamp 1635444444
transform 1 0 28060 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1133_
timestamp 1635444444
transform 1 0 27232 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1635444444
transform 1 0 28428 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_37_313
timestamp 1635444444
transform 1 0 29900 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_319
timestamp 1635444444
transform 1 0 30452 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1635444444
transform -1 0 30820 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_14
timestamp 1635444444
transform 1 0 2392 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_7
timestamp 1635444444
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1635444444
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1697_
timestamp 1635444444
transform 1 0 2116 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1635444444
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1635444444
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1635444444
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1635444444
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1635444444
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1635444444
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1635444444
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1635444444
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1635444444
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1635444444
transform 1 0 8188 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1052_
timestamp 1635444444
transform 1 0 8924 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_38_94
timestamp 1635444444
transform 1 0 9752 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0889_
timestamp 1635444444
transform 1 0 10304 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_38_110
timestamp 1635444444
transform 1 0 11224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_114
timestamp 1635444444
transform 1 0 11592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_123
timestamp 1635444444
transform 1 0 12420 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_129
timestamp 1635444444
transform 1 0 12972 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__or4b_1  _1056_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 11684 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_1  _1536_
timestamp 1635444444
transform 1 0 13064 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1635444444
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_150
timestamp 1635444444
transform 1 0 14904 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1635444444
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1537_
timestamp 1635444444
transform 1 0 14076 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_38_158
timestamp 1635444444
transform 1 0 15640 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_170
timestamp 1635444444
transform 1 0 16744 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1764_
timestamp 1635444444
transform 1 0 15916 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1635444444
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1635444444
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1635444444
transform 1 0 17296 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_200
timestamp 1635444444
transform 1 0 19504 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_211
timestamp 1635444444
transform 1 0 20516 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1389_
timestamp 1635444444
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1390_
timestamp 1635444444
transform 1 0 19872 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_38_228
timestamp 1635444444
transform 1 0 22080 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_235
timestamp 1635444444
transform 1 0 22724 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1385_
timestamp 1635444444
transform 1 0 22448 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1391_
timestamp 1635444444
transform 1 0 21252 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_38_243
timestamp 1635444444
transform 1 0 23460 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1635444444
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_259
timestamp 1635444444
transform 1 0 24932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1635444444
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _1442_
timestamp 1635444444
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1720_
timestamp 1635444444
transform 1 0 23644 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_266
timestamp 1635444444
transform 1 0 25576 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1438_
timestamp 1635444444
transform 1 0 25300 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1635444444
transform 1 0 26128 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_288
timestamp 1635444444
transform 1 0 27600 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_302
timestamp 1635444444
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1130_
timestamp 1635444444
transform 1 0 27968 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_38_312
timestamp 1635444444
transform 1 0 29808 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1635444444
transform -1 0 30820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1635444444
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1710_
timestamp 1635444444
transform 1 0 29532 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1635444444
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1635444444
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1635444444
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1635444444
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1635444444
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1635444444
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1635444444
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1635444444
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1635444444
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1635444444
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1635444444
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1635444444
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1635444444
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1635444444
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_57
timestamp 1635444444
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_65
timestamp 1635444444
transform 1 0 7084 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1635444444
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1635444444
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1635444444
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_83
timestamp 1635444444
transform 1 0 8740 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1635444444
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1635444444
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1635444444
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1058_
timestamp 1635444444
transform 1 0 8924 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1952_
timestamp 1635444444
transform 1 0 7268 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1635444444
transform 1 0 9108 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_39_103
timestamp 1635444444
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_108
timestamp 1635444444
transform 1 0 11040 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_94
timestamp 1635444444
transform 1 0 9752 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1054_
timestamp 1635444444
transform 1 0 10488 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1051_
timestamp 1635444444
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1050_
timestamp 1635444444
transform 1 0 11408 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1635444444
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_116
timestamp 1635444444
transform 1 0 11776 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1635444444
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o211ai_1  _1057_
timestamp 1635444444
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1037_
timestamp 1635444444
transform 1 0 12144 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_40_125
timestamp 1635444444
transform 1 0 12604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_121
timestamp 1635444444
transform 1 0 12236 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1534_
timestamp 1635444444
transform 1 0 12972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_131
timestamp 1635444444
transform 1 0 13156 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _1528_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 13524 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1635444444
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1635444444
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1635444444
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1785_
timestamp 1635444444
transform 1 0 14628 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_149
timestamp 1635444444
transform 1 0 14812 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_141
timestamp 1635444444
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_146
timestamp 1635444444
transform 1 0 14536 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_142
timestamp 1635444444
transform 1 0 14168 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1635444444
transform 1 0 14996 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1525_
timestamp 1635444444
transform 1 0 15916 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_154
timestamp 1635444444
transform 1 0 15272 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_160
timestamp 1635444444
transform 1 0 15824 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_156
timestamp 1635444444
transform 1 0 15456 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1531_
timestamp 1635444444
transform 1 0 16008 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1635444444
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_165
timestamp 1635444444
transform 1 0 16284 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1635444444
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1635444444
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1707_
timestamp 1635444444
transform 1 0 17020 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1696_
timestamp 1635444444
transform 1 0 16928 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_39_179
timestamp 1635444444
transform 1 0 17572 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1635444444
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_192
timestamp 1635444444
transform 1 0 18768 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_180
timestamp 1635444444
transform 1 0 17664 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1635444444
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1635444444
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _1062_
timestamp 1635444444
transform 1 0 18216 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1370_
timestamp 1635444444
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1524_
timestamp 1635444444
transform 1 0 17940 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_39_197
timestamp 1635444444
transform 1 0 19228 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_209
timestamp 1635444444
transform 1 0 20332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1635444444
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_203
timestamp 1635444444
transform 1 0 19780 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_211
timestamp 1635444444
transform 1 0 20516 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1286_
timestamp 1635444444
transform 1 0 20792 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1388_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 19596 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1529_
timestamp 1635444444
transform 1 0 19504 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1387_
timestamp 1635444444
transform 1 0 22172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1635444444
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1635444444
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1635444444
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1787_
timestamp 1635444444
transform 1 0 23092 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1411_
timestamp 1635444444
transform 1 0 22908 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1405_
timestamp 1635444444
transform 1 0 22448 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_235
timestamp 1635444444
transform 1 0 22724 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_231
timestamp 1635444444
transform 1 0 22356 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_233
timestamp 1635444444
transform 1 0 22540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_219
timestamp 1635444444
transform 1 0 21252 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_240
timestamp 1635444444
transform 1 0 23184 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_255
timestamp 1635444444
transform 1 0 24564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1635444444
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_256
timestamp 1635444444
transform 1 0 24656 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1635444444
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1129_
timestamp 1635444444
transform 1 0 25024 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1383_
timestamp 1635444444
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1635444444
transform 1 0 24288 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1635444444
transform 1 0 24932 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1635444444
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1635444444
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_281
timestamp 1635444444
transform 1 0 26956 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_269
timestamp 1635444444
transform 1 0 25852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1635444444
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1131_
timestamp 1635444444
transform 1 0 26588 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_39_285
timestamp 1635444444
transform 1 0 27324 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_302
timestamp 1635444444
transform 1 0 28888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_286
timestamp 1635444444
transform 1 0 27416 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_293
timestamp 1635444444
transform 1 0 28060 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1635444444
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1699_
timestamp 1635444444
transform 1 0 27784 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1635444444
transform 1 0 27416 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1635444444
transform 1 0 28796 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1635444444
transform 1 0 29256 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1635444444
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_309
timestamp 1635444444
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_309
timestamp 1635444444
transform 1 0 29532 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1635444444
transform 1 0 29808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1635444444
transform 1 0 29900 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1635444444
transform -1 0 30820 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1635444444
transform -1 0 30820 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_316
timestamp 1635444444
transform 1 0 30176 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_316
timestamp 1635444444
transform 1 0 30176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_20
timestamp 1635444444
transform 1 0 2944 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1635444444
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_8
timestamp 1635444444
transform 1 0 1840 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1635444444
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1708_
timestamp 1635444444
transform 1 0 1564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_32
timestamp 1635444444
transform 1 0 4048 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_44
timestamp 1635444444
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1635444444
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1635444444
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_69
timestamp 1635444444
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_77
timestamp 1635444444
transform 1 0 8188 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_81
timestamp 1635444444
transform 1 0 8556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1635444444
transform 1 0 8280 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0911_
timestamp 1635444444
transform 1 0 8924 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1635444444
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_90
timestamp 1635444444
transform 1 0 9384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_99
timestamp 1635444444
transform 1 0 10212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0888_
timestamp 1635444444
transform 1 0 9752 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1033_
timestamp 1635444444
transform 1 0 10580 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_41_118
timestamp 1635444444
transform 1 0 11960 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_125
timestamp 1635444444
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1635444444
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0912_
timestamp 1635444444
transform 1 0 12328 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1635444444
transform 1 0 12972 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1035_
timestamp 1635444444
transform 1 0 11500 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_41_132
timestamp 1635444444
transform 1 0 13248 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_139
timestamp 1635444444
transform 1 0 13892 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_148
timestamp 1635444444
transform 1 0 14720 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1635444444
transform 1 0 13616 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1532_
timestamp 1635444444
transform 1 0 15088 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1533_
timestamp 1635444444
transform 1 0 14444 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_156
timestamp 1635444444
transform 1 0 15456 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1635444444
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_169
timestamp 1635444444
transform 1 0 16652 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1635444444
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0914_
timestamp 1635444444
transform 1 0 15824 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1664_
timestamp 1635444444
transform 1 0 16744 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1635444444
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_184
timestamp 1635444444
transform 1 0 18032 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_191
timestamp 1635444444
transform 1 0 18676 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0904_
timestamp 1635444444
transform 1 0 18124 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1262_
timestamp 1635444444
transform 1 0 19044 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_41_200
timestamp 1635444444
transform 1 0 19504 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_208
timestamp 1635444444
transform 1 0 20240 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1357_
timestamp 1635444444
transform 1 0 20424 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1635444444
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_225
timestamp 1635444444
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_229
timestamp 1635444444
transform 1 0 22172 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1635444444
transform 1 0 23092 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1635444444
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1735_
timestamp 1635444444
transform 1 0 22264 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_41_246
timestamp 1635444444
transform 1 0 23736 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_261
timestamp 1635444444
transform 1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1395_
timestamp 1635444444
transform 1 0 23460 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1793_
timestamp 1635444444
transform 1 0 24288 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_41_268
timestamp 1635444444
transform 1 0 25760 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1635444444
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1635444444
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1392_
timestamp 1635444444
transform 1 0 25484 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_293
timestamp 1635444444
transform 1 0 28060 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_297
timestamp 1635444444
transform 1 0 28428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_304
timestamp 1635444444
transform 1 0 29072 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1635444444
transform 1 0 28796 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1635444444
transform 1 0 28152 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_316
timestamp 1635444444
transform 1 0 30176 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1635444444
transform -1 0 30820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1635444444
transform 1 0 29808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_19
timestamp 1635444444
transform 1 0 2852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_7
timestamp 1635444444
transform 1 0 1748 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1635444444
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1635444444
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1635444444
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1635444444
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1635444444
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1635444444
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1635444444
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1635444444
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1635444444
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1635444444
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1635444444
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0892_
timestamp 1635444444
transform 1 0 8924 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_42_101
timestamp 1635444444
transform 1 0 10396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_90
timestamp 1635444444
transform 1 0 9384 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_96
timestamp 1635444444
transform 1 0 9936 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0886_
timestamp 1635444444
transform 1 0 10028 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1794_
timestamp 1635444444
transform 1 0 10764 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_114
timestamp 1635444444
transform 1 0 11592 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_123
timestamp 1635444444
transform 1 0 12420 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_129
timestamp 1635444444
transform 1 0 12972 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0913_
timestamp 1635444444
transform 1 0 11960 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _1064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 13064 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1635444444
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1635444444
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1951_
timestamp 1635444444
transform 1 0 14076 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_42_157
timestamp 1635444444
transform 1 0 15548 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_170
timestamp 1635444444
transform 1 0 16744 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1717_
timestamp 1635444444
transform 1 0 17112 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1798_
timestamp 1635444444
transform 1 0 15916 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_42_181
timestamp 1635444444
transform 1 0 17756 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1635444444
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1635444444
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1255_
timestamp 1635444444
transform 1 0 18308 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_42_203
timestamp 1635444444
transform 1 0 19780 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_207
timestamp 1635444444
transform 1 0 20148 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_214
timestamp 1635444444
transform 1 0 20792 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1277_
timestamp 1635444444
transform 1 0 21160 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1285_
timestamp 1635444444
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1358_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 20240 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_223
timestamp 1635444444
transform 1 0 21620 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_230
timestamp 1635444444
transform 1 0 22264 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_238
timestamp 1635444444
transform 1 0 23000 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1384_
timestamp 1635444444
transform 1 0 21988 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1792_
timestamp 1635444444
transform 1 0 23092 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1635444444
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_256
timestamp 1635444444
transform 1 0 24656 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1635444444
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1403_
timestamp 1635444444
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_268
timestamp 1635444444
transform 1 0 25760 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_274
timestamp 1635444444
transform 1 0 26312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_282
timestamp 1635444444
transform 1 0 27048 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1635444444
transform 1 0 25944 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1126_
timestamp 1635444444
transform 1 0 26680 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_294
timestamp 1635444444
transform 1 0 28152 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_300
timestamp 1635444444
transform 1 0 28704 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1635444444
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1635444444
transform 1 0 28796 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_309
timestamp 1635444444
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_316
timestamp 1635444444
transform 1 0 30176 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1635444444
transform -1 0 30820 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1635444444
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1635444444
transform 1 0 29900 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1635444444
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1635444444
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_8
timestamp 1635444444
transform 1 0 1840 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1635444444
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1718_
timestamp 1635444444
transform 1 0 1564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1728_
timestamp 1635444444
transform 1 0 2208 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1635444444
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1635444444
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1635444444
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1635444444
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1635444444
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1635444444
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1635444444
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_81
timestamp 1635444444
transform 1 0 8556 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_4  _1731_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8740 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1635444444
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_95
timestamp 1635444444
transform 1 0 9844 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1040_
timestamp 1635444444
transform 1 0 10580 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_43_122
timestamp 1635444444
transform 1 0 12328 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1635444444
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__o311a_1  _1065_
timestamp 1635444444
transform 1 0 13064 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1788_
timestamp 1635444444
transform 1 0 11500 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_43_138
timestamp 1635444444
transform 1 0 13800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_146
timestamp 1635444444
transform 1 0 14536 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14168 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_154
timestamp 1635444444
transform 1 0 15272 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1635444444
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 1635444444
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1635444444
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1727_
timestamp 1635444444
transform 1 0 17020 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1797_
timestamp 1635444444
transform 1 0 15364 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_43_180
timestamp 1635444444
transform 1 0 17664 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_188
timestamp 1635444444
transform 1 0 18400 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_192
timestamp 1635444444
transform 1 0 18768 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1122_
timestamp 1635444444
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1298_
timestamp 1635444444
transform 1 0 18860 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_199
timestamp 1635444444
transform 1 0 19412 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_205
timestamp 1635444444
transform 1 0 19964 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_211
timestamp 1635444444
transform 1 0 20516 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_218
timestamp 1635444444
transform 1 0 21160 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1263_
timestamp 1635444444
transform 1 0 20056 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1506_
timestamp 1635444444
transform 1 0 20884 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1635444444
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_233
timestamp 1635444444
transform 1 0 22540 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1635444444
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _1404_
timestamp 1635444444
transform 1 0 21988 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1412_
timestamp 1635444444
transform 1 0 22908 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_243
timestamp 1635444444
transform 1 0 23460 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_247
timestamp 1635444444
transform 1 0 23828 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_257
timestamp 1635444444
transform 1 0 24748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1420_
timestamp 1635444444
transform 1 0 25116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1791_
timestamp 1635444444
transform 1 0 23920 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_43_264
timestamp 1635444444
transform 1 0 25392 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1635444444
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_281
timestamp 1635444444
transform 1 0 26956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1635444444
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_289
timestamp 1635444444
transform 1 0 27692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_301
timestamp 1635444444
transform 1 0 28796 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1117_
timestamp 1635444444
transform 1 0 27324 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_309
timestamp 1635444444
transform 1 0 29532 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_316
timestamp 1635444444
transform 1 0 30176 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1635444444
transform -1 0 30820 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1635444444
transform 1 0 29808 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1635444444
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1635444444
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1635444444
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1635444444
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1635444444
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1635444444
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1635444444
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1635444444
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1635444444
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1635444444
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1635444444
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_85
timestamp 1635444444
transform 1 0 8924 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1635444444
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0893_
timestamp 1635444444
transform 1 0 9016 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_44_107
timestamp 1635444444
transform 1 0 10948 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_96
timestamp 1635444444
transform 1 0 9936 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_2  _0894_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 10304 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_44_119
timestamp 1635444444
transform 1 0 12052 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_123
timestamp 1635444444
transform 1 0 12420 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1635444444
transform 1 0 12144 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 12788 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1635444444
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1635444444
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_141
timestamp 1635444444
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_148
timestamp 1635444444
transform 1 0 14720 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1635444444
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1019_
timestamp 1635444444
transform 1 0 14168 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_157
timestamp 1635444444
transform 1 0 15548 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_164
timestamp 1635444444
transform 1 0 16192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1253_
timestamp 1635444444
transform 1 0 15916 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1371_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 16560 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _1530_
timestamp 1635444444
transform 1 0 15272 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_184
timestamp 1635444444
transform 1 0 18032 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_188
timestamp 1635444444
transform 1 0 18400 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1635444444
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1635444444
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1252_
timestamp 1635444444
transform 1 0 18492 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_197
timestamp 1635444444
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_207
timestamp 1635444444
transform 1 0 20148 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1965_
timestamp 1635444444
transform 1 0 20516 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_wb_clk_i
timestamp 1635444444
transform 1 0 19780 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_227
timestamp 1635444444
transform 1 0 21988 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_231
timestamp 1635444444
transform 1 0 22356 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_238
timestamp 1635444444
transform 1 0 23000 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1394_
timestamp 1635444444
transform 1 0 22448 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1635444444
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1635444444
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1635444444
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_257
timestamp 1635444444
transform 1 0 24748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1635444444
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1413_
timestamp 1635444444
transform 1 0 23368 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1790_
timestamp 1635444444
transform 1 0 24840 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_267
timestamp 1635444444
transform 1 0 25668 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_275
timestamp 1635444444
transform 1 0 26404 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1118_
timestamp 1635444444
transform 1 0 26036 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_287
timestamp 1635444444
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1635444444
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1635444444
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_309
timestamp 1635444444
transform 1 0 29532 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_316
timestamp 1635444444
transform 1 0 30176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1635444444
transform -1 0 30820 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1635444444
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1635444444
transform 1 0 29808 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1635444444
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1635444444
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1635444444
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1635444444
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1635444444
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1635444444
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1635444444
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1635444444
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1635444444
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1635444444
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_81
timestamp 1635444444
transform 1 0 8556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1795_
timestamp 1635444444
transform 1 0 8924 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1635444444
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_94
timestamp 1635444444
transform 1 0 9752 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1366_
timestamp 1635444444
transform 1 0 10120 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1635444444
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_120
timestamp 1635444444
transform 1 0 12144 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_127
timestamp 1635444444
transform 1 0 12788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1635444444
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1635444444
transform 1 0 12512 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1068_
timestamp 1635444444
transform 1 0 13156 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1373_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 11500 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_134
timestamp 1635444444
transform 1 0 13432 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_138
timestamp 1635444444
transform 1 0 13800 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_146
timestamp 1635444444
transform 1 0 14536 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1635444444
transform 1 0 14904 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1060_
timestamp 1635444444
transform 1 0 13892 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_153
timestamp 1635444444
transform 1 0 15180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_157
timestamp 1635444444
transform 1 0 15548 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1635444444
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_169
timestamp 1635444444
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1635444444
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _0884_
timestamp 1635444444
transform 1 0 15640 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1635444444
transform 1 0 16928 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_45_188
timestamp 1635444444
transform 1 0 18400 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1745_
timestamp 1635444444
transform 1 0 18768 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_45_201
timestamp 1635444444
transform 1 0 19596 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_209
timestamp 1635444444
transform 1 0 20332 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _0959_
timestamp 1635444444
transform 1 0 20516 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1635444444
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1635444444
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_233
timestamp 1635444444
transform 1 0 22540 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_240
timestamp 1635444444
transform 1 0 23184 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1635444444
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0957_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 22908 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_wb_clk_i
timestamp 1635444444
transform 1 0 22172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_253
timestamp 1635444444
transform 1 0 24380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1786_
timestamp 1635444444
transform 1 0 23552 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1789_
timestamp 1635444444
transform 1 0 24932 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_268
timestamp 1635444444
transform 1 0 25760 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_275
timestamp 1635444444
transform 1 0 26404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1635444444
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1635444444
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1635444444
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1436_
timestamp 1635444444
transform 1 0 26128 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1635444444
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_305
timestamp 1635444444
transform 1 0 29164 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_311
timestamp 1635444444
transform 1 0 29716 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_316
timestamp 1635444444
transform 1 0 30176 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1635444444
transform -1 0 30820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1635444444
transform 1 0 29808 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_19
timestamp 1635444444
transform 1 0 2852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_7
timestamp 1635444444
transform 1 0 1748 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1635444444
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1635444444
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1635444444
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1635444444
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1635444444
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1635444444
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1635444444
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1635444444
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1635444444
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1635444444
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1635444444
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1635444444
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_65
timestamp 1635444444
transform 1 0 7084 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1635444444
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1635444444
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1635444444
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1635444444
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_73
timestamp 1635444444
transform 1 0 7820 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_78
timestamp 1635444444
transform 1 0 8280 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1635444444
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_69
timestamp 1635444444
transform 1 0 7452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_73
timestamp 1635444444
transform 1 0 7820 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_77
timestamp 1635444444
transform 1 0 8188 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1635444444
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1361_
timestamp 1635444444
transform 1 0 7912 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1362_
timestamp 1635444444
transform 1 0 8004 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_106
timestamp 1635444444
transform 1 0 10856 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_95
timestamp 1635444444
transform 1 0 9844 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1635444444
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_89
timestamp 1635444444
transform 1 0 9292 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_94
timestamp 1635444444
transform 1 0 9752 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0920_
timestamp 1635444444
transform 1 0 9476 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1635444444
transform 1 0 9476 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0972_
timestamp 1635444444
transform 1 0 10120 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_2  _1030_
timestamp 1635444444
transform 1 0 10212 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1635444444
transform 1 0 12052 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0922_
timestamp 1635444444
transform 1 0 11684 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0890_
timestamp 1635444444
transform 1 0 11224 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1635444444
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_119
timestamp 1635444444
transform 1 0 12052 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1635444444
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_115
timestamp 1635444444
transform 1 0 11684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1365_
timestamp 1635444444
transform 1 0 12880 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_124
timestamp 1635444444
transform 1 0 12512 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1950_
timestamp 1635444444
transform 1 0 12420 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_46_132
timestamp 1635444444
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_141
timestamp 1635444444
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_146
timestamp 1635444444
transform 1 0 14536 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_139
timestamp 1635444444
transform 1 0 13892 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1635444444
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14904 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1073_
timestamp 1635444444
transform 1 0 14168 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1635444444
transform 1 0 14260 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_46_159
timestamp 1635444444
transform 1 0 15732 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_168
timestamp 1635444444
transform 1 0 16560 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1635444444
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1635444444
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1635444444
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_173
timestamp 1635444444
transform 1 0 17020 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1635444444
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1128_
timestamp 1635444444
transform 1 0 17112 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1379_
timestamp 1635444444
transform 1 0 16100 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_46_176
timestamp 1635444444
transform 1 0 17296 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1635444444
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1635444444
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_183
timestamp 1635444444
transform 1 0 17940 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1635444444
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1125_
timestamp 1635444444
transform 1 0 17480 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1127_
timestamp 1635444444
transform 1 0 18676 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_46_200
timestamp 1635444444
transform 1 0 19504 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_214
timestamp 1635444444
transform 1 0 20792 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_200
timestamp 1635444444
transform 1 0 19504 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1635444444
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0950_
timestamp 1635444444
transform 1 0 19872 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0956_
timestamp 1635444444
transform 1 0 21068 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0960_
timestamp 1635444444
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1744_
timestamp 1635444444
transform 1 0 19872 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1964_
timestamp 1635444444
transform 1 0 21160 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_46_234
timestamp 1635444444
transform 1 0 22632 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1635444444
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_234
timestamp 1635444444
transform 1 0 22632 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_238
timestamp 1635444444
transform 1 0 23000 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1635444444
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0961_
timestamp 1635444444
transform 1 0 23000 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0963_
timestamp 1635444444
transform 1 0 21804 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1421_
timestamp 1635444444
transform 1 0 23092 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1429_
timestamp 1635444444
transform 1 0 23644 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_245
timestamp 1635444444
transform 1 0 23644 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_241
timestamp 1635444444
transform 1 0 23276 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1422_
timestamp 1635444444
transform 1 0 24380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1393_
timestamp 1635444444
transform 1 0 24012 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1635444444
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_252
timestamp 1635444444
transform 1 0 24288 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1635444444
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1433_
timestamp 1635444444
transform 1 0 24656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1427_
timestamp 1635444444
transform 1 0 25024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_259
timestamp 1635444444
transform 1 0 24932 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_256
timestamp 1635444444
transform 1 0 24656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1439_
timestamp 1635444444
transform 1 0 25668 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1338_
timestamp 1635444444
transform 1 0 25576 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_269
timestamp 1635444444
transform 1 0 25852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_265
timestamp 1635444444
transform 1 0 25484 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_270
timestamp 1635444444
transform 1 0 25944 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_263
timestamp 1635444444
transform 1 0 25300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1444_
timestamp 1635444444
transform 1 0 26312 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1635444444
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 1635444444
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1635444444
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1635444444
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1635444444
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1635444444
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1635444444
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_305
timestamp 1635444444
transform 1 0 29164 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1635444444
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_309
timestamp 1635444444
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_317
timestamp 1635444444
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_311
timestamp 1635444444
transform 1 0 29716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_316
timestamp 1635444444
transform 1 0 30176 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1635444444
transform -1 0 30820 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1635444444
transform -1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1635444444
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1635444444
transform 1 0 29808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1635444444
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1635444444
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1635444444
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1635444444
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1635444444
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1635444444
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1635444444
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1635444444
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_65
timestamp 1635444444
transform 1 0 7084 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_73
timestamp 1635444444
transform 1 0 7820 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1635444444
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1635444444
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1635444444
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1635444444
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1349_
timestamp 1635444444
transform 1 0 7912 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_107
timestamp 1635444444
transform 1 0 10948 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1635444444
transform 1 0 9660 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_98
timestamp 1635444444
transform 1 0 10120 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0973_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 10488 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1635444444
transform 1 0 9844 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_115
timestamp 1635444444
transform 1 0 11684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_123
timestamp 1635444444
transform 1 0 12420 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_130
timestamp 1635444444
transform 1 0 13064 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1635444444
transform 1 0 12788 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0923_
timestamp 1635444444
transform 1 0 12052 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_wb_clk_i
timestamp 1635444444
transform 1 0 11316 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1635444444
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_141
timestamp 1635444444
transform 1 0 14076 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_145
timestamp 1635444444
transform 1 0 14444 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1635444444
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0916_
timestamp 1635444444
transform 1 0 14812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1635444444
transform 1 0 14168 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_153
timestamp 1635444444
transform 1 0 15180 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_167
timestamp 1635444444
transform 1 0 16468 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1380_
timestamp 1635444444
transform 1 0 15548 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1635444444
transform 1 0 16836 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_48_187
timestamp 1635444444
transform 1 0 18308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1635444444
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1635444444
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_213
timestamp 1635444444
transform 1 0 20700 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1635444444
transform 1 0 19228 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_48_219
timestamp 1635444444
transform 1 0 21252 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_229
timestamp 1635444444
transform 1 0 22172 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0967_
timestamp 1635444444
transform 1 0 21344 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1428_
timestamp 1635444444
transform 1 0 22724 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_241
timestamp 1635444444
transform 1 0 23276 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1635444444
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1635444444
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_260
timestamp 1635444444
transform 1 0 25024 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1635444444
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1315_
timestamp 1635444444
transform 1 0 24748 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1341_
timestamp 1635444444
transform 1 0 23644 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_268
timestamp 1635444444
transform 1 0 25760 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1635444444
transform 1 0 25944 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_48_286
timestamp 1635444444
transform 1 0 27416 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_298
timestamp 1635444444
transform 1 0 28520 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1635444444
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_309
timestamp 1635444444
transform 1 0 29532 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_316
timestamp 1635444444
transform 1 0 30176 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1635444444
transform -1 0 30820 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1635444444
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1635444444
transform 1 0 29808 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_19
timestamp 1635444444
transform 1 0 2852 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_7
timestamp 1635444444
transform 1 0 1748 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1635444444
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1635444444
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_31
timestamp 1635444444
transform 1 0 3956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_43
timestamp 1635444444
transform 1 0 5060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1635444444
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1635444444
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1635444444
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_69
timestamp 1635444444
transform 1 0 7452 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_74
timestamp 1635444444
transform 1 0 7912 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1348_
timestamp 1635444444
transform 1 0 7636 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1635444444
transform 1 0 8280 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_49_106
timestamp 1635444444
transform 1 0 10856 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_94
timestamp 1635444444
transform 1 0 9752 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 10120 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_122
timestamp 1635444444
transform 1 0 12328 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1635444444
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_2  _1313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 11500 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1741_
timestamp 1635444444
transform 1 0 12696 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_135
timestamp 1635444444
transform 1 0 13524 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_143
timestamp 1635444444
transform 1 0 14260 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1725_
timestamp 1635444444
transform 1 0 14812 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_wb_clk_i
timestamp 1635444444
transform 1 0 13892 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_154
timestamp 1635444444
transform 1 0 15272 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1635444444
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1635444444
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1650_
timestamp 1635444444
transform 1 0 16652 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _1705_
timestamp 1635444444
transform 1 0 15640 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_179
timestamp 1635444444
transform 1 0 17572 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_188
timestamp 1635444444
transform 1 0 18400 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_195
timestamp 1635444444
transform 1 0 19044 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0965_
timestamp 1635444444
transform 1 0 18768 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1507_
timestamp 1635444444
transform 1 0 18124 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_202
timestamp 1635444444
transform 1 0 19688 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_209
timestamp 1635444444
transform 1 0 20332 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1635444444
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0947_
timestamp 1635444444
transform 1 0 20056 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0964_
timestamp 1635444444
transform 1 0 19412 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1635444444
transform 1 0 20700 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1635444444
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1635444444
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1635444444
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1635444444
transform 1 0 21988 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_49_243
timestamp 1635444444
transform 1 0 23460 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_253
timestamp 1635444444
transform 1 0 24380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1337_
timestamp 1635444444
transform 1 0 24748 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1382_
timestamp 1635444444
transform 1 0 23828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_266
timestamp 1635444444
transform 1 0 25576 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1635444444
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1635444444
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1635444444
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1335_
timestamp 1635444444
transform 1 0 25944 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1336_
timestamp 1635444444
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_284
timestamp 1635444444
transform 1 0 27232 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_291
timestamp 1635444444
transform 1 0 27876 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1339_
timestamp 1635444444
transform 1 0 27600 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1448_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 28612 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_49_306
timestamp 1635444444
transform 1 0 29256 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_316
timestamp 1635444444
transform 1 0 30176 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1635444444
transform -1 0 30820 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1635444444
transform 1 0 29808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1635444444
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1635444444
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1635444444
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1635444444
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1635444444
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1635444444
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1635444444
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1635444444
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1635444444
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1635444444
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1635444444
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1635444444
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1351_
timestamp 1635444444
transform 1 0 8188 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_105
timestamp 1635444444
transform 1 0 10764 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_89
timestamp 1635444444
transform 1 0 9292 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_98
timestamp 1635444444
transform 1 0 10120 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _0975_
timestamp 1635444444
transform 1 0 11132 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1635444444
transform 1 0 10488 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1346_
timestamp 1635444444
transform 1 0 9384 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_118
timestamp 1635444444
transform 1 0 11960 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_126
timestamp 1635444444
transform 1 0 12696 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__a221o_1  _0917_
timestamp 1635444444
transform 1 0 12880 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1635444444
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_144
timestamp 1635444444
transform 1 0 14352 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1635444444
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1635444444
transform 1 0 14076 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1090_
timestamp 1635444444
transform 1 0 14904 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_156
timestamp 1635444444
transform 1 0 15456 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_163
timestamp 1635444444
transform 1 0 16100 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1369_
timestamp 1635444444
transform 1 0 15824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1706_
timestamp 1635444444
transform 1 0 16468 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_50_176
timestamp 1635444444
transform 1 0 17296 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_182
timestamp 1635444444
transform 1 0 17848 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_186
timestamp 1635444444
transform 1 0 18216 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1635444444
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1635444444
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1575_
timestamp 1635444444
transform 1 0 17940 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_197
timestamp 1635444444
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_203
timestamp 1635444444
transform 1 0 19780 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_210
timestamp 1635444444
transform 1 0 20424 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_217
timestamp 1635444444
transform 1 0 21068 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1635444444
transform 1 0 20792 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0945_
timestamp 1635444444
transform 1 0 20148 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0952_
timestamp 1635444444
transform 1 0 19504 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_231
timestamp 1635444444
transform 1 0 22356 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_240
timestamp 1635444444
transform 1 0 23184 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0932_
timestamp 1635444444
transform 1 0 21436 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _1333_
timestamp 1635444444
transform 1 0 22908 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1635444444
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1635444444
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_257
timestamp 1635444444
transform 1 0 24748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1635444444
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1340_
timestamp 1635444444
transform 1 0 24840 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1381_
timestamp 1635444444
transform 1 0 23552 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_267
timestamp 1635444444
transform 1 0 25668 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1635444444
transform 1 0 26036 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_50_287
timestamp 1635444444
transform 1 0 27508 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_295
timestamp 1635444444
transform 1 0 28244 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1635444444
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1446_
timestamp 1635444444
transform 1 0 28428 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_50_309
timestamp 1635444444
transform 1 0 29532 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_316
timestamp 1635444444
transform 1 0 30176 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1635444444
transform -1 0 30820 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1635444444
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1635444444
transform 1 0 29808 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1635444444
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1635444444
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1635444444
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1635444444
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1635444444
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1635444444
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1635444444
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1635444444
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1635444444
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1635444444
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_81
timestamp 1635444444
transform 1 0 8556 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_87
timestamp 1635444444
transform 1 0 9108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1347_
timestamp 1635444444
transform 1 0 8832 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_104
timestamp 1635444444
transform 1 0 10672 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _1345_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9844 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_122
timestamp 1635444444
transform 1 0 12328 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1635444444
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1355_
timestamp 1635444444
transform 1 0 11500 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1740_
timestamp 1635444444
transform 1 0 12696 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_51_135
timestamp 1635444444
transform 1 0 13524 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_143
timestamp 1635444444
transform 1 0 14260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1635444444
transform 1 0 14444 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1635444444
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1635444444
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_169
timestamp 1635444444
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1635444444
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1668_
timestamp 1635444444
transform 1 0 17020 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_182
timestamp 1635444444
transform 1 0 17848 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_195
timestamp 1635444444
transform 1 0 19044 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1726_
timestamp 1635444444
transform 1 0 18216 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_51_203
timestamp 1635444444
transform 1 0 19780 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_211
timestamp 1635444444
transform 1 0 20516 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1635444444
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0946_
timestamp 1635444444
transform 1 0 20700 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1085_
timestamp 1635444444
transform 1 0 19412 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_225
timestamp 1635444444
transform 1 0 21804 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1635444444
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1967_
timestamp 1635444444
transform 1 0 22080 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_51_244
timestamp 1635444444
transform 1 0 23552 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_252
timestamp 1635444444
transform 1 0 24288 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_262
timestamp 1635444444
transform 1 0 25208 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1334_
timestamp 1635444444
transform 1 0 24380 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1635444444
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1635444444
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1314_
timestamp 1635444444
transform 1 0 25576 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1331_
timestamp 1635444444
transform 1 0 26956 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_290
timestamp 1635444444
transform 1 0 27784 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_297
timestamp 1635444444
transform 1 0 28428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1330_
timestamp 1635444444
transform 1 0 28152 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1447_
timestamp 1635444444
transform 1 0 29164 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_308
timestamp 1635444444
transform 1 0 29440 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_316
timestamp 1635444444
transform 1 0 30176 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1635444444
transform -1 0 30820 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1635444444
transform 1 0 29808 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1635444444
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1635444444
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_13
timestamp 1635444444
transform 1 0 2300 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1635444444
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1635444444
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1635444444
transform 1 0 1380 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1635444444
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1635444444
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1635444444
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_25
timestamp 1635444444
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_37
timestamp 1635444444
transform 1 0 4508 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1635444444
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1635444444
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1635444444
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_49
timestamp 1635444444
transform 1 0 5612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1635444444
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1635444444
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1635444444
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1635444444
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1635444444
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1635444444
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_69
timestamp 1635444444
transform 1 0 7452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_73
timestamp 1635444444
transform 1 0 7820 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_77
timestamp 1635444444
transform 1 0 8188 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1635444444
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1342_
timestamp 1635444444
transform 1 0 7912 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1635444444
transform 1 0 8556 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_52_107
timestamp 1635444444
transform 1 0 10948 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_93
timestamp 1635444444
transform 1 0 9660 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_98
timestamp 1635444444
transform 1 0 10120 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1635444444
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_97
timestamp 1635444444
transform 1 0 10028 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0928_
timestamp 1635444444
transform 1 0 10580 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1312_
timestamp 1635444444
transform 1 0 10488 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1344_
timestamp 1635444444
transform 1 0 9844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1635444444
transform 1 0 12144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1354_
timestamp 1635444444
transform 1 0 11592 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1343_
timestamp 1635444444
transform 1 0 11408 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1635444444
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_117
timestamp 1635444444
transform 1 0 11868 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_113
timestamp 1635444444
transform 1 0 11500 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_116
timestamp 1635444444
transform 1 0 11776 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_111
timestamp 1635444444
transform 1 0 11316 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _1742_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 12236 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1635444444
transform 1 0 12880 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_52_124
timestamp 1635444444
transform 1 0 12512 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_130
timestamp 1635444444
transform 1 0 13064 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1635444444
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1635444444
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_142
timestamp 1635444444
transform 1 0 14168 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_150
timestamp 1635444444
transform 1 0 14904 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1635444444
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1972_
timestamp 1635444444
transform 1 0 14076 0 1 30464
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_52_160
timestamp 1635444444
transform 1 0 15824 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_172
timestamp 1635444444
transform 1 0 16928 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_158
timestamp 1635444444
transform 1 0 15640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1635444444
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1635444444
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1635444444
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1656_
timestamp 1635444444
transform 1 0 17020 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1715_
timestamp 1635444444
transform 1 0 15180 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_52_182
timestamp 1635444444
transform 1 0 17848 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1635444444
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_190
timestamp 1635444444
transform 1 0 18584 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1635444444
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_1  _1655_
timestamp 1635444444
transform 1 0 18216 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _1678_
timestamp 1635444444
transform 1 0 18952 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1679_
timestamp 1635444444
transform 1 0 17756 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_52_203
timestamp 1635444444
transform 1 0 19780 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_200
timestamp 1635444444
transform 1 0 19504 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_208
timestamp 1635444444
transform 1 0 20240 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_212
timestamp 1635444444
transform 1 0 20608 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0953_
timestamp 1635444444
transform 1 0 20332 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _1667_
timestamp 1635444444
transform 1 0 19228 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1966_
timestamp 1635444444
transform 1 0 20332 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1635444444
transform 1 0 20976 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_225
timestamp 1635444444
transform 1 0 21804 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_238
timestamp 1635444444
transform 1 0 23000 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1635444444
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_234
timestamp 1635444444
transform 1 0 22632 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1635444444
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0908_
timestamp 1635444444
transform 1 0 23000 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0951_
timestamp 1635444444
transform 1 0 22172 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _0955_
timestamp 1635444444
transform 1 0 21804 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1328_
timestamp 1635444444
transform 1 0 23552 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1320_
timestamp 1635444444
transform 1 0 23920 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_53_247
timestamp 1635444444
transform 1 0 23828 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_241
timestamp 1635444444
transform 1 0 23276 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1635444444
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_247
timestamp 1635444444
transform 1 0 23828 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1635444444
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_258
timestamp 1635444444
transform 1 0 24840 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1635444444
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1635444444
transform 1 0 24564 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_52_271
timestamp 1635444444
transform 1 0 26036 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_278
timestamp 1635444444
transform 1 0 26680 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_274
timestamp 1635444444
transform 1 0 26312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1635444444
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1635444444
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1316_
timestamp 1635444444
transform 1 0 25392 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _1329_
timestamp 1635444444
transform 1 0 26404 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1635444444
transform 1 0 27048 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1635444444
transform 1 0 27140 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_52_298
timestamp 1635444444
transform 1 0 28520 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_299
timestamp 1635444444
transform 1 0 28612 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1450_
timestamp 1635444444
transform 1 0 28980 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1635444444
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_316
timestamp 1635444444
transform 1 0 30176 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_310
timestamp 1635444444
transform 1 0 29624 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_318
timestamp 1635444444
transform 1 0 30360 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1635444444
transform -1 0 30820 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1635444444
transform -1 0 30820 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1635444444
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _1452_
timestamp 1635444444
transform 1 0 29532 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1635444444
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1635444444
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1635444444
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1635444444
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1635444444
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1635444444
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1635444444
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1635444444
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1635444444
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1635444444
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1635444444
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1635444444
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1635444444
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_104
timestamp 1635444444
transform 1 0 10672 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_97
timestamp 1635444444
transform 1 0 10028 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1635444444
transform 1 0 11040 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1523_
timestamp 1635444444
transform 1 0 10120 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_111
timestamp 1635444444
transform 1 0 11316 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_115
timestamp 1635444444
transform 1 0 11684 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_125
timestamp 1635444444
transform 1 0 12604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1737_
timestamp 1635444444
transform 1 0 11776 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_54_137
timestamp 1635444444
transform 1 0 13708 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1635444444
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1635444444
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_153
timestamp 1635444444
transform 1 0 15180 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_162
timestamp 1635444444
transform 1 0 16008 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1666_
timestamp 1635444444
transform 1 0 15732 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1716_
timestamp 1635444444
transform 1 0 16376 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_54_175
timestamp 1635444444
transform 1 0 17204 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_187
timestamp 1635444444
transform 1 0 18308 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1635444444
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1635444444
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1072_
timestamp 1635444444
transform 1 0 18400 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_197
timestamp 1635444444
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_203
timestamp 1635444444
transform 1 0 19780 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_207
timestamp 1635444444
transform 1 0 20148 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_215
timestamp 1635444444
transform 1 0 20884 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0933_
timestamp 1635444444
transform 1 0 21068 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1724_
timestamp 1635444444
transform 1 0 19872 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_227
timestamp 1635444444
transform 1 0 21988 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_240
timestamp 1635444444
transform 1 0 23184 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0939_
timestamp 1635444444
transform 1 0 22356 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_54_244
timestamp 1635444444
transform 1 0 23552 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1635444444
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_259
timestamp 1635444444
transform 1 0 24932 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1635444444
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1332_
timestamp 1635444444
transform 1 0 23644 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1440_
timestamp 1635444444
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_267
timestamp 1635444444
transform 1 0 25668 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_271
timestamp 1635444444
transform 1 0 26036 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1326_
timestamp 1635444444
transform 1 0 25760 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1327_
timestamp 1635444444
transform 1 0 26404 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_54_284
timestamp 1635444444
transform 1 0 27232 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_292
timestamp 1635444444
transform 1 0 27968 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_297
timestamp 1635444444
transform 1 0 28428 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1635444444
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1451_
timestamp 1635444444
transform 1 0 28796 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1453_
timestamp 1635444444
transform 1 0 28152 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_309
timestamp 1635444444
transform 1 0 29532 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_316
timestamp 1635444444
transform 1 0 30176 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1635444444
transform -1 0 30820 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1635444444
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1635444444
transform 1 0 29808 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1635444444
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1635444444
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1635444444
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1635444444
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1635444444
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1635444444
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1635444444
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1635444444
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1635444444
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1635444444
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1635444444
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_104
timestamp 1635444444
transform 1 0 10672 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_93
timestamp 1635444444
transform 1 0 9660 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1734_
timestamp 1635444444
transform 1 0 9844 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_55_113
timestamp 1635444444
transform 1 0 11500 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_117
timestamp 1635444444
transform 1 0 11868 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_130
timestamp 1635444444
transform 1 0 13064 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1635444444
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0924_
timestamp 1635444444
transform 1 0 12236 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1635444444
transform 1 0 11592 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_141
timestamp 1635444444
transform 1 0 14076 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _1044_
timestamp 1635444444
transform 1 0 13432 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1121_
timestamp 1635444444
transform 1 0 14444 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_55_154
timestamp 1635444444
transform 1 0 15272 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1635444444
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_169
timestamp 1635444444
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1635444444
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1113_
timestamp 1635444444
transform 1 0 15824 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1635444444
transform 1 0 17020 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_177
timestamp 1635444444
transform 1 0 17388 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1635444444
transform 1 0 18032 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_196
timestamp 1635444444
transform 1 0 19136 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1651_
timestamp 1635444444
transform 1 0 17756 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_213
timestamp 1635444444
transform 1 0 20700 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0940_
timestamp 1635444444
transform 1 0 21068 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1635444444
transform 1 0 19228 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1635444444
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1635444444
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_237
timestamp 1635444444
transform 1 0 22908 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1635444444
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0935_
timestamp 1635444444
transform 1 0 22080 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_55_244
timestamp 1635444444
transform 1 0 23552 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_252
timestamp 1635444444
transform 1 0 24288 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_260
timestamp 1635444444
transform 1 0 25024 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0936_
timestamp 1635444444
transform 1 0 23276 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1435_
timestamp 1635444444
transform 1 0 24472 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_269
timestamp 1635444444
transform 1 0 25852 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1635444444
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1635444444
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1322_
timestamp 1635444444
transform 1 0 26220 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1324_
timestamp 1635444444
transform 1 0 26956 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1325_
timestamp 1635444444
transform 1 0 25576 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_290
timestamp 1635444444
transform 1 0 27784 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_294
timestamp 1635444444
transform 1 0 28152 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_298
timestamp 1635444444
transform 1 0 28520 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1635444444
transform 1 0 28244 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1455_
timestamp 1635444444
transform 1 0 28888 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_55_309
timestamp 1635444444
transform 1 0 29532 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_316
timestamp 1635444444
transform 1 0 30176 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1635444444
transform -1 0 30820 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1449_
timestamp 1635444444
transform 1 0 29900 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1635444444
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1635444444
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1635444444
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1635444444
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1635444444
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1635444444
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1635444444
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1635444444
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1635444444
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1635444444
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1635444444
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_85
timestamp 1635444444
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1635444444
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_102
timestamp 1635444444
transform 1 0 10488 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_108
timestamp 1635444444
transform 1 0 11040 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_92
timestamp 1635444444
transform 1 0 9568 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_2  _0930_
timestamp 1635444444
transform 1 0 11132 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1222_
timestamp 1635444444
transform 1 0 9292 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1522_
timestamp 1635444444
transform 1 0 9936 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_116
timestamp 1635444444
transform 1 0 11776 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1971_
timestamp 1635444444
transform 1 0 12144 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1635444444
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_141
timestamp 1635444444
transform 1 0 14076 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1635444444
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1635444444
transform 1 0 14168 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_56_158
timestamp 1635444444
transform 1 0 15640 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1635444444
transform 1 0 16376 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_182
timestamp 1635444444
transform 1 0 17848 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1635444444
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1635444444
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1635444444
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1677_
timestamp 1635444444
transform 1 0 18216 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1635444444
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_216
timestamp 1635444444
transform 1 0 20976 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1635444444
transform 1 0 19504 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_56_224
timestamp 1635444444
transform 1 0 21712 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_228
timestamp 1635444444
transform 1 0 22080 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0937_
timestamp 1635444444
transform 1 0 21804 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1635444444
transform 1 0 22448 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1635444444
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_256
timestamp 1635444444
transform 1 0 24656 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1635444444
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1434_
timestamp 1635444444
transform 1 0 25024 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1635444444
transform 1 0 24380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_270
timestamp 1635444444
transform 1 0 25944 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_277
timestamp 1635444444
transform 1 0 26588 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_283
timestamp 1635444444
transform 1 0 27140 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1318_
timestamp 1635444444
transform 1 0 26312 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_300
timestamp 1635444444
transform 1 0 28704 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1635444444
transform 1 0 27232 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_56_309
timestamp 1635444444
transform 1 0 29532 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_316
timestamp 1635444444
transform 1 0 30176 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1635444444
transform -1 0 30820 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1635444444
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1635444444
transform 1 0 29808 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_18
timestamp 1635444444
transform 1 0 2760 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_6
timestamp 1635444444
transform 1 0 1656 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1635444444
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1635444444
transform 1 0 1380 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_30
timestamp 1635444444
transform 1 0 3864 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_42
timestamp 1635444444
transform 1 0 4968 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1635444444
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1635444444
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1635444444
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1635444444
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1635444444
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_102
timestamp 1635444444
transform 1 0 10488 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1758_
timestamp 1635444444
transform 1 0 9660 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1635444444
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_120
timestamp 1635444444
transform 1 0 12144 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_128
timestamp 1635444444
transform 1 0 12880 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1635444444
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_2  _1223_
timestamp 1635444444
transform 1 0 11500 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1635444444
transform 1 0 12512 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_135
timestamp 1635444444
transform 1 0 13524 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_142
timestamp 1635444444
transform 1 0 14168 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_150
timestamp 1635444444
transform 1 0 14904 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0918_
timestamp 1635444444
transform 1 0 13248 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0919_
timestamp 1635444444
transform 1 0 13892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1120_
timestamp 1635444444
transform 1 0 14996 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_57_160
timestamp 1635444444
transform 1 0 15824 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1635444444
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1123_
timestamp 1635444444
transform 1 0 16652 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_178
timestamp 1635444444
transform 1 0 17480 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_182
timestamp 1635444444
transform 1 0 17848 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1944_
timestamp 1635444444
transform 1 0 17940 0 -1 33728
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_57_202
timestamp 1635444444
transform 1 0 19688 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_210
timestamp 1635444444
transform 1 0 20424 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0943_
timestamp 1635444444
transform 1 0 20516 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1635444444
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_225
timestamp 1635444444
transform 1 0 21804 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_231
timestamp 1635444444
transform 1 0 22356 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1635444444
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0925_
timestamp 1635444444
transform 1 0 22080 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1970_
timestamp 1635444444
transform 1 0 22724 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_57_251
timestamp 1635444444
transform 1 0 24196 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_258
timestamp 1635444444
transform 1 0 24840 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1248_
timestamp 1635444444
transform 1 0 24564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1635444444
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1635444444
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_281
timestamp 1635444444
transform 1 0 26956 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1635444444
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1317_
timestamp 1635444444
transform 1 0 25392 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_300
timestamp 1635444444
transform 1 0 28704 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1323_
timestamp 1635444444
transform 1 0 29072 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1635444444
transform 1 0 27232 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_57_307
timestamp 1635444444
transform 1 0 29348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_311
timestamp 1635444444
transform 1 0 29716 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_316
timestamp 1635444444
transform 1 0 30176 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1635444444
transform -1 0 30820 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1635444444
transform 1 0 29808 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1635444444
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1635444444
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1635444444
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1635444444
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1635444444
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1635444444
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1635444444
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1635444444
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1635444444
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1635444444
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1635444444
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1635444444
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1635444444
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_101
timestamp 1635444444
transform 1 0 10396 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_108
timestamp 1635444444
transform 1 0 11040 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_97
timestamp 1635444444
transform 1 0 10028 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1221_
timestamp 1635444444
transform 1 0 10120 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1353_
timestamp 1635444444
transform 1 0 10764 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_115
timestamp 1635444444
transform 1 0 11684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_125
timestamp 1635444444
transform 1 0 12604 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0948_
timestamp 1635444444
transform 1 0 11408 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0966_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 12052 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1635444444
transform 1 0 12972 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1635444444
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1635444444
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_141
timestamp 1635444444
transform 1 0 14076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_147
timestamp 1635444444
transform 1 0 14628 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_151
timestamp 1635444444
transform 1 0 14996 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1635444444
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1690_
timestamp 1635444444
transform 1 0 14720 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_171
timestamp 1635444444
transform 1 0 16836 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1635444444
transform 1 0 15364 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_58_175
timestamp 1635444444
transform 1 0 17204 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_179
timestamp 1635444444
transform 1 0 17572 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1635444444
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1635444444
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1089_
timestamp 1635444444
transform 1 0 17940 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1665_
timestamp 1635444444
transform 1 0 17296 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_197
timestamp 1635444444
transform 1 0 19228 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_207
timestamp 1635444444
transform 1 0 20148 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_214
timestamp 1635444444
transform 1 0 20792 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0941_
timestamp 1635444444
transform 1 0 20516 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1093_
timestamp 1635444444
transform 1 0 19320 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1968_
timestamp 1635444444
transform 1 0 21160 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_234
timestamp 1635444444
transform 1 0 22632 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0926_
timestamp 1635444444
transform 1 0 23000 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_241
timestamp 1635444444
transform 1 0 23276 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_249
timestamp 1635444444
transform 1 0 24012 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1635444444
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_258
timestamp 1635444444
transform 1 0 24840 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1635444444
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1249_
timestamp 1635444444
transform 1 0 24564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1635444444
transform 1 0 25208 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_278
timestamp 1635444444
transform 1 0 26680 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1321_
timestamp 1635444444
transform 1 0 27048 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_58_291
timestamp 1635444444
transform 1 0 27876 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_299
timestamp 1635444444
transform 1 0 28612 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1635444444
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1635444444
transform 1 0 28704 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_316
timestamp 1635444444
transform 1 0 30176 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1635444444
transform -1 0 30820 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1635444444
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _1458_
timestamp 1635444444
transform 1 0 29532 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1635444444
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1635444444
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_18
timestamp 1635444444
transform 1 0 2760 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_6
timestamp 1635444444
transform 1 0 1656 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1635444444
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1635444444
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1635444444
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1635444444
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1635444444
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1635444444
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1635444444
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1635444444
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1635444444
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1635444444
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1635444444
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1635444444
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1635444444
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1635444444
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1635444444
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1635444444
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1635444444
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1635444444
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1635444444
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1635444444
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1635444444
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_101
timestamp 1635444444
transform 1 0 10396 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_106
timestamp 1635444444
transform 1 0 10856 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_93
timestamp 1635444444
transform 1 0 9660 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_105
timestamp 1635444444
transform 1 0 10764 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_109
timestamp 1635444444
transform 1 0 11132 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_97
timestamp 1635444444
transform 1 0 10028 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0921_
timestamp 1635444444
transform 1 0 10488 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1352_
timestamp 1635444444
transform 1 0 10856 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_130
timestamp 1635444444
transform 1 0 13064 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_117
timestamp 1635444444
transform 1 0 11868 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_125
timestamp 1635444444
transform 1 0 12604 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1635444444
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0962_
timestamp 1635444444
transform 1 0 12052 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1828_
timestamp 1635444444
transform 1 0 11500 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_59_150
timestamp 1635444444
transform 1 0 14904 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_136
timestamp 1635444444
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1635444444
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_149
timestamp 1635444444
transform 1 0 14812 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1635444444
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1702_
timestamp 1635444444
transform 1 0 13340 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1635444444
transform 1 0 13432 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_wb_clk_i
timestamp 1635444444
transform 1 0 14444 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_163
timestamp 1635444444
transform 1 0 16100 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1635444444
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_169
timestamp 1635444444
transform 1 0 16652 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_155
timestamp 1635444444
transform 1 0 15364 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_172
timestamp 1635444444
transform 1 0 16928 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1635444444
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1119_
timestamp 1635444444
transform 1 0 15272 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1635444444
transform 1 0 15456 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_59_183
timestamp 1635444444
transform 1 0 17940 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_196
timestamp 1635444444
transform 1 0 19136 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_184
timestamp 1635444444
transform 1 0 18032 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1635444444
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1635444444
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1094_
timestamp 1635444444
transform 1 0 18308 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _1683_
timestamp 1635444444
transform 1 0 17204 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1691_
timestamp 1635444444
transform 1 0 17296 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_wb_clk_i
timestamp 1635444444
transform 1 0 18400 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_209
timestamp 1635444444
transform 1 0 20332 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_213
timestamp 1635444444
transform 1 0 20700 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_218
timestamp 1635444444
transform 1 0 21160 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_207
timestamp 1635444444
transform 1 0 20148 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1092_
timestamp 1635444444
transform 1 0 19504 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1095_
timestamp 1635444444
transform 1 0 19228 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1096_
timestamp 1635444444
transform 1 0 20516 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1635444444
transform 1 0 20792 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_wb_clk_i
timestamp 1635444444
transform 1 0 21712 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1635444444
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_220
timestamp 1635444444
transform 1 0 21344 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_225
timestamp 1635444444
transform 1 0 21804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0944_
timestamp 1635444444
transform 1 0 22356 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_228
timestamp 1635444444
transform 1 0 22080 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1682_
timestamp 1635444444
transform 1 0 23000 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906__1
timestamp 1635444444
transform 1 0 22632 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_237
timestamp 1635444444
transform 1 0 22908 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_234
timestamp 1635444444
transform 1 0 22632 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  net99_2
timestamp 1635444444
transform 1 0 23276 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1240_
timestamp 1635444444
transform 1 0 23736 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1635444444
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_250
timestamp 1635444444
transform 1 0 24104 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_245
timestamp 1635444444
transform 1 0 23644 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_241
timestamp 1635444444
transform 1 0 23276 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1250_
timestamp 1635444444
transform 1 0 24472 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1005_
timestamp 1635444444
transform 1 0 24380 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1635444444
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_257
timestamp 1635444444
transform 1 0 24748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1310_
timestamp 1635444444
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_262
timestamp 1635444444
transform 1 0 25208 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1635444444
transform 1 0 25760 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1311_
timestamp 1635444444
transform 1 0 25760 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_264
timestamp 1635444444
transform 1 0 25392 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0990_
timestamp 1635444444
transform 1 0 26404 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_278
timestamp 1635444444
transform 1 0 26680 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_271
timestamp 1635444444
transform 1 0 26036 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1635444444
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_271
timestamp 1635444444
transform 1 0 26036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1319_
timestamp 1635444444
transform 1 0 26956 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1635444444
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1459_
timestamp 1635444444
transform 1 0 27416 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1456_
timestamp 1635444444
transform 1 0 27600 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_289
timestamp 1635444444
transform 1 0 27692 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_291
timestamp 1635444444
transform 1 0 27876 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_284
timestamp 1635444444
transform 1 0 27232 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1635444444
transform 1 0 28244 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1635444444
transform 1 0 28060 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_296
timestamp 1635444444
transform 1 0 28336 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_299
timestamp 1635444444
transform 1 0 28612 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1635444444
transform 1 0 28704 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1460_
timestamp 1635444444
transform 1 0 28980 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1635444444
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_310
timestamp 1635444444
transform 1 0 29624 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_318
timestamp 1635444444
transform 1 0 30360 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_316
timestamp 1635444444
transform 1 0 30176 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1635444444
transform -1 0 30820 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1635444444
transform -1 0 30820 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1635444444
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _1462_
timestamp 1635444444
transform 1 0 29532 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1635444444
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1635444444
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1635444444
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1635444444
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1635444444
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1635444444
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1635444444
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1635444444
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1635444444
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1635444444
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_81
timestamp 1635444444
transform 1 0 8556 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_85
timestamp 1635444444
transform 1 0 8924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1635444444
transform 1 0 9016 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_61_102
timestamp 1635444444
transform 1 0 10488 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1635444444
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_113
timestamp 1635444444
transform 1 0 11500 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_125
timestamp 1635444444
transform 1 0 12604 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1635444444
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0958_
timestamp 1635444444
transform 1 0 12052 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1945_
timestamp 1635444444
transform 1 0 12972 0 -1 35904
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_61_148
timestamp 1635444444
transform 1 0 14720 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1114_
timestamp 1635444444
transform 1 0 15088 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1635444444
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1635444444
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1635444444
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1106_
timestamp 1635444444
transform 1 0 16652 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_61_179
timestamp 1635444444
transform 1 0 17572 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_186
timestamp 1635444444
transform 1 0 18216 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1091_
timestamp 1635444444
transform 1 0 18584 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1505_
timestamp 1635444444
transform 1 0 17940 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_200
timestamp 1635444444
transform 1 0 19504 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1635444444
transform 1 0 19872 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1635444444
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1635444444
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_231
timestamp 1635444444
transform 1 0 22356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_236
timestamp 1635444444
transform 1 0 22816 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1635444444
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0907_
timestamp 1635444444
transform 1 0 23184 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0980_
timestamp 1635444444
transform 1 0 22448 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_243
timestamp 1635444444
transform 1 0 23460 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_247
timestamp 1635444444
transform 1 0 23828 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1635444444
transform 1 0 23920 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_61_264
timestamp 1635444444
transform 1 0 25392 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_271
timestamp 1635444444
transform 1 0 26036 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1635444444
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1635444444
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0968_
timestamp 1635444444
transform 1 0 25760 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0989_
timestamp 1635444444
transform 1 0 26956 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_284
timestamp 1635444444
transform 1 0 27232 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_291
timestamp 1635444444
transform 1 0 27876 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_300
timestamp 1635444444
transform 1 0 28704 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0992_
timestamp 1635444444
transform 1 0 27600 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1454_
timestamp 1635444444
transform 1 0 28428 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1464_
timestamp 1635444444
transform 1 0 29072 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_61_311
timestamp 1635444444
transform 1 0 29716 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_319
timestamp 1635444444
transform 1 0 30452 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1635444444
transform -1 0 30820 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1635444444
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1635444444
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1635444444
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1635444444
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1635444444
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1635444444
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1635444444
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1635444444
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1635444444
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1635444444
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1635444444
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1635444444
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1635444444
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_97
timestamp 1635444444
transform 1 0 10028 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1821_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 10580 0 1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_62_121
timestamp 1635444444
transform 1 0 12236 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1084_
timestamp 1635444444
transform 1 0 12788 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1635444444
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1635444444
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_145
timestamp 1635444444
transform 1 0 14444 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1635444444
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1635444444
transform 1 0 14536 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_162
timestamp 1635444444
transform 1 0 16008 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_170
timestamp 1635444444
transform 1 0 16744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1635444444
transform 1 0 16836 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_187
timestamp 1635444444
transform 1 0 18308 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1635444444
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1635444444
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_197
timestamp 1635444444
transform 1 0 19228 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_204
timestamp 1635444444
transform 1 0 19872 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1079_
timestamp 1635444444
transform 1 0 19504 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1635444444
transform 1 0 20240 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_62_224
timestamp 1635444444
transform 1 0 21712 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_232
timestamp 1635444444
transform 1 0 22448 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_240
timestamp 1635444444
transform 1 0 23184 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0998_
timestamp 1635444444
transform 1 0 22080 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1083_
timestamp 1635444444
transform 1 0 22816 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1635444444
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1635444444
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1635444444
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_258
timestamp 1635444444
transform 1 0 24840 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1635444444
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1635444444
transform 1 0 24564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1004_
timestamp 1635444444
transform 1 0 23552 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_274
timestamp 1635444444
transform 1 0 26312 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0976_
timestamp 1635444444
transform 1 0 25392 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1958_
timestamp 1635444444
transform 1 0 26864 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_62_296
timestamp 1635444444
transform 1 0 28336 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1635444444
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1635444444
transform 1 0 28704 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_309
timestamp 1635444444
transform 1 0 29532 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_316
timestamp 1635444444
transform 1 0 30176 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1635444444
transform -1 0 30820 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1635444444
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1635444444
transform 1 0 29808 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1635444444
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1635444444
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1635444444
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1635444444
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1635444444
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1635444444
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1635444444
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1635444444
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1635444444
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1635444444
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_81
timestamp 1635444444
transform 1 0 8556 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1078_
timestamp 1635444444
transform 1 0 8648 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_63_104
timestamp 1635444444
transform 1 0 10672 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_91
timestamp 1635444444
transform 1 0 9476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1076_
timestamp 1635444444
transform 1 0 9844 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_63_113
timestamp 1635444444
transform 1 0 11500 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_118
timestamp 1635444444
transform 1 0 11960 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1635444444
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1075_
timestamp 1635444444
transform 1 0 12328 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_wb_clk_i
timestamp 1635444444
transform 1 0 11592 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_132
timestamp 1635444444
transform 1 0 13248 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_146
timestamp 1635444444
transform 1 0 14536 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1074_
timestamp 1635444444
transform 1 0 13616 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1108_
timestamp 1635444444
transform 1 0 14904 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_63_160
timestamp 1635444444
transform 1 0 15824 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_169
timestamp 1635444444
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1635444444
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1107_
timestamp 1635444444
transform 1 0 17020 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_63_182
timestamp 1635444444
transform 1 0 17848 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_190
timestamp 1635444444
transform 1 0 18584 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1088_
timestamp 1635444444
transform 1 0 18768 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_63_202
timestamp 1635444444
transform 1 0 19688 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_216
timestamp 1635444444
transform 1 0 20976 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1099_
timestamp 1635444444
transform 1 0 20056 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1635444444
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_230
timestamp 1635444444
transform 1 0 22264 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1635444444
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1002_
timestamp 1635444444
transform 1 0 22632 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1003_
timestamp 1635444444
transform 1 0 21988 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_243
timestamp 1635444444
transform 1 0 23460 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1635444444
transform 1 0 23828 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_263
timestamp 1635444444
transform 1 0 25300 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1635444444
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1635444444
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0991_
timestamp 1635444444
transform 1 0 25668 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1635444444
transform 1 0 26956 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_63_297
timestamp 1635444444
transform 1 0 28428 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_303
timestamp 1635444444
transform 1 0 28980 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _1467_
timestamp 1635444444
transform 1 0 29072 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_63_311
timestamp 1635444444
transform 1 0 29716 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_319
timestamp 1635444444
transform 1 0 30452 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1635444444
transform -1 0 30820 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_18
timestamp 1635444444
transform 1 0 2760 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_6
timestamp 1635444444
transform 1 0 1656 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1635444444
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1635444444
transform 1 0 1380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1635444444
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1635444444
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1635444444
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1635444444
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1635444444
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1635444444
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1635444444
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1635444444
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1635444444
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1635444444
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_97
timestamp 1635444444
transform 1 0 10028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1635444444
transform 1 0 10396 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_64_117
timestamp 1635444444
transform 1 0 11868 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1080_
timestamp 1635444444
transform 1 0 12420 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_64_132
timestamp 1635444444
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1635444444
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_149
timestamp 1635444444
transform 1 0 14812 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1635444444
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1116_
timestamp 1635444444
transform 1 0 14904 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_64_159
timestamp 1635444444
transform 1 0 15732 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_165
timestamp 1635444444
transform 1 0 16284 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_170
timestamp 1635444444
transform 1 0 16744 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1115_
timestamp 1635444444
transform 1 0 16376 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1714_
timestamp 1635444444
transform 1 0 17112 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_177
timestamp 1635444444
transform 1 0 17388 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1635444444
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1635444444
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1635444444
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1103_
timestamp 1635444444
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_207
timestamp 1635444444
transform 1 0 20148 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_211
timestamp 1635444444
transform 1 0 20516 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1097_
timestamp 1635444444
transform 1 0 19228 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1938_
timestamp 1635444444
transform 1 0 20608 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_64_228
timestamp 1635444444
transform 1 0 22080 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_236
timestamp 1635444444
transform 1 0 22816 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _0999_
timestamp 1635444444
transform 1 0 23000 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1635444444
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1635444444
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_256
timestamp 1635444444
transform 1 0 24656 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_262
timestamp 1635444444
transform 1 0 25208 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1635444444
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1000_
timestamp 1635444444
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_273
timestamp 1635444444
transform 1 0 26220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0978_
timestamp 1635444444
transform 1 0 25300 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _0994_
timestamp 1635444444
transform 1 0 26588 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 1635444444
transform 1 0 27416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 1635444444
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1635444444
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0993_
timestamp 1635444444
transform 1 0 27784 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1474_
timestamp 1635444444
transform 1 0 28428 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_64_316
timestamp 1635444444
transform 1 0 30176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1635444444
transform -1 0 30820 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1635444444
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _1470_
timestamp 1635444444
transform 1 0 29532 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1635444444
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1635444444
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1635444444
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1635444444
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1635444444
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1635444444
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1635444444
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1635444444
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1635444444
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1635444444
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1635444444
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_106
timestamp 1635444444
transform 1 0 10856 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_93
timestamp 1635444444
transform 1 0 9660 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1077_
timestamp 1635444444
transform 1 0 10028 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_65_113
timestamp 1635444444
transform 1 0 11500 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1635444444
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1946_
timestamp 1635444444
transform 1 0 12236 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_65_137
timestamp 1635444444
transform 1 0 13708 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_145
timestamp 1635444444
transform 1 0 14444 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1111_
timestamp 1635444444
transform 1 0 14720 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_65_157
timestamp 1635444444
transform 1 0 15548 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_164
timestamp 1635444444
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_172
timestamp 1635444444
transform 1 0 16928 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1635444444
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1713_
timestamp 1635444444
transform 1 0 16652 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1723_
timestamp 1635444444
transform 1 0 15916 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_65_178
timestamp 1635444444
transform 1 0 17480 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_182
timestamp 1635444444
transform 1 0 17848 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1675_
timestamp 1635444444
transform 1 0 17572 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1635444444
transform 1 0 18216 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_202
timestamp 1635444444
transform 1 0 19688 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_215
timestamp 1635444444
transform 1 0 20884 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1098_
timestamp 1635444444
transform 1 0 20056 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1635444444
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_225
timestamp 1635444444
transform 1 0 21804 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_229
timestamp 1635444444
transform 1 0 22172 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1635444444
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0996_
timestamp 1635444444
transform 1 0 21896 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1635444444
transform 1 0 22540 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_65_249
timestamp 1635444444
transform 1 0 24012 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_258
timestamp 1635444444
transform 1 0 24840 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0981_
timestamp 1635444444
transform 1 0 25208 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1469_
timestamp 1635444444
transform 1 0 24564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_272
timestamp 1635444444
transform 1 0 26128 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1635444444
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0986_
timestamp 1635444444
transform 1 0 26956 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_284
timestamp 1635444444
transform 1 0 27232 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_288
timestamp 1635444444
transform 1 0 27600 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_292
timestamp 1635444444
transform 1 0 27968 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_299
timestamp 1635444444
transform 1 0 28612 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1635444444
transform 1 0 28336 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1465_
timestamp 1635444444
transform 1 0 27692 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1472_
timestamp 1635444444
transform 1 0 28980 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_65_310
timestamp 1635444444
transform 1 0 29624 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_318
timestamp 1635444444
transform 1 0 30360 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1635444444
transform -1 0 30820 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1635444444
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1635444444
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1635444444
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1635444444
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1635444444
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1635444444
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1635444444
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1635444444
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1635444444
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1635444444
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1635444444
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1635444444
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1635444444
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1635444444
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1635444444
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1635444444
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1635444444
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1635444444
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1635444444
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1635444444
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1635444444
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1635444444
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1635444444
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1635444444
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_97
timestamp 1635444444
transform 1 0 10028 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1635444444
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1635444444
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1635444444
transform 1 0 10120 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_114
timestamp 1635444444
transform 1 0 11592 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_126
timestamp 1635444444
transform 1 0 12696 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1635444444
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_113
timestamp 1635444444
transform 1 0 11500 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1635444444
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1635444444
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0954_
timestamp 1635444444
transform 1 0 12052 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_138
timestamp 1635444444
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_137
timestamp 1635444444
transform 1 0 13708 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_145
timestamp 1635444444
transform 1 0 14444 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1635444444
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1635444444
transform 1 0 14076 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1635444444
transform 1 0 14628 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_66_157
timestamp 1635444444
transform 1 0 15548 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_172
timestamp 1635444444
transform 1 0 16928 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_163
timestamp 1635444444
transform 1 0 16100 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1635444444
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1635444444
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1109_
timestamp 1635444444
transform 1 0 16100 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1635444444
transform 1 0 16652 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_66_179
timestamp 1635444444
transform 1 0 17572 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_192
timestamp 1635444444
transform 1 0 18768 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_185
timestamp 1635444444
transform 1 0 18124 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1635444444
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1102_
timestamp 1635444444
transform 1 0 17940 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1649_
timestamp 1635444444
transform 1 0 17296 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1635444444
transform 1 0 18492 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_66_197
timestamp 1635444444
transform 1 0 19228 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_205
timestamp 1635444444
transform 1 0 19964 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_218
timestamp 1635444444
transform 1 0 21160 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1100_
timestamp 1635444444
transform 1 0 20332 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1635444444
transform 1 0 19780 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1703_
timestamp 1635444444
transform 1 0 21620 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1635444444
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_225
timestamp 1635444444
transform 1 0 21804 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_226
timestamp 1635444444
transform 1 0 21896 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_219
timestamp 1635444444
transform 1 0 21252 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1635444444
transform 1 0 22080 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0997_
timestamp 1635444444
transform 1 0 22632 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_231
timestamp 1635444444
transform 1 0 22356 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1477_
timestamp 1635444444
transform 1 0 23000 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_67_237
timestamp 1635444444
transform 1 0 22908 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_237
timestamp 1635444444
transform 1 0 22908 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1473_
timestamp 1635444444
transform 1 0 23644 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1001_
timestamp 1635444444
transform 1 0 23276 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_248
timestamp 1635444444
transform 1 0 23920 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_241
timestamp 1635444444
transform 1 0 23276 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_244
timestamp 1635444444
transform 1 0 23552 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1251_
timestamp 1635444444
transform 1 0 24288 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1635444444
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_261
timestamp 1635444444
transform 1 0 25116 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_66_253
timestamp 1635444444
transform 1 0 24380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1635444444
transform 1 0 24656 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_66_272
timestamp 1635444444
transform 1 0 26128 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_279
timestamp 1635444444
transform 1 0 26772 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1635444444
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 1635444444
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1635444444
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0983_
timestamp 1635444444
transform 1 0 26496 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0985_
timestamp 1635444444
transform 1 0 25668 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1635444444
transform 1 0 27140 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1961_
timestamp 1635444444
transform 1 0 27140 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_66_299
timestamp 1635444444
transform 1 0 28612 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_299
timestamp 1635444444
transform 1 0 28612 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1476_
timestamp 1635444444
transform 1 0 28980 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1635444444
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_309
timestamp 1635444444
transform 1 0 29532 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_316
timestamp 1635444444
transform 1 0 30176 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_310
timestamp 1635444444
transform 1 0 29624 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_318
timestamp 1635444444
transform 1 0 30360 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1635444444
transform -1 0 30820 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1635444444
transform -1 0 30820 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1635444444
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1635444444
transform 1 0 29808 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_18
timestamp 1635444444
transform 1 0 2760 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_6
timestamp 1635444444
transform 1 0 1656 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1635444444
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1635444444
transform 1 0 1380 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_26
timestamp 1635444444
transform 1 0 3496 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1635444444
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1635444444
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1635444444
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1635444444
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1635444444
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1635444444
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1635444444
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1635444444
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1635444444
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1635444444
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1635444444
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1635444444
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1635444444
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1635444444
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1635444444
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1635444444
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_162
timestamp 1635444444
transform 1 0 16008 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_174
timestamp 1635444444
transform 1 0 17112 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1110_
timestamp 1635444444
transform 1 0 15180 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1635444444
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1635444444
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1635444444
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1104_
timestamp 1635444444
transform 1 0 17664 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_68_197
timestamp 1635444444
transform 1 0 19228 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_204
timestamp 1635444444
transform 1 0 19872 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1937_
timestamp 1635444444
transform 1 0 20240 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1635444444
transform 1 0 19596 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_224
timestamp 1635444444
transform 1 0 21712 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_231
timestamp 1635444444
transform 1 0 22356 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_238
timestamp 1635444444
transform 1 0 23000 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0995_
timestamp 1635444444
transform 1 0 22724 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1635444444
transform 1 0 22080 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_244
timestamp 1635444444
transform 1 0 23552 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1635444444
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_262
timestamp 1635444444
transform 1 0 25208 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1635444444
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1635444444
transform 1 0 23644 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1247_
timestamp 1635444444
transform 1 0 24380 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_68_268
timestamp 1635444444
transform 1 0 25760 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_278
timestamp 1635444444
transform 1 0 26680 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0982_
timestamp 1635444444
transform 1 0 25852 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _0988_
timestamp 1635444444
transform 1 0 27048 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_68_291
timestamp 1635444444
transform 1 0 27876 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_299
timestamp 1635444444
transform 1 0 28612 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_304
timestamp 1635444444
transform 1 0 29072 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1635444444
transform 1 0 28704 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_316
timestamp 1635444444
transform 1 0 30176 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1635444444
transform -1 0 30820 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1635444444
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _1479_
timestamp 1635444444
transform 1 0 29532 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1635444444
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1635444444
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1635444444
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1635444444
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1635444444
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1635444444
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1635444444
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1635444444
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1635444444
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1635444444
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1635444444
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1635444444
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1635444444
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1635444444
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_113
timestamp 1635444444
transform 1 0 11500 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1635444444
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1635444444
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0949_
timestamp 1635444444
transform 1 0 12052 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_69_137
timestamp 1635444444
transform 1 0 13708 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_145
timestamp 1635444444
transform 1 0 14444 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_1  _1509_
timestamp 1635444444
transform 1 0 14628 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_153
timestamp 1635444444
transform 1 0 15180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_165
timestamp 1635444444
transform 1 0 16284 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1635444444
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1508_
timestamp 1635444444
transform 1 0 16652 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_175
timestamp 1635444444
transform 1 0 17204 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_187
timestamp 1635444444
transform 1 0 18308 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_208
timestamp 1635444444
transform 1 0 20240 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_216
timestamp 1635444444
transform 1 0 20976 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1101_
timestamp 1635444444
transform 1 0 19412 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1635444444
transform 1 0 21068 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1635444444
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_225
timestamp 1635444444
transform 1 0 21804 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_229
timestamp 1635444444
transform 1 0 22172 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_236
timestamp 1635444444
transform 1 0 22816 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1635444444
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1231_
timestamp 1635444444
transform 1 0 23184 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1489_
timestamp 1635444444
transform 1 0 22540 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1635444444
transform 1 0 21896 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_243
timestamp 1635444444
transform 1 0 23460 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_256
timestamp 1635444444
transform 1 0 24656 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1244_
timestamp 1635444444
transform 1 0 23828 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1245_
timestamp 1635444444
transform 1 0 25024 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_263
timestamp 1635444444
transform 1 0 25300 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_270
timestamp 1635444444
transform 1 0 25944 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_278
timestamp 1635444444
transform 1 0 26680 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1635444444
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1635444444
transform 1 0 25668 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0984_
timestamp 1635444444
transform 1 0 26956 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_284
timestamp 1635444444
transform 1 0 27232 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_292
timestamp 1635444444
transform 1 0 27968 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_297
timestamp 1635444444
transform 1 0 28428 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_304
timestamp 1635444444
transform 1 0 29072 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1466_
timestamp 1635444444
transform 1 0 28796 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1468_
timestamp 1635444444
transform 1 0 28152 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_316
timestamp 1635444444
transform 1 0 30176 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1635444444
transform -1 0 30820 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1635444444
transform 1 0 29808 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1635444444
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1635444444
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1635444444
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1635444444
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1635444444
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1635444444
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1635444444
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1635444444
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1635444444
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1635444444
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1635444444
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1635444444
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1635444444
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1635444444
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1635444444
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1635444444
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1635444444
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1635444444
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_141
timestamp 1635444444
transform 1 0 14076 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1635444444
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1748_
timestamp 1635444444
transform 1 0 14628 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_70_156
timestamp 1635444444
transform 1 0 15456 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_173
timestamp 1635444444
transform 1 0 17020 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1746_
timestamp 1635444444
transform 1 0 16192 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_70_185
timestamp 1635444444
transform 1 0 18124 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_192
timestamp 1635444444
transform 1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1635444444
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1521_
timestamp 1635444444
transform 1 0 18216 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 19412 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_197
timestamp 1635444444
transform 1 0 19228 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_204
timestamp 1635444444
transform 1 0 19872 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_211
timestamp 1635444444
transform 1 0 20516 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_215
timestamp 1635444444
transform 1 0 20884 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1635444444
transform 1 0 20240 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1635444444
transform 1 0 20976 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1635444444
transform 1 0 19596 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_219
timestamp 1635444444
transform 1 0 21252 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_223
timestamp 1635444444
transform 1 0 21620 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_227
timestamp 1635444444
transform 1 0 21988 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_235
timestamp 1635444444
transform 1 0 22724 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_240
timestamp 1635444444
transform 1 0 23184 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1635444444
transform 1 0 21712 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1246_
timestamp 1635444444
transform 1 0 22908 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_247
timestamp 1635444444
transform 1 0 23828 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1635444444
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1635444444
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1243_
timestamp 1635444444
transform 1 0 23552 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1635444444
transform 1 0 24380 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_70_269
timestamp 1635444444
transform 1 0 25852 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_276
timestamp 1635444444
transform 1 0 26496 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_283
timestamp 1635444444
transform 1 0 27140 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0970_
timestamp 1635444444
transform 1 0 26220 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0987_
timestamp 1635444444
transform 1 0 26864 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_289
timestamp 1635444444
transform 1 0 27692 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_293
timestamp 1635444444
transform 1 0 28060 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_304
timestamp 1635444444
transform 1 0 29072 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1471_
timestamp 1635444444
transform 1 0 27784 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1484_
timestamp 1635444444
transform 1 0 28428 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_70_309
timestamp 1635444444
transform 1 0 29532 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_316
timestamp 1635444444
transform 1 0 30176 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1635444444
transform -1 0 30820 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1635444444
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1635444444
transform 1 0 29808 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_18
timestamp 1635444444
transform 1 0 2760 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_6
timestamp 1635444444
transform 1 0 1656 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1635444444
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1635444444
transform 1 0 1380 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_30
timestamp 1635444444
transform 1 0 3864 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_42
timestamp 1635444444
transform 1 0 4968 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_54
timestamp 1635444444
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1635444444
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1635444444
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1635444444
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1635444444
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1635444444
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1635444444
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1635444444
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1635444444
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1635444444
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1635444444
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_137
timestamp 1635444444
transform 1 0 13708 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_143
timestamp 1635444444
transform 1 0 14260 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1747_
timestamp 1635444444
transform 1 0 14352 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_71_153
timestamp 1635444444
transform 1 0 15180 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_163
timestamp 1635444444
transform 1 0 16100 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1635444444
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1635444444
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1254_
timestamp 1635444444
transform 1 0 15548 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1504_
timestamp 1635444444
transform 1 0 16652 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_175
timestamp 1635444444
transform 1 0 17204 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_179
timestamp 1635444444
transform 1 0 17572 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_189
timestamp 1635444444
transform 1 0 18492 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1756_
timestamp 1635444444
transform 1 0 17664 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1757_
timestamp 1635444444
transform 1 0 18860 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_71_202
timestamp 1635444444
transform 1 0 19688 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_208
timestamp 1635444444
transform 1 0 20240 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__or4b_4  _1265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 20332 0 -1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_71_220
timestamp 1635444444
transform 1 0 21344 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_225
timestamp 1635444444
transform 1 0 21804 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_233
timestamp 1635444444
transform 1 0 22540 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1635444444
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1082_
timestamp 1635444444
transform 1 0 22172 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_241
timestamp 1635444444
transform 1 0 23276 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_259
timestamp 1635444444
transform 1 0 24932 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1635444444
transform 1 0 23460 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_71_274
timestamp 1635444444
transform 1 0 26312 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1635444444
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1241_
timestamp 1635444444
transform 1 0 25484 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1962_
timestamp 1635444444
transform 1 0 26956 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_297
timestamp 1635444444
transform 1 0 28428 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1482_
timestamp 1635444444
transform 1 0 28796 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_71_308
timestamp 1635444444
transform 1 0 29440 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_316
timestamp 1635444444
transform 1 0 30176 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1635444444
transform -1 0 30820 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1635444444
transform 1 0 29808 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1635444444
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1635444444
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1635444444
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1635444444
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1635444444
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1635444444
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1635444444
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1635444444
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1635444444
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1635444444
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1635444444
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1635444444
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1635444444
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1635444444
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1635444444
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1635444444
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1635444444
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1635444444
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1635444444
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1635444444
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1635444444
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1635444444
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1635444444
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1635444444
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1635444444
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1635444444
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1635444444
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1635444444
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1635444444
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1635444444
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1635444444
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1635444444
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1635444444
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1635444444
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1635444444
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_141
timestamp 1635444444
transform 1 0 14076 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_152
timestamp 1635444444
transform 1 0 15088 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1635444444
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1635444444
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1510_
timestamp 1635444444
transform 1 0 14812 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1749_
timestamp 1635444444
transform 1 0 14260 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1743_
timestamp 1635444444
transform 1 0 16008 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1502_
timestamp 1635444444
transform 1 0 15824 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_159
timestamp 1635444444
transform 1 0 15732 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_155
timestamp 1635444444
transform 1 0 15364 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_160
timestamp 1635444444
transform 1 0 15824 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1501_
timestamp 1635444444
transform 1 0 16928 0 -1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1635444444
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_169
timestamp 1635444444
transform 1 0 16652 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_164
timestamp 1635444444
transform 1 0 16192 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_171
timestamp 1635444444
transform 1 0 16836 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_185
timestamp 1635444444
transform 1 0 18124 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_182
timestamp 1635444444
transform 1 0 17848 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_192
timestamp 1635444444
transform 1 0 18768 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1635444444
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1356_
timestamp 1635444444
transform 1 0 18676 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1503_
timestamp 1635444444
transform 1 0 17204 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1519_
timestamp 1635444444
transform 1 0 18216 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1733_
timestamp 1635444444
transform 1 0 19136 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1635444444
transform -1 0 19872 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_200
timestamp 1635444444
transform 1 0 19504 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_204
timestamp 1635444444
transform 1 0 19872 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_205
timestamp 1635444444
transform 1 0 19964 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_213
timestamp 1635444444
transform 1 0 20700 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1087_
timestamp 1635444444
transform 1 0 20332 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1359_
timestamp 1635444444
transform 1 0 21068 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1635444444
transform 1 0 20056 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1635444444
transform 1 0 19228 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1378_
timestamp 1635444444
transform 1 0 21804 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1360_
timestamp 1635444444
transform 1 0 21896 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1635444444
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_220
timestamp 1635444444
transform 1 0 21344 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_222
timestamp 1635444444
transform 1 0 21528 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1483_
timestamp 1635444444
transform 1 0 22816 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_228
timestamp 1635444444
transform 1 0 22080 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_230
timestamp 1635444444
transform 1 0 22264 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1242_
timestamp 1635444444
transform 1 0 23000 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_239
timestamp 1635444444
transform 1 0 23092 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_241
timestamp 1635444444
transform 1 0 23276 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_248
timestamp 1635444444
transform 1 0 23920 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_253
timestamp 1635444444
transform 1 0 24380 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_250
timestamp 1635444444
transform 1 0 24104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1635444444
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1225_
timestamp 1635444444
transform 1 0 24656 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1226_
timestamp 1635444444
transform 1 0 24472 0 -1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _1238_
timestamp 1635444444
transform 1 0 23644 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1481_
timestamp 1635444444
transform 1 0 23828 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_266
timestamp 1635444444
transform 1 0 25576 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_264
timestamp 1635444444
transform 1 0 25392 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_271
timestamp 1635444444
transform 1 0 26036 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1635444444
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_281
timestamp 1635444444
transform 1 0 26956 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1635444444
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1235_
timestamp 1635444444
transform 1 0 25760 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1635444444
transform 1 0 25944 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_72_286
timestamp 1635444444
transform 1 0 27416 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_293
timestamp 1635444444
transform 1 0 28060 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_304
timestamp 1635444444
transform 1 0 29072 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_294
timestamp 1635444444
transform 1 0 28152 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_305
timestamp 1635444444
transform 1 0 29164 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1475_
timestamp 1635444444
transform 1 0 27784 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1486_
timestamp 1635444444
transform 1 0 28428 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1488_
timestamp 1635444444
transform 1 0 28520 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1491_
timestamp 1635444444
transform 1 0 27508 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_72_309
timestamp 1635444444
transform 1 0 29532 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_316
timestamp 1635444444
transform 1 0 30176 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_311
timestamp 1635444444
transform 1 0 29716 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_316
timestamp 1635444444
transform 1 0 30176 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1635444444
transform -1 0 30820 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1635444444
transform -1 0 30820 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1635444444
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1635444444
transform 1 0 29808 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1635444444
transform 1 0 29808 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1635444444
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1635444444
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1635444444
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1635444444
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1635444444
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1635444444
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1635444444
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1635444444
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1635444444
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1635444444
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1635444444
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1635444444
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1635444444
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_105
timestamp 1635444444
transform 1 0 10764 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_97
timestamp 1635444444
transform 1 0 10028 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _0942_
timestamp 1635444444
transform 1 0 10856 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_112
timestamp 1635444444
transform 1 0 11408 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_124
timestamp 1635444444
transform 1 0 12512 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_136
timestamp 1635444444
transform 1 0 13616 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_141
timestamp 1635444444
transform 1 0 14076 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_145
timestamp 1635444444
transform 1 0 14444 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_152
timestamp 1635444444
transform 1 0 15088 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1635444444
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1511_
timestamp 1635444444
transform 1 0 14536 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_162
timestamp 1635444444
transform 1 0 16008 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_172
timestamp 1635444444
transform 1 0 16928 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1515_
timestamp 1635444444
transform 1 0 15456 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1517_
timestamp 1635444444
transform 1 0 16376 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_185
timestamp 1635444444
transform 1 0 18124 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_192
timestamp 1635444444
transform 1 0 18768 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1635444444
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1755_
timestamp 1635444444
transform 1 0 17296 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1635444444
transform 1 0 18492 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_197
timestamp 1635444444
transform 1 0 19228 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_204
timestamp 1635444444
transform 1 0 19872 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_210
timestamp 1635444444
transform 1 0 20424 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _1377_
timestamp 1635444444
transform 1 0 19412 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1635444444
transform 1 0 20516 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_74_227
timestamp 1635444444
transform 1 0 21988 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_238
timestamp 1635444444
transform 1 0 23000 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1228_
timestamp 1635444444
transform 1 0 22724 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1635444444
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1635444444
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_253
timestamp 1635444444
transform 1 0 24380 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_257
timestamp 1635444444
transform 1 0 24748 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_261
timestamp 1635444444
transform 1 0 25116 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1635444444
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1233_
timestamp 1635444444
transform 1 0 24840 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1485_
timestamp 1635444444
transform 1 0 23368 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_274
timestamp 1635444444
transform 1 0 26312 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_281
timestamp 1635444444
transform 1 0 26956 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1236_
timestamp 1635444444
transform 1 0 26680 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1237_
timestamp 1635444444
transform 1 0 25484 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_74_288
timestamp 1635444444
transform 1 0 27600 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_295
timestamp 1635444444
transform 1 0 28244 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_302
timestamp 1635444444
transform 1 0 28888 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1239_
timestamp 1635444444
transform 1 0 27324 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1478_
timestamp 1635444444
transform 1 0 28612 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1480_
timestamp 1635444444
transform 1 0 27968 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_74_309
timestamp 1635444444
transform 1 0 29532 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_316
timestamp 1635444444
transform 1 0 30176 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1635444444
transform -1 0 30820 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1635444444
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1635444444
transform 1 0 29808 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_18
timestamp 1635444444
transform 1 0 2760 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_6
timestamp 1635444444
transform 1 0 1656 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1635444444
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1635444444
transform 1 0 1380 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_30
timestamp 1635444444
transform 1 0 3864 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_42
timestamp 1635444444
transform 1 0 4968 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_54
timestamp 1635444444
transform 1 0 6072 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1635444444
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1635444444
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1635444444
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1635444444
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1635444444
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1635444444
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1635444444
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1635444444
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_125
timestamp 1635444444
transform 1 0 12604 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1635444444
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_136
timestamp 1635444444
transform 1 0 13616 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_145
timestamp 1635444444
transform 1 0 14444 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1752_
timestamp 1635444444
transform 1 0 14812 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1635444444
transform 1 0 14168 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1635444444
transform 1 0 13340 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_158
timestamp 1635444444
transform 1 0 15640 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_166
timestamp 1635444444
transform 1 0 16376 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_169
timestamp 1635444444
transform 1 0 16652 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_173
timestamp 1635444444
transform 1 0 17020 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1635444444
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1635444444
transform 1 0 16744 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_187
timestamp 1635444444
transform 1 0 18308 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1513_
timestamp 1635444444
transform 1 0 17388 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1520_
timestamp 1635444444
transform 1 0 18676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_197
timestamp 1635444444
transform 1 0 19228 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_204
timestamp 1635444444
transform 1 0 19872 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_213
timestamp 1635444444
transform 1 0 20700 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1257_
timestamp 1635444444
transform 1 0 20240 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1376_
timestamp 1635444444
transform 1 0 19596 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1490_
timestamp 1635444444
transform 1 0 21068 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_220
timestamp 1635444444
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_225
timestamp 1635444444
transform 1 0 21804 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_231
timestamp 1635444444
transform 1 0 22356 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_238
timestamp 1635444444
transform 1 0 23000 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1635444444
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1219_
timestamp 1635444444
transform 1 0 22724 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1487_
timestamp 1635444444
transform 1 0 22080 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_258
timestamp 1635444444
transform 1 0 24840 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1635444444
transform 1 0 23368 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_75_264
timestamp 1635444444
transform 1 0 25392 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_274
timestamp 1635444444
transform 1 0 26312 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1635444444
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1232_
timestamp 1635444444
transform 1 0 26956 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1234_
timestamp 1635444444
transform 1 0 25484 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_75_284
timestamp 1635444444
transform 1 0 27232 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_290
timestamp 1635444444
transform 1 0 27784 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_298
timestamp 1635444444
transform 1 0 28520 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1499_
timestamp 1635444444
transform 1 0 27876 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1635444444
transform 1 0 29072 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_308
timestamp 1635444444
transform 1 0 29440 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_316
timestamp 1635444444
transform 1 0 30176 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1635444444
transform -1 0 30820 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1635444444
transform 1 0 29808 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_18
timestamp 1635444444
transform 1 0 2760 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_6
timestamp 1635444444
transform 1 0 1656 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1635444444
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1635444444
transform 1 0 1380 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_26
timestamp 1635444444
transform 1 0 3496 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1635444444
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1635444444
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1635444444
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1635444444
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1635444444
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1635444444
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1635444444
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1635444444
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1635444444
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_105
timestamp 1635444444
transform 1 0 10764 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_97
timestamp 1635444444
transform 1 0 10028 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _0934_
timestamp 1635444444
transform 1 0 10856 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_112
timestamp 1635444444
transform 1 0 11408 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_122
timestamp 1635444444
transform 1 0 12328 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_130
timestamp 1635444444
transform 1 0 13064 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__and2_2  _0938_
timestamp 1635444444
transform 1 0 11776 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_135
timestamp 1635444444
transform 1 0 13524 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1635444444
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_141
timestamp 1635444444
transform 1 0 14076 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1635444444
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1751_
timestamp 1635444444
transform 1 0 14628 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1635444444
transform 1 0 13248 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_156
timestamp 1635444444
transform 1 0 15456 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_169
timestamp 1635444444
transform 1 0 16652 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_173
timestamp 1635444444
transform 1 0 17020 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1512_
timestamp 1635444444
transform 1 0 17112 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1753_
timestamp 1635444444
transform 1 0 15824 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_76_184
timestamp 1635444444
transform 1 0 18032 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_192
timestamp 1635444444
transform 1 0 18768 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1635444444
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1017_
timestamp 1635444444
transform 1 0 18400 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_202
timestamp 1635444444
transform 1 0 19688 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_206
timestamp 1635444444
transform 1 0 20056 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_213
timestamp 1635444444
transform 1 0 20700 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1009_
timestamp 1635444444
transform 1 0 20148 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1013_
timestamp 1635444444
transform 1 0 21068 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1016_
timestamp 1635444444
transform 1 0 19228 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_76_222
timestamp 1635444444
transform 1 0 21528 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_230
timestamp 1635444444
transform 1 0 22264 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_235
timestamp 1635444444
transform 1 0 22724 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1220_
timestamp 1635444444
transform 1 0 22448 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1230_
timestamp 1635444444
transform 1 0 23092 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_76_248
timestamp 1635444444
transform 1 0 23920 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_262
timestamp 1635444444
transform 1 0 25208 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1635444444
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1227_
timestamp 1635444444
transform 1 0 24380 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1635444444
transform 1 0 25944 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_76_286
timestamp 1635444444
transform 1 0 27416 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_290
timestamp 1635444444
transform 1 0 27784 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_298
timestamp 1635444444
transform 1 0 28520 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1493_
timestamp 1635444444
transform 1 0 27876 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 1635444444
transform 1 0 29256 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_309
timestamp 1635444444
transform 1 0 29532 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_316
timestamp 1635444444
transform 1 0 30176 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1635444444
transform -1 0 30820 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1635444444
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1635444444
transform 1 0 29808 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_17
timestamp 1635444444
transform 1 0 2668 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_6
timestamp 1635444444
transform 1 0 1656 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1635444444
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0881_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2024 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1635444444
transform 1 0 1380 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_29
timestamp 1635444444
transform 1 0 3772 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_41
timestamp 1635444444
transform 1 0 4876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1635444444
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1635444444
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1635444444
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1635444444
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1635444444
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1635444444
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1635444444
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1635444444
transform -1 0 13248 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1635444444
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1635444444
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_125
timestamp 1635444444
transform 1 0 12604 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_129
timestamp 1635444444
transform 1 0 12972 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1635444444
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_135
timestamp 1635444444
transform 1 0 13524 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_142
timestamp 1635444444
transform 1 0 14168 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1750_
timestamp 1635444444
transform 1 0 14536 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1635444444
transform 1 0 13892 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1635444444
transform 1 0 13248 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_77_155
timestamp 1635444444
transform 1 0 15364 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_164
timestamp 1635444444
transform 1 0 16192 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1635444444
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1635444444
transform 1 0 15916 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1754_
timestamp 1635444444
transform 1 0 16652 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_77_178
timestamp 1635444444
transform 1 0 17480 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_187
timestamp 1635444444
transform 1 0 18308 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1261_
timestamp 1635444444
transform 1 0 17848 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _1372_
timestamp 1635444444
transform 1 0 18676 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_77_204
timestamp 1635444444
transform 1 0 19872 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_216
timestamp 1635444444
transform 1 0 20976 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1256_
timestamp 1635444444
transform 1 0 20240 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_77_230
timestamp 1635444444
transform 1 0 22264 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_236
timestamp 1635444444
transform 1 0 22816 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_240
timestamp 1635444444
transform 1 0 23184 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1635444444
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1014_
timestamp 1635444444
transform 1 0 21804 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _1229_
timestamp 1635444444
transform 1 0 22908 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_260
timestamp 1635444444
transform 1 0 25024 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1635444444
transform 1 0 23552 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_77_274
timestamp 1635444444
transform 1 0 26312 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_281
timestamp 1635444444
transform 1 0 26956 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1635444444
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1635444444
transform 1 0 25392 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1635444444
transform 1 0 27140 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_287
timestamp 1635444444
transform 1 0 27508 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_298
timestamp 1635444444
transform 1 0 28520 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1495_
timestamp 1635444444
transform 1 0 27876 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_77_306
timestamp 1635444444
transform 1 0 29256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_316
timestamp 1635444444
transform 1 0 30176 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1635444444
transform -1 0 30820 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1010_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 29348 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_78_18
timestamp 1635444444
transform 1 0 2760 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_78_3
timestamp 1635444444
transform 1 0 1380 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1635444444
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1932 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_78_26
timestamp 1635444444
transform 1 0 3496 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1635444444
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_41
timestamp 1635444444
transform 1 0 4876 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1635444444
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 1635444444
transform 1 0 4968 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_46
timestamp 1635444444
transform 1 0 5336 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_58
timestamp 1635444444
transform 1 0 6440 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_66
timestamp 1635444444
transform 1 0 7176 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_70
timestamp 1635444444
transform 1 0 7544 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_82
timestamp 1635444444
transform 1 0 8648 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1635444444
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1635444444
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1635444444
transform 1 0 7268 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_104
timestamp 1635444444
transform 1 0 10672 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_97
timestamp 1635444444
transform 1 0 10028 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1635444444
transform 1 0 10304 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_116
timestamp 1635444444
transform 1 0 11776 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_120
timestamp 1635444444
transform 1 0 12144 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_124
timestamp 1635444444
transform 1 0 12512 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_128
timestamp 1635444444
transform 1 0 12880 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1635444444
transform 1 0 11868 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1635444444
transform 1 0 12604 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_78_132
timestamp 1635444444
transform 1 0 13248 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_136
timestamp 1635444444
transform 1 0 13616 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_141
timestamp 1635444444
transform 1 0 14076 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_145
timestamp 1635444444
transform 1 0 14444 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_152
timestamp 1635444444
transform 1 0 15088 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1635444444
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1514_
timestamp 1635444444
transform 1 0 14536 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1635444444
transform 1 0 13340 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_78_162
timestamp 1635444444
transform 1 0 16008 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_174
timestamp 1635444444
transform 1 0 17112 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1258_
timestamp 1635444444
transform 1 0 15456 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1260_
timestamp 1635444444
transform 1 0 16560 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_178
timestamp 1635444444
transform 1 0 17480 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_185
timestamp 1635444444
transform 1 0 18124 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_192
timestamp 1635444444
transform 1 0 18768 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1635444444
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1635444444
transform 1 0 18492 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1259_
timestamp 1635444444
transform 1 0 17572 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_197
timestamp 1635444444
transform 1 0 19228 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_201
timestamp 1635444444
transform 1 0 19596 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_208
timestamp 1635444444
transform 1 0 20240 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1008_
timestamp 1635444444
transform 1 0 20608 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1015_
timestamp 1635444444
transform 1 0 19688 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_220
timestamp 1635444444
transform 1 0 21344 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_227
timestamp 1635444444
transform 1 0 21988 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1635444444
transform 1 0 21712 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1635444444
transform 1 0 22540 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_78_243
timestamp 1635444444
transform 1 0 23460 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1635444444
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1635444444
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1635444444
transform 1 0 24380 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_78_263
timestamp 1635444444
transform 1 0 25300 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1635444444
transform 1 0 25852 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_78_285
timestamp 1635444444
transform 1 0 27324 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_78_298
timestamp 1635444444
transform 1 0 28520 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1497_
timestamp 1635444444
transform 1 0 27876 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_78_306
timestamp 1635444444
transform 1 0 29256 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_78_309
timestamp 1635444444
transform 1 0 29532 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_316
timestamp 1635444444
transform 1 0 30176 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1635444444
transform -1 0 30820 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1635444444
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1635444444
transform 1 0 29808 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_6
timestamp 1635444444
transform 1 0 1656 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1635444444
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1635444444
transform 1 0 1380 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1635444444
transform 1 0 2392 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_79_24
timestamp 1635444444
transform 1 0 3312 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_39
timestamp 1635444444
transform 1 0 4692 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1635444444
transform 1 0 3680 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1635444444
transform 1 0 3772 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 5060 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_49
timestamp 1635444444
transform 1 0 5612 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1635444444
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_60
timestamp 1635444444
transform 1 0 6624 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1635444444
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1635444444
transform 1 0 6348 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1635444444
transform 1 0 6992 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_67
timestamp 1635444444
transform 1 0 7268 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_79_78
timestamp 1635444444
transform 1 0 8280 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1635444444
transform 1 0 8832 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635444444
transform 1 0 8004 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1635444444
transform 1 0 8924 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_79_103
timestamp 1635444444
transform 1 0 10580 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_95
timestamp 1635444444
transform 1 0 9844 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1635444444
transform 1 0 10212 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1635444444
transform 1 0 12512 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1635444444
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_117
timestamp 1635444444
transform 1 0 11868 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_123
timestamp 1635444444
transform 1 0 12420 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_129
timestamp 1635444444
transform 1 0 12972 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1635444444
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1635444444
transform 1 0 12696 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1635444444
transform 1 0 11500 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_136
timestamp 1635444444
transform 1 0 13616 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_141
timestamp 1635444444
transform 1 0 14076 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_148
timestamp 1635444444
transform 1 0 14720 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1635444444
transform 1 0 13984 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1516_
timestamp 1635444444
transform 1 0 15088 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1635444444
transform 1 0 14444 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1635444444
transform 1 0 13340 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_158
timestamp 1635444444
transform 1 0 15640 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_166
timestamp 1635444444
transform 1 0 16376 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_169
timestamp 1635444444
transform 1 0 16652 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1635444444
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1518_
timestamp 1635444444
transform 1 0 16744 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_176
timestamp 1635444444
transform 1 0 17296 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_180
timestamp 1635444444
transform 1 0 17664 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_184
timestamp 1635444444
transform 1 0 18032 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_192
timestamp 1635444444
transform 1 0 18768 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1635444444
transform 1 0 19136 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1635444444
transform 1 0 17756 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1086_
timestamp 1635444444
transform 1 0 18400 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_202
timestamp 1635444444
transform 1 0 19688 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_213
timestamp 1635444444
transform 1 0 20700 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1264_
timestamp 1635444444
transform 1 0 19228 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1635444444
transform 1 0 21068 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 1635444444
transform 1 0 20424 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_220
timestamp 1635444444
transform 1 0 21344 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_235
timestamp 1635444444
transform 1 0 22724 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1635444444
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1635444444
transform 1 0 21804 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_79_243
timestamp 1635444444
transform 1 0 23460 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_248
timestamp 1635444444
transform 1 0 23920 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1635444444
transform 1 0 24288 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1494_
timestamp 1635444444
transform 1 0 23644 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1635444444
transform 1 0 24380 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_79_263
timestamp 1635444444
transform 1 0 25300 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_271
timestamp 1635444444
transform 1 0 26036 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_276
timestamp 1635444444
transform 1 0 26496 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_281
timestamp 1635444444
transform 1 0 26956 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1635444444
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1635444444
transform 1 0 26128 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_285
timestamp 1635444444
transform 1 0 27324 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_292
timestamp 1635444444
transform 1 0 27968 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_301
timestamp 1635444444
transform 1 0 28796 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 1635444444
transform 1 0 27416 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1635444444
transform 1 0 28336 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_79_307
timestamp 1635444444
transform 1 0 29348 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_309
timestamp 1635444444
transform 1 0 29532 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_316
timestamp 1635444444
transform 1 0 30176 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1635444444
transform -1 0 30820 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1635444444
transform 1 0 29440 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1635444444
transform 1 0 29808 0 -1 45696
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 4904 800 5024 6 hb_clk_o
port 0 nsew signal tristate
rlabel metal3 s 0 6944 800 7064 6 hb_clkn_o
port 1 nsew signal tristate
rlabel metal3 s 0 2864 800 2984 6 hb_csn_o
port 2 nsew signal tristate
rlabel metal3 s 0 32920 800 33040 6 hb_dq_i[0]
port 3 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 hb_dq_i[1]
port 4 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 hb_dq_i[2]
port 5 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 hb_dq_i[3]
port 6 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 hb_dq_i[4]
port 7 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 hb_dq_i[5]
port 8 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 hb_dq_i[6]
port 9 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 hb_dq_i[7]
port 10 nsew signal input
rlabel metal3 s 0 14832 800 14952 6 hb_dq_o[0]
port 11 nsew signal tristate
rlabel metal3 s 0 16872 800 16992 6 hb_dq_o[1]
port 12 nsew signal tristate
rlabel metal3 s 0 18912 800 19032 6 hb_dq_o[2]
port 13 nsew signal tristate
rlabel metal3 s 0 20952 800 21072 6 hb_dq_o[3]
port 14 nsew signal tristate
rlabel metal3 s 0 22856 800 22976 6 hb_dq_o[4]
port 15 nsew signal tristate
rlabel metal3 s 0 24896 800 25016 6 hb_dq_o[5]
port 16 nsew signal tristate
rlabel metal3 s 0 26936 800 27056 6 hb_dq_o[6]
port 17 nsew signal tristate
rlabel metal3 s 0 28840 800 28960 6 hb_dq_o[7]
port 18 nsew signal tristate
rlabel metal3 s 0 12928 800 13048 6 hb_dq_oen
port 19 nsew signal tristate
rlabel metal3 s 0 960 800 1080 6 hb_rstn_o
port 20 nsew signal tristate
rlabel metal3 s 0 30880 800 31000 6 hb_rwds_i
port 21 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 hb_rwds_o
port 22 nsew signal tristate
rlabel metal3 s 0 10888 800 11008 6 hb_rwds_oen
port 23 nsew signal tristate
rlabel metal2 s 386 47200 442 48000 6 rst_i
port 24 nsew signal input
rlabel metal4 s 5909 2128 6229 45744 6 vccd1
port 25 nsew power input
rlabel metal4 s 15839 2128 16159 45744 6 vccd1
port 25 nsew power input
rlabel metal4 s 25770 2128 26090 45744 6 vccd1
port 25 nsew power input
rlabel metal4 s 10874 2128 11194 45744 6 vssd1
port 26 nsew ground input
rlabel metal4 s 20805 2128 21125 45744 6 vssd1
port 26 nsew ground input
rlabel metal2 s 1122 47200 1178 48000 6 wb_clk_i
port 27 nsew signal input
rlabel metal2 s 1858 47200 1914 48000 6 wb_rst_i
port 28 nsew signal input
rlabel metal3 s 31200 47472 32000 47592 6 wbs_ack_o
port 29 nsew signal tristate
rlabel metal2 s 7930 47200 7986 48000 6 wbs_adr_i[0]
port 30 nsew signal input
rlabel metal2 s 15566 47200 15622 48000 6 wbs_adr_i[10]
port 31 nsew signal input
rlabel metal2 s 16394 47200 16450 48000 6 wbs_adr_i[11]
port 32 nsew signal input
rlabel metal2 s 17130 47200 17186 48000 6 wbs_adr_i[12]
port 33 nsew signal input
rlabel metal2 s 17866 47200 17922 48000 6 wbs_adr_i[13]
port 34 nsew signal input
rlabel metal2 s 18602 47200 18658 48000 6 wbs_adr_i[14]
port 35 nsew signal input
rlabel metal2 s 19430 47200 19486 48000 6 wbs_adr_i[15]
port 36 nsew signal input
rlabel metal2 s 20166 47200 20222 48000 6 wbs_adr_i[16]
port 37 nsew signal input
rlabel metal2 s 20902 47200 20958 48000 6 wbs_adr_i[17]
port 38 nsew signal input
rlabel metal2 s 21730 47200 21786 48000 6 wbs_adr_i[18]
port 39 nsew signal input
rlabel metal2 s 22466 47200 22522 48000 6 wbs_adr_i[19]
port 40 nsew signal input
rlabel metal2 s 8758 47200 8814 48000 6 wbs_adr_i[1]
port 41 nsew signal input
rlabel metal2 s 23202 47200 23258 48000 6 wbs_adr_i[20]
port 42 nsew signal input
rlabel metal2 s 23938 47200 23994 48000 6 wbs_adr_i[21]
port 43 nsew signal input
rlabel metal2 s 24766 47200 24822 48000 6 wbs_adr_i[22]
port 44 nsew signal input
rlabel metal2 s 25502 47200 25558 48000 6 wbs_adr_i[23]
port 45 nsew signal input
rlabel metal2 s 26238 47200 26294 48000 6 wbs_adr_i[24]
port 46 nsew signal input
rlabel metal2 s 27066 47200 27122 48000 6 wbs_adr_i[25]
port 47 nsew signal input
rlabel metal2 s 27802 47200 27858 48000 6 wbs_adr_i[26]
port 48 nsew signal input
rlabel metal2 s 28538 47200 28594 48000 6 wbs_adr_i[27]
port 49 nsew signal input
rlabel metal2 s 29274 47200 29330 48000 6 wbs_adr_i[28]
port 50 nsew signal input
rlabel metal2 s 30102 47200 30158 48000 6 wbs_adr_i[29]
port 51 nsew signal input
rlabel metal2 s 9494 47200 9550 48000 6 wbs_adr_i[2]
port 52 nsew signal input
rlabel metal2 s 30838 47200 30894 48000 6 wbs_adr_i[30]
port 53 nsew signal input
rlabel metal2 s 31574 47200 31630 48000 6 wbs_adr_i[31]
port 54 nsew signal input
rlabel metal2 s 10230 47200 10286 48000 6 wbs_adr_i[3]
port 55 nsew signal input
rlabel metal2 s 11058 47200 11114 48000 6 wbs_adr_i[4]
port 56 nsew signal input
rlabel metal2 s 11794 47200 11850 48000 6 wbs_adr_i[5]
port 57 nsew signal input
rlabel metal2 s 12530 47200 12586 48000 6 wbs_adr_i[6]
port 58 nsew signal input
rlabel metal2 s 13266 47200 13322 48000 6 wbs_adr_i[7]
port 59 nsew signal input
rlabel metal2 s 14094 47200 14150 48000 6 wbs_adr_i[8]
port 60 nsew signal input
rlabel metal2 s 14830 47200 14886 48000 6 wbs_adr_i[9]
port 61 nsew signal input
rlabel metal2 s 3422 47200 3478 48000 6 wbs_cyc_i
port 62 nsew signal input
rlabel metal3 s 31200 280 32000 400 6 wbs_dat_i[0]
port 63 nsew signal input
rlabel metal3 s 31200 7624 32000 7744 6 wbs_dat_i[10]
port 64 nsew signal input
rlabel metal3 s 31200 8304 32000 8424 6 wbs_dat_i[11]
port 65 nsew signal input
rlabel metal3 s 31200 9120 32000 9240 6 wbs_dat_i[12]
port 66 nsew signal input
rlabel metal3 s 31200 9800 32000 9920 6 wbs_dat_i[13]
port 67 nsew signal input
rlabel metal3 s 31200 10616 32000 10736 6 wbs_dat_i[14]
port 68 nsew signal input
rlabel metal3 s 31200 11296 32000 11416 6 wbs_dat_i[15]
port 69 nsew signal input
rlabel metal3 s 31200 11976 32000 12096 6 wbs_dat_i[16]
port 70 nsew signal input
rlabel metal3 s 31200 12792 32000 12912 6 wbs_dat_i[17]
port 71 nsew signal input
rlabel metal3 s 31200 13472 32000 13592 6 wbs_dat_i[18]
port 72 nsew signal input
rlabel metal3 s 31200 14288 32000 14408 6 wbs_dat_i[19]
port 73 nsew signal input
rlabel metal3 s 31200 960 32000 1080 6 wbs_dat_i[1]
port 74 nsew signal input
rlabel metal3 s 31200 14968 32000 15088 6 wbs_dat_i[20]
port 75 nsew signal input
rlabel metal3 s 31200 15784 32000 15904 6 wbs_dat_i[21]
port 76 nsew signal input
rlabel metal3 s 31200 16464 32000 16584 6 wbs_dat_i[22]
port 77 nsew signal input
rlabel metal3 s 31200 17144 32000 17264 6 wbs_dat_i[23]
port 78 nsew signal input
rlabel metal3 s 31200 17960 32000 18080 6 wbs_dat_i[24]
port 79 nsew signal input
rlabel metal3 s 31200 18640 32000 18760 6 wbs_dat_i[25]
port 80 nsew signal input
rlabel metal3 s 31200 19456 32000 19576 6 wbs_dat_i[26]
port 81 nsew signal input
rlabel metal3 s 31200 20136 32000 20256 6 wbs_dat_i[27]
port 82 nsew signal input
rlabel metal3 s 31200 20952 32000 21072 6 wbs_dat_i[28]
port 83 nsew signal input
rlabel metal3 s 31200 21632 32000 21752 6 wbs_dat_i[29]
port 84 nsew signal input
rlabel metal3 s 31200 1640 32000 1760 6 wbs_dat_i[2]
port 85 nsew signal input
rlabel metal3 s 31200 22312 32000 22432 6 wbs_dat_i[30]
port 86 nsew signal input
rlabel metal3 s 31200 23128 32000 23248 6 wbs_dat_i[31]
port 87 nsew signal input
rlabel metal3 s 31200 2456 32000 2576 6 wbs_dat_i[3]
port 88 nsew signal input
rlabel metal3 s 31200 3136 32000 3256 6 wbs_dat_i[4]
port 89 nsew signal input
rlabel metal3 s 31200 3952 32000 4072 6 wbs_dat_i[5]
port 90 nsew signal input
rlabel metal3 s 31200 4632 32000 4752 6 wbs_dat_i[6]
port 91 nsew signal input
rlabel metal3 s 31200 5448 32000 5568 6 wbs_dat_i[7]
port 92 nsew signal input
rlabel metal3 s 31200 6128 32000 6248 6 wbs_dat_i[8]
port 93 nsew signal input
rlabel metal3 s 31200 6808 32000 6928 6 wbs_dat_i[9]
port 94 nsew signal input
rlabel metal3 s 31200 23808 32000 23928 6 wbs_dat_o[0]
port 95 nsew signal tristate
rlabel metal3 s 31200 31288 32000 31408 6 wbs_dat_o[10]
port 96 nsew signal tristate
rlabel metal3 s 31200 31968 32000 32088 6 wbs_dat_o[11]
port 97 nsew signal tristate
rlabel metal3 s 31200 32648 32000 32768 6 wbs_dat_o[12]
port 98 nsew signal tristate
rlabel metal3 s 31200 33464 32000 33584 6 wbs_dat_o[13]
port 99 nsew signal tristate
rlabel metal3 s 31200 34144 32000 34264 6 wbs_dat_o[14]
port 100 nsew signal tristate
rlabel metal3 s 31200 34960 32000 35080 6 wbs_dat_o[15]
port 101 nsew signal tristate
rlabel metal3 s 31200 35640 32000 35760 6 wbs_dat_o[16]
port 102 nsew signal tristate
rlabel metal3 s 31200 36456 32000 36576 6 wbs_dat_o[17]
port 103 nsew signal tristate
rlabel metal3 s 31200 37136 32000 37256 6 wbs_dat_o[18]
port 104 nsew signal tristate
rlabel metal3 s 31200 37816 32000 37936 6 wbs_dat_o[19]
port 105 nsew signal tristate
rlabel metal3 s 31200 24624 32000 24744 6 wbs_dat_o[1]
port 106 nsew signal tristate
rlabel metal3 s 31200 38632 32000 38752 6 wbs_dat_o[20]
port 107 nsew signal tristate
rlabel metal3 s 31200 39312 32000 39432 6 wbs_dat_o[21]
port 108 nsew signal tristate
rlabel metal3 s 31200 40128 32000 40248 6 wbs_dat_o[22]
port 109 nsew signal tristate
rlabel metal3 s 31200 40808 32000 40928 6 wbs_dat_o[23]
port 110 nsew signal tristate
rlabel metal3 s 31200 41624 32000 41744 6 wbs_dat_o[24]
port 111 nsew signal tristate
rlabel metal3 s 31200 42304 32000 42424 6 wbs_dat_o[25]
port 112 nsew signal tristate
rlabel metal3 s 31200 42984 32000 43104 6 wbs_dat_o[26]
port 113 nsew signal tristate
rlabel metal3 s 31200 43800 32000 43920 6 wbs_dat_o[27]
port 114 nsew signal tristate
rlabel metal3 s 31200 44480 32000 44600 6 wbs_dat_o[28]
port 115 nsew signal tristate
rlabel metal3 s 31200 45296 32000 45416 6 wbs_dat_o[29]
port 116 nsew signal tristate
rlabel metal3 s 31200 25304 32000 25424 6 wbs_dat_o[2]
port 117 nsew signal tristate
rlabel metal3 s 31200 45976 32000 46096 6 wbs_dat_o[30]
port 118 nsew signal tristate
rlabel metal3 s 31200 46792 32000 46912 6 wbs_dat_o[31]
port 119 nsew signal tristate
rlabel metal3 s 31200 26120 32000 26240 6 wbs_dat_o[3]
port 120 nsew signal tristate
rlabel metal3 s 31200 26800 32000 26920 6 wbs_dat_o[4]
port 121 nsew signal tristate
rlabel metal3 s 31200 27480 32000 27600 6 wbs_dat_o[5]
port 122 nsew signal tristate
rlabel metal3 s 31200 28296 32000 28416 6 wbs_dat_o[6]
port 123 nsew signal tristate
rlabel metal3 s 31200 28976 32000 29096 6 wbs_dat_o[7]
port 124 nsew signal tristate
rlabel metal3 s 31200 29792 32000 29912 6 wbs_dat_o[8]
port 125 nsew signal tristate
rlabel metal3 s 31200 30472 32000 30592 6 wbs_dat_o[9]
port 126 nsew signal tristate
rlabel metal2 s 4894 47200 4950 48000 6 wbs_sel_i[0]
port 127 nsew signal input
rlabel metal2 s 5722 47200 5778 48000 6 wbs_sel_i[1]
port 128 nsew signal input
rlabel metal2 s 6458 47200 6514 48000 6 wbs_sel_i[2]
port 129 nsew signal input
rlabel metal2 s 7194 47200 7250 48000 6 wbs_sel_i[3]
port 130 nsew signal input
rlabel metal2 s 2594 47200 2650 48000 6 wbs_stb_i
port 131 nsew signal input
rlabel metal2 s 4158 47200 4214 48000 6 wbs_we_i
port 132 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32000 48000
<< end >>
