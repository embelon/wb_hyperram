`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  reg [0:0] PI_wb_clk_i;
  reg [0:0] PI_rst_i;
  reg [0:0] PI_wb_rst_i;
  reg [0:0] PI_wbs_we_i;
  reg [0:0] PI_wbs_stb_i;
  reg [31:0] PI_wbs_dat_i;
  reg [31:0] PI_wbs_addr_i;
  reg [0:0] PI_hb_rwds_i;
  reg [7:0] PI_hb_dq_i;
  reg [3:0] PI_wbs_sel_i;
  reg [0:0] PI_wbs_cyc_i;
  wb_hyperram UUT (
    .wb_clk_i(PI_wb_clk_i),
    .rst_i(PI_rst_i),
    .wb_rst_i(PI_wb_rst_i),
    .wbs_we_i(PI_wbs_we_i),
    .wbs_stb_i(PI_wbs_stb_i),
    .wbs_dat_i(PI_wbs_dat_i),
    .wbs_addr_i(PI_wbs_addr_i),
    .hb_rwds_i(PI_hb_rwds_i),
    .hb_dq_i(PI_hb_dq_i),
    .wbs_sel_i(PI_wbs_sel_i),
    .wbs_cyc_i(PI_wbs_cyc_i)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    // UUT.$and$wb_hyperram.\v:0$461_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$470_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$474_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$492_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$505_Y  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:156:execute$4351  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:156:execute$4361  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:168:execute$4353  = 1'b1;
    // UUT.$auto$clk2fflogic.\cc:192:execute$4357  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:192:execute$4367  = 1'b0;
    // UUT.$eq$wb_hyperram.\v:419$652_Y  = 1'b0;
    // UUT.$eq$wb_hyperram.\v:528$794_Y  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:254$128_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:254$128_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:256$129_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:256$129_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:260$130_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:260$130_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:265$131_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:265$131_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:267$132_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:267$132_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:272$133_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:272$133_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:274$134_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:274$134_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:306$135_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:306$135_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:307$136_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:311$137_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:311$137_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:312$138_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:313$139_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:314$140_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:315$141_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:316$142_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:320$143_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:320$143_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:321$144_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:322$145_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:323$146_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:324$147_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:333$148_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:334$149_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:335$150_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:336$151_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:340$152_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:343$153_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:346$154_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:349$155_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:354$156_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:370$157_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:384$158_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:399$159_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:413$160_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:429$161_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:445$162_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:458$163_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:474$164_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:494$165_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:508$166_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:508$166_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:515$167_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:515$167_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:517$168_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:517$168_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:519$169_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:519$169_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:521$170_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:521$170_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:523$171_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:523$171_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:530$172_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:530$172_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:532$173_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:532$173_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:534$174_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:534$174_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:536$175_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:536$175_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:543$176_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:543$176_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:545$177_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:545$177_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:551$178_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:551$178_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:553$179_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:553$179_EN  = 1'b0;
    // UUT.$past$wb_hyperram.\v:314$17$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:315$18$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:316$19$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:317$20$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:333$25$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:334$26$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:335$28$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:358$30$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:359$31$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:365$36$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:365$37$0  = 6'b000000;
    // UUT.$past$wb_hyperram.\v:374$40$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:377$42$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:388$48$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:391$50$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:392$51$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:403$58$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:406$60$0  = 5'b00000;
    // UUT.$past$wb_hyperram.\v:431$72$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:432$73$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:438$77$0  = 3'b000;
    // UUT.$past$wb_hyperram.\v:476$91$0  = 1'b0;
    UUT.f_past_valid = 1'b0;
    // UUT.hram.$and$hyperram.\v:0$1506_Y  = 1'b0;
    // UUT.hram.$and$hyperram.\v:0$1515_Y  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4151  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4161  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4171  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4181  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4191  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4201  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4211  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4221  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4231  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4241  = 5'b00001;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4251  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4261  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4271  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4281  = 48'b000000000000000000000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4291  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4301  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4311  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4321  = 3'b010;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4331  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4341  = 6'b100000;
    // UUT.hram.$auto$clk2fflogic.\cc:168:execute$4153  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:168:execute$4203  = 1'b1;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4157  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4167  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4177  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4187  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4197  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4207  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4217  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4227  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4237  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4247  = 5'b00000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4257  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4267  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4277  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4287  = 48'b000000000000000000000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4297  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4307  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4317  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4327  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4337  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4347  = 6'b000000;
    // UUT.hram.$formal$hyperram.\v:1001$1139_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1001$1139_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1004$1140_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1004$1140_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1007$1141_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1007$1141_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1012$1142_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1015$1143_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1015$1143_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1018$1144_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1018$1144_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1021$1145_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1021$1145_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1024$1146_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1024$1146_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1029$1147_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1033$1148_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1033$1148_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1035$1149_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1035$1149_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1039$1150_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1039$1150_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1047$1152_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1047$1152_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1052$1153_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1052$1153_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1055$1154_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1055$1154_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1056$1155_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1056$1155_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1057$1156_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1057$1156_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1058$1157_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1058$1157_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1066$1158_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1066$1158_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1067$1159_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1068$1160_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1069$1161_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:395$1084_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:395$1084_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:398$1085_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:398$1085_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:848$1086_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:848$1086_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:854$1087_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:855$1088_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:861$1089_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:861$1089_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:862$1090_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:863$1091_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:866$1092_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:866$1092_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:868$1093_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:868$1093_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:871$1094_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:871$1094_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:873$1095_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:873$1095_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:873$1096_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:875$1097_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:883$1098_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:883$1098_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:885$1099_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:885$1099_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:889$1100_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:889$1100_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:890$1101_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:890$1101_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:891$1102_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:891$1102_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:892$1103_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:892$1103_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:893$1104_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:893$1104_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:894$1105_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:894$1105_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:900$1106_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:900$1106_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:901$1107_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:901$1107_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:902$1108_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:902$1108_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:903$1109_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:903$1109_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:911$1110_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:911$1110_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:913$1111_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:913$1111_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:917$1112_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:917$1112_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:919$1113_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:919$1113_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:926$1114_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:926$1114_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:927$1115_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:928$1116_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:929$1117_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:931$1118_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:931$1118_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:937$1119_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:937$1119_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:941$1120_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:941$1120_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:944$1121_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:944$1121_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:947$1122_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:947$1122_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:950$1123_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:950$1123_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:953$1124_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:953$1124_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:956$1125_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:956$1125_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:959$1126_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:959$1126_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:962$1127_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:962$1127_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:965$1128_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:965$1128_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:968$1129_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:968$1129_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:974$1130_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:974$1130_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:977$1131_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:977$1131_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:980$1132_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:980$1132_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:983$1133_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:983$1133_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:987$1134_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:987$1134_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:989$1135_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:989$1135_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:993$1136_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:993$1136_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:995$1137_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:995$1137_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:997$1138_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:997$1138_EN  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1014$1049$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1014$1050$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1046$1061$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1046$1062$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1051$1066$0  = 8'b00000000;
    // UUT.hram.$past$hyperram.\v:1066$1076$0  = 32'b00000000000000000000000000000000;
    // UUT.hram.$past$hyperram.\v:1067$1077$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:1068$1078$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1069$1079$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:861$998$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:862$999$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:863$1000$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:865$1001$0  = 5'b00000;
    // UUT.hram.$past$hyperram.\v:870$1003$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:875$1005$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:876$1006$0  = 1'b0;
    UUT.hram.f_past_valid = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4131  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4133  = 1'b1;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4137  = 6'b000000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4111  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4113  = 1'b1;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4117  = 4'b0000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4121  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4123  = 1'b1;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4127  = 8'b00000000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4141  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4143  = 1'b1;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4147  = 5'b00000;
    UUT.wb_state = 2'b00;

    // state 0
    PI_wb_clk_i = 1'b0;
    PI_rst_i = 1'b1;
    PI_wb_rst_i = 1'b1;
    PI_wbs_we_i = 1'b0;
    PI_wbs_stb_i = 1'b0;
    PI_wbs_dat_i = 32'b10000000000000000000000000000000;
    PI_wbs_addr_i = 32'b00000000000000000000000010000000;
    PI_hb_rwds_i = 1'b0;
    PI_hb_dq_i = 8'b00000000;
    PI_wbs_sel_i = 4'b1000;
    PI_wbs_cyc_i = 1'b0;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      PI_wb_clk_i <= 1'b1;
      PI_rst_i <= 1'b1;
      PI_wb_rst_i <= 1'b1;
      PI_wbs_we_i <= 1'b0;
      PI_wbs_stb_i <= 1'b0;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
      PI_hb_rwds_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_sel_i <= 4'b0000;
      PI_wbs_cyc_i <= 1'b0;
    end

    // state 2
    if (cycle == 1) begin
      PI_wb_clk_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_we_i <= 1'b0;
      PI_wbs_stb_i <= 1'b0;
      PI_wbs_dat_i <= 32'b10000000000000000000000000000000;
      PI_wbs_addr_i <= 32'b00000000000000000000000010000000;
      PI_hb_rwds_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_sel_i <= 4'b1000;
      PI_wbs_cyc_i <= 1'b0;
    end

    // state 3
    if (cycle == 2) begin
      PI_wb_clk_i <= 1'b1;
      PI_rst_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_we_i <= 1'b0;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
      PI_hb_rwds_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_sel_i <= 4'b0000;
      PI_wbs_cyc_i <= 1'b1;
    end

    // state 4
    if (cycle == 3) begin
      PI_wb_clk_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_we_i <= 1'b1;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_dat_i <= 32'b00000000000000000000000000001001;
      PI_wbs_addr_i <= 32'b00110100000000100000000000001000;
      PI_hb_rwds_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_sel_i <= 4'b1001;
      PI_wbs_cyc_i <= 1'b1;
    end

    // state 5
    if (cycle == 4) begin
      PI_wb_clk_i <= 1'b1;
      PI_rst_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_we_i <= 1'b1;
      PI_wbs_stb_i <= 1'b1;
      PI_wbs_dat_i <= 32'b00000000000000000000000000001001;
      PI_wbs_addr_i <= 32'b00110100000000100000000000001000;
      PI_hb_rwds_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_sel_i <= 4'b1001;
      PI_wbs_cyc_i <= 1'b1;
    end

    // state 6
    if (cycle == 5) begin
      PI_wb_clk_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_we_i <= 1'b0;
      PI_wbs_stb_i <= 1'b0;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
      PI_hb_rwds_i <= 1'b0;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_sel_i <= 4'b0000;
      PI_wbs_cyc_i <= 1'b0;
    end

    genclock <= cycle < 6;
    cycle <= cycle + 1;
  end
endmodule
