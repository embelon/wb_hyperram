module dump();
    initial begin
        $dumpfile ("wb_hyperram.vcd");
        $dumpvars (0, test_top);
        #1;
    end
endmodule
