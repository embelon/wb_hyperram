VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_hyperram
  CLASS BLOCK ;
  FOREIGN wb_hyperram ;
  ORIGIN 0.000 0.000 ;
  SIZE 160.000 BY 240.000 ;
  PIN hb_clk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 24.520 160.000 25.120 ;
    END
  END hb_clk_o
  PIN hb_clkn_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 34.720 160.000 35.320 ;
    END
  END hb_clkn_o
  PIN hb_csn_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 14.320 160.000 14.920 ;
    END
  END hb_csn_o
  PIN hb_dq_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 164.600 160.000 165.200 ;
    END
  END hb_dq_i[0]
  PIN hb_dq_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 174.800 160.000 175.400 ;
    END
  END hb_dq_i[1]
  PIN hb_dq_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 184.320 160.000 184.920 ;
    END
  END hb_dq_i[2]
  PIN hb_dq_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 194.520 160.000 195.120 ;
    END
  END hb_dq_i[3]
  PIN hb_dq_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 204.720 160.000 205.320 ;
    END
  END hb_dq_i[4]
  PIN hb_dq_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 214.240 160.000 214.840 ;
    END
  END hb_dq_i[5]
  PIN hb_dq_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 224.440 160.000 225.040 ;
    END
  END hb_dq_i[6]
  PIN hb_dq_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 234.640 160.000 235.240 ;
    END
  END hb_dq_i[7]
  PIN hb_dq_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 74.160 160.000 74.760 ;
    END
  END hb_dq_o[0]
  PIN hb_dq_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 84.360 160.000 84.960 ;
    END
  END hb_dq_o[1]
  PIN hb_dq_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 94.560 160.000 95.160 ;
    END
  END hb_dq_o[2]
  PIN hb_dq_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 104.760 160.000 105.360 ;
    END
  END hb_dq_o[3]
  PIN hb_dq_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 114.280 160.000 114.880 ;
    END
  END hb_dq_o[4]
  PIN hb_dq_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 124.480 160.000 125.080 ;
    END
  END hb_dq_o[5]
  PIN hb_dq_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 134.680 160.000 135.280 ;
    END
  END hb_dq_o[6]
  PIN hb_dq_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 144.200 160.000 144.800 ;
    END
  END hb_dq_o[7]
  PIN hb_dq_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 64.640 160.000 65.240 ;
    END
  END hb_dq_oen
  PIN hb_rstn_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 4.800 160.000 5.400 ;
    END
  END hb_rstn_o
  PIN hb_rwds_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 154.400 160.000 155.000 ;
    END
  END hb_rwds_i
  PIN hb_rwds_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 44.240 160.000 44.840 ;
    END
  END hb_rwds_o
  PIN hb_rwds_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 54.440 160.000 55.040 ;
    END
  END hb_rwds_oen
  PIN rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END rst_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.545 10.640 31.145 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.195 10.640 80.795 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.850 10.640 130.450 228.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 54.370 10.640 55.970 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.025 10.640 105.625 228.720 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 154.875 228.565 ;
      LAYER met1 ;
        RECT 1.910 6.840 158.170 228.720 ;
      LAYER met2 ;
        RECT 1.940 4.280 158.140 237.845 ;
        RECT 2.490 1.515 5.330 4.280 ;
        RECT 6.170 1.515 9.010 4.280 ;
        RECT 9.850 1.515 12.690 4.280 ;
        RECT 13.530 1.515 16.830 4.280 ;
        RECT 17.670 1.515 20.510 4.280 ;
        RECT 21.350 1.515 24.190 4.280 ;
        RECT 25.030 1.515 28.330 4.280 ;
        RECT 29.170 1.515 32.010 4.280 ;
        RECT 32.850 1.515 35.690 4.280 ;
        RECT 36.530 1.515 39.370 4.280 ;
        RECT 40.210 1.515 43.510 4.280 ;
        RECT 44.350 1.515 47.190 4.280 ;
        RECT 48.030 1.515 50.870 4.280 ;
        RECT 51.710 1.515 55.010 4.280 ;
        RECT 55.850 1.515 58.690 4.280 ;
        RECT 59.530 1.515 62.370 4.280 ;
        RECT 63.210 1.515 66.050 4.280 ;
        RECT 66.890 1.515 70.190 4.280 ;
        RECT 71.030 1.515 73.870 4.280 ;
        RECT 74.710 1.515 77.550 4.280 ;
        RECT 78.390 1.515 81.690 4.280 ;
        RECT 82.530 1.515 85.370 4.280 ;
        RECT 86.210 1.515 89.050 4.280 ;
        RECT 89.890 1.515 92.730 4.280 ;
        RECT 93.570 1.515 96.870 4.280 ;
        RECT 97.710 1.515 100.550 4.280 ;
        RECT 101.390 1.515 104.230 4.280 ;
        RECT 105.070 1.515 108.370 4.280 ;
        RECT 109.210 1.515 112.050 4.280 ;
        RECT 112.890 1.515 115.730 4.280 ;
        RECT 116.570 1.515 119.410 4.280 ;
        RECT 120.250 1.515 123.550 4.280 ;
        RECT 124.390 1.515 127.230 4.280 ;
        RECT 128.070 1.515 130.910 4.280 ;
        RECT 131.750 1.515 135.050 4.280 ;
        RECT 135.890 1.515 138.730 4.280 ;
        RECT 139.570 1.515 142.410 4.280 ;
        RECT 143.250 1.515 146.090 4.280 ;
        RECT 146.930 1.515 150.230 4.280 ;
        RECT 151.070 1.515 153.910 4.280 ;
        RECT 154.750 1.515 157.590 4.280 ;
      LAYER met3 ;
        RECT 4.400 236.960 156.000 237.825 ;
        RECT 4.000 235.640 156.000 236.960 ;
        RECT 4.000 234.960 155.600 235.640 ;
        RECT 4.400 234.240 155.600 234.960 ;
        RECT 4.400 233.560 156.000 234.240 ;
        RECT 4.000 230.880 156.000 233.560 ;
        RECT 4.400 229.480 156.000 230.880 ;
        RECT 4.000 227.480 156.000 229.480 ;
        RECT 4.400 226.080 156.000 227.480 ;
        RECT 4.000 225.440 156.000 226.080 ;
        RECT 4.000 224.040 155.600 225.440 ;
        RECT 4.000 223.400 156.000 224.040 ;
        RECT 4.400 222.000 156.000 223.400 ;
        RECT 4.000 220.000 156.000 222.000 ;
        RECT 4.400 218.600 156.000 220.000 ;
        RECT 4.000 215.920 156.000 218.600 ;
        RECT 4.400 215.240 156.000 215.920 ;
        RECT 4.400 214.520 155.600 215.240 ;
        RECT 4.000 213.840 155.600 214.520 ;
        RECT 4.000 212.520 156.000 213.840 ;
        RECT 4.400 211.120 156.000 212.520 ;
        RECT 4.000 209.120 156.000 211.120 ;
        RECT 4.400 207.720 156.000 209.120 ;
        RECT 4.000 205.720 156.000 207.720 ;
        RECT 4.000 205.040 155.600 205.720 ;
        RECT 4.400 204.320 155.600 205.040 ;
        RECT 4.400 203.640 156.000 204.320 ;
        RECT 4.000 201.640 156.000 203.640 ;
        RECT 4.400 200.240 156.000 201.640 ;
        RECT 4.000 197.560 156.000 200.240 ;
        RECT 4.400 196.160 156.000 197.560 ;
        RECT 4.000 195.520 156.000 196.160 ;
        RECT 4.000 194.160 155.600 195.520 ;
        RECT 4.400 194.120 155.600 194.160 ;
        RECT 4.400 192.760 156.000 194.120 ;
        RECT 4.000 190.080 156.000 192.760 ;
        RECT 4.400 188.680 156.000 190.080 ;
        RECT 4.000 186.680 156.000 188.680 ;
        RECT 4.400 185.320 156.000 186.680 ;
        RECT 4.400 185.280 155.600 185.320 ;
        RECT 4.000 183.920 155.600 185.280 ;
        RECT 4.000 183.280 156.000 183.920 ;
        RECT 4.400 181.880 156.000 183.280 ;
        RECT 4.000 179.200 156.000 181.880 ;
        RECT 4.400 177.800 156.000 179.200 ;
        RECT 4.000 175.800 156.000 177.800 ;
        RECT 4.400 174.400 155.600 175.800 ;
        RECT 4.000 171.720 156.000 174.400 ;
        RECT 4.400 170.320 156.000 171.720 ;
        RECT 4.000 168.320 156.000 170.320 ;
        RECT 4.400 166.920 156.000 168.320 ;
        RECT 4.000 165.600 156.000 166.920 ;
        RECT 4.000 164.240 155.600 165.600 ;
        RECT 4.400 164.200 155.600 164.240 ;
        RECT 4.400 162.840 156.000 164.200 ;
        RECT 4.000 160.840 156.000 162.840 ;
        RECT 4.400 159.440 156.000 160.840 ;
        RECT 4.000 157.440 156.000 159.440 ;
        RECT 4.400 156.040 156.000 157.440 ;
        RECT 4.000 155.400 156.000 156.040 ;
        RECT 4.000 154.000 155.600 155.400 ;
        RECT 4.000 153.360 156.000 154.000 ;
        RECT 4.400 151.960 156.000 153.360 ;
        RECT 4.000 149.960 156.000 151.960 ;
        RECT 4.400 148.560 156.000 149.960 ;
        RECT 4.000 145.880 156.000 148.560 ;
        RECT 4.400 145.200 156.000 145.880 ;
        RECT 4.400 144.480 155.600 145.200 ;
        RECT 4.000 143.800 155.600 144.480 ;
        RECT 4.000 142.480 156.000 143.800 ;
        RECT 4.400 141.080 156.000 142.480 ;
        RECT 4.000 138.400 156.000 141.080 ;
        RECT 4.400 137.000 156.000 138.400 ;
        RECT 4.000 135.680 156.000 137.000 ;
        RECT 4.000 135.000 155.600 135.680 ;
        RECT 4.400 134.280 155.600 135.000 ;
        RECT 4.400 133.600 156.000 134.280 ;
        RECT 4.000 131.600 156.000 133.600 ;
        RECT 4.400 130.200 156.000 131.600 ;
        RECT 4.000 127.520 156.000 130.200 ;
        RECT 4.400 126.120 156.000 127.520 ;
        RECT 4.000 125.480 156.000 126.120 ;
        RECT 4.000 124.120 155.600 125.480 ;
        RECT 4.400 124.080 155.600 124.120 ;
        RECT 4.400 122.720 156.000 124.080 ;
        RECT 4.000 120.040 156.000 122.720 ;
        RECT 4.400 118.640 156.000 120.040 ;
        RECT 4.000 116.640 156.000 118.640 ;
        RECT 4.400 115.280 156.000 116.640 ;
        RECT 4.400 115.240 155.600 115.280 ;
        RECT 4.000 113.880 155.600 115.240 ;
        RECT 4.000 112.560 156.000 113.880 ;
        RECT 4.400 111.160 156.000 112.560 ;
        RECT 4.000 109.160 156.000 111.160 ;
        RECT 4.400 107.760 156.000 109.160 ;
        RECT 4.000 105.760 156.000 107.760 ;
        RECT 4.400 104.360 155.600 105.760 ;
        RECT 4.000 101.680 156.000 104.360 ;
        RECT 4.400 100.280 156.000 101.680 ;
        RECT 4.000 98.280 156.000 100.280 ;
        RECT 4.400 96.880 156.000 98.280 ;
        RECT 4.000 95.560 156.000 96.880 ;
        RECT 4.000 94.200 155.600 95.560 ;
        RECT 4.400 94.160 155.600 94.200 ;
        RECT 4.400 92.800 156.000 94.160 ;
        RECT 4.000 90.800 156.000 92.800 ;
        RECT 4.400 89.400 156.000 90.800 ;
        RECT 4.000 86.720 156.000 89.400 ;
        RECT 4.400 85.360 156.000 86.720 ;
        RECT 4.400 85.320 155.600 85.360 ;
        RECT 4.000 83.960 155.600 85.320 ;
        RECT 4.000 83.320 156.000 83.960 ;
        RECT 4.400 81.920 156.000 83.320 ;
        RECT 4.000 79.920 156.000 81.920 ;
        RECT 4.400 78.520 156.000 79.920 ;
        RECT 4.000 75.840 156.000 78.520 ;
        RECT 4.400 75.160 156.000 75.840 ;
        RECT 4.400 74.440 155.600 75.160 ;
        RECT 4.000 73.760 155.600 74.440 ;
        RECT 4.000 72.440 156.000 73.760 ;
        RECT 4.400 71.040 156.000 72.440 ;
        RECT 4.000 68.360 156.000 71.040 ;
        RECT 4.400 66.960 156.000 68.360 ;
        RECT 4.000 65.640 156.000 66.960 ;
        RECT 4.000 64.960 155.600 65.640 ;
        RECT 4.400 64.240 155.600 64.960 ;
        RECT 4.400 63.560 156.000 64.240 ;
        RECT 4.000 60.880 156.000 63.560 ;
        RECT 4.400 59.480 156.000 60.880 ;
        RECT 4.000 57.480 156.000 59.480 ;
        RECT 4.400 56.080 156.000 57.480 ;
        RECT 4.000 55.440 156.000 56.080 ;
        RECT 4.000 54.080 155.600 55.440 ;
        RECT 4.400 54.040 155.600 54.080 ;
        RECT 4.400 52.680 156.000 54.040 ;
        RECT 4.000 50.000 156.000 52.680 ;
        RECT 4.400 48.600 156.000 50.000 ;
        RECT 4.000 46.600 156.000 48.600 ;
        RECT 4.400 45.240 156.000 46.600 ;
        RECT 4.400 45.200 155.600 45.240 ;
        RECT 4.000 43.840 155.600 45.200 ;
        RECT 4.000 42.520 156.000 43.840 ;
        RECT 4.400 41.120 156.000 42.520 ;
        RECT 4.000 39.120 156.000 41.120 ;
        RECT 4.400 37.720 156.000 39.120 ;
        RECT 4.000 35.720 156.000 37.720 ;
        RECT 4.000 35.040 155.600 35.720 ;
        RECT 4.400 34.320 155.600 35.040 ;
        RECT 4.400 33.640 156.000 34.320 ;
        RECT 4.000 31.640 156.000 33.640 ;
        RECT 4.400 30.240 156.000 31.640 ;
        RECT 4.000 28.240 156.000 30.240 ;
        RECT 4.400 26.840 156.000 28.240 ;
        RECT 4.000 25.520 156.000 26.840 ;
        RECT 4.000 24.160 155.600 25.520 ;
        RECT 4.400 24.120 155.600 24.160 ;
        RECT 4.400 22.760 156.000 24.120 ;
        RECT 4.000 20.760 156.000 22.760 ;
        RECT 4.400 19.360 156.000 20.760 ;
        RECT 4.000 16.680 156.000 19.360 ;
        RECT 4.400 15.320 156.000 16.680 ;
        RECT 4.400 15.280 155.600 15.320 ;
        RECT 4.000 13.920 155.600 15.280 ;
        RECT 4.000 13.280 156.000 13.920 ;
        RECT 4.400 11.880 156.000 13.280 ;
        RECT 4.000 9.200 156.000 11.880 ;
        RECT 4.400 7.800 156.000 9.200 ;
        RECT 4.000 5.800 156.000 7.800 ;
        RECT 4.400 4.400 155.600 5.800 ;
        RECT 4.000 2.400 156.000 4.400 ;
        RECT 4.400 1.535 156.000 2.400 ;
      LAYER met4 ;
        RECT 39.855 10.640 53.970 228.720 ;
        RECT 56.370 10.640 78.795 228.720 ;
        RECT 81.195 10.640 88.025 228.720 ;
  END
END wb_hyperram
END LIBRARY

