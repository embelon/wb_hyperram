`ifndef VERILATOR
module testbench;
  reg [4095:0] vcdfile;
  reg clock;
`else
module testbench(input clock, output reg genclock);
  initial genclock = 1;
`endif
  reg genclock = 1;
  reg [31:0] cycle = 0;
  reg [0:0] PI_wbs_stb_i;
  reg [0:0] PI_wb_clk_i;
  reg [0:0] PI_wb_rst_i;
  reg [3:0] PI_wbs_sel_i;
  reg [31:0] PI_wbs_addr_i;
  reg [7:0] PI_hb_dq_i;
  reg [31:0] PI_wbs_dat_i;
  reg [0:0] PI_hb_rwds_i;
  reg [0:0] PI_wbs_cyc_i;
  reg [0:0] PI_rst_i;
  reg [0:0] PI_wbs_we_i;
  wb_hyperram UUT (
    .wbs_stb_i(PI_wbs_stb_i),
    .wb_clk_i(PI_wb_clk_i),
    .wb_rst_i(PI_wb_rst_i),
    .wbs_sel_i(PI_wbs_sel_i),
    .wbs_addr_i(PI_wbs_addr_i),
    .hb_dq_i(PI_hb_dq_i),
    .wbs_dat_i(PI_wbs_dat_i),
    .hb_rwds_i(PI_hb_rwds_i),
    .wbs_cyc_i(PI_wbs_cyc_i),
    .rst_i(PI_rst_i),
    .wbs_we_i(PI_wbs_we_i)
  );
`ifndef VERILATOR
  initial begin
    if ($value$plusargs("vcd=%s", vcdfile)) begin
      $dumpfile(vcdfile);
      $dumpvars(0, testbench);
    end
    #5 clock = 0;
    while (genclock) begin
      #5 clock = 0;
      #5 clock = 1;
    end
  end
`endif
  initial begin
`ifndef VERILATOR
    #1;
`endif
    // UUT.$and$wb_hyperram.\v:0$463_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$472_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$476_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$494_Y  = 1'b0;
    // UUT.$and$wb_hyperram.\v:0$507_Y  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:156:execute$5077  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:156:execute$5087  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:156:execute$5097  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:168:execute$5079  = 1'b1;
    // UUT.$auto$clk2fflogic.\cc:192:execute$5083  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:192:execute$5093  = 1'b0;
    // UUT.$auto$clk2fflogic.\cc:192:execute$5103  = 1'b0;
    // UUT.$eq$wb_hyperram.\v:435$654_Y  = 1'b0;
    // UUT.$eq$wb_hyperram.\v:544$796_Y  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:270$128_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:270$128_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:272$129_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:272$129_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:276$130_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:276$130_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:281$131_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:281$131_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:283$132_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:283$132_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:288$133_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:288$133_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:290$134_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:290$134_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:322$135_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:322$135_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:323$136_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:327$137_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:327$137_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:328$138_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:329$139_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:330$140_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:331$141_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:332$142_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:336$143_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:336$143_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:337$144_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:338$145_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:339$146_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:340$147_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:349$148_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:350$149_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:351$150_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:352$151_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:356$152_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:359$153_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:362$154_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:365$155_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:370$156_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:386$157_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:400$158_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:415$159_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:429$160_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:445$161_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:461$162_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:474$163_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:490$164_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:510$165_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:524$166_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:524$166_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:531$167_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:531$167_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:533$168_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:533$168_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:535$169_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:535$169_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:537$170_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:537$170_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:539$171_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:539$171_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:546$172_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:546$172_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:548$173_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:548$173_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:550$174_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:550$174_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:552$175_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:552$175_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:559$176_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:559$176_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:561$177_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:561$177_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:567$178_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:567$178_EN  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:569$179_CHECK  = 1'b0;
    // UUT.$formal$wb_hyperram.\v:569$179_EN  = 1'b0;
    // UUT.$past$wb_hyperram.\v:330$17$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:331$18$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:332$19$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:333$20$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:349$25$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:350$26$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:351$28$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:374$30$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:375$31$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:381$36$0  = 32'b00000000000000000000000000000000;
    // UUT.$past$wb_hyperram.\v:381$37$0  = 6'b000000;
    // UUT.$past$wb_hyperram.\v:390$40$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:393$42$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:404$48$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:407$50$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:408$51$0  = 4'b0000;
    // UUT.$past$wb_hyperram.\v:419$58$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:422$60$0  = 5'b00000;
    // UUT.$past$wb_hyperram.\v:447$72$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:448$73$0  = 1'b0;
    // UUT.$past$wb_hyperram.\v:454$77$0  = 3'b000;
    // UUT.$past$wb_hyperram.\v:492$91$0  = 1'b0;
    UUT.f_past_valid = 1'b0;
    // UUT.hram.$and$hyperram.\v:0$1484_Y  = 1'b0;
    // UUT.hram.$and$hyperram.\v:0$1493_Y  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4877  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4887  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4897  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4907  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4917  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4927  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4937  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4947  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4957  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4967  = 5'b00000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4977  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4987  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$4997  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$5007  = 48'b000000000000000000000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$5017  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$5027  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$5037  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$5047  = 3'b010;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$5057  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:156:execute$5067  = 6'b100000;
    // UUT.hram.$auto$clk2fflogic.\cc:168:execute$4879  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:168:execute$4929  = 1'b1;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4883  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4893  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4903  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4913  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4923  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4933  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4943  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4953  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4963  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4973  = 5'b00000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4983  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$4993  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$5003  = 32'b00000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$5013  = 48'b000000000000000000000000000000000000000000000000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$5023  = 4'b0000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$5033  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$5043  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$5053  = 3'b000;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$5063  = 1'b0;
    // UUT.hram.$auto$clk2fflogic.\cc:192:execute$5073  = 6'b000000;
    // UUT.hram.$formal$hyperram.\v:1001$1128_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1001$1128_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1005$1129_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1005$1129_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1007$1130_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1007$1130_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1011$1131_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1011$1131_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1013$1132_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1013$1132_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1015$1133_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1015$1133_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1019$1134_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1019$1134_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1022$1135_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1022$1135_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1025$1136_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1025$1136_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1030$1137_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1033$1138_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1033$1138_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1036$1139_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1036$1139_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1039$1140_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1039$1140_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1042$1141_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1042$1141_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1047$1142_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1051$1143_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1051$1143_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1053$1144_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1053$1144_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1057$1145_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1057$1145_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1065$1147_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1065$1147_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1068$1148_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1068$1148_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1077$1149_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1077$1149_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1078$1150_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1078$1150_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1079$1151_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1079$1151_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1080$1152_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1080$1152_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1088$1153_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1088$1153_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1089$1154_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1090$1155_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:1091$1156_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:402$1085_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:402$1085_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:405$1086_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:405$1086_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:854$1087_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:854$1087_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:860$1088_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:861$1089_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:867$1090_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:867$1090_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:868$1091_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:869$1092_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:872$1093_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:872$1093_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:874$1094_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:874$1094_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:877$1095_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:877$1095_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:879$1096_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:879$1096_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:879$1097_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:881$1098_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:889$1099_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:889$1099_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:891$1100_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:891$1100_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:893$1101_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:893$1101_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:907$1102_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:907$1102_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:923$1103_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:923$1103_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:925$1104_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:925$1104_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:929$1105_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:929$1105_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:931$1106_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:931$1106_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:937$1107_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:937$1107_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:939$1108_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:939$1108_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:944$1109_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:944$1109_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:945$1110_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:946$1111_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:947$1112_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:949$1113_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:949$1113_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:955$1114_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:955$1114_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:959$1115_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:959$1115_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:962$1116_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:962$1116_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:965$1117_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:965$1117_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:968$1118_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:968$1118_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:971$1119_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:971$1119_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:974$1120_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:974$1120_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:977$1121_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:977$1121_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:980$1122_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:980$1122_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:983$1123_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:983$1123_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:986$1124_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:986$1124_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:992$1125_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:992$1125_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:995$1126_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:995$1126_EN  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:998$1127_CHECK  = 1'b0;
    // UUT.hram.$formal$hyperram.\v:998$1127_EN  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1032$1051$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1032$1052$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1064$1062$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1067$1064$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1067$1065$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1077$1069$0  = 8'b00000000;
    // UUT.hram.$past$hyperram.\v:1088$1077$0  = 32'b00000000000000000000000000000000;
    // UUT.hram.$past$hyperram.\v:1089$1078$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:1090$1079$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:1091$1080$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:867$1000$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:868$1001$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:869$1002$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:871$1003$0  = 5'b00000;
    // UUT.hram.$past$hyperram.\v:876$1005$0  = 4'b0000;
    // UUT.hram.$past$hyperram.\v:881$1007$0  = 1'b0;
    // UUT.hram.$past$hyperram.\v:882$1008$0  = 1'b0;
    UUT.hram.f_past_valid = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4487  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4497  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4507  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4517  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4527  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4537  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4547  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4557  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4567  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4577  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4587  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4597  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4607  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4489  = 1'b1;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4493  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4513  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4523  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4533  = 6'b000000;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4543  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4553  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4563  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4573  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4583  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4593  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4603  = 1'b0;
    // UUT.latency_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4613  = 6'b000000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4357  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4367  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4377  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4387  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4397  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4407  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4417  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4427  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4437  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4447  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4457  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4467  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4477  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4359  = 1'b1;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4363  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4383  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4393  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4403  = 4'b0000;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4413  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4423  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4433  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4443  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4453  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4463  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4473  = 1'b0;
    // UUT.tcsh_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4483  = 4'b0000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4617  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4627  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4637  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4647  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4657  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4667  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4677  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4687  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4697  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4707  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4717  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4727  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4737  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4619  = 1'b1;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4623  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4643  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4653  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4663  = 8'b00000000;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4673  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4683  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4693  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4703  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4713  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4723  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4733  = 1'b0;
    // UUT.tpre_tpost_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4743  = 8'b00000000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4747  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4757  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4767  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4777  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4787  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4797  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4807  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4817  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4827  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4837  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4847  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4857  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:156:execute$4867  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:168:execute$4749  = 1'b1;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4753  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4773  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4783  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4793  = 5'b00000;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4803  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4813  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4823  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4833  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4843  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4853  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4863  = 1'b0;
    // UUT.trmax_shadow_reg.$auto$clk2fflogic.\cc:192:execute$4873  = 5'b00000;
    UUT.wb_state = 2'b00;

    // state 0
    PI_wbs_stb_i = 1'b0;
    PI_wb_clk_i = 1'b0;
    PI_wb_rst_i = 1'b1;
    PI_wbs_sel_i = 4'b1000;
    PI_wbs_addr_i = 32'b00000000001000000000000000000000;
    PI_hb_dq_i = 8'b00000000;
    PI_wbs_dat_i = 32'b10000000000000000000000000000000;
    PI_hb_rwds_i = 1'b0;
    PI_wbs_cyc_i = 1'b0;
    PI_rst_i = 1'b1;
    PI_wbs_we_i = 1'b0;
  end
  always @(posedge clock) begin
    // state 1
    if (cycle == 0) begin
      PI_wbs_stb_i <= 1'b0;
      PI_wb_clk_i <= 1'b1;
      PI_wb_rst_i <= 1'b1;
      PI_wbs_sel_i <= 4'b0000;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_cyc_i <= 1'b0;
      PI_rst_i <= 1'b1;
      PI_wbs_we_i <= 1'b0;
    end

    // state 2
    if (cycle == 1) begin
      PI_wbs_stb_i <= 1'b0;
      PI_wb_clk_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_sel_i <= 4'b1000;
      PI_wbs_addr_i <= 32'b00000000001000000000000000000000;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b10000000000000000000000000000000;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_cyc_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_wbs_we_i <= 1'b0;
    end

    // state 3
    if (cycle == 2) begin
      PI_wbs_stb_i <= 1'b1;
      PI_wb_clk_i <= 1'b1;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_sel_i <= 4'b0000;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_cyc_i <= 1'b1;
      PI_rst_i <= 1'b0;
      PI_wbs_we_i <= 1'b0;
    end

    // state 4
    if (cycle == 3) begin
      PI_wbs_stb_i <= 1'b1;
      PI_wb_clk_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_sel_i <= 4'b1001;
      PI_wbs_addr_i <= 32'b00110000110000000000000000000100;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000010101101;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_cyc_i <= 1'b1;
      PI_rst_i <= 1'b0;
      PI_wbs_we_i <= 1'b1;
    end

    // state 5
    if (cycle == 4) begin
      PI_wbs_stb_i <= 1'b1;
      PI_wb_clk_i <= 1'b1;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_sel_i <= 4'b1001;
      PI_wbs_addr_i <= 32'b00110000110000000000000000000100;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000010101101;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_cyc_i <= 1'b1;
      PI_rst_i <= 1'b0;
      PI_wbs_we_i <= 1'b1;
    end

    // state 6
    if (cycle == 5) begin
      PI_wbs_stb_i <= 1'b0;
      PI_wb_clk_i <= 1'b0;
      PI_wb_rst_i <= 1'b0;
      PI_wbs_sel_i <= 4'b0000;
      PI_wbs_addr_i <= 32'b00000000000000000000000000000000;
      PI_hb_dq_i <= 8'b00000000;
      PI_wbs_dat_i <= 32'b00000000000000000000000000000000;
      PI_hb_rwds_i <= 1'b0;
      PI_wbs_cyc_i <= 1'b0;
      PI_rst_i <= 1'b0;
      PI_wbs_we_i <= 1'b0;
    end

    genclock <= cycle < 6;
    cycle <= cycle + 1;
  end
endmodule
