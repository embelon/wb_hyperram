VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_hyperram
  CLASS BLOCK ;
  FOREIGN wb_hyperram ;
  ORIGIN 0.000 0.000 ;
  SIZE 160.000 BY 240.000 ;
  PIN hb_clk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END hb_clk_o
  PIN hb_clkn_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END hb_clkn_o
  PIN hb_csn_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END hb_csn_o
  PIN hb_dq_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END hb_dq_i[0]
  PIN hb_dq_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END hb_dq_i[1]
  PIN hb_dq_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END hb_dq_i[2]
  PIN hb_dq_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END hb_dq_i[3]
  PIN hb_dq_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END hb_dq_i[4]
  PIN hb_dq_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END hb_dq_i[5]
  PIN hb_dq_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END hb_dq_i[6]
  PIN hb_dq_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END hb_dq_i[7]
  PIN hb_dq_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END hb_dq_o[0]
  PIN hb_dq_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END hb_dq_o[1]
  PIN hb_dq_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END hb_dq_o[2]
  PIN hb_dq_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END hb_dq_o[3]
  PIN hb_dq_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END hb_dq_o[4]
  PIN hb_dq_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END hb_dq_o[5]
  PIN hb_dq_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END hb_dq_o[6]
  PIN hb_dq_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END hb_dq_o[7]
  PIN hb_dq_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END hb_dq_oen
  PIN hb_rstn_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END hb_rstn_o
  PIN hb_rwds_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END hb_rwds_i
  PIN hb_rwds_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END hb_rwds_o
  PIN hb_rwds_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END hb_rwds_oen
  PIN rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 236.000 2.210 240.000 ;
    END
  END rst_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.545 10.640 31.145 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.195 10.640 80.795 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.850 10.640 130.450 228.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 54.370 10.640 55.970 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.025 10.640 105.625 228.720 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 236.000 5.890 240.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 236.000 9.570 240.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 237.360 160.000 237.960 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 236.000 39.930 240.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 236.000 78.110 240.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 236.000 82.250 240.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 236.000 85.930 240.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 236.000 89.610 240.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 236.000 93.290 240.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 236.000 97.430 240.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 236.000 101.110 240.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 236.000 104.790 240.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 236.000 108.930 240.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 236.000 112.610 240.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 236.000 44.070 240.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 236.000 116.290 240.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 236.000 119.970 240.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 236.000 124.110 240.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 236.000 127.790 240.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 236.000 131.470 240.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 236.000 135.610 240.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 236.000 139.290 240.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 236.000 142.970 240.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 236.000 146.650 240.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 236.000 150.790 240.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 236.000 47.750 240.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 236.000 154.470 240.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 236.000 158.150 240.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 236.000 51.430 240.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 236.000 55.570 240.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 236.000 59.250 240.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 236.000 62.930 240.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 236.000 66.610 240.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 236.000 70.750 240.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 236.000 74.430 240.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 236.000 17.390 240.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 1.400 160.000 2.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 38.120 160.000 38.720 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 41.520 160.000 42.120 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 45.600 160.000 46.200 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 49.000 160.000 49.600 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 53.080 160.000 53.680 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 56.480 160.000 57.080 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 59.880 160.000 60.480 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 63.960 160.000 64.560 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 67.360 160.000 67.960 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 71.440 160.000 72.040 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 4.800 160.000 5.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 74.840 160.000 75.440 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 78.920 160.000 79.520 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 82.320 160.000 82.920 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 85.720 160.000 86.320 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 89.800 160.000 90.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 93.200 160.000 93.800 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 97.280 160.000 97.880 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 100.680 160.000 101.280 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 104.760 160.000 105.360 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 108.160 160.000 108.760 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 8.200 160.000 8.800 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 111.560 160.000 112.160 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 115.640 160.000 116.240 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 12.280 160.000 12.880 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 15.680 160.000 16.280 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 19.760 160.000 20.360 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 23.160 160.000 23.760 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 27.240 160.000 27.840 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 30.640 160.000 31.240 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 34.040 160.000 34.640 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 119.040 160.000 119.640 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 156.440 160.000 157.040 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 159.840 160.000 160.440 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 163.240 160.000 163.840 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 167.320 160.000 167.920 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 170.720 160.000 171.320 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 174.800 160.000 175.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 178.200 160.000 178.800 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 182.280 160.000 182.880 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 185.680 160.000 186.280 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 189.080 160.000 189.680 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 123.120 160.000 123.720 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 193.160 160.000 193.760 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 196.560 160.000 197.160 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 200.640 160.000 201.240 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 204.040 160.000 204.640 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 208.120 160.000 208.720 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 211.520 160.000 212.120 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 214.920 160.000 215.520 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 219.000 160.000 219.600 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 222.400 160.000 223.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 226.480 160.000 227.080 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 126.520 160.000 127.120 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 229.880 160.000 230.480 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 233.960 160.000 234.560 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 130.600 160.000 131.200 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 134.000 160.000 134.600 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 137.400 160.000 138.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 141.480 160.000 142.080 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 144.880 160.000 145.480 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 148.960 160.000 149.560 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.000 152.360 160.000 152.960 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 236.000 24.750 240.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 236.000 28.890 240.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 236.000 32.570 240.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 236.000 36.250 240.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 236.000 13.250 240.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 236.000 21.070 240.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 158.095 228.565 ;
      LAYER met1 ;
        RECT 1.910 10.640 158.170 229.120 ;
      LAYER met2 ;
        RECT 2.490 235.720 5.330 237.845 ;
        RECT 6.170 235.720 9.010 237.845 ;
        RECT 9.850 235.720 12.690 237.845 ;
        RECT 13.530 235.720 16.830 237.845 ;
        RECT 17.670 235.720 20.510 237.845 ;
        RECT 21.350 235.720 24.190 237.845 ;
        RECT 25.030 235.720 28.330 237.845 ;
        RECT 29.170 235.720 32.010 237.845 ;
        RECT 32.850 235.720 35.690 237.845 ;
        RECT 36.530 235.720 39.370 237.845 ;
        RECT 40.210 235.720 43.510 237.845 ;
        RECT 44.350 235.720 47.190 237.845 ;
        RECT 48.030 235.720 50.870 237.845 ;
        RECT 51.710 235.720 55.010 237.845 ;
        RECT 55.850 235.720 58.690 237.845 ;
        RECT 59.530 235.720 62.370 237.845 ;
        RECT 63.210 235.720 66.050 237.845 ;
        RECT 66.890 235.720 70.190 237.845 ;
        RECT 71.030 235.720 73.870 237.845 ;
        RECT 74.710 235.720 77.550 237.845 ;
        RECT 78.390 235.720 81.690 237.845 ;
        RECT 82.530 235.720 85.370 237.845 ;
        RECT 86.210 235.720 89.050 237.845 ;
        RECT 89.890 235.720 92.730 237.845 ;
        RECT 93.570 235.720 96.870 237.845 ;
        RECT 97.710 235.720 100.550 237.845 ;
        RECT 101.390 235.720 104.230 237.845 ;
        RECT 105.070 235.720 108.370 237.845 ;
        RECT 109.210 235.720 112.050 237.845 ;
        RECT 112.890 235.720 115.730 237.845 ;
        RECT 116.570 235.720 119.410 237.845 ;
        RECT 120.250 235.720 123.550 237.845 ;
        RECT 124.390 235.720 127.230 237.845 ;
        RECT 128.070 235.720 130.910 237.845 ;
        RECT 131.750 235.720 135.050 237.845 ;
        RECT 135.890 235.720 138.730 237.845 ;
        RECT 139.570 235.720 142.410 237.845 ;
        RECT 143.250 235.720 146.090 237.845 ;
        RECT 146.930 235.720 150.230 237.845 ;
        RECT 151.070 235.720 153.910 237.845 ;
        RECT 154.750 235.720 157.590 237.845 ;
        RECT 1.940 1.515 158.140 235.720 ;
      LAYER met3 ;
        RECT 4.000 236.960 155.600 237.825 ;
        RECT 4.000 235.640 156.000 236.960 ;
        RECT 4.400 234.960 156.000 235.640 ;
        RECT 4.400 234.240 155.600 234.960 ;
        RECT 4.000 233.560 155.600 234.240 ;
        RECT 4.000 230.880 156.000 233.560 ;
        RECT 4.000 229.480 155.600 230.880 ;
        RECT 4.000 227.480 156.000 229.480 ;
        RECT 4.000 226.080 155.600 227.480 ;
        RECT 4.000 225.440 156.000 226.080 ;
        RECT 4.400 224.040 156.000 225.440 ;
        RECT 4.000 223.400 156.000 224.040 ;
        RECT 4.000 222.000 155.600 223.400 ;
        RECT 4.000 220.000 156.000 222.000 ;
        RECT 4.000 218.600 155.600 220.000 ;
        RECT 4.000 215.920 156.000 218.600 ;
        RECT 4.000 215.240 155.600 215.920 ;
        RECT 4.400 214.520 155.600 215.240 ;
        RECT 4.400 213.840 156.000 214.520 ;
        RECT 4.000 212.520 156.000 213.840 ;
        RECT 4.000 211.120 155.600 212.520 ;
        RECT 4.000 209.120 156.000 211.120 ;
        RECT 4.000 207.720 155.600 209.120 ;
        RECT 4.000 205.720 156.000 207.720 ;
        RECT 4.400 205.040 156.000 205.720 ;
        RECT 4.400 204.320 155.600 205.040 ;
        RECT 4.000 203.640 155.600 204.320 ;
        RECT 4.000 201.640 156.000 203.640 ;
        RECT 4.000 200.240 155.600 201.640 ;
        RECT 4.000 197.560 156.000 200.240 ;
        RECT 4.000 196.160 155.600 197.560 ;
        RECT 4.000 195.520 156.000 196.160 ;
        RECT 4.400 194.160 156.000 195.520 ;
        RECT 4.400 194.120 155.600 194.160 ;
        RECT 4.000 192.760 155.600 194.120 ;
        RECT 4.000 190.080 156.000 192.760 ;
        RECT 4.000 188.680 155.600 190.080 ;
        RECT 4.000 186.680 156.000 188.680 ;
        RECT 4.000 185.320 155.600 186.680 ;
        RECT 4.400 185.280 155.600 185.320 ;
        RECT 4.400 183.920 156.000 185.280 ;
        RECT 4.000 183.280 156.000 183.920 ;
        RECT 4.000 181.880 155.600 183.280 ;
        RECT 4.000 179.200 156.000 181.880 ;
        RECT 4.000 177.800 155.600 179.200 ;
        RECT 4.000 175.800 156.000 177.800 ;
        RECT 4.400 174.400 155.600 175.800 ;
        RECT 4.000 171.720 156.000 174.400 ;
        RECT 4.000 170.320 155.600 171.720 ;
        RECT 4.000 168.320 156.000 170.320 ;
        RECT 4.000 166.920 155.600 168.320 ;
        RECT 4.000 165.600 156.000 166.920 ;
        RECT 4.400 164.240 156.000 165.600 ;
        RECT 4.400 164.200 155.600 164.240 ;
        RECT 4.000 162.840 155.600 164.200 ;
        RECT 4.000 160.840 156.000 162.840 ;
        RECT 4.000 159.440 155.600 160.840 ;
        RECT 4.000 157.440 156.000 159.440 ;
        RECT 4.000 156.040 155.600 157.440 ;
        RECT 4.000 155.400 156.000 156.040 ;
        RECT 4.400 154.000 156.000 155.400 ;
        RECT 4.000 153.360 156.000 154.000 ;
        RECT 4.000 151.960 155.600 153.360 ;
        RECT 4.000 149.960 156.000 151.960 ;
        RECT 4.000 148.560 155.600 149.960 ;
        RECT 4.000 145.880 156.000 148.560 ;
        RECT 4.000 145.200 155.600 145.880 ;
        RECT 4.400 144.480 155.600 145.200 ;
        RECT 4.400 143.800 156.000 144.480 ;
        RECT 4.000 142.480 156.000 143.800 ;
        RECT 4.000 141.080 155.600 142.480 ;
        RECT 4.000 138.400 156.000 141.080 ;
        RECT 4.000 137.000 155.600 138.400 ;
        RECT 4.000 135.680 156.000 137.000 ;
        RECT 4.400 135.000 156.000 135.680 ;
        RECT 4.400 134.280 155.600 135.000 ;
        RECT 4.000 133.600 155.600 134.280 ;
        RECT 4.000 131.600 156.000 133.600 ;
        RECT 4.000 130.200 155.600 131.600 ;
        RECT 4.000 127.520 156.000 130.200 ;
        RECT 4.000 126.120 155.600 127.520 ;
        RECT 4.000 125.480 156.000 126.120 ;
        RECT 4.400 124.120 156.000 125.480 ;
        RECT 4.400 124.080 155.600 124.120 ;
        RECT 4.000 122.720 155.600 124.080 ;
        RECT 4.000 120.040 156.000 122.720 ;
        RECT 4.000 118.640 155.600 120.040 ;
        RECT 4.000 116.640 156.000 118.640 ;
        RECT 4.000 115.280 155.600 116.640 ;
        RECT 4.400 115.240 155.600 115.280 ;
        RECT 4.400 113.880 156.000 115.240 ;
        RECT 4.000 112.560 156.000 113.880 ;
        RECT 4.000 111.160 155.600 112.560 ;
        RECT 4.000 109.160 156.000 111.160 ;
        RECT 4.000 107.760 155.600 109.160 ;
        RECT 4.000 105.760 156.000 107.760 ;
        RECT 4.400 104.360 155.600 105.760 ;
        RECT 4.000 101.680 156.000 104.360 ;
        RECT 4.000 100.280 155.600 101.680 ;
        RECT 4.000 98.280 156.000 100.280 ;
        RECT 4.000 96.880 155.600 98.280 ;
        RECT 4.000 95.560 156.000 96.880 ;
        RECT 4.400 94.200 156.000 95.560 ;
        RECT 4.400 94.160 155.600 94.200 ;
        RECT 4.000 92.800 155.600 94.160 ;
        RECT 4.000 90.800 156.000 92.800 ;
        RECT 4.000 89.400 155.600 90.800 ;
        RECT 4.000 86.720 156.000 89.400 ;
        RECT 4.000 85.360 155.600 86.720 ;
        RECT 4.400 85.320 155.600 85.360 ;
        RECT 4.400 83.960 156.000 85.320 ;
        RECT 4.000 83.320 156.000 83.960 ;
        RECT 4.000 81.920 155.600 83.320 ;
        RECT 4.000 79.920 156.000 81.920 ;
        RECT 4.000 78.520 155.600 79.920 ;
        RECT 4.000 75.840 156.000 78.520 ;
        RECT 4.000 75.160 155.600 75.840 ;
        RECT 4.400 74.440 155.600 75.160 ;
        RECT 4.400 73.760 156.000 74.440 ;
        RECT 4.000 72.440 156.000 73.760 ;
        RECT 4.000 71.040 155.600 72.440 ;
        RECT 4.000 68.360 156.000 71.040 ;
        RECT 4.000 66.960 155.600 68.360 ;
        RECT 4.000 65.640 156.000 66.960 ;
        RECT 4.400 64.960 156.000 65.640 ;
        RECT 4.400 64.240 155.600 64.960 ;
        RECT 4.000 63.560 155.600 64.240 ;
        RECT 4.000 60.880 156.000 63.560 ;
        RECT 4.000 59.480 155.600 60.880 ;
        RECT 4.000 57.480 156.000 59.480 ;
        RECT 4.000 56.080 155.600 57.480 ;
        RECT 4.000 55.440 156.000 56.080 ;
        RECT 4.400 54.080 156.000 55.440 ;
        RECT 4.400 54.040 155.600 54.080 ;
        RECT 4.000 52.680 155.600 54.040 ;
        RECT 4.000 50.000 156.000 52.680 ;
        RECT 4.000 48.600 155.600 50.000 ;
        RECT 4.000 46.600 156.000 48.600 ;
        RECT 4.000 45.240 155.600 46.600 ;
        RECT 4.400 45.200 155.600 45.240 ;
        RECT 4.400 43.840 156.000 45.200 ;
        RECT 4.000 42.520 156.000 43.840 ;
        RECT 4.000 41.120 155.600 42.520 ;
        RECT 4.000 39.120 156.000 41.120 ;
        RECT 4.000 37.720 155.600 39.120 ;
        RECT 4.000 35.720 156.000 37.720 ;
        RECT 4.400 35.040 156.000 35.720 ;
        RECT 4.400 34.320 155.600 35.040 ;
        RECT 4.000 33.640 155.600 34.320 ;
        RECT 4.000 31.640 156.000 33.640 ;
        RECT 4.000 30.240 155.600 31.640 ;
        RECT 4.000 28.240 156.000 30.240 ;
        RECT 4.000 26.840 155.600 28.240 ;
        RECT 4.000 25.520 156.000 26.840 ;
        RECT 4.400 24.160 156.000 25.520 ;
        RECT 4.400 24.120 155.600 24.160 ;
        RECT 4.000 22.760 155.600 24.120 ;
        RECT 4.000 20.760 156.000 22.760 ;
        RECT 4.000 19.360 155.600 20.760 ;
        RECT 4.000 16.680 156.000 19.360 ;
        RECT 4.000 15.320 155.600 16.680 ;
        RECT 4.400 15.280 155.600 15.320 ;
        RECT 4.400 13.920 156.000 15.280 ;
        RECT 4.000 13.280 156.000 13.920 ;
        RECT 4.000 11.880 155.600 13.280 ;
        RECT 4.000 9.200 156.000 11.880 ;
        RECT 4.000 7.800 155.600 9.200 ;
        RECT 4.000 5.800 156.000 7.800 ;
        RECT 4.400 4.400 155.600 5.800 ;
        RECT 4.000 2.400 156.000 4.400 ;
        RECT 4.000 1.535 155.600 2.400 ;
      LAYER met4 ;
        RECT 81.195 10.640 103.625 228.720 ;
        RECT 106.025 10.640 107.345 228.720 ;
  END
END wb_hyperram
END LIBRARY

