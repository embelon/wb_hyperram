magic
tech sky130A
magscale 1 2
timestamp 1636583420
<< locali >>
rect 7757 35683 7791 35785
rect 12909 31195 12943 31433
rect 3617 28407 3651 28509
rect 6377 25687 6411 25857
rect 6377 24599 6411 24769
rect 8953 15487 8987 15657
rect 16221 9979 16255 10217
rect 6377 8415 6411 8517
rect 15853 2975 15887 3145
rect 20269 2907 20303 3009
rect 30941 2839 30975 4573
<< viali >>
rect 7113 45577 7147 45611
rect 1685 45441 1719 45475
rect 2421 45441 2455 45475
rect 3157 45441 3191 45475
rect 3985 45441 4019 45475
rect 4629 45441 4663 45475
rect 5273 45441 5307 45475
rect 6469 45441 6503 45475
rect 7297 45441 7331 45475
rect 30113 45441 30147 45475
rect 2237 45305 2271 45339
rect 2973 45305 3007 45339
rect 5089 45305 5123 45339
rect 1501 45237 1535 45271
rect 3801 45237 3835 45271
rect 4445 45237 4479 45271
rect 6653 45237 6687 45271
rect 29929 45237 29963 45271
rect 2237 45033 2271 45067
rect 5089 45033 5123 45067
rect 5273 45033 5307 45067
rect 1685 44829 1719 44863
rect 2421 44829 2455 44863
rect 3065 44829 3099 44863
rect 4077 44829 4111 44863
rect 4721 44829 4755 44863
rect 5733 44829 5767 44863
rect 7021 44829 7055 44863
rect 7205 44829 7239 44863
rect 7297 44829 7331 44863
rect 7389 44829 7423 44863
rect 7573 44829 7607 44863
rect 8217 44829 8251 44863
rect 30113 44829 30147 44863
rect 1501 44693 1535 44727
rect 2881 44693 2915 44727
rect 4261 44693 4295 44727
rect 5089 44693 5123 44727
rect 5917 44693 5951 44727
rect 6837 44693 6871 44727
rect 8033 44693 8067 44727
rect 29929 44693 29963 44727
rect 4445 44489 4479 44523
rect 4905 44489 4939 44523
rect 5089 44489 5123 44523
rect 8125 44489 8159 44523
rect 4261 44421 4295 44455
rect 6990 44421 7024 44455
rect 1685 44353 1719 44387
rect 2329 44353 2363 44387
rect 2973 44353 3007 44387
rect 6745 44353 6779 44387
rect 8769 44353 8803 44387
rect 8953 44353 8987 44387
rect 9149 44359 9183 44393
rect 9321 44353 9355 44387
rect 3893 44285 3927 44319
rect 9045 44285 9079 44319
rect 5457 44217 5491 44251
rect 1501 44149 1535 44183
rect 2145 44149 2179 44183
rect 2789 44149 2823 44183
rect 4261 44149 4295 44183
rect 5089 44149 5123 44183
rect 8585 44149 8619 44183
rect 5273 43945 5307 43979
rect 5457 43945 5491 43979
rect 20085 43945 20119 43979
rect 2329 43877 2363 43911
rect 8401 43877 8435 43911
rect 5917 43809 5951 43843
rect 8953 43809 8987 43843
rect 20453 43809 20487 43843
rect 21373 43809 21407 43843
rect 1685 43741 1719 43775
rect 2145 43741 2179 43775
rect 2973 43741 3007 43775
rect 3985 43741 4019 43775
rect 4905 43741 4939 43775
rect 8217 43741 8251 43775
rect 20269 43741 20303 43775
rect 21189 43741 21223 43775
rect 6184 43673 6218 43707
rect 9198 43673 9232 43707
rect 21005 43673 21039 43707
rect 1501 43605 1535 43639
rect 2789 43605 2823 43639
rect 3801 43605 3835 43639
rect 5273 43605 5307 43639
rect 7297 43605 7331 43639
rect 10333 43605 10367 43639
rect 6377 43401 6411 43435
rect 8125 43401 8159 43435
rect 9965 43401 9999 43435
rect 10425 43401 10459 43435
rect 8830 43333 8864 43367
rect 1685 43265 1719 43299
rect 2329 43265 2363 43299
rect 2789 43265 2823 43299
rect 3617 43265 3651 43299
rect 4261 43265 4295 43299
rect 4905 43265 4939 43299
rect 5641 43265 5675 43299
rect 6561 43265 6595 43299
rect 7389 43265 7423 43299
rect 7573 43265 7607 43299
rect 7941 43265 7975 43299
rect 10609 43265 10643 43299
rect 30113 43265 30147 43299
rect 7665 43197 7699 43231
rect 7757 43197 7791 43231
rect 8585 43197 8619 43231
rect 4721 43129 4755 43163
rect 5825 43129 5859 43163
rect 1501 43061 1535 43095
rect 2145 43061 2179 43095
rect 2973 43061 3007 43095
rect 3433 43061 3467 43095
rect 4077 43061 4111 43095
rect 29929 43061 29963 43095
rect 2513 42857 2547 42891
rect 4721 42857 4755 42891
rect 6653 42857 6687 42891
rect 8401 42857 8435 42891
rect 7021 42721 7055 42755
rect 1685 42653 1719 42687
rect 2145 42653 2179 42687
rect 3985 42653 4019 42687
rect 5089 42653 5123 42687
rect 6009 42653 6043 42687
rect 6837 42653 6871 42687
rect 7113 42653 7147 42687
rect 7205 42653 7239 42687
rect 7389 42653 7423 42687
rect 8217 42653 8251 42687
rect 9137 42653 9171 42687
rect 19809 42653 19843 42687
rect 19993 42653 20027 42687
rect 2513 42585 2547 42619
rect 1501 42517 1535 42551
rect 2697 42517 2731 42551
rect 3801 42517 3835 42551
rect 4537 42517 4571 42551
rect 4721 42517 4755 42551
rect 6193 42517 6227 42551
rect 8953 42517 8987 42551
rect 19625 42517 19659 42551
rect 3709 42313 3743 42347
rect 2513 42245 2547 42279
rect 1685 42177 1719 42211
rect 3525 42177 3559 42211
rect 4721 42177 4755 42211
rect 5641 42177 5675 42211
rect 6745 42177 6779 42211
rect 6929 42177 6963 42211
rect 7297 42177 7331 42211
rect 7941 42177 7975 42211
rect 7021 42109 7055 42143
rect 7113 42109 7147 42143
rect 2145 42041 2179 42075
rect 5825 42041 5859 42075
rect 1501 41973 1535 42007
rect 2513 41973 2547 42007
rect 2697 41973 2731 42007
rect 4905 41973 4939 42007
rect 7481 41973 7515 42007
rect 8125 41973 8159 42007
rect 2513 41769 2547 41803
rect 2697 41769 2731 41803
rect 7021 41769 7055 41803
rect 3801 41633 3835 41667
rect 5917 41633 5951 41667
rect 8401 41633 8435 41667
rect 1685 41565 1719 41599
rect 2145 41565 2179 41599
rect 5641 41565 5675 41599
rect 9137 41565 9171 41599
rect 2513 41497 2547 41531
rect 4068 41497 4102 41531
rect 8134 41497 8168 41531
rect 1501 41429 1535 41463
rect 5181 41429 5215 41463
rect 8953 41429 8987 41463
rect 2513 41225 2547 41259
rect 3985 41225 4019 41259
rect 6745 41225 6779 41259
rect 8815 41225 8849 41259
rect 16129 41225 16163 41259
rect 2329 41157 2363 41191
rect 1961 41089 1995 41123
rect 3249 41089 3283 41123
rect 3433 41089 3467 41123
rect 3812 41089 3846 41123
rect 5558 41089 5592 41123
rect 7858 41089 7892 41123
rect 8125 41089 8159 41123
rect 15945 41089 15979 41123
rect 16773 41089 16807 41123
rect 30113 41089 30147 41123
rect 3525 41021 3559 41055
rect 3617 41021 3651 41055
rect 5825 41021 5859 41055
rect 8585 41021 8619 41055
rect 2329 40885 2363 40919
rect 4445 40885 4479 40919
rect 16773 40885 16807 40919
rect 29929 40885 29963 40919
rect 2513 40681 2547 40715
rect 2697 40681 2731 40715
rect 4353 40681 4387 40715
rect 2145 40613 2179 40647
rect 4813 40545 4847 40579
rect 7205 40545 7239 40579
rect 15117 40545 15151 40579
rect 15393 40545 15427 40579
rect 15669 40545 15703 40579
rect 1685 40477 1719 40511
rect 4537 40477 4571 40511
rect 4721 40477 4755 40511
rect 4905 40477 4939 40511
rect 5089 40477 5123 40511
rect 6101 40477 6135 40511
rect 6377 40477 6411 40511
rect 6929 40477 6963 40511
rect 9137 40477 9171 40511
rect 9597 40477 9631 40511
rect 12357 40477 12391 40511
rect 13001 40477 13035 40511
rect 14473 40477 14507 40511
rect 14657 40477 14691 40511
rect 15510 40477 15544 40511
rect 16957 40477 16991 40511
rect 17693 40477 17727 40511
rect 2513 40409 2547 40443
rect 16773 40409 16807 40443
rect 17601 40409 17635 40443
rect 1501 40341 1535 40375
rect 8953 40341 8987 40375
rect 9781 40341 9815 40375
rect 12541 40341 12575 40375
rect 13185 40341 13219 40375
rect 16313 40341 16347 40375
rect 17141 40341 17175 40375
rect 4537 40137 4571 40171
rect 5181 40137 5215 40171
rect 7941 40137 7975 40171
rect 12173 40137 12207 40171
rect 15669 40137 15703 40171
rect 15301 40069 15335 40103
rect 1685 40001 1719 40035
rect 2513 40001 2547 40035
rect 3424 40001 3458 40035
rect 4997 40001 5031 40035
rect 5641 40001 5675 40035
rect 6377 40001 6411 40035
rect 6561 40001 6595 40035
rect 6929 40001 6963 40035
rect 7113 40001 7147 40035
rect 7757 40001 7791 40035
rect 8401 40001 8435 40035
rect 10158 40001 10192 40035
rect 10425 40001 10459 40035
rect 11989 40001 12023 40035
rect 12633 40001 12667 40035
rect 14473 40001 14507 40035
rect 16681 40001 16715 40035
rect 16865 40001 16899 40035
rect 17601 40001 17635 40035
rect 19165 40001 19199 40035
rect 22293 40001 22327 40035
rect 3157 39933 3191 39967
rect 6653 39933 6687 39967
rect 6745 39933 6779 39967
rect 12817 39933 12851 39967
rect 13553 39933 13587 39967
rect 13670 39933 13704 39967
rect 13829 39933 13863 39967
rect 15025 39933 15059 39967
rect 15209 39933 15243 39967
rect 17325 39933 17359 39967
rect 17718 39933 17752 39967
rect 17877 39933 17911 39967
rect 21833 39933 21867 39967
rect 22385 39933 22419 39967
rect 13277 39865 13311 39899
rect 1501 39797 1535 39831
rect 2697 39797 2731 39831
rect 5825 39797 5859 39831
rect 8585 39797 8619 39831
rect 9045 39797 9079 39831
rect 18521 39797 18555 39831
rect 18981 39797 19015 39831
rect 2329 39593 2363 39627
rect 2513 39593 2547 39627
rect 3065 39593 3099 39627
rect 3801 39593 3835 39627
rect 5733 39593 5767 39627
rect 13001 39593 13035 39627
rect 1961 39525 1995 39559
rect 4997 39525 5031 39559
rect 12173 39525 12207 39559
rect 15117 39525 15151 39559
rect 17509 39525 17543 39559
rect 4169 39457 4203 39491
rect 6745 39457 6779 39491
rect 7665 39457 7699 39491
rect 9045 39457 9079 39491
rect 14657 39457 14691 39491
rect 15393 39457 15427 39491
rect 15510 39457 15544 39491
rect 15669 39457 15703 39491
rect 16865 39457 16899 39491
rect 17049 39457 17083 39491
rect 3249 39389 3283 39423
rect 3985 39389 4019 39423
rect 4258 39389 4292 39423
rect 4353 39389 4387 39423
rect 4537 39389 4571 39423
rect 5181 39389 5215 39423
rect 5917 39389 5951 39423
rect 6377 39389 6411 39423
rect 6561 39389 6595 39423
rect 6653 39389 6687 39423
rect 6929 39389 6963 39423
rect 7757 39389 7791 39423
rect 8401 39389 8435 39423
rect 11989 39389 12023 39423
rect 14473 39389 14507 39423
rect 18153 39389 18187 39423
rect 19809 39389 19843 39423
rect 30113 39389 30147 39423
rect 2329 39321 2363 39355
rect 9312 39321 9346 39355
rect 12633 39321 12667 39355
rect 12817 39321 12851 39355
rect 16313 39321 16347 39355
rect 17141 39321 17175 39355
rect 19625 39321 19659 39355
rect 7113 39253 7147 39287
rect 8217 39253 8251 39287
rect 10425 39253 10459 39287
rect 17969 39253 18003 39287
rect 19993 39253 20027 39287
rect 29929 39253 29963 39287
rect 2605 39049 2639 39083
rect 5181 39049 5215 39083
rect 7941 39049 7975 39083
rect 9321 39049 9355 39083
rect 14381 39049 14415 39083
rect 16129 39049 16163 39083
rect 16865 39049 16899 39083
rect 17693 39049 17727 39083
rect 17785 39049 17819 39083
rect 18797 39049 18831 39083
rect 18889 39049 18923 39083
rect 19993 39049 20027 39083
rect 21925 39049 21959 39083
rect 2421 38981 2455 39015
rect 15761 38981 15795 39015
rect 1409 38913 1443 38947
rect 2053 38913 2087 38947
rect 3249 38913 3283 38947
rect 3985 38913 4019 38947
rect 4997 38913 5031 38947
rect 5641 38913 5675 38947
rect 6561 38913 6595 38947
rect 6828 38913 6862 38947
rect 8585 38913 8619 38947
rect 8769 38913 8803 38947
rect 9137 38913 9171 38947
rect 10333 38913 10367 38947
rect 12541 38913 12575 38947
rect 13461 38913 13495 38947
rect 15117 38913 15151 38947
rect 15209 38913 15243 38947
rect 15945 38913 15979 38947
rect 16681 38913 16715 38947
rect 20085 38913 20119 38947
rect 22109 38913 22143 38947
rect 8861 38845 8895 38879
rect 8953 38845 8987 38879
rect 12725 38845 12759 38879
rect 13578 38845 13612 38879
rect 13737 38845 13771 38879
rect 17969 38845 18003 38879
rect 18613 38845 18647 38879
rect 19809 38845 19843 38879
rect 22293 38845 22327 38879
rect 13185 38777 13219 38811
rect 1593 38709 1627 38743
rect 2421 38709 2455 38743
rect 3065 38709 3099 38743
rect 4169 38709 4203 38743
rect 5733 38709 5767 38743
rect 10517 38709 10551 38743
rect 17325 38709 17359 38743
rect 19257 38709 19291 38743
rect 20453 38709 20487 38743
rect 2329 38505 2363 38539
rect 2513 38505 2547 38539
rect 6975 38505 7009 38539
rect 8401 38505 8435 38539
rect 9689 38505 9723 38539
rect 14105 38505 14139 38539
rect 18245 38505 18279 38539
rect 19625 38505 19659 38539
rect 20085 38505 20119 38539
rect 1961 38437 1995 38471
rect 12357 38437 12391 38471
rect 4169 38369 4203 38403
rect 5733 38369 5767 38403
rect 6745 38369 6779 38403
rect 9229 38369 9263 38403
rect 13093 38369 13127 38403
rect 13461 38369 13495 38403
rect 15025 38369 15059 38403
rect 2973 38301 3007 38335
rect 3985 38301 4019 38335
rect 4261 38301 4295 38335
rect 4353 38301 4387 38335
rect 4537 38301 4571 38335
rect 5457 38301 5491 38335
rect 8217 38301 8251 38335
rect 8953 38301 8987 38335
rect 9137 38301 9171 38335
rect 9321 38301 9355 38335
rect 9505 38301 9539 38335
rect 10425 38301 10459 38335
rect 11069 38301 11103 38335
rect 12173 38301 12207 38335
rect 13369 38301 13403 38335
rect 14289 38301 14323 38335
rect 14473 38301 14507 38335
rect 14933 38301 14967 38335
rect 15117 38301 15151 38335
rect 17877 38301 17911 38335
rect 19257 38301 19291 38335
rect 20269 38301 20303 38335
rect 2329 38233 2363 38267
rect 12817 38233 12851 38267
rect 18061 38233 18095 38267
rect 19441 38233 19475 38267
rect 3157 38165 3191 38199
rect 3801 38165 3835 38199
rect 10609 38165 10643 38199
rect 11253 38165 11287 38199
rect 2329 37961 2363 37995
rect 7573 37961 7607 37995
rect 13369 37961 13403 37995
rect 14565 37961 14599 37995
rect 3464 37893 3498 37927
rect 11774 37893 11808 37927
rect 17877 37893 17911 37927
rect 1685 37825 1719 37859
rect 4169 37825 4203 37859
rect 4436 37825 4470 37859
rect 6561 37825 6595 37859
rect 6745 37825 6779 37859
rect 6929 37825 6963 37859
rect 7113 37825 7147 37859
rect 7757 37825 7791 37859
rect 8217 37825 8251 37859
rect 8484 37825 8518 37859
rect 10057 37825 10091 37859
rect 10241 37825 10275 37859
rect 10609 37825 10643 37859
rect 11529 37825 11563 37859
rect 13645 37825 13679 37859
rect 14105 37825 14139 37859
rect 14381 37825 14415 37859
rect 15025 37825 15059 37859
rect 17693 37825 17727 37859
rect 18061 37825 18095 37859
rect 18705 37825 18739 37859
rect 3709 37757 3743 37791
rect 6837 37757 6871 37791
rect 10333 37757 10367 37791
rect 10425 37757 10459 37791
rect 13369 37757 13403 37791
rect 15117 37757 15151 37791
rect 14197 37689 14231 37723
rect 1501 37621 1535 37655
rect 5549 37621 5583 37655
rect 6377 37621 6411 37655
rect 9597 37621 9631 37655
rect 10793 37621 10827 37655
rect 12909 37621 12943 37655
rect 13553 37621 13587 37655
rect 18521 37621 18555 37655
rect 2329 37417 2363 37451
rect 7481 37417 7515 37451
rect 8953 37417 8987 37451
rect 12725 37417 12759 37451
rect 13093 37417 13127 37451
rect 2513 37349 2547 37383
rect 5365 37281 5399 37315
rect 5641 37281 5675 37315
rect 9413 37281 9447 37315
rect 15761 37281 15795 37315
rect 16037 37281 16071 37315
rect 16154 37281 16188 37315
rect 16313 37281 16347 37315
rect 17969 37281 18003 37315
rect 1961 37213 1995 37247
rect 2973 37213 3007 37247
rect 3985 37213 4019 37247
rect 6101 37213 6135 37247
rect 6368 37213 6402 37247
rect 8401 37213 8435 37247
rect 9137 37213 9171 37247
rect 9321 37213 9355 37247
rect 9505 37213 9539 37247
rect 9689 37213 9723 37247
rect 10609 37213 10643 37247
rect 10876 37213 10910 37247
rect 13001 37213 13035 37247
rect 13093 37213 13127 37247
rect 14105 37213 14139 37247
rect 14289 37213 14323 37247
rect 14657 37213 14691 37247
rect 15117 37213 15151 37247
rect 15301 37213 15335 37247
rect 18061 37213 18095 37247
rect 18153 37213 18187 37247
rect 19441 37213 19475 37247
rect 30113 37213 30147 37247
rect 2329 37145 2363 37179
rect 14565 37145 14599 37179
rect 3157 37077 3191 37111
rect 3801 37077 3835 37111
rect 8217 37077 8251 37111
rect 11989 37077 12023 37111
rect 16957 37077 16991 37111
rect 18521 37077 18555 37111
rect 19257 37077 19291 37111
rect 29929 37077 29963 37111
rect 1593 36873 1627 36907
rect 2605 36873 2639 36907
rect 3617 36873 3651 36907
rect 5457 36873 5491 36907
rect 10885 36873 10919 36907
rect 11529 36873 11563 36907
rect 14933 36873 14967 36907
rect 17233 36873 17267 36907
rect 17601 36873 17635 36907
rect 18797 36873 18831 36907
rect 2421 36805 2455 36839
rect 4077 36805 4111 36839
rect 1409 36737 1443 36771
rect 2053 36737 2087 36771
rect 3433 36737 3467 36771
rect 4261 36737 4295 36771
rect 4629 36737 4663 36771
rect 4813 36737 4847 36771
rect 5641 36737 5675 36771
rect 7389 36737 7423 36771
rect 8033 36737 8067 36771
rect 9045 36737 9079 36771
rect 10149 36737 10183 36771
rect 10333 36737 10367 36771
rect 10517 36737 10551 36771
rect 10701 36737 10735 36771
rect 11713 36737 11747 36771
rect 12449 36737 12483 36771
rect 13185 36737 13219 36771
rect 13829 36737 13863 36771
rect 14105 36737 14139 36771
rect 14197 36737 14231 36771
rect 14841 36737 14875 36771
rect 15025 36737 15059 36771
rect 18613 36737 18647 36771
rect 19257 36737 19291 36771
rect 19524 36737 19558 36771
rect 22109 36737 22143 36771
rect 4445 36669 4479 36703
rect 4537 36669 4571 36703
rect 10425 36669 10459 36703
rect 13277 36669 13311 36703
rect 14381 36669 14415 36703
rect 16957 36669 16991 36703
rect 17141 36669 17175 36703
rect 22293 36669 22327 36703
rect 6929 36601 6963 36635
rect 2421 36533 2455 36567
rect 7205 36533 7239 36567
rect 7849 36533 7883 36567
rect 9229 36533 9263 36567
rect 12633 36533 12667 36567
rect 13921 36533 13955 36567
rect 20637 36533 20671 36567
rect 21925 36533 21959 36567
rect 3985 36329 4019 36363
rect 5273 36329 5307 36363
rect 7205 36329 7239 36363
rect 16957 36329 16991 36363
rect 9781 36261 9815 36295
rect 6009 36193 6043 36227
rect 10241 36193 10275 36227
rect 15301 36193 15335 36227
rect 15761 36193 15795 36227
rect 16037 36193 16071 36227
rect 16154 36193 16188 36227
rect 20269 36193 20303 36227
rect 1685 36125 1719 36159
rect 2421 36125 2455 36159
rect 3065 36125 3099 36159
rect 3801 36125 3835 36159
rect 4629 36125 4663 36159
rect 5089 36125 5123 36159
rect 5733 36125 5767 36159
rect 7481 36125 7515 36159
rect 8125 36125 8159 36159
rect 9137 36125 9171 36159
rect 9597 36125 9631 36159
rect 12812 36125 12846 36159
rect 13184 36125 13218 36159
rect 13277 36125 13311 36159
rect 15117 36125 15151 36159
rect 16313 36125 16347 36159
rect 17601 36125 17635 36159
rect 18429 36125 18463 36159
rect 20821 36125 20855 36159
rect 21097 36125 21131 36159
rect 10508 36057 10542 36091
rect 12909 36057 12943 36091
rect 13001 36057 13035 36091
rect 19993 36057 20027 36091
rect 20085 36057 20119 36091
rect 21281 36057 21315 36091
rect 1501 35989 1535 36023
rect 2237 35989 2271 36023
rect 2881 35989 2915 36023
rect 4445 35989 4479 36023
rect 7021 35989 7055 36023
rect 7941 35989 7975 36023
rect 8953 35989 8987 36023
rect 11621 35989 11655 36023
rect 12633 35989 12667 36023
rect 17785 35989 17819 36023
rect 18245 35989 18279 36023
rect 19625 35989 19659 36023
rect 20913 35989 20947 36023
rect 2237 35785 2271 35819
rect 5549 35785 5583 35819
rect 6837 35785 6871 35819
rect 7757 35785 7791 35819
rect 9229 35785 9263 35819
rect 10701 35785 10735 35819
rect 19533 35785 19567 35819
rect 20361 35785 20395 35819
rect 12909 35717 12943 35751
rect 1869 35649 1903 35683
rect 2881 35649 2915 35683
rect 3525 35649 3559 35683
rect 4905 35649 4939 35683
rect 5733 35649 5767 35683
rect 6377 35649 6411 35683
rect 7757 35649 7791 35683
rect 7849 35649 7883 35683
rect 8116 35649 8150 35683
rect 9965 35649 9999 35683
rect 10149 35649 10183 35683
rect 10241 35649 10275 35683
rect 10517 35649 10551 35683
rect 11805 35649 11839 35683
rect 12633 35649 12667 35683
rect 12781 35649 12815 35683
rect 13001 35649 13035 35683
rect 13098 35649 13132 35683
rect 17049 35649 17083 35683
rect 18153 35649 18187 35683
rect 18420 35649 18454 35683
rect 20269 35649 20303 35683
rect 20453 35649 20487 35683
rect 10333 35581 10367 35615
rect 16773 35581 16807 35615
rect 16957 35581 16991 35615
rect 3065 35513 3099 35547
rect 2237 35445 2271 35479
rect 2421 35445 2455 35479
rect 3709 35445 3743 35479
rect 4721 35445 4755 35479
rect 6469 35445 6503 35479
rect 11897 35445 11931 35479
rect 13277 35445 13311 35479
rect 17417 35445 17451 35479
rect 2237 35241 2271 35275
rect 2421 35241 2455 35275
rect 5825 35241 5859 35275
rect 8401 35241 8435 35275
rect 10609 35241 10643 35275
rect 16589 35241 16623 35275
rect 20453 35241 20487 35275
rect 1869 35173 1903 35207
rect 3801 35105 3835 35139
rect 7941 35105 7975 35139
rect 9597 35105 9631 35139
rect 15393 35105 15427 35139
rect 15786 35105 15820 35139
rect 17141 35105 17175 35139
rect 17325 35105 17359 35139
rect 2881 35037 2915 35071
rect 6009 35037 6043 35071
rect 6561 35037 6595 35071
rect 6653 35037 6687 35071
rect 7665 35037 7699 35071
rect 7849 35031 7883 35065
rect 8033 35037 8067 35071
rect 8200 35037 8234 35071
rect 9321 35037 9355 35071
rect 10793 35037 10827 35071
rect 11713 35037 11747 35071
rect 14749 35037 14783 35071
rect 14933 35037 14967 35071
rect 15669 35037 15703 35071
rect 15945 35037 15979 35071
rect 18245 35037 18279 35071
rect 20269 35037 20303 35071
rect 20545 35037 20579 35071
rect 21005 35037 21039 35071
rect 21189 35037 21223 35071
rect 22109 35037 22143 35071
rect 22293 35037 22327 35071
rect 30113 35037 30147 35071
rect 2237 34969 2271 35003
rect 4068 34969 4102 35003
rect 11980 34969 12014 35003
rect 18429 34969 18463 35003
rect 21097 34969 21131 35003
rect 3065 34901 3099 34935
rect 5181 34901 5215 34935
rect 13093 34901 13127 34935
rect 17417 34901 17451 34935
rect 17785 34901 17819 34935
rect 18613 34901 18647 34935
rect 20085 34901 20119 34935
rect 21925 34901 21959 34935
rect 29929 34901 29963 34935
rect 2421 34697 2455 34731
rect 3985 34697 4019 34731
rect 4445 34697 4479 34731
rect 6377 34697 6411 34731
rect 7021 34697 7055 34731
rect 8769 34697 8803 34731
rect 13737 34697 13771 34731
rect 16129 34697 16163 34731
rect 17049 34697 17083 34731
rect 18889 34697 18923 34731
rect 19533 34697 19567 34731
rect 20545 34697 20579 34731
rect 20729 34697 20763 34731
rect 20821 34697 20855 34731
rect 2237 34629 2271 34663
rect 11621 34629 11655 34663
rect 12624 34629 12658 34663
rect 20637 34629 20671 34663
rect 1869 34561 1903 34595
rect 3249 34561 3283 34595
rect 3433 34561 3467 34595
rect 3525 34561 3559 34595
rect 3801 34561 3835 34595
rect 5569 34561 5603 34595
rect 5825 34561 5859 34595
rect 6561 34561 6595 34595
rect 7205 34561 7239 34595
rect 7849 34561 7883 34595
rect 8677 34561 8711 34595
rect 11529 34561 11563 34595
rect 14473 34561 14507 34595
rect 15326 34561 15360 34595
rect 16865 34561 16899 34595
rect 17776 34561 17810 34595
rect 19530 34561 19564 34595
rect 21005 34561 21039 34595
rect 3617 34493 3651 34527
rect 9873 34493 9907 34527
rect 10149 34493 10183 34527
rect 12357 34493 12391 34527
rect 14289 34493 14323 34527
rect 15209 34493 15243 34527
rect 15485 34493 15519 34527
rect 17509 34493 17543 34527
rect 19993 34493 20027 34527
rect 14933 34425 14967 34459
rect 2237 34357 2271 34391
rect 7665 34357 7699 34391
rect 19349 34357 19383 34391
rect 19901 34357 19935 34391
rect 2237 34153 2271 34187
rect 2421 34153 2455 34187
rect 5641 34153 5675 34187
rect 7205 34153 7239 34187
rect 18061 34153 18095 34187
rect 18613 34153 18647 34187
rect 1869 34085 1903 34119
rect 15485 34085 15519 34119
rect 20729 34085 20763 34119
rect 6101 34017 6135 34051
rect 8033 34017 8067 34051
rect 12081 34017 12115 34051
rect 19993 34017 20027 34051
rect 20085 34017 20119 34051
rect 3157 33949 3191 33983
rect 3801 33949 3835 33983
rect 5825 33949 5859 33983
rect 6009 33949 6043 33983
rect 6193 33949 6227 33983
rect 6377 33949 6411 33983
rect 7021 33949 7055 33983
rect 7849 33949 7883 33983
rect 8125 33949 8159 33983
rect 8217 33949 8251 33983
rect 8401 33949 8435 33983
rect 9321 33949 9355 33983
rect 11345 33949 11379 33983
rect 11805 33949 11839 33983
rect 14105 33949 14139 33983
rect 17877 33949 17911 33983
rect 18061 33949 18095 33983
rect 18705 33949 18739 33983
rect 21281 33949 21315 33983
rect 21741 33949 21775 33983
rect 22385 33949 22419 33983
rect 2237 33881 2271 33915
rect 4046 33881 4080 33915
rect 11100 33881 11134 33915
rect 14372 33881 14406 33915
rect 20913 33881 20947 33915
rect 21833 33881 21867 33915
rect 2973 33813 3007 33847
rect 5181 33813 5215 33847
rect 7665 33813 7699 33847
rect 9505 33813 9539 33847
rect 9965 33813 9999 33847
rect 19533 33813 19567 33847
rect 19901 33813 19935 33847
rect 21005 33813 21039 33847
rect 21097 33813 21131 33847
rect 22569 33813 22603 33847
rect 2605 33609 2639 33643
rect 5549 33609 5583 33643
rect 10977 33609 11011 33643
rect 12081 33609 12115 33643
rect 15669 33609 15703 33643
rect 18337 33609 18371 33643
rect 18889 33609 18923 33643
rect 19073 33609 19107 33643
rect 21281 33609 21315 33643
rect 20913 33541 20947 33575
rect 1685 33473 1719 33507
rect 2421 33473 2455 33507
rect 3249 33473 3283 33507
rect 3801 33473 3835 33507
rect 3985 33473 4019 33507
rect 4353 33473 4387 33507
rect 4537 33473 4571 33507
rect 5733 33473 5767 33507
rect 6469 33473 6503 33507
rect 7297 33473 7331 33507
rect 8125 33473 8159 33507
rect 8309 33473 8343 33507
rect 8493 33473 8527 33507
rect 8677 33473 8711 33507
rect 9781 33473 9815 33507
rect 9965 33473 9999 33507
rect 10149 33473 10183 33507
rect 10333 33473 10367 33507
rect 10793 33473 10827 33507
rect 11529 33473 11563 33507
rect 11805 33473 11839 33507
rect 11897 33473 11931 33507
rect 12081 33473 12115 33507
rect 14298 33473 14332 33507
rect 14565 33473 14599 33507
rect 15485 33473 15519 33507
rect 16681 33473 16715 33507
rect 18245 33473 18279 33507
rect 18429 33473 18463 33507
rect 19070 33473 19104 33507
rect 19441 33473 19475 33507
rect 22385 33473 22419 33507
rect 30113 33473 30147 33507
rect 4169 33405 4203 33439
rect 4261 33405 4295 33439
rect 8401 33405 8435 33439
rect 10057 33405 10091 33439
rect 19533 33405 19567 33439
rect 20637 33405 20671 33439
rect 20821 33405 20855 33439
rect 3065 33337 3099 33371
rect 1501 33269 1535 33303
rect 6653 33269 6687 33303
rect 7113 33269 7147 33303
rect 7941 33269 7975 33303
rect 9597 33269 9631 33303
rect 11621 33269 11655 33303
rect 13185 33269 13219 33303
rect 16865 33269 16899 33303
rect 22569 33269 22603 33303
rect 29929 33269 29963 33303
rect 4721 33065 4755 33099
rect 8401 33065 8435 33099
rect 10517 33065 10551 33099
rect 16497 33065 16531 33099
rect 20361 33065 20395 33099
rect 20729 33065 20763 33099
rect 5733 32997 5767 33031
rect 10057 32929 10091 32963
rect 10149 32929 10183 32963
rect 15117 32929 15151 32963
rect 17049 32929 17083 32963
rect 20453 32929 20487 32963
rect 1409 32861 1443 32895
rect 2329 32861 2363 32895
rect 3157 32861 3191 32895
rect 4077 32861 4111 32895
rect 4905 32861 4939 32895
rect 6377 32861 6411 32895
rect 7021 32861 7055 32895
rect 7288 32861 7322 32895
rect 9045 32861 9079 32895
rect 9781 32861 9815 32895
rect 9965 32861 9999 32895
rect 10333 32861 10367 32895
rect 11161 32861 11195 32895
rect 11621 32861 11655 32895
rect 19717 32861 19751 32895
rect 20361 32861 20395 32895
rect 22293 32861 22327 32895
rect 22477 32861 22511 32895
rect 5549 32793 5583 32827
rect 11888 32793 11922 32827
rect 15384 32793 15418 32827
rect 17316 32793 17350 32827
rect 1593 32725 1627 32759
rect 2145 32725 2179 32759
rect 2973 32725 3007 32759
rect 4261 32725 4295 32759
rect 6561 32725 6595 32759
rect 9229 32725 9263 32759
rect 10977 32725 11011 32759
rect 13001 32725 13035 32759
rect 18429 32725 18463 32759
rect 19809 32725 19843 32759
rect 22109 32725 22143 32759
rect 2237 32521 2271 32555
rect 4261 32521 4295 32555
rect 6929 32521 6963 32555
rect 8769 32521 8803 32555
rect 9597 32521 9631 32555
rect 15761 32521 15795 32555
rect 17969 32521 18003 32555
rect 18613 32521 18647 32555
rect 20561 32521 20595 32555
rect 7656 32453 7690 32487
rect 10710 32453 10744 32487
rect 15485 32453 15519 32487
rect 20361 32453 20395 32487
rect 1869 32385 1903 32419
rect 3148 32385 3182 32419
rect 5365 32385 5399 32419
rect 6745 32385 6779 32419
rect 7389 32385 7423 32419
rect 10977 32385 11011 32419
rect 11888 32385 11922 32419
rect 15117 32385 15151 32419
rect 15265 32385 15299 32419
rect 15393 32385 15427 32419
rect 15623 32385 15657 32419
rect 17233 32385 17267 32419
rect 17417 32385 17451 32419
rect 17509 32385 17543 32419
rect 17785 32385 17819 32419
rect 18521 32385 18555 32419
rect 19625 32385 19659 32419
rect 19809 32385 19843 32419
rect 2881 32317 2915 32351
rect 5641 32317 5675 32351
rect 11621 32317 11655 32351
rect 17601 32317 17635 32351
rect 18705 32317 18739 32351
rect 2237 32181 2271 32215
rect 2421 32181 2455 32215
rect 13001 32181 13035 32215
rect 19073 32181 19107 32215
rect 19625 32181 19659 32215
rect 20545 32181 20579 32215
rect 20729 32181 20763 32215
rect 2789 31977 2823 32011
rect 3801 31977 3835 32011
rect 9781 31977 9815 32011
rect 16037 31977 16071 32011
rect 17233 31977 17267 32011
rect 19257 31977 19291 32011
rect 19625 31977 19659 32011
rect 19809 31977 19843 32011
rect 7113 31909 7147 31943
rect 8401 31909 8435 31943
rect 10609 31909 10643 31943
rect 19717 31909 19751 31943
rect 20637 31909 20671 31943
rect 4169 31841 4203 31875
rect 5549 31841 5583 31875
rect 9413 31841 9447 31875
rect 11253 31841 11287 31875
rect 14105 31841 14139 31875
rect 22017 31841 22051 31875
rect 1685 31773 1719 31807
rect 2605 31773 2639 31807
rect 3985 31773 4019 31807
rect 4261 31773 4295 31807
rect 4353 31773 4387 31807
rect 4537 31773 4571 31807
rect 5825 31773 5859 31807
rect 6469 31773 6503 31807
rect 6929 31773 6963 31807
rect 7573 31773 7607 31807
rect 8217 31773 8251 31807
rect 9873 31773 9907 31807
rect 10425 31773 10459 31807
rect 11529 31773 11563 31807
rect 15945 31773 15979 31807
rect 17417 31773 17451 31807
rect 18521 31773 18555 31807
rect 18613 31773 18647 31807
rect 19533 31773 19567 31807
rect 19993 31773 20027 31807
rect 20453 31773 20487 31807
rect 21741 31773 21775 31807
rect 14350 31705 14384 31739
rect 17601 31705 17635 31739
rect 1501 31637 1535 31671
rect 6377 31637 6411 31671
rect 7757 31637 7791 31671
rect 15485 31637 15519 31671
rect 1409 31433 1443 31467
rect 3065 31433 3099 31467
rect 10793 31433 10827 31467
rect 12265 31433 12299 31467
rect 12909 31433 12943 31467
rect 13645 31433 13679 31467
rect 15393 31433 15427 31467
rect 17877 31433 17911 31467
rect 19441 31433 19475 31467
rect 2421 31365 2455 31399
rect 1593 31297 1627 31331
rect 3249 31297 3283 31331
rect 3893 31297 3927 31331
rect 4077 31297 4111 31331
rect 4261 31297 4295 31331
rect 4445 31297 4479 31331
rect 7490 31297 7524 31331
rect 7757 31297 7791 31331
rect 8309 31297 8343 31331
rect 9505 31297 9539 31331
rect 10885 31297 10919 31331
rect 11529 31297 11563 31331
rect 11713 31297 11747 31331
rect 12081 31297 12115 31331
rect 2053 31229 2087 31263
rect 4169 31229 4203 31263
rect 5457 31229 5491 31263
rect 5733 31229 5767 31263
rect 11805 31229 11839 31263
rect 11897 31229 11931 31263
rect 13369 31365 13403 31399
rect 14381 31365 14415 31399
rect 17785 31365 17819 31399
rect 13001 31297 13035 31331
rect 13094 31297 13128 31331
rect 13277 31297 13311 31331
rect 13507 31297 13541 31331
rect 14105 31297 14139 31331
rect 14253 31297 14287 31331
rect 14473 31297 14507 31331
rect 14570 31297 14604 31331
rect 15761 31297 15795 31331
rect 15853 31297 15887 31331
rect 16681 31297 16715 31331
rect 18705 31297 18739 31331
rect 18889 31297 18923 31331
rect 18981 31297 19015 31331
rect 19257 31297 19291 31331
rect 19901 31297 19935 31331
rect 20729 31297 20763 31331
rect 21115 31297 21149 31331
rect 21281 31297 21315 31331
rect 29837 31297 29871 31331
rect 16037 31229 16071 31263
rect 17601 31229 17635 31263
rect 19073 31229 19107 31263
rect 20913 31229 20947 31263
rect 21005 31229 21039 31263
rect 21833 31229 21867 31263
rect 22109 31229 22143 31263
rect 30113 31229 30147 31263
rect 2605 31161 2639 31195
rect 8769 31161 8803 31195
rect 12909 31161 12943 31195
rect 20545 31161 20579 31195
rect 2421 31093 2455 31127
rect 3709 31093 3743 31127
rect 6377 31093 6411 31127
rect 8585 31093 8619 31127
rect 9781 31093 9815 31127
rect 9965 31093 9999 31127
rect 14749 31093 14783 31127
rect 16773 31093 16807 31127
rect 18245 31093 18279 31127
rect 19993 31093 20027 31127
rect 2421 30889 2455 30923
rect 3065 30889 3099 30923
rect 5917 30889 5951 30923
rect 9321 30889 9355 30923
rect 9873 30889 9907 30923
rect 15393 30889 15427 30923
rect 18521 30889 18555 30923
rect 19993 30889 20027 30923
rect 20177 30889 20211 30923
rect 1593 30821 1627 30855
rect 2053 30821 2087 30855
rect 2605 30821 2639 30855
rect 7113 30821 7147 30855
rect 11989 30821 12023 30855
rect 14105 30821 14139 30855
rect 17417 30821 17451 30855
rect 18613 30821 18647 30855
rect 20913 30821 20947 30855
rect 5089 30753 5123 30787
rect 5181 30753 5215 30787
rect 6377 30753 6411 30787
rect 7573 30753 7607 30787
rect 11529 30753 11563 30787
rect 18429 30753 18463 30787
rect 21189 30753 21223 30787
rect 23305 30753 23339 30787
rect 1409 30685 1443 30719
rect 3249 30685 3283 30719
rect 3801 30685 3835 30719
rect 4905 30685 4939 30719
rect 5273 30685 5307 30719
rect 5457 30685 5491 30719
rect 6101 30685 6135 30719
rect 6285 30685 6319 30719
rect 6469 30685 6503 30719
rect 6653 30685 6687 30719
rect 7297 30685 7331 30719
rect 7481 30685 7515 30719
rect 7665 30685 7699 30719
rect 7849 30685 7883 30719
rect 9413 30685 9447 30719
rect 10057 30685 10091 30719
rect 10701 30685 10735 30719
rect 11253 30685 11287 30719
rect 11437 30685 11471 30719
rect 11621 30685 11655 30719
rect 11805 30685 11839 30719
rect 13001 30685 13035 30719
rect 13277 30685 13311 30719
rect 14243 30685 14277 30719
rect 14473 30685 14507 30719
rect 14601 30685 14635 30719
rect 14749 30685 14783 30719
rect 15301 30685 15335 30719
rect 16037 30685 16071 30719
rect 17141 30685 17175 30719
rect 17233 30685 17267 30719
rect 17509 30685 17543 30719
rect 18705 30685 18739 30719
rect 21281 30685 21315 30719
rect 21649 30685 21683 30719
rect 21833 30685 21867 30719
rect 22017 30685 22051 30719
rect 23213 30685 23247 30719
rect 14381 30617 14415 30651
rect 16221 30617 16255 30651
rect 19809 30617 19843 30651
rect 20009 30617 20043 30651
rect 22477 30617 22511 30651
rect 22661 30617 22695 30651
rect 2421 30549 2455 30583
rect 3985 30549 4019 30583
rect 4721 30549 4755 30583
rect 8953 30549 8987 30583
rect 10517 30549 10551 30583
rect 16957 30549 16991 30583
rect 2329 30345 2363 30379
rect 4629 30345 4663 30379
rect 7757 30345 7791 30379
rect 16681 30345 16715 30379
rect 17877 30345 17911 30379
rect 3516 30277 3550 30311
rect 6644 30277 6678 30311
rect 18337 30277 18371 30311
rect 21833 30277 21867 30311
rect 1961 30209 1995 30243
rect 5641 30209 5675 30243
rect 8677 30209 8711 30243
rect 9597 30209 9631 30243
rect 9864 30209 9898 30243
rect 11805 30209 11839 30243
rect 12357 30209 12391 30243
rect 12633 30209 12667 30243
rect 14197 30209 14231 30243
rect 14464 30209 14498 30243
rect 17049 30209 17083 30243
rect 18245 30209 18279 30243
rect 19165 30209 19199 30243
rect 19993 30209 20027 30243
rect 20269 30209 20303 30243
rect 22017 30209 22051 30243
rect 22201 30209 22235 30243
rect 22653 30209 22687 30243
rect 3249 30141 3283 30175
rect 6377 30141 6411 30175
rect 17141 30141 17175 30175
rect 17233 30141 17267 30175
rect 18429 30141 18463 30175
rect 10977 30073 11011 30107
rect 15577 30073 15611 30107
rect 19349 30073 19383 30107
rect 2329 30005 2363 30039
rect 2513 30005 2547 30039
rect 5825 30005 5859 30039
rect 8217 30005 8251 30039
rect 8585 30005 8619 30039
rect 11713 30005 11747 30039
rect 22753 30005 22787 30039
rect 2421 29801 2455 29835
rect 2605 29801 2639 29835
rect 6193 29801 6227 29835
rect 7389 29801 7423 29835
rect 10701 29801 10735 29835
rect 11069 29801 11103 29835
rect 17509 29801 17543 29835
rect 2053 29733 2087 29767
rect 21373 29733 21407 29767
rect 10609 29665 10643 29699
rect 14105 29665 14139 29699
rect 16957 29665 16991 29699
rect 22109 29665 22143 29699
rect 1409 29597 1443 29631
rect 3065 29597 3099 29631
rect 4169 29597 4203 29631
rect 4436 29597 4470 29631
rect 6009 29597 6043 29631
rect 8217 29597 8251 29631
rect 9689 29597 9723 29631
rect 10885 29597 10919 29631
rect 12633 29597 12667 29631
rect 12909 29597 12943 29631
rect 16313 29597 16347 29631
rect 17969 29597 18003 29631
rect 19993 29597 20027 29631
rect 20361 29597 20395 29631
rect 21189 29597 21223 29631
rect 21833 29597 21867 29631
rect 22201 29597 22235 29631
rect 2421 29529 2455 29563
rect 7297 29529 7331 29563
rect 12081 29529 12115 29563
rect 14350 29529 14384 29563
rect 16221 29529 16255 29563
rect 19809 29529 19843 29563
rect 20821 29529 20855 29563
rect 22318 29529 22352 29563
rect 1593 29461 1627 29495
rect 3249 29461 3283 29495
rect 5549 29461 5583 29495
rect 8033 29461 8067 29495
rect 9505 29461 9539 29495
rect 11989 29461 12023 29495
rect 15485 29461 15519 29495
rect 17049 29461 17083 29495
rect 17141 29461 17175 29495
rect 18153 29461 18187 29495
rect 20085 29461 20119 29495
rect 20177 29461 20211 29495
rect 21005 29461 21039 29495
rect 21097 29461 21131 29495
rect 22477 29461 22511 29495
rect 2329 29257 2363 29291
rect 3433 29257 3467 29291
rect 5273 29257 5307 29291
rect 8769 29257 8803 29291
rect 9137 29257 9171 29291
rect 11897 29257 11931 29291
rect 13185 29257 13219 29291
rect 14657 29257 14691 29291
rect 21005 29257 21039 29291
rect 22385 29257 22419 29291
rect 12633 29189 12667 29223
rect 13553 29189 13587 29223
rect 16037 29189 16071 29223
rect 23090 29189 23124 29223
rect 1685 29121 1719 29155
rect 2145 29121 2179 29155
rect 3617 29121 3651 29155
rect 4261 29121 4295 29155
rect 5089 29121 5123 29155
rect 7021 29121 7055 29155
rect 8033 29121 8067 29155
rect 10149 29121 10183 29155
rect 11989 29121 12023 29155
rect 13323 29121 13357 29155
rect 13461 29121 13495 29155
rect 13681 29121 13715 29155
rect 13829 29121 13863 29155
rect 14749 29121 14783 29155
rect 15945 29121 15979 29155
rect 16681 29121 16715 29155
rect 16865 29121 16899 29155
rect 17049 29121 17083 29155
rect 17233 29121 17267 29155
rect 18061 29121 18095 29155
rect 18245 29121 18279 29155
rect 18337 29121 18371 29155
rect 20729 29121 20763 29155
rect 22201 29121 22235 29155
rect 22845 29121 22879 29155
rect 29837 29121 29871 29155
rect 7113 29053 7147 29087
rect 7205 29053 7239 29087
rect 9229 29053 9263 29087
rect 9321 29053 9355 29087
rect 16957 29053 16991 29087
rect 17417 29053 17451 29087
rect 17969 29053 18003 29087
rect 20545 29053 20579 29087
rect 20637 29053 20671 29087
rect 20821 29053 20855 29087
rect 1501 28985 1535 29019
rect 7849 28985 7883 29019
rect 9965 28985 9999 29019
rect 12449 28985 12483 29019
rect 17877 28985 17911 29019
rect 24225 28985 24259 29019
rect 30021 28985 30055 29019
rect 4077 28917 4111 28951
rect 6653 28917 6687 28951
rect 3985 28713 4019 28747
rect 5181 28713 5215 28747
rect 5825 28713 5859 28747
rect 11345 28713 11379 28747
rect 16497 28713 16531 28747
rect 22661 28713 22695 28747
rect 12081 28645 12115 28679
rect 14749 28645 14783 28679
rect 2697 28577 2731 28611
rect 7021 28577 7055 28611
rect 8125 28577 8159 28611
rect 9965 28577 9999 28611
rect 16957 28577 16991 28611
rect 17141 28577 17175 28611
rect 18061 28577 18095 28611
rect 18245 28577 18279 28611
rect 21281 28577 21315 28611
rect 1685 28509 1719 28543
rect 2605 28509 2639 28543
rect 2789 28509 2823 28543
rect 3617 28509 3651 28543
rect 3801 28509 3835 28543
rect 4997 28509 5031 28543
rect 5641 28509 5675 28543
rect 6745 28509 6779 28543
rect 7941 28509 7975 28543
rect 9137 28509 9171 28543
rect 12725 28509 12759 28543
rect 12818 28509 12852 28543
rect 13001 28509 13035 28543
rect 13190 28509 13224 28543
rect 15393 28509 15427 28543
rect 19901 28509 19935 28543
rect 20453 28509 20487 28543
rect 10232 28441 10266 28475
rect 11897 28441 11931 28475
rect 13093 28441 13127 28475
rect 14565 28441 14599 28475
rect 15209 28441 15243 28475
rect 15577 28441 15611 28475
rect 21526 28441 21560 28475
rect 1501 28373 1535 28407
rect 3617 28373 3651 28407
rect 6377 28373 6411 28407
rect 6837 28373 6871 28407
rect 7573 28373 7607 28407
rect 8033 28373 8067 28407
rect 9045 28373 9079 28407
rect 13369 28373 13403 28407
rect 16865 28373 16899 28407
rect 18337 28373 18371 28407
rect 18705 28373 18739 28407
rect 19901 28373 19935 28407
rect 20637 28373 20671 28407
rect 4721 28169 4755 28203
rect 6837 28169 6871 28203
rect 7481 28169 7515 28203
rect 9229 28169 9263 28203
rect 10333 28169 10367 28203
rect 14473 28169 14507 28203
rect 16129 28169 16163 28203
rect 17049 28169 17083 28203
rect 20545 28169 20579 28203
rect 30021 28169 30055 28203
rect 3893 28101 3927 28135
rect 4077 28101 4111 28135
rect 5457 28101 5491 28135
rect 10885 28101 10919 28135
rect 12357 28101 12391 28135
rect 17509 28101 17543 28135
rect 20637 28101 20671 28135
rect 22017 28101 22051 28135
rect 1685 28033 1719 28067
rect 2145 28033 2179 28067
rect 2329 28033 2363 28067
rect 3065 28033 3099 28067
rect 4629 28033 4663 28067
rect 4813 28033 4847 28067
rect 7021 28033 7055 28067
rect 7665 28033 7699 28067
rect 7757 28033 7791 28067
rect 8033 28033 8067 28067
rect 8493 28033 8527 28067
rect 8677 28033 8711 28067
rect 9045 28033 9079 28067
rect 9689 28033 9723 28067
rect 9782 28033 9816 28067
rect 9965 28033 9999 28067
rect 10057 28033 10091 28067
rect 10195 28033 10229 28067
rect 10977 28033 11011 28067
rect 11529 28033 11563 28067
rect 13093 28033 13127 28067
rect 13360 28033 13394 28067
rect 14933 28033 14967 28067
rect 15761 28033 15795 28067
rect 15945 28033 15979 28067
rect 17417 28033 17451 28067
rect 18613 28033 18647 28067
rect 18705 28033 18739 28067
rect 18981 28033 19015 28067
rect 20361 28033 20395 28067
rect 20453 28033 20487 28067
rect 20729 28033 20763 28067
rect 20821 28033 20855 28067
rect 21833 28033 21867 28067
rect 22201 28033 22235 28067
rect 29837 28033 29871 28067
rect 2237 27965 2271 27999
rect 8769 27965 8803 27999
rect 8861 27965 8895 27999
rect 17601 27965 17635 27999
rect 5641 27897 5675 27931
rect 12173 27897 12207 27931
rect 1501 27829 1535 27863
rect 2881 27829 2915 27863
rect 7941 27829 7975 27863
rect 11621 27829 11655 27863
rect 15025 27829 15059 27863
rect 18429 27829 18463 27863
rect 18889 27829 18923 27863
rect 5825 27625 5859 27659
rect 7297 27625 7331 27659
rect 7481 27625 7515 27659
rect 16129 27625 16163 27659
rect 19257 27625 19291 27659
rect 21097 27625 21131 27659
rect 6561 27557 6595 27591
rect 8309 27557 8343 27591
rect 9781 27557 9815 27591
rect 10793 27557 10827 27591
rect 14473 27557 14507 27591
rect 21649 27557 21683 27591
rect 10701 27489 10735 27523
rect 14841 27489 14875 27523
rect 15393 27489 15427 27523
rect 15577 27489 15611 27523
rect 16681 27489 16715 27523
rect 18245 27489 18279 27523
rect 19809 27489 19843 27523
rect 20821 27489 20855 27523
rect 2605 27421 2639 27455
rect 2789 27421 2823 27455
rect 4445 27421 4479 27455
rect 7757 27421 7791 27455
rect 8401 27421 8435 27455
rect 9137 27421 9171 27455
rect 9285 27421 9319 27455
rect 9643 27421 9677 27455
rect 10885 27421 10919 27455
rect 10977 27421 11011 27455
rect 11437 27421 11471 27455
rect 14381 27421 14415 27455
rect 14657 27421 14691 27455
rect 15301 27421 15335 27455
rect 16497 27421 16531 27455
rect 17325 27421 17359 27455
rect 17969 27421 18003 27455
rect 18153 27421 18187 27455
rect 18337 27421 18371 27455
rect 18521 27421 18555 27455
rect 20453 27421 20487 27455
rect 20637 27421 20671 27455
rect 20729 27421 20763 27455
rect 20913 27421 20947 27455
rect 21557 27421 21591 27455
rect 29837 27421 29871 27455
rect 4712 27353 4746 27387
rect 6745 27353 6779 27387
rect 9413 27353 9447 27387
rect 9505 27353 9539 27387
rect 11682 27353 11716 27387
rect 19717 27353 19751 27387
rect 2697 27285 2731 27319
rect 12817 27285 12851 27319
rect 15577 27285 15611 27319
rect 16589 27285 16623 27319
rect 17417 27285 17451 27319
rect 18705 27285 18739 27319
rect 19625 27285 19659 27319
rect 30021 27285 30055 27319
rect 5825 27081 5859 27115
rect 10885 27081 10919 27115
rect 16681 27081 16715 27115
rect 20545 27081 20579 27115
rect 8493 27013 8527 27047
rect 8677 27013 8711 27047
rect 15945 27013 15979 27047
rect 22017 27013 22051 27047
rect 1685 26945 1719 26979
rect 3341 26945 3375 26979
rect 3608 26945 3642 26979
rect 5365 26945 5399 26979
rect 5641 26945 5675 26979
rect 6653 26945 6687 26979
rect 7481 26945 7515 26979
rect 7849 26945 7883 26979
rect 8033 26945 8067 26979
rect 9505 26945 9539 26979
rect 9772 26945 9806 26979
rect 11529 26945 11563 26979
rect 12797 26945 12831 26979
rect 14749 26945 14783 26979
rect 15025 26945 15059 26979
rect 15117 26945 15151 26979
rect 15301 26945 15335 26979
rect 15761 26945 15795 26979
rect 16129 26945 16163 26979
rect 16865 26945 16899 26979
rect 17509 26945 17543 26979
rect 17969 26945 18003 26979
rect 18153 26945 18187 26979
rect 18245 26945 18279 26979
rect 18429 26945 18463 26979
rect 18613 26945 18647 26979
rect 19441 26945 19475 26979
rect 20177 26945 20211 26979
rect 20361 26945 20395 26979
rect 22201 26945 22235 26979
rect 5457 26877 5491 26911
rect 7665 26877 7699 26911
rect 7757 26877 7791 26911
rect 12541 26877 12575 26911
rect 20085 26877 20119 26911
rect 1501 26809 1535 26843
rect 5549 26809 5583 26843
rect 6745 26809 6779 26843
rect 11621 26809 11655 26843
rect 14841 26809 14875 26843
rect 18337 26809 18371 26843
rect 4721 26741 4755 26775
rect 7297 26741 7331 26775
rect 13921 26741 13955 26775
rect 17417 26741 17451 26775
rect 19533 26741 19567 26775
rect 21833 26741 21867 26775
rect 4905 26537 4939 26571
rect 9873 26537 9907 26571
rect 10425 26537 10459 26571
rect 14289 26537 14323 26571
rect 14657 26537 14691 26571
rect 15209 26537 15243 26571
rect 17509 26537 17543 26571
rect 17969 26537 18003 26571
rect 20821 26537 20855 26571
rect 6009 26469 6043 26503
rect 6101 26469 6135 26503
rect 7021 26469 7055 26503
rect 11161 26469 11195 26503
rect 12633 26469 12667 26503
rect 20637 26469 20671 26503
rect 23029 26469 23063 26503
rect 7481 26401 7515 26435
rect 7573 26401 7607 26435
rect 18521 26401 18555 26435
rect 21649 26401 21683 26435
rect 21925 26401 21959 26435
rect 1685 26333 1719 26367
rect 2697 26333 2731 26367
rect 2881 26333 2915 26367
rect 4261 26333 4295 26367
rect 4354 26333 4388 26367
rect 4629 26333 4663 26367
rect 4767 26333 4801 26367
rect 5917 26333 5951 26367
rect 6193 26333 6227 26367
rect 7389 26333 7423 26367
rect 8309 26333 8343 26367
rect 8401 26333 8435 26367
rect 9229 26333 9263 26367
rect 9322 26333 9356 26367
rect 9505 26333 9539 26367
rect 9735 26333 9769 26367
rect 10517 26333 10551 26367
rect 11253 26333 11287 26367
rect 11897 26333 11931 26367
rect 12081 26333 12115 26367
rect 12173 26333 12207 26367
rect 12265 26333 12299 26367
rect 12449 26333 12483 26367
rect 13277 26333 13311 26367
rect 14289 26333 14323 26367
rect 14473 26333 14507 26367
rect 15117 26333 15151 26367
rect 15761 26333 15795 26367
rect 15945 26333 15979 26367
rect 19257 26333 19291 26367
rect 20913 26333 20947 26367
rect 21005 26333 21039 26367
rect 23121 26333 23155 26367
rect 4537 26265 4571 26299
rect 6377 26265 6411 26299
rect 9597 26265 9631 26299
rect 13093 26265 13127 26299
rect 15853 26265 15887 26299
rect 17141 26265 17175 26299
rect 17325 26265 17359 26299
rect 18429 26265 18463 26299
rect 19349 26265 19383 26299
rect 1501 26197 1535 26231
rect 2789 26197 2823 26231
rect 18337 26197 18371 26231
rect 2789 25993 2823 26027
rect 3801 25993 3835 26027
rect 7757 25993 7791 26027
rect 8953 25993 8987 26027
rect 9321 25993 9355 26027
rect 9413 25993 9447 26027
rect 11529 25993 11563 26027
rect 14933 25993 14967 26027
rect 16681 25993 16715 26027
rect 17141 25993 17175 26027
rect 18337 25993 18371 26027
rect 4169 25925 4203 25959
rect 5733 25925 5767 25959
rect 10241 25925 10275 25959
rect 15761 25925 15795 25959
rect 15945 25925 15979 25959
rect 18705 25925 18739 25959
rect 1685 25857 1719 25891
rect 2697 25857 2731 25891
rect 2881 25857 2915 25891
rect 3980 25857 4014 25891
rect 4077 25857 4111 25891
rect 4297 25857 4331 25891
rect 4445 25857 4479 25891
rect 4905 25857 4939 25891
rect 6377 25857 6411 25891
rect 6929 25857 6963 25891
rect 7941 25857 7975 25891
rect 8033 25857 8067 25891
rect 8309 25857 8343 25891
rect 10333 25857 10367 25891
rect 10977 25857 11011 25891
rect 11713 25857 11747 25891
rect 11989 25857 12023 25891
rect 12081 25857 12115 25891
rect 12265 25857 12299 25891
rect 13930 25857 13964 25891
rect 14841 25857 14875 25891
rect 17049 25857 17083 25891
rect 19625 25857 19659 25891
rect 20545 25857 20579 25891
rect 20729 25857 20763 25891
rect 20821 25857 20855 25891
rect 21097 25857 21131 25891
rect 22089 25857 22123 25891
rect 4997 25721 5031 25755
rect 7021 25789 7055 25823
rect 7205 25789 7239 25823
rect 9505 25789 9539 25823
rect 11897 25789 11931 25823
rect 14197 25789 14231 25823
rect 17325 25789 17359 25823
rect 18797 25789 18831 25823
rect 18889 25789 18923 25823
rect 19901 25789 19935 25823
rect 19993 25789 20027 25823
rect 20913 25789 20947 25823
rect 21833 25789 21867 25823
rect 10885 25721 10919 25755
rect 1501 25653 1535 25687
rect 5641 25653 5675 25687
rect 6377 25653 6411 25687
rect 6561 25653 6595 25687
rect 8217 25653 8251 25687
rect 12817 25653 12851 25687
rect 16129 25653 16163 25687
rect 19717 25653 19751 25687
rect 20085 25653 20119 25687
rect 21281 25653 21315 25687
rect 23213 25653 23247 25687
rect 11069 25449 11103 25483
rect 12817 25449 12851 25483
rect 17785 25449 17819 25483
rect 19625 25449 19659 25483
rect 21373 25449 21407 25483
rect 23213 25449 23247 25483
rect 5641 25381 5675 25415
rect 7573 25381 7607 25415
rect 10793 25381 10827 25415
rect 14841 25381 14875 25415
rect 9413 25313 9447 25347
rect 10701 25313 10735 25347
rect 12357 25313 12391 25347
rect 12449 25313 12483 25347
rect 16681 25313 16715 25347
rect 18337 25313 18371 25347
rect 19901 25313 19935 25347
rect 21005 25313 21039 25347
rect 21833 25313 21867 25347
rect 4261 25245 4295 25279
rect 6193 25245 6227 25279
rect 8309 25245 8343 25279
rect 9137 25245 9171 25279
rect 9229 25245 9263 25279
rect 9505 25245 9539 25279
rect 10609 25245 10643 25279
rect 10885 25245 10919 25279
rect 12081 25245 12115 25279
rect 12265 25245 12299 25279
rect 12633 25245 12667 25279
rect 13277 25245 13311 25279
rect 13369 25245 13403 25279
rect 15301 25245 15335 25279
rect 19533 25245 19567 25279
rect 19993 25245 20027 25279
rect 20637 25245 20671 25279
rect 20821 25245 20855 25279
rect 20913 25245 20947 25279
rect 21189 25245 21223 25279
rect 22089 25245 22123 25279
rect 29837 25245 29871 25279
rect 4528 25177 4562 25211
rect 6460 25177 6494 25211
rect 14657 25177 14691 25211
rect 16957 25177 16991 25211
rect 18245 25177 18279 25211
rect 8217 25109 8251 25143
rect 8953 25109 8987 25143
rect 15393 25109 15427 25143
rect 16865 25109 16899 25143
rect 17325 25109 17359 25143
rect 18153 25109 18187 25143
rect 20177 25109 20211 25143
rect 30021 25109 30055 25143
rect 4813 24905 4847 24939
rect 7665 24905 7699 24939
rect 9321 24905 9355 24939
rect 12909 24905 12943 24939
rect 17877 24905 17911 24939
rect 19901 24905 19935 24939
rect 21005 24905 21039 24939
rect 15209 24837 15243 24871
rect 20361 24837 20395 24871
rect 1685 24769 1719 24803
rect 2697 24769 2731 24803
rect 2881 24769 2915 24803
rect 4077 24769 4111 24803
rect 4261 24769 4295 24803
rect 4629 24769 4663 24803
rect 5733 24769 5767 24803
rect 6377 24769 6411 24803
rect 6745 24769 6779 24803
rect 8585 24769 8619 24803
rect 8769 24769 8803 24803
rect 8953 24769 8987 24803
rect 9137 24769 9171 24803
rect 10241 24769 10275 24803
rect 10425 24769 10459 24803
rect 10517 24769 10551 24803
rect 10793 24769 10827 24803
rect 11529 24769 11563 24803
rect 11785 24769 11819 24803
rect 14749 24769 14783 24803
rect 14841 24769 14875 24803
rect 15025 24769 15059 24803
rect 15669 24769 15703 24803
rect 19073 24769 19107 24803
rect 19625 24769 19659 24803
rect 19717 24769 19751 24803
rect 20821 24769 20855 24803
rect 2789 24701 2823 24735
rect 4353 24701 4387 24735
rect 4445 24701 4479 24735
rect 1501 24633 1535 24667
rect 5549 24633 5583 24667
rect 7757 24701 7791 24735
rect 7849 24701 7883 24735
rect 8861 24701 8895 24735
rect 10609 24701 10643 24735
rect 10977 24701 11011 24735
rect 17601 24701 17635 24735
rect 17785 24701 17819 24735
rect 19901 24701 19935 24735
rect 20637 24701 20671 24735
rect 7297 24633 7331 24667
rect 6377 24565 6411 24599
rect 6653 24565 6687 24599
rect 15761 24565 15795 24599
rect 18245 24565 18279 24599
rect 18981 24565 19015 24599
rect 20453 24565 20487 24599
rect 6377 24361 6411 24395
rect 8125 24361 8159 24395
rect 14289 24361 14323 24395
rect 17877 24361 17911 24395
rect 19809 24361 19843 24395
rect 2789 24225 2823 24259
rect 4261 24225 4295 24259
rect 6009 24225 6043 24259
rect 7665 24225 7699 24259
rect 9781 24225 9815 24259
rect 12357 24225 12391 24259
rect 12449 24225 12483 24259
rect 16037 24225 16071 24259
rect 17325 24225 17359 24259
rect 22293 24225 22327 24259
rect 22477 24225 22511 24259
rect 1685 24157 1719 24191
rect 2697 24157 2731 24191
rect 2881 24157 2915 24191
rect 3985 24157 4019 24191
rect 4169 24157 4203 24191
rect 4353 24157 4387 24191
rect 4537 24157 4571 24191
rect 4997 24157 5031 24191
rect 5641 24157 5675 24191
rect 5825 24157 5859 24191
rect 5917 24157 5951 24191
rect 6193 24157 6227 24191
rect 7389 24157 7423 24191
rect 7573 24157 7607 24191
rect 7757 24157 7791 24191
rect 7941 24157 7975 24191
rect 9045 24157 9079 24191
rect 9137 24157 9171 24191
rect 12081 24157 12115 24191
rect 12265 24157 12299 24191
rect 12633 24157 12667 24191
rect 14197 24157 14231 24191
rect 14381 24157 14415 24191
rect 14841 24157 14875 24191
rect 14989 24157 15023 24191
rect 15209 24157 15243 24191
rect 15306 24157 15340 24191
rect 17509 24157 17543 24191
rect 18429 24157 18463 24191
rect 18613 24157 18647 24191
rect 19901 24157 19935 24191
rect 20361 24157 20395 24191
rect 5089 24089 5123 24123
rect 10026 24089 10060 24123
rect 15117 24089 15151 24123
rect 16221 24089 16255 24123
rect 22201 24089 22235 24123
rect 1501 24021 1535 24055
rect 3801 24021 3835 24055
rect 11161 24021 11195 24055
rect 12817 24021 12851 24055
rect 15485 24021 15519 24055
rect 16313 24021 16347 24055
rect 16681 24021 16715 24055
rect 17417 24021 17451 24055
rect 18521 24021 18555 24055
rect 20453 24021 20487 24055
rect 21833 24021 21867 24055
rect 4169 23817 4203 23851
rect 7665 23817 7699 23851
rect 9873 23817 9907 23851
rect 14289 23817 14323 23851
rect 18521 23817 18555 23851
rect 20085 23817 20119 23851
rect 11713 23749 11747 23783
rect 11897 23749 11931 23783
rect 13176 23749 13210 23783
rect 21925 23749 21959 23783
rect 2789 23681 2823 23715
rect 3056 23681 3090 23715
rect 4813 23681 4847 23715
rect 5181 23681 5215 23715
rect 5365 23681 5399 23715
rect 6377 23681 6411 23715
rect 6561 23681 6595 23715
rect 6653 23681 6687 23715
rect 6929 23681 6963 23715
rect 7849 23681 7883 23715
rect 7941 23681 7975 23715
rect 8217 23681 8251 23715
rect 9137 23681 9171 23715
rect 9321 23681 9355 23715
rect 9505 23681 9539 23715
rect 9689 23681 9723 23715
rect 10517 23681 10551 23715
rect 12909 23681 12943 23715
rect 14749 23681 14783 23715
rect 15761 23681 15795 23715
rect 16681 23681 16715 23715
rect 17141 23681 17175 23715
rect 17509 23681 17543 23715
rect 20269 23681 20303 23715
rect 20453 23681 20487 23715
rect 21097 23681 21131 23715
rect 22109 23681 22143 23715
rect 1409 23613 1443 23647
rect 1685 23613 1719 23647
rect 4997 23613 5031 23647
rect 5089 23613 5123 23647
rect 6745 23613 6779 23647
rect 9413 23613 9447 23647
rect 10425 23613 10459 23647
rect 15485 23613 15519 23647
rect 15669 23613 15703 23647
rect 17233 23613 17267 23647
rect 17417 23613 17451 23647
rect 18613 23613 18647 23647
rect 18797 23613 18831 23647
rect 21189 23613 21223 23647
rect 22661 23613 22695 23647
rect 22937 23613 22971 23647
rect 14841 23545 14875 23579
rect 4629 23477 4663 23511
rect 7113 23477 7147 23511
rect 8125 23477 8159 23511
rect 16129 23477 16163 23511
rect 16773 23477 16807 23511
rect 18153 23477 18187 23511
rect 20269 23477 20303 23511
rect 5457 23273 5491 23307
rect 7297 23273 7331 23307
rect 14933 23273 14967 23307
rect 15485 23273 15519 23307
rect 16773 23273 16807 23307
rect 19533 23273 19567 23307
rect 22569 23273 22603 23307
rect 4077 23137 4111 23171
rect 5917 23137 5951 23171
rect 9597 23137 9631 23171
rect 11253 23137 11287 23171
rect 12357 23137 12391 23171
rect 12449 23137 12483 23171
rect 16405 23137 16439 23171
rect 21465 23137 21499 23171
rect 21925 23137 21959 23171
rect 1409 23069 1443 23103
rect 2053 23069 2087 23103
rect 4344 23069 4378 23103
rect 6184 23069 6218 23103
rect 7757 23069 7791 23103
rect 9229 23069 9263 23103
rect 9413 23069 9447 23103
rect 9505 23069 9539 23103
rect 9781 23069 9815 23103
rect 10885 23069 10919 23103
rect 11069 23069 11103 23103
rect 11161 23069 11195 23103
rect 11437 23069 11471 23103
rect 12081 23069 12115 23103
rect 12265 23069 12299 23103
rect 12633 23069 12667 23103
rect 15393 23069 15427 23103
rect 16037 23069 16071 23103
rect 16221 23069 16255 23103
rect 16313 23069 16347 23103
rect 16589 23069 16623 23103
rect 18153 23069 18187 23103
rect 19441 23069 19475 23103
rect 20085 23069 20119 23103
rect 20269 23069 20303 23103
rect 20361 23069 20395 23103
rect 20453 23069 20487 23103
rect 21373 23069 21407 23103
rect 23581 23069 23615 23103
rect 29837 23069 29871 23103
rect 14565 23001 14599 23035
rect 14749 23001 14783 23035
rect 22753 23001 22787 23035
rect 22937 23001 22971 23035
rect 1593 22933 1627 22967
rect 2237 22933 2271 22967
rect 7849 22933 7883 22967
rect 9965 22933 9999 22967
rect 11621 22933 11655 22967
rect 12817 22933 12851 22967
rect 18337 22933 18371 22967
rect 20729 22933 20763 22967
rect 21741 22933 21775 22967
rect 23397 22933 23431 22967
rect 30021 22933 30055 22967
rect 7665 22729 7699 22763
rect 13829 22729 13863 22763
rect 14289 22729 14323 22763
rect 16957 22729 16991 22763
rect 17417 22729 17451 22763
rect 18981 22729 19015 22763
rect 19809 22729 19843 22763
rect 22201 22729 22235 22763
rect 15402 22661 15436 22695
rect 18153 22661 18187 22695
rect 20361 22661 20395 22695
rect 21833 22661 21867 22695
rect 22845 22661 22879 22695
rect 23029 22661 23063 22695
rect 1409 22593 1443 22627
rect 2237 22593 2271 22627
rect 2697 22593 2731 22627
rect 4997 22593 5031 22627
rect 6653 22593 6687 22627
rect 7849 22593 7883 22627
rect 8217 22593 8251 22627
rect 8401 22593 8435 22627
rect 9965 22593 9999 22627
rect 12449 22593 12483 22627
rect 12705 22593 12739 22627
rect 15669 22593 15703 22627
rect 17049 22593 17083 22627
rect 18337 22593 18371 22627
rect 19165 22593 19199 22627
rect 19901 22593 19935 22627
rect 20729 22593 20763 22627
rect 22006 22593 22040 22627
rect 5273 22525 5307 22559
rect 6377 22525 6411 22559
rect 8033 22525 8067 22559
rect 8125 22525 8159 22559
rect 10241 22525 10275 22559
rect 16865 22525 16899 22559
rect 20545 22525 20579 22559
rect 22661 22525 22695 22559
rect 20729 22457 20763 22491
rect 1593 22389 1627 22423
rect 2053 22389 2087 22423
rect 2881 22389 2915 22423
rect 18521 22389 18555 22423
rect 11161 22185 11195 22219
rect 13001 22185 13035 22219
rect 17969 22185 18003 22219
rect 20913 22185 20947 22219
rect 22569 22185 22603 22219
rect 4629 22049 4663 22083
rect 6653 22049 6687 22083
rect 9045 22049 9079 22083
rect 15393 22049 15427 22083
rect 16589 22049 16623 22083
rect 16957 22049 16991 22083
rect 18429 22049 18463 22083
rect 18613 22049 18647 22083
rect 19717 22049 19751 22083
rect 19901 22049 19935 22083
rect 20545 22049 20579 22083
rect 1869 21981 1903 22015
rect 4721 21981 4755 22015
rect 6561 21981 6595 22015
rect 7389 21981 7423 22015
rect 9781 21981 9815 22015
rect 10048 21981 10082 22015
rect 11621 21981 11655 22015
rect 15490 21981 15524 22015
rect 16497 21981 16531 22015
rect 16681 21981 16715 22015
rect 16773 21981 16807 22015
rect 17049 21981 17083 22015
rect 20453 21981 20487 22015
rect 20729 21981 20763 22015
rect 21833 21981 21867 22015
rect 22477 21981 22511 22015
rect 2136 21913 2170 21947
rect 8033 21913 8067 21947
rect 8217 21913 8251 21947
rect 8401 21913 8435 21947
rect 9229 21913 9263 21947
rect 11888 21913 11922 21947
rect 15117 21913 15151 21947
rect 15301 21913 15335 21947
rect 15393 21913 15427 21947
rect 18337 21913 18371 21947
rect 19625 21913 19659 21947
rect 21649 21913 21683 21947
rect 22017 21913 22051 21947
rect 3249 21845 3283 21879
rect 7481 21845 7515 21879
rect 19257 21845 19291 21879
rect 7665 21641 7699 21675
rect 8953 21641 8987 21675
rect 10793 21641 10827 21675
rect 12265 21641 12299 21675
rect 14933 21641 14967 21675
rect 17417 21641 17451 21675
rect 17877 21641 17911 21675
rect 18337 21641 18371 21675
rect 21005 21641 21039 21675
rect 6745 21573 6779 21607
rect 8585 21573 8619 21607
rect 9669 21573 9703 21607
rect 15393 21573 15427 21607
rect 20085 21573 20119 21607
rect 1961 21505 1995 21539
rect 2228 21505 2262 21539
rect 3801 21505 3835 21539
rect 6556 21505 6590 21539
rect 6653 21505 6687 21539
rect 6873 21505 6907 21539
rect 7021 21505 7055 21539
rect 7757 21505 7791 21539
rect 8316 21505 8350 21539
rect 8402 21505 8436 21539
rect 8685 21505 8719 21539
rect 8815 21505 8849 21539
rect 11529 21505 11563 21539
rect 11713 21505 11747 21539
rect 11805 21505 11839 21539
rect 12081 21505 12115 21539
rect 15301 21505 15335 21539
rect 16681 21505 16715 21539
rect 16865 21505 16899 21539
rect 16957 21505 16991 21539
rect 17233 21505 17267 21539
rect 18245 21505 18279 21539
rect 19073 21505 19107 21539
rect 19246 21505 19280 21539
rect 19349 21505 19383 21539
rect 19625 21505 19659 21539
rect 20269 21505 20303 21539
rect 21097 21505 21131 21539
rect 29837 21505 29871 21539
rect 9413 21437 9447 21471
rect 11897 21437 11931 21471
rect 15485 21437 15519 21471
rect 17049 21437 17083 21471
rect 18429 21437 18463 21471
rect 3341 21301 3375 21335
rect 3893 21301 3927 21335
rect 6377 21301 6411 21335
rect 19073 21301 19107 21335
rect 19533 21301 19567 21335
rect 20453 21301 20487 21335
rect 30021 21301 30055 21335
rect 2329 21097 2363 21131
rect 5457 21097 5491 21131
rect 7389 21097 7423 21131
rect 8217 21097 8251 21131
rect 8401 21097 8435 21131
rect 16773 21097 16807 21131
rect 17233 21097 17267 21131
rect 19257 21097 19291 21131
rect 19717 21097 19751 21131
rect 10425 21029 10459 21063
rect 21741 21029 21775 21063
rect 1961 20961 1995 20995
rect 4169 20961 4203 20995
rect 9689 20961 9723 20995
rect 15485 20961 15519 20995
rect 16221 20961 16255 20995
rect 17785 20961 17819 20995
rect 21097 20961 21131 20995
rect 1593 20893 1627 20927
rect 1777 20893 1811 20927
rect 1869 20893 1903 20927
rect 2145 20893 2179 20927
rect 3065 20893 3099 20927
rect 3801 20893 3835 20927
rect 3985 20893 4019 20927
rect 4077 20893 4111 20927
rect 4353 20893 4387 20927
rect 6570 20893 6604 20927
rect 6837 20893 6871 20927
rect 7481 20893 7515 20927
rect 7941 20893 7975 20927
rect 9965 20893 9999 20927
rect 13369 20893 13403 20927
rect 13461 20893 13495 20927
rect 16313 20893 16347 20927
rect 17693 20893 17727 20927
rect 18429 20893 18463 20927
rect 18613 20893 18647 20927
rect 19441 20893 19475 20927
rect 19533 20893 19567 20927
rect 19809 20893 19843 20927
rect 21005 20893 21039 20927
rect 21925 20893 21959 20927
rect 22109 20893 22143 20927
rect 10609 20825 10643 20859
rect 15209 20825 15243 20859
rect 16405 20825 16439 20859
rect 3157 20757 3191 20791
rect 4537 20757 4571 20791
rect 14841 20757 14875 20791
rect 15301 20757 15335 20791
rect 17601 20757 17635 20791
rect 18521 20757 18555 20791
rect 20545 20757 20579 20791
rect 20913 20757 20947 20791
rect 2237 20553 2271 20587
rect 5181 20553 5215 20587
rect 8033 20553 8067 20587
rect 9321 20553 9355 20587
rect 15393 20553 15427 20587
rect 16865 20553 16899 20587
rect 19165 20553 19199 20587
rect 19257 20553 19291 20587
rect 20269 20553 20303 20587
rect 20729 20553 20763 20587
rect 22293 20553 22327 20587
rect 4068 20485 4102 20519
rect 8493 20485 8527 20519
rect 9689 20485 9723 20519
rect 11713 20485 11747 20519
rect 12265 20485 12299 20519
rect 14933 20485 14967 20519
rect 17325 20485 17359 20519
rect 22201 20485 22235 20519
rect 1501 20417 1535 20451
rect 1685 20417 1719 20451
rect 1777 20417 1811 20451
rect 2053 20417 2087 20451
rect 2881 20417 2915 20451
rect 5641 20417 5675 20451
rect 6920 20417 6954 20451
rect 8677 20417 8711 20451
rect 8861 20417 8895 20451
rect 9505 20417 9539 20451
rect 10149 20417 10183 20451
rect 12449 20417 12483 20451
rect 13461 20417 13495 20451
rect 13921 20417 13955 20451
rect 15025 20417 15059 20451
rect 15853 20417 15887 20451
rect 16129 20417 16163 20451
rect 17233 20417 17267 20451
rect 18061 20417 18095 20451
rect 18245 20417 18279 20451
rect 20637 20417 20671 20451
rect 1869 20349 1903 20383
rect 3801 20349 3835 20383
rect 6653 20349 6687 20383
rect 10241 20349 10275 20383
rect 14841 20349 14875 20383
rect 17417 20349 17451 20383
rect 19073 20349 19107 20383
rect 20821 20349 20855 20383
rect 22385 20349 22419 20383
rect 13553 20281 13587 20315
rect 21833 20281 21867 20315
rect 2697 20213 2731 20247
rect 5733 20213 5767 20247
rect 11621 20213 11655 20247
rect 13645 20213 13679 20247
rect 13783 20213 13817 20247
rect 18429 20213 18463 20247
rect 19625 20213 19659 20247
rect 7113 20009 7147 20043
rect 7573 20009 7607 20043
rect 7941 20009 7975 20043
rect 9413 20009 9447 20043
rect 12909 20009 12943 20043
rect 16681 20009 16715 20043
rect 20453 20009 20487 20043
rect 3249 19941 3283 19975
rect 9873 19941 9907 19975
rect 10425 19941 10459 19975
rect 14381 19941 14415 19975
rect 14473 19941 14507 19975
rect 19349 19941 19383 19975
rect 21741 19941 21775 19975
rect 4445 19873 4479 19907
rect 6653 19873 6687 19907
rect 6745 19873 6779 19907
rect 10609 19873 10643 19907
rect 11529 19873 11563 19907
rect 15761 19873 15795 19907
rect 16037 19873 16071 19907
rect 17969 19873 18003 19907
rect 1869 19805 1903 19839
rect 4077 19805 4111 19839
rect 4261 19805 4295 19839
rect 4353 19805 4387 19839
rect 4629 19805 4663 19839
rect 5365 19805 5399 19839
rect 6377 19805 6411 19839
rect 6561 19805 6595 19839
rect 6929 19805 6963 19839
rect 8033 19805 8067 19839
rect 9597 19805 9631 19839
rect 9689 19805 9723 19839
rect 9965 19805 9999 19839
rect 10701 19805 10735 19839
rect 10977 19805 11011 19839
rect 11069 19805 11103 19839
rect 13553 19805 13587 19839
rect 14105 19805 14139 19839
rect 14289 19805 14323 19839
rect 14565 19805 14599 19839
rect 15853 19805 15887 19839
rect 15945 19805 15979 19839
rect 16865 19805 16899 19839
rect 17693 19805 17727 19839
rect 19441 19805 19475 19839
rect 20177 19805 20211 19839
rect 20269 19805 20303 19839
rect 20545 19805 20579 19839
rect 21925 19805 21959 19839
rect 22109 19805 22143 19839
rect 2136 19737 2170 19771
rect 11796 19737 11830 19771
rect 13461 19737 13495 19771
rect 4813 19669 4847 19703
rect 5457 19669 5491 19703
rect 14749 19669 14783 19703
rect 15577 19669 15611 19703
rect 17325 19669 17359 19703
rect 17785 19669 17819 19703
rect 19993 19669 20027 19703
rect 13185 19465 13219 19499
rect 14105 19465 14139 19499
rect 16037 19465 16071 19499
rect 17601 19465 17635 19499
rect 18797 19465 18831 19499
rect 4620 19397 4654 19431
rect 8677 19397 8711 19431
rect 9321 19397 9355 19431
rect 10057 19397 10091 19431
rect 10241 19397 10275 19431
rect 11897 19397 11931 19431
rect 15218 19397 15252 19431
rect 19165 19397 19199 19431
rect 19257 19397 19291 19431
rect 23213 19397 23247 19431
rect 1409 19329 1443 19363
rect 2237 19329 2271 19363
rect 2504 19329 2538 19363
rect 4353 19329 4387 19363
rect 6377 19329 6411 19363
rect 6469 19329 6503 19363
rect 8769 19329 8803 19363
rect 9413 19329 9447 19363
rect 9873 19329 9907 19363
rect 10977 19329 11011 19363
rect 15485 19329 15519 19363
rect 15945 19329 15979 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 17969 19329 18003 19363
rect 19993 19329 20027 19363
rect 20269 19329 20303 19363
rect 20361 19329 20395 19363
rect 20545 19329 20579 19363
rect 21005 19329 21039 19363
rect 21189 19329 21223 19363
rect 22477 19329 22511 19363
rect 22569 19329 22603 19363
rect 22753 19329 22787 19363
rect 29837 19329 29871 19363
rect 18061 19261 18095 19295
rect 18245 19261 18279 19295
rect 19349 19261 19383 19295
rect 1593 19193 1627 19227
rect 5733 19193 5767 19227
rect 10793 19193 10827 19227
rect 3617 19125 3651 19159
rect 16773 19125 16807 19159
rect 20085 19125 20119 19159
rect 20177 19125 20211 19159
rect 21005 19125 21039 19159
rect 30021 19125 30055 19159
rect 2237 18921 2271 18955
rect 12265 18921 12299 18955
rect 18245 18921 18279 18955
rect 19349 18921 19383 18955
rect 29929 18921 29963 18955
rect 4031 18853 4065 18887
rect 11069 18853 11103 18887
rect 14289 18853 14323 18887
rect 21649 18853 21683 18887
rect 1777 18785 1811 18819
rect 1869 18785 1903 18819
rect 6469 18785 6503 18819
rect 7849 18785 7883 18819
rect 7941 18785 7975 18819
rect 9229 18785 9263 18819
rect 11897 18785 11931 18819
rect 15025 18785 15059 18819
rect 17325 18785 17359 18819
rect 20453 18785 20487 18819
rect 20545 18785 20579 18819
rect 22201 18785 22235 18819
rect 1501 18717 1535 18751
rect 1685 18717 1719 18751
rect 2053 18717 2087 18751
rect 3801 18717 3835 18751
rect 5457 18717 5491 18751
rect 6193 18717 6227 18751
rect 7665 18717 7699 18751
rect 8033 18717 8067 18751
rect 8217 18717 8251 18751
rect 8953 18717 8987 18751
rect 9137 18717 9171 18751
rect 9321 18717 9355 18751
rect 9505 18717 9539 18751
rect 11529 18717 11563 18751
rect 11713 18717 11747 18751
rect 11805 18717 11839 18751
rect 12081 18717 12115 18751
rect 12725 18717 12759 18751
rect 14197 18717 14231 18751
rect 16313 18717 16347 18751
rect 17601 18717 17635 18751
rect 18429 18717 18463 18751
rect 19257 18717 19291 18751
rect 20361 18717 20395 18751
rect 22017 18717 22051 18751
rect 22109 18717 22143 18751
rect 29929 18717 29963 18751
rect 30113 18717 30147 18751
rect 3157 18649 3191 18683
rect 10885 18649 10919 18683
rect 15117 18649 15151 18683
rect 15209 18649 15243 18683
rect 16037 18649 16071 18683
rect 3065 18581 3099 18615
rect 5549 18581 5583 18615
rect 7481 18581 7515 18615
rect 9689 18581 9723 18615
rect 12909 18581 12943 18615
rect 15577 18581 15611 18615
rect 19993 18581 20027 18615
rect 2421 18377 2455 18411
rect 4169 18377 4203 18411
rect 4813 18377 4847 18411
rect 5733 18377 5767 18411
rect 8309 18377 8343 18411
rect 8861 18377 8895 18411
rect 12081 18377 12115 18411
rect 15393 18377 15427 18411
rect 18981 18377 19015 18411
rect 19349 18377 19383 18411
rect 20545 18377 20579 18411
rect 20913 18377 20947 18411
rect 21833 18377 21867 18411
rect 30021 18377 30055 18411
rect 5641 18309 5675 18343
rect 7196 18309 7230 18343
rect 12817 18309 12851 18343
rect 15301 18309 15335 18343
rect 19441 18309 19475 18343
rect 1685 18241 1719 18275
rect 1869 18241 1903 18275
rect 2237 18241 2271 18275
rect 3065 18241 3099 18275
rect 3433 18241 3467 18275
rect 3617 18241 3651 18275
rect 4261 18241 4295 18275
rect 4997 18241 5031 18275
rect 6929 18241 6963 18275
rect 9974 18241 10008 18275
rect 10241 18241 10275 18275
rect 10977 18241 11011 18275
rect 11989 18241 12023 18275
rect 12909 18241 12943 18275
rect 16865 18241 16899 18275
rect 21005 18241 21039 18275
rect 22017 18241 22051 18275
rect 29929 18241 29963 18275
rect 30113 18241 30147 18275
rect 1961 18173 1995 18207
rect 2053 18173 2087 18207
rect 3249 18173 3283 18207
rect 3341 18173 3375 18207
rect 15577 18173 15611 18207
rect 17141 18173 17175 18207
rect 19533 18173 19567 18207
rect 21097 18173 21131 18207
rect 10793 18105 10827 18139
rect 2881 18037 2915 18071
rect 14933 18037 14967 18071
rect 6009 17833 6043 17867
rect 7941 17833 7975 17867
rect 11345 17833 11379 17867
rect 15485 17833 15519 17867
rect 16773 17833 16807 17867
rect 19717 17833 19751 17867
rect 20637 17833 20671 17867
rect 13277 17765 13311 17799
rect 14473 17765 14507 17799
rect 18429 17765 18463 17799
rect 21833 17765 21867 17799
rect 3801 17697 3835 17731
rect 13369 17697 13403 17731
rect 13553 17697 13587 17731
rect 14289 17697 14323 17731
rect 14381 17697 14415 17731
rect 15393 17697 15427 17731
rect 15577 17697 15611 17731
rect 16221 17697 16255 17731
rect 19257 17697 19291 17731
rect 1593 17629 1627 17663
rect 1860 17629 1894 17663
rect 4077 17629 4111 17663
rect 5273 17629 5307 17663
rect 6101 17629 6135 17663
rect 6561 17629 6595 17663
rect 9965 17629 9999 17663
rect 12449 17629 12483 17663
rect 12633 17629 12667 17663
rect 13277 17629 13311 17663
rect 14105 17629 14139 17663
rect 14565 17629 14599 17663
rect 15301 17629 15335 17663
rect 16405 17629 16439 17663
rect 17877 17629 17911 17663
rect 18153 17629 18187 17663
rect 18705 17629 18739 17663
rect 19441 17629 19475 17663
rect 19533 17629 19567 17663
rect 19809 17629 19843 17663
rect 20269 17629 20303 17663
rect 20453 17629 20487 17663
rect 21097 17629 21131 17663
rect 21741 17629 21775 17663
rect 6828 17561 6862 17595
rect 10210 17561 10244 17595
rect 21189 17561 21223 17595
rect 2973 17493 3007 17527
rect 5089 17493 5123 17527
rect 12541 17493 12575 17527
rect 14749 17493 14783 17527
rect 16313 17493 16347 17527
rect 7481 17289 7515 17323
rect 9137 17289 9171 17323
rect 9597 17289 9631 17323
rect 14841 17289 14875 17323
rect 16957 17289 16991 17323
rect 20453 17289 20487 17323
rect 21925 17289 21959 17323
rect 11980 17221 12014 17255
rect 14197 17221 14231 17255
rect 17601 17221 17635 17255
rect 18429 17221 18463 17255
rect 1409 17153 1443 17187
rect 2605 17153 2639 17187
rect 4160 17153 4194 17187
rect 6745 17153 6779 17187
rect 6929 17153 6963 17187
rect 7297 17153 7331 17187
rect 8401 17153 8435 17187
rect 8585 17153 8619 17187
rect 8677 17153 8711 17187
rect 8953 17153 8987 17187
rect 10721 17153 10755 17187
rect 14013 17153 14047 17187
rect 14749 17153 14783 17187
rect 17141 17153 17175 17187
rect 18061 17153 18095 17187
rect 18245 17153 18279 17187
rect 19257 17153 19291 17187
rect 19441 17153 19475 17187
rect 19671 17153 19705 17187
rect 19809 17153 19843 17187
rect 20729 17153 20763 17187
rect 21833 17153 21867 17187
rect 29837 17153 29871 17187
rect 2881 17085 2915 17119
rect 3893 17085 3927 17119
rect 7021 17085 7055 17119
rect 7113 17085 7147 17119
rect 8769 17085 8803 17119
rect 10977 17085 11011 17119
rect 11713 17085 11747 17119
rect 13829 17085 13863 17119
rect 17233 17085 17267 17119
rect 19533 17085 19567 17119
rect 20453 17085 20487 17119
rect 20637 17085 20671 17119
rect 1593 16949 1627 16983
rect 5273 16949 5307 16983
rect 13093 16949 13127 16983
rect 19993 16949 20027 16983
rect 30021 16949 30055 16983
rect 10977 16745 11011 16779
rect 13277 16745 13311 16779
rect 14105 16745 14139 16779
rect 17233 16745 17267 16779
rect 21741 16745 21775 16779
rect 14381 16677 14415 16711
rect 15117 16677 15151 16711
rect 4353 16609 4387 16643
rect 9505 16609 9539 16643
rect 10517 16609 10551 16643
rect 13185 16609 13219 16643
rect 14473 16609 14507 16643
rect 1409 16541 1443 16575
rect 2973 16541 3007 16575
rect 3249 16541 3283 16575
rect 6193 16541 6227 16575
rect 6837 16541 6871 16575
rect 9781 16541 9815 16575
rect 10241 16541 10275 16575
rect 10425 16541 10459 16575
rect 10609 16541 10643 16575
rect 10793 16541 10827 16575
rect 11989 16541 12023 16575
rect 13406 16541 13440 16575
rect 13553 16541 13587 16575
rect 14289 16541 14323 16575
rect 14565 16541 14599 16575
rect 15301 16541 15335 16575
rect 16221 16541 16255 16575
rect 16405 16541 16439 16575
rect 17049 16541 17083 16575
rect 17233 16541 17267 16575
rect 19441 16541 19475 16575
rect 20361 16541 20395 16575
rect 20617 16541 20651 16575
rect 4598 16473 4632 16507
rect 12357 16473 12391 16507
rect 16589 16473 16623 16507
rect 1593 16405 1627 16439
rect 5733 16405 5767 16439
rect 6285 16405 6319 16439
rect 6929 16405 6963 16439
rect 12909 16405 12943 16439
rect 17417 16405 17451 16439
rect 19349 16405 19383 16439
rect 4261 16201 4295 16235
rect 7205 16201 7239 16235
rect 10977 16201 11011 16235
rect 13737 16201 13771 16235
rect 18337 16201 18371 16235
rect 30021 16201 30055 16235
rect 7113 16133 7147 16167
rect 12725 16133 12759 16167
rect 20269 16133 20303 16167
rect 1941 16065 1975 16099
rect 3525 16065 3559 16099
rect 3709 16065 3743 16099
rect 4077 16065 4111 16099
rect 4997 16065 5031 16099
rect 5641 16065 5675 16099
rect 6377 16065 6411 16099
rect 9045 16065 9079 16099
rect 9597 16065 9631 16099
rect 9864 16065 9898 16099
rect 12817 16065 12851 16099
rect 13553 16065 13587 16099
rect 14473 16065 14507 16099
rect 16957 16065 16991 16099
rect 17224 16065 17258 16099
rect 18889 16065 18923 16099
rect 19073 16065 19107 16099
rect 19257 16065 19291 16099
rect 19441 16065 19475 16099
rect 20453 16065 20487 16099
rect 21189 16065 21223 16099
rect 29929 16065 29963 16099
rect 30113 16065 30147 16099
rect 1685 15997 1719 16031
rect 3801 15997 3835 16031
rect 3893 15997 3927 16031
rect 8769 15997 8803 16031
rect 13277 15997 13311 16031
rect 14749 15997 14783 16031
rect 19165 15997 19199 16031
rect 3065 15929 3099 15963
rect 20085 15929 20119 15963
rect 5089 15861 5123 15895
rect 5733 15861 5767 15895
rect 6469 15861 6503 15895
rect 13369 15861 13403 15895
rect 15853 15861 15887 15895
rect 19625 15861 19659 15895
rect 21005 15861 21039 15895
rect 1777 15657 1811 15691
rect 4537 15657 4571 15691
rect 8953 15657 8987 15691
rect 9781 15657 9815 15691
rect 14565 15657 14599 15691
rect 16129 15657 16163 15691
rect 17417 15657 17451 15691
rect 20821 15657 20855 15691
rect 29929 15657 29963 15691
rect 2145 15521 2179 15555
rect 4169 15521 4203 15555
rect 6009 15521 6043 15555
rect 9413 15521 9447 15555
rect 10333 15521 10367 15555
rect 13461 15521 13495 15555
rect 15025 15521 15059 15555
rect 16957 15521 16991 15555
rect 1961 15453 1995 15487
rect 2237 15453 2271 15487
rect 2329 15453 2363 15487
rect 2513 15453 2547 15487
rect 3157 15453 3191 15487
rect 3801 15453 3835 15487
rect 3985 15453 4019 15487
rect 4077 15453 4111 15487
rect 4353 15453 4387 15487
rect 5089 15453 5123 15487
rect 5733 15453 5767 15487
rect 5917 15453 5951 15487
rect 6101 15453 6135 15487
rect 6285 15453 6319 15487
rect 7573 15453 7607 15487
rect 7666 15453 7700 15487
rect 8079 15453 8113 15487
rect 8953 15453 8987 15487
rect 9045 15453 9079 15487
rect 9229 15453 9263 15487
rect 9321 15453 9355 15487
rect 9597 15453 9631 15487
rect 10241 15453 10275 15487
rect 12633 15453 12667 15487
rect 13093 15453 13127 15487
rect 13277 15453 13311 15487
rect 14749 15453 14783 15487
rect 14933 15453 14967 15487
rect 15113 15451 15147 15485
rect 15301 15453 15335 15487
rect 16681 15453 16715 15487
rect 16853 15453 16887 15487
rect 17049 15453 17083 15487
rect 17233 15453 17267 15487
rect 18613 15453 18647 15487
rect 19441 15453 19475 15487
rect 19708 15453 19742 15487
rect 21281 15453 21315 15487
rect 29929 15453 29963 15487
rect 30113 15453 30147 15487
rect 7849 15385 7883 15419
rect 7941 15385 7975 15419
rect 16037 15385 16071 15419
rect 2973 15317 3007 15351
rect 5181 15317 5215 15351
rect 6469 15317 6503 15351
rect 8217 15317 8251 15351
rect 12449 15317 12483 15351
rect 18521 15317 18555 15351
rect 21465 15317 21499 15351
rect 7665 15113 7699 15147
rect 17693 15113 17727 15147
rect 3525 15045 3559 15079
rect 4230 15045 4264 15079
rect 8778 15045 8812 15079
rect 9750 15045 9784 15079
rect 11805 15045 11839 15079
rect 18429 15045 18463 15079
rect 19533 15045 19567 15079
rect 1777 14977 1811 15011
rect 1961 14977 1995 15011
rect 2145 14977 2179 15011
rect 2329 14977 2363 15011
rect 2789 14977 2823 15011
rect 2973 14977 3007 15011
rect 3157 14977 3191 15011
rect 3341 14977 3375 15011
rect 6377 14977 6411 15011
rect 6561 14977 6595 15011
rect 6653 14977 6687 15011
rect 6929 14977 6963 15011
rect 9045 14977 9079 15011
rect 9505 14977 9539 15011
rect 12265 14977 12299 15011
rect 12403 14977 12437 15011
rect 12541 14977 12575 15011
rect 13277 14977 13311 15011
rect 13461 14977 13495 15011
rect 14473 14977 14507 15011
rect 14729 14977 14763 15011
rect 17141 14977 17175 15011
rect 17417 14977 17451 15011
rect 17509 14977 17543 15011
rect 18153 14977 18187 15011
rect 18301 14977 18335 15011
rect 18521 14977 18555 15011
rect 18618 14977 18652 15011
rect 19349 14977 19383 15011
rect 20453 14977 20487 15011
rect 20729 14977 20763 15011
rect 20821 14977 20855 15011
rect 21833 14977 21867 15011
rect 22109 14977 22143 15011
rect 29193 14977 29227 15011
rect 29377 14977 29411 15011
rect 29837 14977 29871 15011
rect 2053 14909 2087 14943
rect 3065 14909 3099 14943
rect 3985 14909 4019 14943
rect 6745 14909 6779 14943
rect 7113 14841 7147 14875
rect 20545 14841 20579 14875
rect 21005 14841 21039 14875
rect 29193 14841 29227 14875
rect 30021 14841 30055 14875
rect 1593 14773 1627 14807
rect 5365 14773 5399 14807
rect 10885 14773 10919 14807
rect 13277 14773 13311 14807
rect 15853 14773 15887 14807
rect 17233 14773 17267 14807
rect 18797 14773 18831 14807
rect 1593 14569 1627 14603
rect 5181 14569 5215 14603
rect 8125 14569 8159 14603
rect 9597 14569 9631 14603
rect 14473 14569 14507 14603
rect 18429 14569 18463 14603
rect 29929 14569 29963 14603
rect 13553 14501 13587 14535
rect 19901 14501 19935 14535
rect 20361 14501 20395 14535
rect 2789 14433 2823 14467
rect 5917 14433 5951 14467
rect 6377 14433 6411 14467
rect 7113 14433 7147 14467
rect 12173 14433 12207 14467
rect 14933 14433 14967 14467
rect 16313 14433 16347 14467
rect 17417 14433 17451 14467
rect 17877 14433 17911 14467
rect 1409 14365 1443 14399
rect 2513 14365 2547 14399
rect 2697 14365 2731 14399
rect 2881 14365 2915 14399
rect 3065 14365 3099 14399
rect 3801 14365 3835 14399
rect 5641 14365 5675 14399
rect 5825 14365 5859 14399
rect 6009 14365 6043 14399
rect 6193 14365 6227 14399
rect 6837 14365 6871 14399
rect 7021 14365 7055 14399
rect 7205 14365 7239 14399
rect 7389 14365 7423 14399
rect 8953 14365 8987 14399
rect 9046 14365 9080 14399
rect 9321 14365 9355 14399
rect 9418 14365 9452 14399
rect 10793 14365 10827 14399
rect 10977 14365 11011 14399
rect 11529 14365 11563 14399
rect 12440 14365 12474 14399
rect 14657 14365 14691 14399
rect 14841 14365 14875 14399
rect 15025 14365 15059 14399
rect 15209 14365 15243 14399
rect 16221 14365 16255 14399
rect 16497 14365 16531 14399
rect 16589 14365 16623 14399
rect 17325 14365 17359 14399
rect 17601 14365 17635 14399
rect 17693 14365 17727 14399
rect 18337 14365 18371 14399
rect 19809 14365 19843 14399
rect 20085 14365 20119 14399
rect 20177 14365 20211 14399
rect 20821 14365 20855 14399
rect 29929 14365 29963 14399
rect 30113 14365 30147 14399
rect 3249 14297 3283 14331
rect 4046 14297 4080 14331
rect 8217 14297 8251 14331
rect 8401 14297 8435 14331
rect 9229 14297 9263 14331
rect 10149 14297 10183 14331
rect 10333 14297 10367 14331
rect 16773 14297 16807 14331
rect 7573 14229 7607 14263
rect 10885 14229 10919 14263
rect 11713 14229 11747 14263
rect 21051 14229 21085 14263
rect 2789 14025 2823 14059
rect 5733 14025 5767 14059
rect 7113 14025 7147 14059
rect 11713 14025 11747 14059
rect 19165 14025 19199 14059
rect 30021 14025 30055 14059
rect 12817 13957 12851 13991
rect 15577 13957 15611 13991
rect 1409 13889 1443 13923
rect 1665 13889 1699 13923
rect 3617 13889 3651 13923
rect 4905 13889 4939 13923
rect 4997 13889 5031 13923
rect 5641 13889 5675 13923
rect 6365 13889 6399 13923
rect 6561 13889 6595 13923
rect 6653 13889 6687 13923
rect 6929 13889 6963 13923
rect 8309 13889 8343 13923
rect 8953 13889 8987 13923
rect 10057 13889 10091 13923
rect 10609 13889 10643 13923
rect 11897 13889 11931 13923
rect 12633 13889 12667 13923
rect 13553 13889 13587 13923
rect 15117 13889 15151 13923
rect 16865 13889 16899 13923
rect 17141 13889 17175 13923
rect 17601 13889 17635 13923
rect 17785 13889 17819 13923
rect 18613 13889 18647 13923
rect 19349 13889 19383 13923
rect 20269 13889 20303 13923
rect 20545 13889 20579 13923
rect 20637 13889 20671 13923
rect 29929 13889 29963 13923
rect 30113 13889 30147 13923
rect 3341 13821 3375 13855
rect 6745 13821 6779 13855
rect 9137 13821 9171 13855
rect 12081 13821 12115 13855
rect 16957 13821 16991 13855
rect 20821 13821 20855 13855
rect 8125 13753 8159 13787
rect 20361 13753 20395 13787
rect 9873 13685 9907 13719
rect 10793 13685 10827 13719
rect 13461 13685 13495 13719
rect 16681 13685 16715 13719
rect 17141 13685 17175 13719
rect 17877 13685 17911 13719
rect 18521 13685 18555 13719
rect 4169 13481 4203 13515
rect 9689 13481 9723 13515
rect 9873 13481 9907 13515
rect 11713 13481 11747 13515
rect 18245 13481 18279 13515
rect 19717 13481 19751 13515
rect 6469 13413 6503 13447
rect 14473 13413 14507 13447
rect 15761 13413 15795 13447
rect 2237 13345 2271 13379
rect 6009 13345 6043 13379
rect 7205 13345 7239 13379
rect 13093 13345 13127 13379
rect 20453 13345 20487 13379
rect 1409 13277 1443 13311
rect 2513 13277 2547 13311
rect 4077 13277 4111 13311
rect 5733 13277 5767 13311
rect 5917 13277 5951 13311
rect 6101 13277 6135 13311
rect 6285 13277 6319 13311
rect 6929 13277 6963 13311
rect 8401 13277 8435 13311
rect 10333 13277 10367 13311
rect 10600 13277 10634 13311
rect 14933 13277 14967 13311
rect 15301 13277 15335 13311
rect 16129 13277 16163 13311
rect 17141 13277 17175 13311
rect 17233 13277 17267 13311
rect 17509 13277 17543 13311
rect 17785 13277 17819 13311
rect 18245 13277 18279 13311
rect 18337 13277 18371 13311
rect 19809 13277 19843 13311
rect 20361 13277 20395 13311
rect 20637 13277 20671 13311
rect 20729 13277 20763 13311
rect 29837 13277 29871 13311
rect 5181 13209 5215 13243
rect 9505 13209 9539 13243
rect 12817 13209 12851 13243
rect 14289 13209 14323 13243
rect 15117 13209 15151 13243
rect 15945 13209 15979 13243
rect 16957 13209 16991 13243
rect 20913 13209 20947 13243
rect 1593 13141 1627 13175
rect 5089 13141 5123 13175
rect 8309 13141 8343 13175
rect 9715 13141 9749 13175
rect 18613 13141 18647 13175
rect 30021 13141 30055 13175
rect 5641 12937 5675 12971
rect 16129 12937 16163 12971
rect 18337 12937 18371 12971
rect 30021 12937 30055 12971
rect 5733 12869 5767 12903
rect 10609 12869 10643 12903
rect 13093 12869 13127 12903
rect 15301 12869 15335 12903
rect 19450 12869 19484 12903
rect 20177 12869 20211 12903
rect 1409 12801 1443 12835
rect 2789 12801 2823 12835
rect 3065 12801 3099 12835
rect 3873 12801 3907 12835
rect 6377 12801 6411 12835
rect 6561 12801 6595 12835
rect 6653 12801 6687 12835
rect 6929 12801 6963 12835
rect 7113 12801 7147 12835
rect 9505 12801 9539 12835
rect 9689 12801 9723 12835
rect 11897 12801 11931 12835
rect 12081 12801 12115 12835
rect 12449 12801 12483 12835
rect 13277 12801 13311 12835
rect 15025 12801 15059 12835
rect 15761 12801 15795 12835
rect 15945 12801 15979 12835
rect 16865 12801 16899 12835
rect 17049 12801 17083 12835
rect 17325 12801 17359 12835
rect 19717 12801 19751 12835
rect 20269 12801 20303 12835
rect 29929 12801 29963 12835
rect 30113 12801 30147 12835
rect 3617 12733 3651 12767
rect 6745 12733 6779 12767
rect 8493 12733 8527 12767
rect 8769 12733 8803 12767
rect 10793 12733 10827 12767
rect 12173 12733 12207 12767
rect 12265 12733 12299 12767
rect 16681 12733 16715 12767
rect 1593 12597 1627 12631
rect 4997 12597 5031 12631
rect 9321 12597 9355 12631
rect 12633 12597 12667 12631
rect 15761 12597 15795 12631
rect 5733 12393 5767 12427
rect 6469 12393 6503 12427
rect 14197 12393 14231 12427
rect 17877 12393 17911 12427
rect 18429 12325 18463 12359
rect 2881 12257 2915 12291
rect 3801 12257 3835 12291
rect 7389 12257 7423 12291
rect 7481 12257 7515 12291
rect 15485 12257 15519 12291
rect 18521 12257 18555 12291
rect 20545 12257 20579 12291
rect 21005 12257 21039 12291
rect 1409 12189 1443 12223
rect 2513 12189 2547 12223
rect 2697 12189 2731 12223
rect 2789 12189 2823 12223
rect 3065 12189 3099 12223
rect 5641 12189 5675 12223
rect 6561 12189 6595 12223
rect 7113 12189 7147 12223
rect 7297 12189 7331 12223
rect 7665 12189 7699 12223
rect 10333 12189 10367 12223
rect 10977 12189 11011 12223
rect 14841 12189 14875 12223
rect 15761 12189 15795 12223
rect 18002 12189 18036 12223
rect 19441 12189 19475 12223
rect 19625 12189 19659 12223
rect 20453 12189 20487 12223
rect 20729 12189 20763 12223
rect 20821 12189 20855 12223
rect 21465 12189 21499 12223
rect 3249 12121 3283 12155
rect 4046 12121 4080 12155
rect 7849 12121 7883 12155
rect 10066 12121 10100 12155
rect 11244 12121 11278 12155
rect 14289 12121 14323 12155
rect 21649 12121 21683 12155
rect 1593 12053 1627 12087
rect 5181 12053 5215 12087
rect 8953 12053 8987 12087
rect 12357 12053 12391 12087
rect 14933 12053 14967 12087
rect 18061 12053 18095 12087
rect 19809 12053 19843 12087
rect 21833 12053 21867 12087
rect 3341 11849 3375 11883
rect 4813 11849 4847 11883
rect 5733 11849 5767 11883
rect 8861 11849 8895 11883
rect 10977 11849 11011 11883
rect 13645 11849 13679 11883
rect 17785 11849 17819 11883
rect 17969 11849 18003 11883
rect 20637 11849 20671 11883
rect 4721 11781 4755 11815
rect 12532 11781 12566 11815
rect 19073 11781 19107 11815
rect 19257 11781 19291 11815
rect 1409 11713 1443 11747
rect 2605 11713 2639 11747
rect 2789 11713 2823 11747
rect 2973 11713 3007 11747
rect 3157 11713 3191 11747
rect 5641 11713 5675 11747
rect 7205 11713 7239 11747
rect 7389 11713 7423 11747
rect 7481 11713 7515 11747
rect 7757 11713 7791 11747
rect 8677 11713 8711 11747
rect 8999 11713 9033 11747
rect 9321 11713 9355 11747
rect 10241 11713 10275 11747
rect 10425 11713 10459 11747
rect 10517 11713 10551 11747
rect 10793 11713 10827 11747
rect 12265 11713 12299 11747
rect 14105 11713 14139 11747
rect 14372 11713 14406 11747
rect 15945 11713 15979 11747
rect 16681 11713 16715 11747
rect 17910 11713 17944 11747
rect 18337 11713 18371 11747
rect 19901 11713 19935 11747
rect 20085 11713 20119 11747
rect 20453 11713 20487 11747
rect 22201 11713 22235 11747
rect 2881 11645 2915 11679
rect 7573 11645 7607 11679
rect 10609 11645 10643 11679
rect 18429 11645 18463 11679
rect 20177 11645 20211 11679
rect 20269 11645 20303 11679
rect 22477 11645 22511 11679
rect 16037 11577 16071 11611
rect 1593 11509 1627 11543
rect 7941 11509 7975 11543
rect 9091 11509 9125 11543
rect 15485 11509 15519 11543
rect 16773 11509 16807 11543
rect 19441 11509 19475 11543
rect 8401 11305 8435 11339
rect 17877 11305 17911 11339
rect 18429 11305 18463 11339
rect 19901 11305 19935 11339
rect 21189 11305 21223 11339
rect 2789 11237 2823 11271
rect 15485 11237 15519 11271
rect 4169 11169 4203 11203
rect 5457 11169 5491 11203
rect 7021 11169 7055 11203
rect 9137 11169 9171 11203
rect 13185 11169 13219 11203
rect 14105 11169 14139 11203
rect 16313 11169 16347 11203
rect 17509 11169 17543 11203
rect 20361 11169 20395 11203
rect 1409 11101 1443 11135
rect 3801 11101 3835 11135
rect 3985 11101 4019 11135
rect 4077 11101 4111 11135
rect 4353 11101 4387 11135
rect 5549 11101 5583 11135
rect 5677 11101 5711 11135
rect 7288 11101 7322 11135
rect 9413 11101 9447 11135
rect 10149 11101 10183 11135
rect 12817 11101 12851 11135
rect 13001 11101 13035 11135
rect 13093 11101 13127 11135
rect 13369 11101 13403 11135
rect 15945 11101 15979 11135
rect 16129 11101 16163 11135
rect 16221 11101 16255 11135
rect 16497 11101 16531 11135
rect 16681 11101 16715 11135
rect 17141 11101 17175 11135
rect 17325 11101 17359 11135
rect 17417 11101 17451 11135
rect 17693 11101 17727 11135
rect 18521 11101 18555 11135
rect 20085 11101 20119 11135
rect 20269 11101 20303 11135
rect 20453 11101 20487 11135
rect 20637 11101 20671 11135
rect 21281 11101 21315 11135
rect 29837 11101 29871 11135
rect 1676 11033 1710 11067
rect 5273 11033 5307 11067
rect 5457 11033 5491 11067
rect 10416 11033 10450 11067
rect 13553 11033 13587 11067
rect 14350 11033 14384 11067
rect 4537 10965 4571 10999
rect 11529 10965 11563 10999
rect 30021 10965 30055 10999
rect 10701 10761 10735 10795
rect 13737 10761 13771 10795
rect 18061 10761 18095 10795
rect 20545 10761 20579 10795
rect 21097 10761 21131 10795
rect 2145 10693 2179 10727
rect 3056 10693 3090 10727
rect 5365 10693 5399 10727
rect 5549 10693 5583 10727
rect 5641 10693 5675 10727
rect 6837 10693 6871 10727
rect 15853 10693 15887 10727
rect 17417 10693 17451 10727
rect 1409 10625 1443 10659
rect 1593 10625 1627 10659
rect 1685 10625 1719 10659
rect 1961 10625 1995 10659
rect 2789 10625 2823 10659
rect 5769 10625 5803 10659
rect 6433 10625 6467 10659
rect 6561 10625 6595 10659
rect 6653 10625 6687 10659
rect 8217 10625 8251 10659
rect 8953 10625 8987 10659
rect 9965 10625 9999 10659
rect 10149 10625 10183 10659
rect 10517 10625 10551 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 11805 10625 11839 10659
rect 12081 10625 12115 10659
rect 13001 10625 13035 10659
rect 13185 10625 13219 10659
rect 13553 10625 13587 10659
rect 15025 10625 15059 10659
rect 15209 10625 15243 10659
rect 15669 10625 15703 10659
rect 15945 10625 15979 10659
rect 16073 10625 16107 10659
rect 16681 10625 16715 10659
rect 16865 10625 16899 10659
rect 16957 10625 16991 10659
rect 17233 10625 17267 10659
rect 17969 10625 18003 10659
rect 18889 10625 18923 10659
rect 19809 10625 19843 10659
rect 19993 10625 20027 10659
rect 20361 10625 20395 10659
rect 21189 10625 21223 10659
rect 1777 10557 1811 10591
rect 5365 10557 5399 10591
rect 10241 10557 10275 10591
rect 10333 10557 10367 10591
rect 11897 10557 11931 10591
rect 13277 10557 13311 10591
rect 13369 10557 13403 10591
rect 15761 10557 15795 10591
rect 17049 10557 17083 10591
rect 19349 10557 19383 10591
rect 20085 10557 20119 10591
rect 20177 10557 20211 10591
rect 4169 10489 4203 10523
rect 6837 10489 6871 10523
rect 8769 10489 8803 10523
rect 8125 10421 8159 10455
rect 12265 10421 12299 10455
rect 19073 10421 19107 10455
rect 9229 10217 9263 10251
rect 10333 10217 10367 10251
rect 16221 10217 16255 10251
rect 20453 10217 20487 10251
rect 2881 10149 2915 10183
rect 12633 10149 12667 10183
rect 14473 10081 14507 10115
rect 1685 10013 1719 10047
rect 1869 10013 1903 10047
rect 1955 10013 1989 10047
rect 2099 10013 2133 10047
rect 2237 10013 2271 10047
rect 3065 10013 3099 10047
rect 3893 10013 3927 10047
rect 5917 10013 5951 10047
rect 6101 10013 6135 10047
rect 6193 10013 6227 10047
rect 6285 10013 6319 10047
rect 6469 10013 6503 10047
rect 7113 10013 7147 10047
rect 7849 10013 7883 10047
rect 11253 10013 11287 10047
rect 14105 10013 14139 10047
rect 14289 10013 14323 10047
rect 14381 10013 14415 10047
rect 14657 10013 14691 10047
rect 16589 10081 16623 10115
rect 17417 10081 17451 10115
rect 18521 10081 18555 10115
rect 16497 10013 16531 10047
rect 16717 10013 16751 10047
rect 17289 10013 17323 10047
rect 17693 10013 17727 10047
rect 18337 10013 18371 10047
rect 18613 10013 18647 10047
rect 20361 10013 20395 10047
rect 21281 10013 21315 10047
rect 4160 9945 4194 9979
rect 6929 9945 6963 9979
rect 7665 9945 7699 9979
rect 9413 9945 9447 9979
rect 9597 9945 9631 9979
rect 10057 9945 10091 9979
rect 10241 9945 10275 9979
rect 11520 9945 11554 9979
rect 13185 9945 13219 9979
rect 13369 9945 13403 9979
rect 15393 9945 15427 9979
rect 15577 9945 15611 9979
rect 16221 9945 16255 9979
rect 16313 9945 16347 9979
rect 16589 9945 16623 9979
rect 17417 9945 17451 9979
rect 17509 9945 17543 9979
rect 21526 9945 21560 9979
rect 2421 9877 2455 9911
rect 5273 9877 5307 9911
rect 5733 9877 5767 9911
rect 14841 9877 14875 9911
rect 18153 9877 18187 9911
rect 22661 9877 22695 9911
rect 3525 9673 3559 9707
rect 17325 9673 17359 9707
rect 19257 9673 19291 9707
rect 19809 9673 19843 9707
rect 2412 9605 2446 9639
rect 6745 9605 6779 9639
rect 6837 9605 6871 9639
rect 7665 9605 7699 9639
rect 10701 9605 10735 9639
rect 10885 9605 10919 9639
rect 16037 9605 16071 9639
rect 18144 9605 18178 9639
rect 1409 9537 1443 9571
rect 4077 9537 4111 9571
rect 4261 9537 4295 9571
rect 4629 9537 4663 9571
rect 5641 9537 5675 9571
rect 6617 9537 6651 9571
rect 7021 9537 7055 9571
rect 11529 9537 11563 9571
rect 12449 9537 12483 9571
rect 13461 9537 13495 9571
rect 14749 9537 14783 9571
rect 14933 9537 14967 9571
rect 15117 9537 15151 9571
rect 15301 9537 15335 9571
rect 15945 9537 15979 9571
rect 17233 9537 17267 9571
rect 19717 9537 19751 9571
rect 2145 9469 2179 9503
rect 4353 9469 4387 9503
rect 4445 9469 4479 9503
rect 8217 9469 8251 9503
rect 8493 9469 8527 9503
rect 12173 9469 12207 9503
rect 13737 9469 13771 9503
rect 15025 9469 15059 9503
rect 17877 9469 17911 9503
rect 5457 9401 5491 9435
rect 7021 9401 7055 9435
rect 1593 9333 1627 9367
rect 4813 9333 4847 9367
rect 7573 9333 7607 9367
rect 9597 9333 9631 9367
rect 11621 9333 11655 9367
rect 15485 9333 15519 9367
rect 6469 9129 6503 9163
rect 9689 9129 9723 9163
rect 10241 9129 10275 9163
rect 17141 9129 17175 9163
rect 19809 9129 19843 9163
rect 21097 9129 21131 9163
rect 15577 9061 15611 9095
rect 2881 8993 2915 9027
rect 3801 8993 3835 9027
rect 5089 8993 5123 9027
rect 9229 8993 9263 9027
rect 10885 8993 10919 9027
rect 20637 8993 20671 9027
rect 21557 8993 21591 9027
rect 1409 8925 1443 8959
rect 2605 8925 2639 8959
rect 4077 8925 4111 8959
rect 5356 8925 5390 8959
rect 8309 8925 8343 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9321 8925 9355 8959
rect 9505 8925 9539 8959
rect 10609 8925 10643 8959
rect 11621 8925 11655 8959
rect 13286 8925 13320 8959
rect 13553 8925 13587 8959
rect 14197 8925 14231 8959
rect 16405 8925 16439 8959
rect 17049 8925 17083 8959
rect 17785 8925 17819 8959
rect 17969 8923 18003 8957
rect 18055 8925 18089 8959
rect 18199 8925 18233 8959
rect 18337 8925 18371 8959
rect 19717 8925 19751 8959
rect 20361 8925 20395 8959
rect 20545 8925 20579 8959
rect 20729 8925 20763 8959
rect 20913 8925 20947 8959
rect 29837 8925 29871 8959
rect 8042 8857 8076 8891
rect 14464 8857 14498 8891
rect 21824 8857 21858 8891
rect 1593 8789 1627 8823
rect 6929 8789 6963 8823
rect 10701 8789 10735 8823
rect 11529 8789 11563 8823
rect 12173 8789 12207 8823
rect 16313 8789 16347 8823
rect 18521 8789 18555 8823
rect 22937 8789 22971 8823
rect 30021 8789 30055 8823
rect 3065 8585 3099 8619
rect 3617 8585 3651 8619
rect 5641 8585 5675 8619
rect 10793 8585 10827 8619
rect 11529 8585 11563 8619
rect 19809 8585 19843 8619
rect 21833 8585 21867 8619
rect 30021 8585 30055 8619
rect 6377 8517 6411 8551
rect 10885 8517 10919 8551
rect 1685 8449 1719 8483
rect 1952 8449 1986 8483
rect 3801 8449 3835 8483
rect 4261 8449 4295 8483
rect 4528 8449 4562 8483
rect 8309 8449 8343 8483
rect 9965 8449 9999 8483
rect 10241 8449 10275 8483
rect 11897 8449 11931 8483
rect 13093 8449 13127 8483
rect 14381 8449 14415 8483
rect 14648 8449 14682 8483
rect 17141 8449 17175 8483
rect 17417 8449 17451 8483
rect 18429 8449 18463 8483
rect 18705 8449 18739 8483
rect 20729 8449 20763 8483
rect 21097 8449 21131 8483
rect 21281 8449 21315 8483
rect 22017 8449 22051 8483
rect 22201 8449 22235 8483
rect 22385 8449 22419 8483
rect 22569 8449 22603 8483
rect 29929 8449 29963 8483
rect 30113 8449 30147 8483
rect 6377 8381 6411 8415
rect 6469 8381 6503 8415
rect 6745 8381 6779 8415
rect 8585 8381 8619 8415
rect 10149 8381 10183 8415
rect 11989 8381 12023 8415
rect 12081 8381 12115 8415
rect 13369 8381 13403 8415
rect 20913 8381 20947 8415
rect 21005 8381 21039 8415
rect 22293 8381 22327 8415
rect 9781 8313 9815 8347
rect 15761 8313 15795 8347
rect 10149 8245 10183 8279
rect 20545 8245 20579 8279
rect 2237 8041 2271 8075
rect 5089 8041 5123 8075
rect 7297 8041 7331 8075
rect 9505 8041 9539 8075
rect 10057 8041 10091 8075
rect 10517 8041 10551 8075
rect 12265 8041 12299 8075
rect 12909 8041 12943 8075
rect 17417 8041 17451 8075
rect 21281 8041 21315 8075
rect 18521 7973 18555 8007
rect 1869 7905 1903 7939
rect 4077 7905 4111 7939
rect 6929 7905 6963 7939
rect 9413 7905 9447 7939
rect 11713 7905 11747 7939
rect 14197 7905 14231 7939
rect 15117 7905 15151 7939
rect 1501 7837 1535 7871
rect 1685 7837 1719 7871
rect 1777 7837 1811 7871
rect 2053 7837 2087 7871
rect 3801 7837 3835 7871
rect 5273 7837 5307 7871
rect 5457 7837 5491 7871
rect 5549 7837 5583 7871
rect 5641 7837 5675 7871
rect 5825 7837 5859 7871
rect 6561 7837 6595 7871
rect 6745 7837 6779 7871
rect 6837 7837 6871 7871
rect 7113 7837 7147 7871
rect 9505 7837 9539 7871
rect 10241 7837 10275 7871
rect 10333 7837 10367 7871
rect 12725 7837 12759 7871
rect 12909 7837 12943 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 14841 7839 14875 7873
rect 15025 7837 15059 7871
rect 15209 7837 15243 7871
rect 15393 7837 15427 7871
rect 16037 7837 16071 7871
rect 19901 7837 19935 7871
rect 20168 7837 20202 7871
rect 7849 7769 7883 7803
rect 8033 7769 8067 7803
rect 10517 7769 10551 7803
rect 15577 7769 15611 7803
rect 16282 7769 16316 7803
rect 18337 7769 18371 7803
rect 9137 7701 9171 7735
rect 11805 7701 11839 7735
rect 11897 7701 11931 7735
rect 2237 7497 2271 7531
rect 6469 7497 6503 7531
rect 10149 7497 10183 7531
rect 12173 7497 12207 7531
rect 14749 7497 14783 7531
rect 17969 7497 18003 7531
rect 23213 7497 23247 7531
rect 2789 7429 2823 7463
rect 2973 7429 3007 7463
rect 5641 7429 5675 7463
rect 5825 7429 5859 7463
rect 10517 7429 10551 7463
rect 11621 7429 11655 7463
rect 17325 7429 17359 7463
rect 19993 7429 20027 7463
rect 21281 7429 21315 7463
rect 22078 7429 22112 7463
rect 1409 7361 1443 7395
rect 2053 7361 2087 7395
rect 4537 7361 4571 7395
rect 6561 7361 6595 7395
rect 7021 7361 7055 7395
rect 7205 7361 7239 7395
rect 7573 7361 7607 7395
rect 8493 7361 8527 7395
rect 8677 7361 8711 7395
rect 9045 7361 9079 7395
rect 10333 7361 10367 7395
rect 11529 7361 11563 7395
rect 11713 7361 11747 7395
rect 12541 7361 12575 7395
rect 13185 7361 13219 7395
rect 14013 7361 14047 7395
rect 14197 7361 14231 7395
rect 14289 7361 14323 7395
rect 14565 7361 14599 7395
rect 15209 7361 15243 7395
rect 15393 7361 15427 7395
rect 15485 7361 15519 7395
rect 15761 7361 15795 7395
rect 19082 7361 19116 7395
rect 20545 7361 20579 7395
rect 20729 7361 20763 7395
rect 20913 7361 20947 7395
rect 21097 7361 21131 7395
rect 21833 7361 21867 7395
rect 29837 7361 29871 7395
rect 4261 7293 4295 7327
rect 7297 7293 7331 7327
rect 7389 7293 7423 7327
rect 8769 7293 8803 7327
rect 8861 7293 8895 7327
rect 12449 7293 12483 7327
rect 13461 7293 13495 7327
rect 14381 7293 14415 7327
rect 15577 7293 15611 7327
rect 19349 7293 19383 7327
rect 20821 7293 20855 7327
rect 1593 7225 1627 7259
rect 17509 7225 17543 7259
rect 7757 7157 7791 7191
rect 9229 7157 9263 7191
rect 12541 7157 12575 7191
rect 13001 7157 13035 7191
rect 13369 7157 13403 7191
rect 15945 7157 15979 7191
rect 19901 7157 19935 7191
rect 30021 7157 30055 7191
rect 6561 6953 6595 6987
rect 7021 6953 7055 6987
rect 11713 6953 11747 6987
rect 12817 6885 12851 6919
rect 18061 6885 18095 6919
rect 1777 6817 1811 6851
rect 12081 6817 12115 6851
rect 13461 6817 13495 6851
rect 15025 6817 15059 6851
rect 16865 6817 16899 6851
rect 19533 6817 19567 6851
rect 1409 6749 1443 6783
rect 1593 6749 1627 6783
rect 1685 6749 1719 6783
rect 1961 6749 1995 6783
rect 2605 6749 2639 6783
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 4261 6749 4295 6783
rect 4353 6749 4387 6783
rect 4537 6749 4571 6783
rect 5733 6749 5767 6783
rect 6009 6749 6043 6783
rect 6377 6749 6411 6783
rect 6561 6749 6595 6783
rect 8134 6749 8168 6783
rect 8401 6749 8435 6783
rect 10057 6749 10091 6783
rect 10333 6749 10367 6783
rect 10977 6749 11011 6783
rect 11897 6749 11931 6783
rect 12173 6749 12207 6783
rect 13185 6749 13219 6783
rect 15301 6749 15335 6783
rect 15945 6749 15979 6783
rect 16497 6749 16531 6783
rect 16681 6749 16715 6783
rect 16782 6749 16816 6783
rect 17049 6749 17083 6783
rect 19441 6749 19475 6783
rect 20085 6749 20119 6783
rect 5181 6681 5215 6715
rect 13277 6681 13311 6715
rect 17877 6681 17911 6715
rect 20352 6681 20386 6715
rect 2145 6613 2179 6647
rect 2789 6613 2823 6647
rect 3801 6613 3835 6647
rect 5089 6613 5123 6647
rect 10885 6613 10919 6647
rect 15761 6613 15795 6647
rect 17233 6613 17267 6647
rect 21465 6613 21499 6647
rect 2881 6409 2915 6443
rect 8953 6409 8987 6443
rect 9689 6409 9723 6443
rect 1768 6341 1802 6375
rect 10425 6341 10459 6375
rect 10793 6341 10827 6375
rect 1501 6273 1535 6307
rect 3341 6273 3375 6307
rect 3525 6273 3559 6307
rect 3893 6273 3927 6307
rect 5089 6273 5123 6307
rect 5273 6273 5307 6307
rect 5641 6273 5675 6307
rect 5825 6273 5859 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 6745 6273 6779 6307
rect 6929 6273 6963 6307
rect 7573 6273 7607 6307
rect 7840 6273 7874 6307
rect 10057 6273 10091 6307
rect 10517 6273 10551 6307
rect 12449 6273 12483 6307
rect 13277 6273 13311 6307
rect 13461 6273 13495 6307
rect 13737 6273 13771 6307
rect 14289 6273 14323 6307
rect 14556 6273 14590 6307
rect 17794 6273 17828 6307
rect 18061 6273 18095 6307
rect 18705 6273 18739 6307
rect 19625 6273 19659 6307
rect 19901 6273 19935 6307
rect 3617 6205 3651 6239
rect 3709 6205 3743 6239
rect 6653 6205 6687 6239
rect 12173 6205 12207 6239
rect 12357 6205 12391 6239
rect 18521 6205 18555 6239
rect 5641 6137 5675 6171
rect 9505 6137 9539 6171
rect 12817 6137 12851 6171
rect 15669 6137 15703 6171
rect 16681 6137 16715 6171
rect 4077 6069 4111 6103
rect 7113 6069 7147 6103
rect 13645 6069 13679 6103
rect 3249 5865 3283 5899
rect 9413 5865 9447 5899
rect 10793 5865 10827 5899
rect 13461 5865 13495 5899
rect 16957 5865 16991 5899
rect 18245 5865 18279 5899
rect 20729 5865 20763 5899
rect 5549 5797 5583 5831
rect 6469 5797 6503 5831
rect 19257 5797 19291 5831
rect 1869 5729 1903 5763
rect 4169 5729 4203 5763
rect 11437 5729 11471 5763
rect 12817 5729 12851 5763
rect 13001 5729 13035 5763
rect 14381 5729 14415 5763
rect 17877 5729 17911 5763
rect 20269 5729 20303 5763
rect 20361 5729 20395 5763
rect 4436 5661 4470 5695
rect 6009 5661 6043 5695
rect 6285 5661 6319 5695
rect 6653 5661 6687 5695
rect 6837 5661 6871 5695
rect 9505 5661 9539 5695
rect 11989 5661 12023 5695
rect 14105 5661 14139 5695
rect 15577 5661 15611 5695
rect 17509 5661 17543 5695
rect 17693 5661 17727 5695
rect 17785 5661 17819 5695
rect 18061 5661 18095 5695
rect 19441 5661 19475 5695
rect 19993 5661 20027 5695
rect 20177 5661 20211 5695
rect 20545 5661 20579 5695
rect 2136 5593 2170 5627
rect 11161 5593 11195 5627
rect 12081 5593 12115 5627
rect 15822 5593 15856 5627
rect 11253 5525 11287 5559
rect 13093 5525 13127 5559
rect 4997 5321 5031 5355
rect 11529 5321 11563 5355
rect 13277 5321 13311 5355
rect 14933 5321 14967 5355
rect 19901 5321 19935 5355
rect 1685 5185 1719 5219
rect 3617 5185 3651 5219
rect 3884 5185 3918 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 6929 5185 6963 5219
rect 7021 5185 7055 5219
rect 8401 5185 8435 5219
rect 8585 5185 8619 5219
rect 8769 5185 8803 5219
rect 8953 5185 8987 5219
rect 10793 5185 10827 5219
rect 11713 5185 11747 5219
rect 13093 5185 13127 5219
rect 13921 5185 13955 5219
rect 15117 5185 15151 5219
rect 15393 5185 15427 5219
rect 15485 5185 15519 5219
rect 15669 5185 15703 5219
rect 16865 5185 16899 5219
rect 18061 5185 18095 5219
rect 21014 5185 21048 5219
rect 21281 5185 21315 5219
rect 29837 5185 29871 5219
rect 1409 5117 1443 5151
rect 8677 5117 8711 5151
rect 11989 5117 12023 5151
rect 12817 5117 12851 5151
rect 15301 5117 15335 5151
rect 17785 5117 17819 5151
rect 6377 5049 6411 5083
rect 10977 5049 11011 5083
rect 13737 5049 13771 5083
rect 9137 4981 9171 5015
rect 11897 4981 11931 5015
rect 12909 4981 12943 5015
rect 16681 4981 16715 5015
rect 17877 4981 17911 5015
rect 18245 4981 18279 5015
rect 30021 4981 30055 5015
rect 6561 4777 6595 4811
rect 11253 4777 11287 4811
rect 14105 4777 14139 4811
rect 15301 4777 15335 4811
rect 19349 4777 19383 4811
rect 20637 4777 20671 4811
rect 12449 4709 12483 4743
rect 1409 4641 1443 4675
rect 1685 4641 1719 4675
rect 5733 4641 5767 4675
rect 7941 4641 7975 4675
rect 9321 4641 9355 4675
rect 13553 4641 13587 4675
rect 14565 4641 14599 4675
rect 14749 4641 14783 4675
rect 15853 4641 15887 4675
rect 16865 4641 16899 4675
rect 18245 4641 18279 4675
rect 18337 4641 18371 4675
rect 5549 4573 5583 4607
rect 5825 4573 5859 4607
rect 5917 4573 5951 4607
rect 6101 4573 6135 4607
rect 8953 4573 8987 4607
rect 9137 4573 9171 4607
rect 9229 4573 9263 4607
rect 9505 4573 9539 4607
rect 10609 4573 10643 4607
rect 10701 4573 10735 4607
rect 12541 4573 12575 4607
rect 13369 4573 13403 4607
rect 16681 4573 16715 4607
rect 16957 4573 16991 4607
rect 17969 4573 18003 4607
rect 18153 4573 18187 4607
rect 18521 4573 18555 4607
rect 19441 4573 19475 4607
rect 19901 4573 19935 4607
rect 20085 4573 20119 4607
rect 20177 4573 20211 4607
rect 20269 4573 20303 4607
rect 20453 4573 20487 4607
rect 30113 4573 30147 4607
rect 30941 4573 30975 4607
rect 7674 4505 7708 4539
rect 11437 4505 11471 4539
rect 11621 4505 11655 4539
rect 12265 4505 12299 4539
rect 14473 4505 14507 4539
rect 18705 4505 18739 4539
rect 5365 4437 5399 4471
rect 9689 4437 9723 4471
rect 12541 4437 12575 4471
rect 15669 4437 15703 4471
rect 15761 4437 15795 4471
rect 16497 4437 16531 4471
rect 29929 4437 29963 4471
rect 7113 4233 7147 4267
rect 9689 4233 9723 4267
rect 15577 4233 15611 4267
rect 16681 4233 16715 4267
rect 18337 4233 18371 4267
rect 1869 4165 1903 4199
rect 8576 4165 8610 4199
rect 17049 4165 17083 4199
rect 2789 4097 2823 4131
rect 3617 4097 3651 4131
rect 5181 4097 5215 4131
rect 5365 4097 5399 4131
rect 5549 4097 5583 4131
rect 5733 4097 5767 4131
rect 6377 4097 6411 4131
rect 6561 4097 6595 4131
rect 6653 4097 6687 4131
rect 6745 4097 6779 4131
rect 6929 4097 6963 4131
rect 8309 4097 8343 4131
rect 10149 4097 10183 4131
rect 10333 4097 10367 4131
rect 10425 4097 10459 4131
rect 10701 4097 10735 4131
rect 11989 4097 12023 4131
rect 13829 4097 13863 4131
rect 14289 4097 14323 4131
rect 15761 4097 15795 4131
rect 15945 4097 15979 4131
rect 16037 4097 16071 4131
rect 17141 4097 17175 4131
rect 19450 4097 19484 4131
rect 19717 4097 19751 4131
rect 20177 4097 20211 4131
rect 20361 4097 20395 4131
rect 20729 4097 20763 4131
rect 22017 4097 22051 4131
rect 29285 4097 29319 4131
rect 30113 4097 30147 4131
rect 5457 4029 5491 4063
rect 10517 4029 10551 4063
rect 11897 4029 11931 4063
rect 13553 4029 13587 4063
rect 14565 4029 14599 4063
rect 17233 4029 17267 4063
rect 20453 4029 20487 4063
rect 20545 4029 20579 4063
rect 3065 3961 3099 3995
rect 3801 3961 3835 3995
rect 11621 3961 11655 3995
rect 21833 3961 21867 3995
rect 2145 3893 2179 3927
rect 4997 3893 5031 3927
rect 10885 3893 10919 3927
rect 11989 3893 12023 3927
rect 20913 3893 20947 3927
rect 29469 3893 29503 3927
rect 29929 3893 29963 3927
rect 1593 3689 1627 3723
rect 2421 3689 2455 3723
rect 4445 3689 4479 3723
rect 6653 3689 6687 3723
rect 10793 3689 10827 3723
rect 11437 3689 11471 3723
rect 13185 3689 13219 3723
rect 15577 3689 15611 3723
rect 16773 3689 16807 3723
rect 17969 3689 18003 3723
rect 19257 3689 19291 3723
rect 21281 3689 21315 3723
rect 22845 3689 22879 3723
rect 11621 3621 11655 3655
rect 5273 3553 5307 3587
rect 9413 3553 9447 3587
rect 14105 3553 14139 3587
rect 14381 3553 14415 3587
rect 16129 3553 16163 3587
rect 17417 3553 17451 3587
rect 18521 3553 18555 3587
rect 20637 3553 20671 3587
rect 21465 3553 21499 3587
rect 1409 3485 1443 3519
rect 2513 3485 2547 3519
rect 5540 3485 5574 3519
rect 9680 3485 9714 3519
rect 11253 3485 11287 3519
rect 11345 3485 11379 3519
rect 12081 3485 12115 3519
rect 12541 3485 12575 3519
rect 12909 3485 12943 3519
rect 15945 3485 15979 3519
rect 20381 3485 20415 3519
rect 21281 3485 21315 3519
rect 22385 3485 22419 3519
rect 23029 3485 23063 3519
rect 28089 3485 28123 3519
rect 28825 3485 28859 3519
rect 29745 3485 29779 3519
rect 2697 3417 2731 3451
rect 4353 3417 4387 3451
rect 16037 3417 16071 3451
rect 18429 3417 18463 3451
rect 21741 3417 21775 3451
rect 17141 3349 17175 3383
rect 17233 3349 17267 3383
rect 18337 3349 18371 3383
rect 21097 3349 21131 3383
rect 22201 3349 22235 3383
rect 27905 3349 27939 3383
rect 28641 3349 28675 3383
rect 29561 3349 29595 3383
rect 3801 3145 3835 3179
rect 8677 3145 8711 3179
rect 10609 3145 10643 3179
rect 11529 3145 11563 3179
rect 14473 3145 14507 3179
rect 15853 3145 15887 3179
rect 15945 3145 15979 3179
rect 16865 3145 16899 3179
rect 17785 3145 17819 3179
rect 18153 3145 18187 3179
rect 19441 3145 19475 3179
rect 23581 3145 23615 3179
rect 27353 3145 27387 3179
rect 29377 3145 29411 3179
rect 1869 3077 1903 3111
rect 3157 3077 3191 3111
rect 4712 3077 4746 3111
rect 9496 3077 9530 3111
rect 11989 3077 12023 3111
rect 2789 3009 2823 3043
rect 3617 3009 3651 3043
rect 4445 3009 4479 3043
rect 6561 3009 6595 3043
rect 7297 3009 7331 3043
rect 7941 3009 7975 3043
rect 8585 3009 8619 3043
rect 9229 3009 9263 3043
rect 11713 3009 11747 3043
rect 12541 3009 12575 3043
rect 13001 3009 13035 3043
rect 13093 3009 13127 3043
rect 14105 3009 14139 3043
rect 15117 3009 15151 3043
rect 15393 3009 15427 3043
rect 17325 3077 17359 3111
rect 20453 3077 20487 3111
rect 27813 3077 27847 3111
rect 28273 3077 28307 3111
rect 28457 3077 28491 3111
rect 16129 3009 16163 3043
rect 17049 3009 17083 3043
rect 18245 3009 18279 3043
rect 19257 3009 19291 3043
rect 20269 3009 20303 3043
rect 20637 3009 20671 3043
rect 20729 3009 20763 3043
rect 22017 3009 22051 3043
rect 22109 3009 22143 3043
rect 22477 3009 22511 3043
rect 23121 3009 23155 3043
rect 23765 3009 23799 3043
rect 27537 3009 27571 3043
rect 29561 3009 29595 3043
rect 29929 3009 29963 3043
rect 30021 3009 30055 3043
rect 11897 2941 11931 2975
rect 13829 2941 13863 2975
rect 14013 2941 14047 2975
rect 15301 2941 15335 2975
rect 15853 2941 15887 2975
rect 17141 2941 17175 2975
rect 18337 2941 18371 2975
rect 18981 2941 19015 2975
rect 27629 2941 27663 2975
rect 5825 2873 5859 2907
rect 6745 2873 6779 2907
rect 7481 2873 7515 2907
rect 14933 2873 14967 2907
rect 20269 2873 20303 2907
rect 2145 2805 2179 2839
rect 8125 2805 8159 2839
rect 11713 2805 11747 2839
rect 15209 2805 15243 2839
rect 17325 2805 17359 2839
rect 19073 2805 19107 2839
rect 20453 2805 20487 2839
rect 20913 2805 20947 2839
rect 21833 2805 21867 2839
rect 22293 2805 22327 2839
rect 22937 2805 22971 2839
rect 27813 2805 27847 2839
rect 28641 2805 28675 2839
rect 29653 2805 29687 2839
rect 30941 2805 30975 2839
rect 2881 2601 2915 2635
rect 4445 2601 4479 2635
rect 7665 2601 7699 2635
rect 9137 2601 9171 2635
rect 14105 2601 14139 2635
rect 15025 2601 15059 2635
rect 15945 2601 15979 2635
rect 17601 2601 17635 2635
rect 18521 2601 18555 2635
rect 20453 2601 20487 2635
rect 21097 2601 21131 2635
rect 21925 2601 21959 2635
rect 25697 2601 25731 2635
rect 27169 2601 27203 2635
rect 27629 2601 27663 2635
rect 30021 2601 30055 2635
rect 6561 2533 6595 2567
rect 14473 2533 14507 2567
rect 16773 2533 16807 2567
rect 19257 2533 19291 2567
rect 24409 2533 24443 2567
rect 25053 2533 25087 2567
rect 2237 2465 2271 2499
rect 8401 2465 8435 2499
rect 9873 2465 9907 2499
rect 11805 2465 11839 2499
rect 14565 2465 14599 2499
rect 15485 2465 15519 2499
rect 16681 2465 16715 2499
rect 17141 2465 17175 2499
rect 20361 2465 20395 2499
rect 21189 2465 21223 2499
rect 1961 2397 1995 2431
rect 3065 2397 3099 2431
rect 4997 2397 5031 2431
rect 5273 2397 5307 2431
rect 6377 2397 6411 2431
rect 7481 2397 7515 2431
rect 8953 2397 8987 2431
rect 9597 2397 9631 2431
rect 11529 2397 11563 2431
rect 13369 2397 13403 2431
rect 14289 2397 14323 2431
rect 15209 2397 15243 2431
rect 15393 2397 15427 2431
rect 16129 2397 16163 2431
rect 16957 2397 16991 2431
rect 17785 2397 17819 2431
rect 17969 2397 18003 2431
rect 18061 2397 18095 2431
rect 18705 2397 18739 2431
rect 19441 2397 19475 2431
rect 20453 2397 20487 2431
rect 21281 2397 21315 2431
rect 22845 2397 22879 2431
rect 23489 2397 23523 2431
rect 24593 2397 24627 2431
rect 25237 2397 25271 2431
rect 25881 2397 25915 2431
rect 26985 2397 27019 2431
rect 27813 2397 27847 2431
rect 28733 2397 28767 2431
rect 29837 2397 29871 2431
rect 4169 2329 4203 2363
rect 8217 2329 8251 2363
rect 13553 2329 13587 2363
rect 22017 2329 22051 2363
rect 22201 2329 22235 2363
rect 20085 2261 20119 2295
rect 20913 2261 20947 2295
rect 22661 2261 22695 2295
rect 23305 2261 23339 2295
rect 28917 2261 28951 2295
<< metal1 >>
rect 1104 45722 30820 45744
rect 1104 45670 10880 45722
rect 10932 45670 10944 45722
rect 10996 45670 11008 45722
rect 11060 45670 11072 45722
rect 11124 45670 11136 45722
rect 11188 45670 20811 45722
rect 20863 45670 20875 45722
rect 20927 45670 20939 45722
rect 20991 45670 21003 45722
rect 21055 45670 21067 45722
rect 21119 45670 30820 45722
rect 1104 45648 30820 45670
rect 7101 45611 7159 45617
rect 7101 45577 7113 45611
rect 7147 45577 7159 45611
rect 7101 45571 7159 45577
rect 7116 45540 7144 45571
rect 3160 45512 7144 45540
rect 1670 45472 1676 45484
rect 1631 45444 1676 45472
rect 1670 45432 1676 45444
rect 1728 45432 1734 45484
rect 3160 45481 3188 45512
rect 2409 45475 2467 45481
rect 2409 45441 2421 45475
rect 2455 45441 2467 45475
rect 2409 45435 2467 45441
rect 3145 45475 3203 45481
rect 3145 45441 3157 45475
rect 3191 45441 3203 45475
rect 3145 45435 3203 45441
rect 3973 45475 4031 45481
rect 3973 45441 3985 45475
rect 4019 45472 4031 45475
rect 4522 45472 4528 45484
rect 4019 45444 4528 45472
rect 4019 45441 4031 45444
rect 3973 45435 4031 45441
rect 2424 45404 2452 45435
rect 4522 45432 4528 45444
rect 4580 45432 4586 45484
rect 4617 45475 4675 45481
rect 4617 45441 4629 45475
rect 4663 45472 4675 45475
rect 4890 45472 4896 45484
rect 4663 45444 4896 45472
rect 4663 45441 4675 45444
rect 4617 45435 4675 45441
rect 4890 45432 4896 45444
rect 4948 45432 4954 45484
rect 5261 45475 5319 45481
rect 5261 45441 5273 45475
rect 5307 45472 5319 45475
rect 5442 45472 5448 45484
rect 5307 45444 5448 45472
rect 5307 45441 5319 45444
rect 5261 45435 5319 45441
rect 5442 45432 5448 45444
rect 5500 45432 5506 45484
rect 6454 45472 6460 45484
rect 6415 45444 6460 45472
rect 6454 45432 6460 45444
rect 6512 45432 6518 45484
rect 7282 45472 7288 45484
rect 7243 45444 7288 45472
rect 7282 45432 7288 45444
rect 7340 45432 7346 45484
rect 30098 45472 30104 45484
rect 30059 45444 30104 45472
rect 30098 45432 30104 45444
rect 30156 45432 30162 45484
rect 2424 45376 5120 45404
rect 2222 45336 2228 45348
rect 2183 45308 2228 45336
rect 2222 45296 2228 45308
rect 2280 45296 2286 45348
rect 2958 45336 2964 45348
rect 2919 45308 2964 45336
rect 2958 45296 2964 45308
rect 3016 45296 3022 45348
rect 5092 45345 5120 45376
rect 5077 45339 5135 45345
rect 5077 45305 5089 45339
rect 5123 45305 5135 45339
rect 5077 45299 5135 45305
rect 1489 45271 1547 45277
rect 1489 45237 1501 45271
rect 1535 45268 1547 45271
rect 2774 45268 2780 45280
rect 1535 45240 2780 45268
rect 1535 45237 1547 45240
rect 1489 45231 1547 45237
rect 2774 45228 2780 45240
rect 2832 45228 2838 45280
rect 3786 45268 3792 45280
rect 3747 45240 3792 45268
rect 3786 45228 3792 45240
rect 3844 45228 3850 45280
rect 4430 45268 4436 45280
rect 4391 45240 4436 45268
rect 4430 45228 4436 45240
rect 4488 45228 4494 45280
rect 6641 45271 6699 45277
rect 6641 45237 6653 45271
rect 6687 45268 6699 45271
rect 6730 45268 6736 45280
rect 6687 45240 6736 45268
rect 6687 45237 6699 45240
rect 6641 45231 6699 45237
rect 6730 45228 6736 45240
rect 6788 45228 6794 45280
rect 28994 45228 29000 45280
rect 29052 45268 29058 45280
rect 29917 45271 29975 45277
rect 29917 45268 29929 45271
rect 29052 45240 29929 45268
rect 29052 45228 29058 45240
rect 29917 45237 29929 45240
rect 29963 45237 29975 45271
rect 29917 45231 29975 45237
rect 1104 45178 30820 45200
rect 1104 45126 5915 45178
rect 5967 45126 5979 45178
rect 6031 45126 6043 45178
rect 6095 45126 6107 45178
rect 6159 45126 6171 45178
rect 6223 45126 15846 45178
rect 15898 45126 15910 45178
rect 15962 45126 15974 45178
rect 16026 45126 16038 45178
rect 16090 45126 16102 45178
rect 16154 45126 25776 45178
rect 25828 45126 25840 45178
rect 25892 45126 25904 45178
rect 25956 45126 25968 45178
rect 26020 45126 26032 45178
rect 26084 45126 30820 45178
rect 1104 45104 30820 45126
rect 2225 45067 2283 45073
rect 2225 45033 2237 45067
rect 2271 45064 2283 45067
rect 2866 45064 2872 45076
rect 2271 45036 2872 45064
rect 2271 45033 2283 45036
rect 2225 45027 2283 45033
rect 2866 45024 2872 45036
rect 2924 45024 2930 45076
rect 4246 45024 4252 45076
rect 4304 45064 4310 45076
rect 5077 45067 5135 45073
rect 5077 45064 5089 45067
rect 4304 45036 5089 45064
rect 4304 45024 4310 45036
rect 5077 45033 5089 45036
rect 5123 45033 5135 45067
rect 5077 45027 5135 45033
rect 5261 45067 5319 45073
rect 5261 45033 5273 45067
rect 5307 45064 5319 45067
rect 7282 45064 7288 45076
rect 5307 45036 7288 45064
rect 5307 45033 5319 45036
rect 5261 45027 5319 45033
rect 7282 45024 7288 45036
rect 7340 45024 7346 45076
rect 7374 44956 7380 45008
rect 7432 44996 7438 45008
rect 7432 44968 7604 44996
rect 7432 44956 7438 44968
rect 4430 44928 4436 44940
rect 1688 44900 4436 44928
rect 1688 44869 1716 44900
rect 4430 44888 4436 44900
rect 4488 44888 4494 44940
rect 1673 44863 1731 44869
rect 1673 44829 1685 44863
rect 1719 44829 1731 44863
rect 2406 44860 2412 44872
rect 2367 44832 2412 44860
rect 1673 44823 1731 44829
rect 2406 44820 2412 44832
rect 2464 44820 2470 44872
rect 3053 44863 3111 44869
rect 3053 44829 3065 44863
rect 3099 44860 3111 44863
rect 3142 44860 3148 44872
rect 3099 44832 3148 44860
rect 3099 44829 3111 44832
rect 3053 44823 3111 44829
rect 3142 44820 3148 44832
rect 3200 44820 3206 44872
rect 4062 44860 4068 44872
rect 4023 44832 4068 44860
rect 4062 44820 4068 44832
rect 4120 44820 4126 44872
rect 4709 44863 4767 44869
rect 4709 44829 4721 44863
rect 4755 44860 4767 44863
rect 5350 44860 5356 44872
rect 4755 44832 5356 44860
rect 4755 44829 4767 44832
rect 4709 44823 4767 44829
rect 5350 44820 5356 44832
rect 5408 44820 5414 44872
rect 5718 44860 5724 44872
rect 5679 44832 5724 44860
rect 5718 44820 5724 44832
rect 5776 44820 5782 44872
rect 6638 44820 6644 44872
rect 6696 44860 6702 44872
rect 7009 44863 7067 44869
rect 7009 44860 7021 44863
rect 6696 44832 7021 44860
rect 6696 44820 6702 44832
rect 7009 44829 7021 44832
rect 7055 44829 7067 44863
rect 7190 44860 7196 44872
rect 7151 44832 7196 44860
rect 7009 44823 7067 44829
rect 7190 44820 7196 44832
rect 7248 44820 7254 44872
rect 7285 44863 7343 44869
rect 7285 44829 7297 44863
rect 7331 44829 7343 44863
rect 7285 44823 7343 44829
rect 7377 44863 7435 44869
rect 7377 44829 7389 44863
rect 7423 44860 7435 44863
rect 7466 44860 7472 44872
rect 7423 44832 7472 44860
rect 7423 44829 7435 44832
rect 7377 44823 7435 44829
rect 1486 44724 1492 44736
rect 1447 44696 1492 44724
rect 1486 44684 1492 44696
rect 1544 44684 1550 44736
rect 2866 44724 2872 44736
rect 2827 44696 2872 44724
rect 2866 44684 2872 44696
rect 2924 44684 2930 44736
rect 4246 44724 4252 44736
rect 4207 44696 4252 44724
rect 4246 44684 4252 44696
rect 4304 44684 4310 44736
rect 5077 44727 5135 44733
rect 5077 44693 5089 44727
rect 5123 44724 5135 44727
rect 5534 44724 5540 44736
rect 5123 44696 5540 44724
rect 5123 44693 5135 44696
rect 5077 44687 5135 44693
rect 5534 44684 5540 44696
rect 5592 44684 5598 44736
rect 5810 44684 5816 44736
rect 5868 44724 5874 44736
rect 5905 44727 5963 44733
rect 5905 44724 5917 44727
rect 5868 44696 5917 44724
rect 5868 44684 5874 44696
rect 5905 44693 5917 44696
rect 5951 44693 5963 44727
rect 6822 44724 6828 44736
rect 6783 44696 6828 44724
rect 5905 44687 5963 44693
rect 6822 44684 6828 44696
rect 6880 44684 6886 44736
rect 7300 44724 7328 44823
rect 7466 44820 7472 44832
rect 7524 44820 7530 44872
rect 7576 44869 7604 44968
rect 7561 44863 7619 44869
rect 7561 44829 7573 44863
rect 7607 44829 7619 44863
rect 8202 44860 8208 44872
rect 8163 44832 8208 44860
rect 7561 44823 7619 44829
rect 8202 44820 8208 44832
rect 8260 44820 8266 44872
rect 30006 44820 30012 44872
rect 30064 44860 30070 44872
rect 30101 44863 30159 44869
rect 30101 44860 30113 44863
rect 30064 44832 30113 44860
rect 30064 44820 30070 44832
rect 30101 44829 30113 44832
rect 30147 44829 30159 44863
rect 30101 44823 30159 44829
rect 7650 44724 7656 44736
rect 7300 44696 7656 44724
rect 7650 44684 7656 44696
rect 7708 44684 7714 44736
rect 8018 44724 8024 44736
rect 7979 44696 8024 44724
rect 8018 44684 8024 44696
rect 8076 44684 8082 44736
rect 29914 44724 29920 44736
rect 29875 44696 29920 44724
rect 29914 44684 29920 44696
rect 29972 44684 29978 44736
rect 1104 44634 30820 44656
rect 1104 44582 10880 44634
rect 10932 44582 10944 44634
rect 10996 44582 11008 44634
rect 11060 44582 11072 44634
rect 11124 44582 11136 44634
rect 11188 44582 20811 44634
rect 20863 44582 20875 44634
rect 20927 44582 20939 44634
rect 20991 44582 21003 44634
rect 21055 44582 21067 44634
rect 21119 44582 30820 44634
rect 1104 44560 30820 44582
rect 4430 44520 4436 44532
rect 4391 44492 4436 44520
rect 4430 44480 4436 44492
rect 4488 44480 4494 44532
rect 4890 44520 4896 44532
rect 4851 44492 4896 44520
rect 4890 44480 4896 44492
rect 4948 44480 4954 44532
rect 5077 44523 5135 44529
rect 5077 44489 5089 44523
rect 5123 44520 5135 44523
rect 6638 44520 6644 44532
rect 5123 44492 6644 44520
rect 5123 44489 5135 44492
rect 5077 44483 5135 44489
rect 6638 44480 6644 44492
rect 6696 44520 6702 44532
rect 8113 44523 8171 44529
rect 8113 44520 8125 44523
rect 6696 44492 8125 44520
rect 6696 44480 6702 44492
rect 8113 44489 8125 44492
rect 8159 44489 8171 44523
rect 8113 44483 8171 44489
rect 3786 44452 3792 44464
rect 1688 44424 3792 44452
rect 1688 44393 1716 44424
rect 3786 44412 3792 44424
rect 3844 44412 3850 44464
rect 4249 44455 4307 44461
rect 4249 44421 4261 44455
rect 4295 44421 4307 44455
rect 4249 44415 4307 44421
rect 1673 44387 1731 44393
rect 1673 44353 1685 44387
rect 1719 44353 1731 44387
rect 2314 44384 2320 44396
rect 2275 44356 2320 44384
rect 1673 44347 1731 44353
rect 2314 44344 2320 44356
rect 2372 44344 2378 44396
rect 2958 44384 2964 44396
rect 2919 44356 2964 44384
rect 2958 44344 2964 44356
rect 3016 44344 3022 44396
rect 4264 44384 4292 44415
rect 6822 44412 6828 44464
rect 6880 44452 6886 44464
rect 6978 44455 7036 44461
rect 6978 44452 6990 44455
rect 6880 44424 6990 44452
rect 6880 44412 6886 44424
rect 6978 44421 6990 44424
rect 7024 44421 7036 44455
rect 6978 44415 7036 44421
rect 7190 44412 7196 44464
rect 7248 44452 7254 44464
rect 7248 44424 8984 44452
rect 7248 44412 7254 44424
rect 6730 44384 6736 44396
rect 4264 44356 6592 44384
rect 6691 44356 6736 44384
rect 3881 44319 3939 44325
rect 3881 44285 3893 44319
rect 3927 44316 3939 44319
rect 6564 44316 6592 44356
rect 6730 44344 6736 44356
rect 6788 44344 6794 44396
rect 8956 44393 8984 44424
rect 9137 44393 9195 44399
rect 8757 44387 8815 44393
rect 8757 44384 8769 44387
rect 6840 44356 8769 44384
rect 6840 44316 6868 44356
rect 8757 44353 8769 44356
rect 8803 44353 8815 44387
rect 8757 44347 8815 44353
rect 8941 44387 8999 44393
rect 8941 44353 8953 44387
rect 8987 44353 8999 44387
rect 9137 44359 9149 44393
rect 9183 44390 9195 44393
rect 9183 44362 9260 44390
rect 9183 44359 9195 44362
rect 9137 44353 9195 44359
rect 8941 44347 8999 44353
rect 3927 44288 5396 44316
rect 6564 44288 6868 44316
rect 3927 44285 3939 44288
rect 3881 44279 3939 44285
rect 5368 44260 5396 44288
rect 4264 44220 5120 44248
rect 4264 44192 4292 44220
rect 1486 44180 1492 44192
rect 1447 44152 1492 44180
rect 1486 44140 1492 44152
rect 1544 44140 1550 44192
rect 1762 44140 1768 44192
rect 1820 44180 1826 44192
rect 2133 44183 2191 44189
rect 2133 44180 2145 44183
rect 1820 44152 2145 44180
rect 1820 44140 1826 44152
rect 2133 44149 2145 44152
rect 2179 44149 2191 44183
rect 2133 44143 2191 44149
rect 2777 44183 2835 44189
rect 2777 44149 2789 44183
rect 2823 44180 2835 44183
rect 3050 44180 3056 44192
rect 2823 44152 3056 44180
rect 2823 44149 2835 44152
rect 2777 44143 2835 44149
rect 3050 44140 3056 44152
rect 3108 44140 3114 44192
rect 4246 44180 4252 44192
rect 4207 44152 4252 44180
rect 4246 44140 4252 44152
rect 4304 44140 4310 44192
rect 5092 44189 5120 44220
rect 5350 44208 5356 44260
rect 5408 44248 5414 44260
rect 5445 44251 5503 44257
rect 5445 44248 5457 44251
rect 5408 44220 5457 44248
rect 5408 44208 5414 44220
rect 5445 44217 5457 44220
rect 5491 44217 5503 44251
rect 8772 44248 8800 44347
rect 8846 44276 8852 44328
rect 8904 44316 8910 44328
rect 9033 44319 9091 44325
rect 9033 44316 9045 44319
rect 8904 44288 9045 44316
rect 8904 44276 8910 44288
rect 9033 44285 9045 44288
rect 9079 44285 9091 44319
rect 9232 44316 9260 44362
rect 9309 44387 9367 44393
rect 9309 44353 9321 44387
rect 9355 44384 9367 44387
rect 9858 44384 9864 44396
rect 9355 44356 9864 44384
rect 9355 44353 9367 44356
rect 9309 44347 9367 44353
rect 9858 44344 9864 44356
rect 9916 44344 9922 44396
rect 20070 44384 20076 44396
rect 16546 44356 20076 44384
rect 9490 44316 9496 44328
rect 9232 44288 9496 44316
rect 9033 44279 9091 44285
rect 9490 44276 9496 44288
rect 9548 44316 9554 44328
rect 16546 44316 16574 44356
rect 20070 44344 20076 44356
rect 20128 44344 20134 44396
rect 9548 44288 16574 44316
rect 9548 44276 9554 44288
rect 9950 44248 9956 44260
rect 8772 44220 9956 44248
rect 5445 44211 5503 44217
rect 9950 44208 9956 44220
rect 10008 44208 10014 44260
rect 5077 44183 5135 44189
rect 5077 44149 5089 44183
rect 5123 44180 5135 44183
rect 5258 44180 5264 44192
rect 5123 44152 5264 44180
rect 5123 44149 5135 44152
rect 5077 44143 5135 44149
rect 5258 44140 5264 44152
rect 5316 44140 5322 44192
rect 8570 44180 8576 44192
rect 8531 44152 8576 44180
rect 8570 44140 8576 44152
rect 8628 44140 8634 44192
rect 1104 44090 30820 44112
rect 1104 44038 5915 44090
rect 5967 44038 5979 44090
rect 6031 44038 6043 44090
rect 6095 44038 6107 44090
rect 6159 44038 6171 44090
rect 6223 44038 15846 44090
rect 15898 44038 15910 44090
rect 15962 44038 15974 44090
rect 16026 44038 16038 44090
rect 16090 44038 16102 44090
rect 16154 44038 25776 44090
rect 25828 44038 25840 44090
rect 25892 44038 25904 44090
rect 25956 44038 25968 44090
rect 26020 44038 26032 44090
rect 26084 44038 30820 44090
rect 1104 44016 30820 44038
rect 4062 43936 4068 43988
rect 4120 43976 4126 43988
rect 4982 43976 4988 43988
rect 4120 43948 4988 43976
rect 4120 43936 4126 43948
rect 4982 43936 4988 43948
rect 5040 43936 5046 43988
rect 5258 43976 5264 43988
rect 5219 43948 5264 43976
rect 5258 43936 5264 43948
rect 5316 43936 5322 43988
rect 5442 43976 5448 43988
rect 5403 43948 5448 43976
rect 5442 43936 5448 43948
rect 5500 43936 5506 43988
rect 7650 43936 7656 43988
rect 7708 43976 7714 43988
rect 8846 43976 8852 43988
rect 7708 43948 8852 43976
rect 7708 43936 7714 43948
rect 8846 43936 8852 43948
rect 8904 43936 8910 43988
rect 20070 43976 20076 43988
rect 20031 43948 20076 43976
rect 20070 43936 20076 43948
rect 20128 43936 20134 43988
rect 2317 43911 2375 43917
rect 2317 43877 2329 43911
rect 2363 43908 2375 43911
rect 3326 43908 3332 43920
rect 2363 43880 3332 43908
rect 2363 43877 2375 43880
rect 2317 43871 2375 43877
rect 3326 43868 3332 43880
rect 3384 43868 3390 43920
rect 2866 43840 2872 43852
rect 1688 43812 2872 43840
rect 1688 43781 1716 43812
rect 2866 43800 2872 43812
rect 2924 43800 2930 43852
rect 4080 43840 4108 43936
rect 8389 43911 8447 43917
rect 8389 43877 8401 43911
rect 8435 43877 8447 43911
rect 8389 43871 8447 43877
rect 2976 43812 4108 43840
rect 1673 43775 1731 43781
rect 1673 43741 1685 43775
rect 1719 43741 1731 43775
rect 1673 43735 1731 43741
rect 2133 43775 2191 43781
rect 2133 43741 2145 43775
rect 2179 43772 2191 43775
rect 2590 43772 2596 43784
rect 2179 43744 2596 43772
rect 2179 43741 2191 43744
rect 2133 43735 2191 43741
rect 2590 43732 2596 43744
rect 2648 43732 2654 43784
rect 2976 43781 3004 43812
rect 5810 43800 5816 43852
rect 5868 43840 5874 43852
rect 5905 43843 5963 43849
rect 5905 43840 5917 43843
rect 5868 43812 5917 43840
rect 5868 43800 5874 43812
rect 5905 43809 5917 43812
rect 5951 43809 5963 43843
rect 8404 43840 8432 43871
rect 8941 43843 8999 43849
rect 8941 43840 8953 43843
rect 8404 43812 8953 43840
rect 5905 43803 5963 43809
rect 8941 43809 8953 43812
rect 8987 43809 8999 43843
rect 8941 43803 8999 43809
rect 20441 43843 20499 43849
rect 20441 43809 20453 43843
rect 20487 43840 20499 43843
rect 21361 43843 21419 43849
rect 20487 43812 21312 43840
rect 20487 43809 20499 43812
rect 20441 43803 20499 43809
rect 2961 43775 3019 43781
rect 2961 43741 2973 43775
rect 3007 43741 3019 43775
rect 3970 43772 3976 43784
rect 3931 43744 3976 43772
rect 2961 43735 3019 43741
rect 3970 43732 3976 43744
rect 4028 43732 4034 43784
rect 4893 43775 4951 43781
rect 4893 43741 4905 43775
rect 4939 43772 4951 43775
rect 5350 43772 5356 43784
rect 4939 43744 5356 43772
rect 4939 43741 4951 43744
rect 4893 43735 4951 43741
rect 5350 43732 5356 43744
rect 5408 43732 5414 43784
rect 8205 43775 8263 43781
rect 8205 43741 8217 43775
rect 8251 43772 8263 43775
rect 10410 43772 10416 43784
rect 8251 43744 10416 43772
rect 8251 43741 8263 43744
rect 8205 43735 8263 43741
rect 10410 43732 10416 43744
rect 10468 43732 10474 43784
rect 20162 43732 20168 43784
rect 20220 43772 20226 43784
rect 20257 43775 20315 43781
rect 20257 43772 20269 43775
rect 20220 43744 20269 43772
rect 20220 43732 20226 43744
rect 20257 43741 20269 43744
rect 20303 43772 20315 43775
rect 21177 43775 21235 43781
rect 21177 43772 21189 43775
rect 20303 43744 21189 43772
rect 20303 43741 20315 43744
rect 20257 43735 20315 43741
rect 21177 43741 21189 43744
rect 21223 43741 21235 43775
rect 21284 43772 21312 43812
rect 21361 43809 21373 43843
rect 21407 43840 21419 43843
rect 28994 43840 29000 43852
rect 21407 43812 29000 43840
rect 21407 43809 21419 43812
rect 21361 43803 21419 43809
rect 28994 43800 29000 43812
rect 29052 43800 29058 43852
rect 29914 43772 29920 43784
rect 21284 43744 29920 43772
rect 21177 43735 21235 43741
rect 29914 43732 29920 43744
rect 29972 43732 29978 43784
rect 6172 43707 6230 43713
rect 6172 43673 6184 43707
rect 6218 43704 6230 43707
rect 6638 43704 6644 43716
rect 6218 43676 6644 43704
rect 6218 43673 6230 43676
rect 6172 43667 6230 43673
rect 6638 43664 6644 43676
rect 6696 43664 6702 43716
rect 8110 43664 8116 43716
rect 8168 43704 8174 43716
rect 9186 43707 9244 43713
rect 9186 43704 9198 43707
rect 8168 43676 9198 43704
rect 8168 43664 8174 43676
rect 9186 43673 9198 43676
rect 9232 43673 9244 43707
rect 9186 43667 9244 43673
rect 9766 43664 9772 43716
rect 9824 43704 9830 43716
rect 20993 43707 21051 43713
rect 20993 43704 21005 43707
rect 9824 43676 21005 43704
rect 9824 43664 9830 43676
rect 20993 43673 21005 43676
rect 21039 43673 21051 43707
rect 20993 43667 21051 43673
rect 1486 43636 1492 43648
rect 1447 43608 1492 43636
rect 1486 43596 1492 43608
rect 1544 43596 1550 43648
rect 2498 43596 2504 43648
rect 2556 43636 2562 43648
rect 2777 43639 2835 43645
rect 2777 43636 2789 43639
rect 2556 43608 2789 43636
rect 2556 43596 2562 43608
rect 2777 43605 2789 43608
rect 2823 43605 2835 43639
rect 3786 43636 3792 43648
rect 3747 43608 3792 43636
rect 2777 43599 2835 43605
rect 3786 43596 3792 43608
rect 3844 43596 3850 43648
rect 5261 43639 5319 43645
rect 5261 43605 5273 43639
rect 5307 43636 5319 43639
rect 6822 43636 6828 43648
rect 5307 43608 6828 43636
rect 5307 43605 5319 43608
rect 5261 43599 5319 43605
rect 6822 43596 6828 43608
rect 6880 43636 6886 43648
rect 7285 43639 7343 43645
rect 7285 43636 7297 43639
rect 6880 43608 7297 43636
rect 6880 43596 6886 43608
rect 7285 43605 7297 43608
rect 7331 43605 7343 43639
rect 7285 43599 7343 43605
rect 8018 43596 8024 43648
rect 8076 43636 8082 43648
rect 10321 43639 10379 43645
rect 10321 43636 10333 43639
rect 8076 43608 10333 43636
rect 8076 43596 8082 43608
rect 10321 43605 10333 43608
rect 10367 43605 10379 43639
rect 10321 43599 10379 43605
rect 1104 43546 30820 43568
rect 1104 43494 10880 43546
rect 10932 43494 10944 43546
rect 10996 43494 11008 43546
rect 11060 43494 11072 43546
rect 11124 43494 11136 43546
rect 11188 43494 20811 43546
rect 20863 43494 20875 43546
rect 20927 43494 20939 43546
rect 20991 43494 21003 43546
rect 21055 43494 21067 43546
rect 21119 43494 30820 43546
rect 1104 43472 30820 43494
rect 5718 43392 5724 43444
rect 5776 43432 5782 43444
rect 6365 43435 6423 43441
rect 6365 43432 6377 43435
rect 5776 43404 6377 43432
rect 5776 43392 5782 43404
rect 6365 43401 6377 43404
rect 6411 43401 6423 43435
rect 8110 43432 8116 43444
rect 8071 43404 8116 43432
rect 6365 43395 6423 43401
rect 8110 43392 8116 43404
rect 8168 43392 8174 43444
rect 9950 43432 9956 43444
rect 9911 43404 9956 43432
rect 9950 43392 9956 43404
rect 10008 43392 10014 43444
rect 10410 43432 10416 43444
rect 10371 43404 10416 43432
rect 10410 43392 10416 43404
rect 10468 43392 10474 43444
rect 5534 43324 5540 43376
rect 5592 43364 5598 43376
rect 8018 43364 8024 43376
rect 5592 43336 8024 43364
rect 5592 43324 5598 43336
rect 8018 43324 8024 43336
rect 8076 43364 8082 43376
rect 8076 43336 8169 43364
rect 8076 43324 8082 43336
rect 8570 43324 8576 43376
rect 8628 43364 8634 43376
rect 8818 43367 8876 43373
rect 8818 43364 8830 43367
rect 8628 43336 8830 43364
rect 8628 43324 8634 43336
rect 8818 43333 8830 43336
rect 8864 43333 8876 43367
rect 8818 43327 8876 43333
rect 1673 43299 1731 43305
rect 1673 43265 1685 43299
rect 1719 43265 1731 43299
rect 1673 43259 1731 43265
rect 1688 43228 1716 43259
rect 1854 43256 1860 43308
rect 1912 43296 1918 43308
rect 2317 43299 2375 43305
rect 2317 43296 2329 43299
rect 1912 43268 2329 43296
rect 1912 43256 1918 43268
rect 2317 43265 2329 43268
rect 2363 43265 2375 43299
rect 2317 43259 2375 43265
rect 2774 43256 2780 43308
rect 2832 43296 2838 43308
rect 3602 43296 3608 43308
rect 2832 43268 2877 43296
rect 3563 43268 3608 43296
rect 2832 43256 2838 43268
rect 3602 43256 3608 43268
rect 3660 43256 3666 43308
rect 3878 43256 3884 43308
rect 3936 43296 3942 43308
rect 4249 43299 4307 43305
rect 4249 43296 4261 43299
rect 3936 43268 4261 43296
rect 3936 43256 3942 43268
rect 4249 43265 4261 43268
rect 4295 43265 4307 43299
rect 4249 43259 4307 43265
rect 4338 43256 4344 43308
rect 4396 43296 4402 43308
rect 4893 43299 4951 43305
rect 4893 43296 4905 43299
rect 4396 43268 4905 43296
rect 4396 43256 4402 43268
rect 4893 43265 4905 43268
rect 4939 43265 4951 43299
rect 4893 43259 4951 43265
rect 5629 43299 5687 43305
rect 5629 43265 5641 43299
rect 5675 43296 5687 43299
rect 5718 43296 5724 43308
rect 5675 43268 5724 43296
rect 5675 43265 5687 43268
rect 5629 43259 5687 43265
rect 5718 43256 5724 43268
rect 5776 43296 5782 43308
rect 6549 43299 6607 43305
rect 6549 43296 6561 43299
rect 5776 43268 6561 43296
rect 5776 43256 5782 43268
rect 6549 43265 6561 43268
rect 6595 43265 6607 43299
rect 7374 43296 7380 43308
rect 7335 43268 7380 43296
rect 6549 43259 6607 43265
rect 7374 43256 7380 43268
rect 7432 43256 7438 43308
rect 7561 43299 7619 43305
rect 7561 43265 7573 43299
rect 7607 43296 7619 43299
rect 7929 43299 7987 43305
rect 7607 43268 7889 43296
rect 7607 43265 7619 43268
rect 7561 43259 7619 43265
rect 1688 43200 2774 43228
rect 2746 43160 2774 43200
rect 7006 43188 7012 43240
rect 7064 43228 7070 43240
rect 7650 43228 7656 43240
rect 7064 43200 7656 43228
rect 7064 43188 7070 43200
rect 7650 43188 7656 43200
rect 7708 43188 7714 43240
rect 7745 43231 7803 43237
rect 7745 43197 7757 43231
rect 7791 43197 7803 43231
rect 7861 43228 7889 43268
rect 7929 43265 7941 43299
rect 7975 43296 7987 43299
rect 8036 43296 8064 43324
rect 7975 43268 8064 43296
rect 7975 43265 7987 43268
rect 7929 43259 7987 43265
rect 9122 43256 9128 43308
rect 9180 43296 9186 43308
rect 10597 43299 10655 43305
rect 10597 43296 10609 43299
rect 9180 43268 10609 43296
rect 9180 43256 9186 43268
rect 10597 43265 10609 43268
rect 10643 43265 10655 43299
rect 30098 43296 30104 43308
rect 30059 43268 30104 43296
rect 10597 43259 10655 43265
rect 30098 43256 30104 43268
rect 30156 43256 30162 43308
rect 8018 43228 8024 43240
rect 7861 43200 8024 43228
rect 7745 43191 7803 43197
rect 4709 43163 4767 43169
rect 4709 43160 4721 43163
rect 2746 43132 4721 43160
rect 4709 43129 4721 43132
rect 4755 43129 4767 43163
rect 4709 43123 4767 43129
rect 5813 43163 5871 43169
rect 5813 43129 5825 43163
rect 5859 43160 5871 43163
rect 6454 43160 6460 43172
rect 5859 43132 6460 43160
rect 5859 43129 5871 43132
rect 5813 43123 5871 43129
rect 6454 43120 6460 43132
rect 6512 43120 6518 43172
rect 7190 43120 7196 43172
rect 7248 43160 7254 43172
rect 7760 43160 7788 43191
rect 8018 43188 8024 43200
rect 8076 43188 8082 43240
rect 8570 43228 8576 43240
rect 8531 43200 8576 43228
rect 8570 43188 8576 43200
rect 8628 43188 8634 43240
rect 7248 43132 7788 43160
rect 7248 43120 7254 43132
rect 1394 43052 1400 43104
rect 1452 43092 1458 43104
rect 1489 43095 1547 43101
rect 1489 43092 1501 43095
rect 1452 43064 1501 43092
rect 1452 43052 1458 43064
rect 1489 43061 1501 43064
rect 1535 43061 1547 43095
rect 2130 43092 2136 43104
rect 2091 43064 2136 43092
rect 1489 43055 1547 43061
rect 2130 43052 2136 43064
rect 2188 43052 2194 43104
rect 2958 43092 2964 43104
rect 2919 43064 2964 43092
rect 2958 43052 2964 43064
rect 3016 43052 3022 43104
rect 3418 43092 3424 43104
rect 3379 43064 3424 43092
rect 3418 43052 3424 43064
rect 3476 43052 3482 43104
rect 3510 43052 3516 43104
rect 3568 43092 3574 43104
rect 4065 43095 4123 43101
rect 4065 43092 4077 43095
rect 3568 43064 4077 43092
rect 3568 43052 3574 43064
rect 4065 43061 4077 43064
rect 4111 43061 4123 43095
rect 29914 43092 29920 43104
rect 29875 43064 29920 43092
rect 4065 43055 4123 43061
rect 29914 43052 29920 43064
rect 29972 43052 29978 43104
rect 1104 43002 30820 43024
rect 1104 42950 5915 43002
rect 5967 42950 5979 43002
rect 6031 42950 6043 43002
rect 6095 42950 6107 43002
rect 6159 42950 6171 43002
rect 6223 42950 15846 43002
rect 15898 42950 15910 43002
rect 15962 42950 15974 43002
rect 16026 42950 16038 43002
rect 16090 42950 16102 43002
rect 16154 42950 25776 43002
rect 25828 42950 25840 43002
rect 25892 42950 25904 43002
rect 25956 42950 25968 43002
rect 26020 42950 26032 43002
rect 26084 42950 30820 43002
rect 1104 42928 30820 42950
rect 2498 42888 2504 42900
rect 2459 42860 2504 42888
rect 2498 42848 2504 42860
rect 2556 42848 2562 42900
rect 4709 42891 4767 42897
rect 4709 42857 4721 42891
rect 4755 42888 4767 42891
rect 5258 42888 5264 42900
rect 4755 42860 5264 42888
rect 4755 42857 4767 42860
rect 4709 42851 4767 42857
rect 5258 42848 5264 42860
rect 5316 42848 5322 42900
rect 6638 42888 6644 42900
rect 6599 42860 6644 42888
rect 6638 42848 6644 42860
rect 6696 42848 6702 42900
rect 8389 42891 8447 42897
rect 8389 42857 8401 42891
rect 8435 42888 8447 42891
rect 8570 42888 8576 42900
rect 8435 42860 8576 42888
rect 8435 42857 8447 42860
rect 8389 42851 8447 42857
rect 8570 42848 8576 42860
rect 8628 42848 8634 42900
rect 7190 42820 7196 42832
rect 7024 42792 7196 42820
rect 3786 42752 3792 42764
rect 1688 42724 3792 42752
rect 1688 42693 1716 42724
rect 3786 42712 3792 42724
rect 3844 42712 3850 42764
rect 7024 42761 7052 42792
rect 7190 42780 7196 42792
rect 7248 42780 7254 42832
rect 8018 42780 8024 42832
rect 8076 42820 8082 42832
rect 9766 42820 9772 42832
rect 8076 42792 9772 42820
rect 8076 42780 8082 42792
rect 9766 42780 9772 42792
rect 9824 42780 9830 42832
rect 7009 42755 7067 42761
rect 7009 42721 7021 42755
rect 7055 42721 7067 42755
rect 9858 42752 9864 42764
rect 7009 42715 7067 42721
rect 7392 42724 9864 42752
rect 7392 42696 7420 42724
rect 9858 42712 9864 42724
rect 9916 42712 9922 42764
rect 1673 42687 1731 42693
rect 1673 42653 1685 42687
rect 1719 42653 1731 42687
rect 1673 42647 1731 42653
rect 2133 42687 2191 42693
rect 2133 42653 2145 42687
rect 2179 42684 2191 42687
rect 2222 42684 2228 42696
rect 2179 42656 2228 42684
rect 2179 42653 2191 42656
rect 2133 42647 2191 42653
rect 2222 42644 2228 42656
rect 2280 42644 2286 42696
rect 3694 42644 3700 42696
rect 3752 42684 3758 42696
rect 3973 42687 4031 42693
rect 3973 42684 3985 42687
rect 3752 42656 3985 42684
rect 3752 42644 3758 42656
rect 3973 42653 3985 42656
rect 4019 42653 4031 42687
rect 5074 42684 5080 42696
rect 5035 42656 5080 42684
rect 3973 42647 4031 42653
rect 5074 42644 5080 42656
rect 5132 42644 5138 42696
rect 5718 42644 5724 42696
rect 5776 42684 5782 42696
rect 5997 42687 6055 42693
rect 5997 42684 6009 42687
rect 5776 42656 6009 42684
rect 5776 42644 5782 42656
rect 5997 42653 6009 42656
rect 6043 42653 6055 42687
rect 6822 42684 6828 42696
rect 6783 42656 6828 42684
rect 5997 42647 6055 42653
rect 6822 42644 6828 42656
rect 6880 42644 6886 42696
rect 7101 42687 7159 42693
rect 7101 42684 7113 42687
rect 7024 42656 7113 42684
rect 7024 42628 7052 42656
rect 7101 42653 7113 42656
rect 7147 42653 7159 42687
rect 7101 42647 7159 42653
rect 7193 42687 7251 42693
rect 7193 42653 7205 42687
rect 7239 42653 7251 42687
rect 7193 42647 7251 42653
rect 2501 42619 2559 42625
rect 2501 42585 2513 42619
rect 2547 42616 2559 42619
rect 6730 42616 6736 42628
rect 2547 42588 6736 42616
rect 2547 42585 2559 42588
rect 2501 42579 2559 42585
rect 6730 42576 6736 42588
rect 6788 42576 6794 42628
rect 7006 42576 7012 42628
rect 7064 42576 7070 42628
rect 7208 42616 7236 42647
rect 7374 42644 7380 42696
rect 7432 42684 7438 42696
rect 8205 42687 8263 42693
rect 7432 42656 7525 42684
rect 7432 42644 7438 42656
rect 8205 42653 8217 42687
rect 8251 42684 8263 42687
rect 9122 42684 9128 42696
rect 8251 42656 8984 42684
rect 9083 42656 9128 42684
rect 8251 42653 8263 42656
rect 8205 42647 8263 42653
rect 7650 42616 7656 42628
rect 7208 42588 7656 42616
rect 7650 42576 7656 42588
rect 7708 42576 7714 42628
rect 1486 42548 1492 42560
rect 1447 42520 1492 42548
rect 1486 42508 1492 42520
rect 1544 42508 1550 42560
rect 2685 42551 2743 42557
rect 2685 42517 2697 42551
rect 2731 42548 2743 42551
rect 3142 42548 3148 42560
rect 2731 42520 3148 42548
rect 2731 42517 2743 42520
rect 2685 42511 2743 42517
rect 3142 42508 3148 42520
rect 3200 42508 3206 42560
rect 3786 42548 3792 42560
rect 3747 42520 3792 42548
rect 3786 42508 3792 42520
rect 3844 42508 3850 42560
rect 4522 42548 4528 42560
rect 4483 42520 4528 42548
rect 4522 42508 4528 42520
rect 4580 42508 4586 42560
rect 4706 42548 4712 42560
rect 4667 42520 4712 42548
rect 4706 42508 4712 42520
rect 4764 42508 4770 42560
rect 6181 42551 6239 42557
rect 6181 42517 6193 42551
rect 6227 42548 6239 42551
rect 6546 42548 6552 42560
rect 6227 42520 6552 42548
rect 6227 42517 6239 42520
rect 6181 42511 6239 42517
rect 6546 42508 6552 42520
rect 6604 42508 6610 42560
rect 8956 42557 8984 42656
rect 9122 42644 9128 42656
rect 9180 42644 9186 42696
rect 19797 42687 19855 42693
rect 19797 42653 19809 42687
rect 19843 42653 19855 42687
rect 19797 42647 19855 42653
rect 19981 42687 20039 42693
rect 19981 42653 19993 42687
rect 20027 42684 20039 42687
rect 29914 42684 29920 42696
rect 20027 42656 29920 42684
rect 20027 42653 20039 42656
rect 19981 42647 20039 42653
rect 19812 42616 19840 42647
rect 29914 42644 29920 42656
rect 29972 42644 29978 42696
rect 20162 42616 20168 42628
rect 19812 42588 20168 42616
rect 20162 42576 20168 42588
rect 20220 42576 20226 42628
rect 8941 42551 8999 42557
rect 8941 42517 8953 42551
rect 8987 42517 8999 42551
rect 8941 42511 8999 42517
rect 10226 42508 10232 42560
rect 10284 42548 10290 42560
rect 19613 42551 19671 42557
rect 19613 42548 19625 42551
rect 10284 42520 19625 42548
rect 10284 42508 10290 42520
rect 19613 42517 19625 42520
rect 19659 42517 19671 42551
rect 19613 42511 19671 42517
rect 1104 42458 30820 42480
rect 1104 42406 10880 42458
rect 10932 42406 10944 42458
rect 10996 42406 11008 42458
rect 11060 42406 11072 42458
rect 11124 42406 11136 42458
rect 11188 42406 20811 42458
rect 20863 42406 20875 42458
rect 20927 42406 20939 42458
rect 20991 42406 21003 42458
rect 21055 42406 21067 42458
rect 21119 42406 30820 42458
rect 1104 42384 30820 42406
rect 3050 42344 3056 42356
rect 1688 42316 3056 42344
rect 1688 42217 1716 42316
rect 3050 42304 3056 42316
rect 3108 42304 3114 42356
rect 3694 42344 3700 42356
rect 3655 42316 3700 42344
rect 3694 42304 3700 42316
rect 3752 42304 3758 42356
rect 7282 42344 7288 42356
rect 6932 42316 7288 42344
rect 2501 42279 2559 42285
rect 2501 42245 2513 42279
rect 2547 42245 2559 42279
rect 2501 42239 2559 42245
rect 1673 42211 1731 42217
rect 1673 42177 1685 42211
rect 1719 42177 1731 42211
rect 1673 42171 1731 42177
rect 2133 42075 2191 42081
rect 2133 42041 2145 42075
rect 2179 42072 2191 42075
rect 2222 42072 2228 42084
rect 2179 42044 2228 42072
rect 2179 42041 2191 42044
rect 2133 42035 2191 42041
rect 2222 42032 2228 42044
rect 2280 42032 2286 42084
rect 2516 42072 2544 42239
rect 3234 42168 3240 42220
rect 3292 42208 3298 42220
rect 3513 42211 3571 42217
rect 3513 42208 3525 42211
rect 3292 42180 3525 42208
rect 3292 42168 3298 42180
rect 3513 42177 3525 42180
rect 3559 42208 3571 42211
rect 4709 42211 4767 42217
rect 4709 42208 4721 42211
rect 3559 42180 4721 42208
rect 3559 42177 3571 42180
rect 3513 42171 3571 42177
rect 4709 42177 4721 42180
rect 4755 42177 4767 42211
rect 4709 42171 4767 42177
rect 5629 42211 5687 42217
rect 5629 42177 5641 42211
rect 5675 42208 5687 42211
rect 5718 42208 5724 42220
rect 5675 42180 5724 42208
rect 5675 42177 5687 42180
rect 5629 42171 5687 42177
rect 5718 42168 5724 42180
rect 5776 42168 5782 42220
rect 6454 42168 6460 42220
rect 6512 42208 6518 42220
rect 6932 42217 6960 42316
rect 7282 42304 7288 42316
rect 7340 42344 7346 42356
rect 7340 42316 16574 42344
rect 7340 42304 7346 42316
rect 6733 42211 6791 42217
rect 6733 42208 6745 42211
rect 6512 42180 6745 42208
rect 6512 42168 6518 42180
rect 6733 42177 6745 42180
rect 6779 42177 6791 42211
rect 6733 42171 6791 42177
rect 6917 42211 6975 42217
rect 6917 42177 6929 42211
rect 6963 42177 6975 42211
rect 6917 42171 6975 42177
rect 7285 42211 7343 42217
rect 7285 42177 7297 42211
rect 7331 42208 7343 42211
rect 7742 42208 7748 42220
rect 7331 42180 7748 42208
rect 7331 42177 7343 42180
rect 7285 42171 7343 42177
rect 7742 42168 7748 42180
rect 7800 42168 7806 42220
rect 7929 42211 7987 42217
rect 7929 42177 7941 42211
rect 7975 42177 7987 42211
rect 16546 42208 16574 42316
rect 21910 42208 21916 42220
rect 16546 42180 21916 42208
rect 7929 42171 7987 42177
rect 2682 42100 2688 42152
rect 2740 42140 2746 42152
rect 5074 42140 5080 42152
rect 2740 42112 5080 42140
rect 2740 42100 2746 42112
rect 5074 42100 5080 42112
rect 5132 42100 5138 42152
rect 7006 42140 7012 42152
rect 6967 42112 7012 42140
rect 7006 42100 7012 42112
rect 7064 42100 7070 42152
rect 7101 42143 7159 42149
rect 7101 42109 7113 42143
rect 7147 42140 7159 42143
rect 7190 42140 7196 42152
rect 7147 42112 7196 42140
rect 7147 42109 7159 42112
rect 7101 42103 7159 42109
rect 7190 42100 7196 42112
rect 7248 42100 7254 42152
rect 5813 42075 5871 42081
rect 2516 42044 5028 42072
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 1489 42007 1547 42013
rect 1489 42004 1501 42007
rect 1452 41976 1501 42004
rect 1452 41964 1458 41976
rect 1489 41973 1501 41976
rect 1535 41973 1547 42007
rect 2498 42004 2504 42016
rect 2459 41976 2504 42004
rect 1489 41967 1547 41973
rect 2498 41964 2504 41976
rect 2556 41964 2562 42016
rect 2685 42007 2743 42013
rect 2685 41973 2697 42007
rect 2731 42004 2743 42007
rect 4338 42004 4344 42016
rect 2731 41976 4344 42004
rect 2731 41973 2743 41976
rect 2685 41967 2743 41973
rect 4338 41964 4344 41976
rect 4396 41964 4402 42016
rect 4890 42004 4896 42016
rect 4851 41976 4896 42004
rect 4890 41964 4896 41976
rect 4948 41964 4954 42016
rect 5000 42004 5028 42044
rect 5813 42041 5825 42075
rect 5859 42072 5871 42075
rect 7944 42072 7972 42171
rect 21910 42168 21916 42180
rect 21968 42168 21974 42220
rect 5859 42044 7972 42072
rect 5859 42041 5871 42044
rect 5813 42035 5871 42041
rect 6914 42004 6920 42016
rect 5000 41976 6920 42004
rect 6914 41964 6920 41976
rect 6972 41964 6978 42016
rect 7466 42004 7472 42016
rect 7427 41976 7472 42004
rect 7466 41964 7472 41976
rect 7524 41964 7530 42016
rect 8113 42007 8171 42013
rect 8113 41973 8125 42007
rect 8159 42004 8171 42007
rect 8386 42004 8392 42016
rect 8159 41976 8392 42004
rect 8159 41973 8171 41976
rect 8113 41967 8171 41973
rect 8386 41964 8392 41976
rect 8444 41964 8450 42016
rect 1104 41914 30820 41936
rect 1104 41862 5915 41914
rect 5967 41862 5979 41914
rect 6031 41862 6043 41914
rect 6095 41862 6107 41914
rect 6159 41862 6171 41914
rect 6223 41862 15846 41914
rect 15898 41862 15910 41914
rect 15962 41862 15974 41914
rect 16026 41862 16038 41914
rect 16090 41862 16102 41914
rect 16154 41862 25776 41914
rect 25828 41862 25840 41914
rect 25892 41862 25904 41914
rect 25956 41862 25968 41914
rect 26020 41862 26032 41914
rect 26084 41862 30820 41914
rect 1104 41840 30820 41862
rect 2498 41800 2504 41812
rect 2459 41772 2504 41800
rect 2498 41760 2504 41772
rect 2556 41760 2562 41812
rect 2685 41803 2743 41809
rect 2685 41769 2697 41803
rect 2731 41800 2743 41803
rect 3970 41800 3976 41812
rect 2731 41772 3976 41800
rect 2731 41769 2743 41772
rect 2685 41763 2743 41769
rect 3970 41760 3976 41772
rect 4028 41760 4034 41812
rect 4706 41760 4712 41812
rect 4764 41800 4770 41812
rect 7009 41803 7067 41809
rect 7009 41800 7021 41803
rect 4764 41772 7021 41800
rect 4764 41760 4770 41772
rect 7009 41769 7021 41772
rect 7055 41800 7067 41803
rect 7742 41800 7748 41812
rect 7055 41772 7748 41800
rect 7055 41769 7067 41772
rect 7009 41763 7067 41769
rect 7742 41760 7748 41772
rect 7800 41760 7806 41812
rect 3510 41664 3516 41676
rect 1688 41636 3516 41664
rect 1688 41605 1716 41636
rect 3510 41624 3516 41636
rect 3568 41624 3574 41676
rect 3786 41664 3792 41676
rect 3747 41636 3792 41664
rect 3786 41624 3792 41636
rect 3844 41624 3850 41676
rect 5074 41624 5080 41676
rect 5132 41664 5138 41676
rect 5905 41667 5963 41673
rect 5905 41664 5917 41667
rect 5132 41636 5917 41664
rect 5132 41624 5138 41636
rect 5905 41633 5917 41636
rect 5951 41633 5963 41667
rect 8386 41664 8392 41676
rect 8347 41636 8392 41664
rect 5905 41627 5963 41633
rect 8386 41624 8392 41636
rect 8444 41624 8450 41676
rect 1673 41599 1731 41605
rect 1673 41565 1685 41599
rect 1719 41565 1731 41599
rect 1673 41559 1731 41565
rect 2133 41599 2191 41605
rect 2133 41565 2145 41599
rect 2179 41596 2191 41599
rect 2222 41596 2228 41608
rect 2179 41568 2228 41596
rect 2179 41565 2191 41568
rect 2133 41559 2191 41565
rect 2222 41556 2228 41568
rect 2280 41596 2286 41608
rect 2682 41596 2688 41608
rect 2280 41568 2688 41596
rect 2280 41556 2286 41568
rect 2682 41556 2688 41568
rect 2740 41556 2746 41608
rect 5626 41596 5632 41608
rect 3988 41568 4292 41596
rect 5587 41568 5632 41596
rect 2501 41531 2559 41537
rect 2501 41497 2513 41531
rect 2547 41528 2559 41531
rect 3988 41528 4016 41568
rect 4062 41537 4068 41540
rect 2547 41500 4016 41528
rect 2547 41497 2559 41500
rect 2501 41491 2559 41497
rect 4056 41491 4068 41537
rect 4120 41528 4126 41540
rect 4264 41528 4292 41568
rect 5626 41556 5632 41568
rect 5684 41556 5690 41608
rect 6546 41556 6552 41608
rect 6604 41596 6610 41608
rect 9125 41599 9183 41605
rect 9125 41596 9137 41599
rect 6604 41568 9137 41596
rect 6604 41556 6610 41568
rect 9125 41565 9137 41568
rect 9171 41565 9183 41599
rect 9125 41559 9183 41565
rect 6270 41528 6276 41540
rect 4120 41500 4156 41528
rect 4264 41500 6276 41528
rect 4062 41488 4068 41491
rect 4120 41488 4126 41500
rect 6270 41488 6276 41500
rect 6328 41488 6334 41540
rect 7466 41488 7472 41540
rect 7524 41528 7530 41540
rect 8122 41531 8180 41537
rect 8122 41528 8134 41531
rect 7524 41500 8134 41528
rect 7524 41488 7530 41500
rect 8122 41497 8134 41500
rect 8168 41497 8180 41531
rect 10226 41528 10232 41540
rect 8122 41491 8180 41497
rect 8220 41500 10232 41528
rect 1302 41420 1308 41472
rect 1360 41460 1366 41472
rect 1489 41463 1547 41469
rect 1489 41460 1501 41463
rect 1360 41432 1501 41460
rect 1360 41420 1366 41432
rect 1489 41429 1501 41432
rect 1535 41429 1547 41463
rect 1489 41423 1547 41429
rect 3786 41420 3792 41472
rect 3844 41460 3850 41472
rect 5169 41463 5227 41469
rect 5169 41460 5181 41463
rect 3844 41432 5181 41460
rect 3844 41420 3850 41432
rect 5169 41429 5181 41432
rect 5215 41429 5227 41463
rect 5169 41423 5227 41429
rect 7650 41420 7656 41472
rect 7708 41460 7714 41472
rect 8220 41460 8248 41500
rect 10226 41488 10232 41500
rect 10284 41488 10290 41540
rect 8938 41460 8944 41472
rect 7708 41432 8248 41460
rect 8899 41432 8944 41460
rect 7708 41420 7714 41432
rect 8938 41420 8944 41432
rect 8996 41420 9002 41472
rect 1104 41370 30820 41392
rect 1104 41318 10880 41370
rect 10932 41318 10944 41370
rect 10996 41318 11008 41370
rect 11060 41318 11072 41370
rect 11124 41318 11136 41370
rect 11188 41318 20811 41370
rect 20863 41318 20875 41370
rect 20927 41318 20939 41370
rect 20991 41318 21003 41370
rect 21055 41318 21067 41370
rect 21119 41318 30820 41370
rect 1104 41296 30820 41318
rect 2501 41259 2559 41265
rect 2501 41225 2513 41259
rect 2547 41256 2559 41259
rect 3878 41256 3884 41268
rect 2547 41228 3884 41256
rect 2547 41225 2559 41228
rect 2501 41219 2559 41225
rect 3878 41216 3884 41228
rect 3936 41216 3942 41268
rect 3973 41259 4031 41265
rect 3973 41225 3985 41259
rect 4019 41256 4031 41259
rect 4062 41256 4068 41268
rect 4019 41228 4068 41256
rect 4019 41225 4031 41228
rect 3973 41219 4031 41225
rect 4062 41216 4068 41228
rect 4120 41216 4126 41268
rect 6730 41256 6736 41268
rect 6691 41228 6736 41256
rect 6730 41216 6736 41228
rect 6788 41216 6794 41268
rect 7006 41216 7012 41268
rect 7064 41256 7070 41268
rect 8803 41259 8861 41265
rect 8803 41256 8815 41259
rect 7064 41228 8815 41256
rect 7064 41216 7070 41228
rect 8803 41225 8815 41228
rect 8849 41225 8861 41259
rect 8803 41219 8861 41225
rect 16117 41259 16175 41265
rect 16117 41225 16129 41259
rect 16163 41225 16175 41259
rect 16117 41219 16175 41225
rect 2317 41191 2375 41197
rect 2317 41157 2329 41191
rect 2363 41188 2375 41191
rect 16132 41188 16160 41219
rect 2363 41160 3832 41188
rect 16132 41160 16804 41188
rect 2363 41157 2375 41160
rect 2317 41151 2375 41157
rect 3804 41132 3832 41160
rect 1949 41123 2007 41129
rect 1949 41089 1961 41123
rect 1995 41120 2007 41123
rect 2130 41120 2136 41132
rect 1995 41092 2136 41120
rect 1995 41089 2007 41092
rect 1949 41083 2007 41089
rect 2130 41080 2136 41092
rect 2188 41080 2194 41132
rect 3237 41123 3295 41129
rect 3237 41089 3249 41123
rect 3283 41089 3295 41123
rect 3237 41083 3295 41089
rect 3421 41123 3479 41129
rect 3421 41089 3433 41123
rect 3467 41120 3479 41123
rect 3694 41120 3700 41132
rect 3467 41092 3700 41120
rect 3467 41089 3479 41092
rect 3421 41083 3479 41089
rect 2317 40919 2375 40925
rect 2317 40885 2329 40919
rect 2363 40916 2375 40919
rect 2406 40916 2412 40928
rect 2363 40888 2412 40916
rect 2363 40885 2375 40888
rect 2317 40879 2375 40885
rect 2406 40876 2412 40888
rect 2464 40876 2470 40928
rect 3252 40916 3280 41083
rect 3694 41080 3700 41092
rect 3752 41080 3758 41132
rect 3786 41080 3792 41132
rect 3844 41129 3850 41132
rect 3844 41123 3858 41129
rect 3846 41120 3858 41123
rect 3846 41092 3889 41120
rect 3846 41089 3858 41092
rect 3844 41083 3858 41089
rect 3844 41080 3850 41083
rect 4338 41080 4344 41132
rect 4396 41120 4402 41132
rect 5546 41123 5604 41129
rect 5546 41120 5558 41123
rect 4396 41092 5558 41120
rect 4396 41080 4402 41092
rect 5546 41089 5558 41092
rect 5592 41089 5604 41123
rect 5546 41083 5604 41089
rect 7098 41080 7104 41132
rect 7156 41120 7162 41132
rect 7846 41123 7904 41129
rect 7846 41120 7858 41123
rect 7156 41092 7858 41120
rect 7156 41080 7162 41092
rect 7846 41089 7858 41092
rect 7892 41089 7904 41123
rect 7846 41083 7904 41089
rect 8113 41123 8171 41129
rect 8113 41089 8125 41123
rect 8159 41120 8171 41123
rect 8938 41120 8944 41132
rect 8159 41092 8944 41120
rect 8159 41089 8171 41092
rect 8113 41083 8171 41089
rect 8938 41080 8944 41092
rect 8996 41080 9002 41132
rect 15933 41123 15991 41129
rect 15933 41089 15945 41123
rect 15979 41120 15991 41123
rect 16206 41120 16212 41132
rect 15979 41092 16212 41120
rect 15979 41089 15991 41092
rect 15933 41083 15991 41089
rect 16206 41080 16212 41092
rect 16264 41080 16270 41132
rect 16776 41129 16804 41160
rect 16761 41123 16819 41129
rect 16761 41089 16773 41123
rect 16807 41120 16819 41123
rect 16850 41120 16856 41132
rect 16807 41092 16856 41120
rect 16807 41089 16819 41092
rect 16761 41083 16819 41089
rect 16850 41080 16856 41092
rect 16908 41080 16914 41132
rect 30098 41120 30104 41132
rect 30059 41092 30104 41120
rect 30098 41080 30104 41092
rect 30156 41080 30162 41132
rect 3510 41052 3516 41064
rect 3471 41024 3516 41052
rect 3510 41012 3516 41024
rect 3568 41012 3574 41064
rect 3605 41055 3663 41061
rect 3605 41021 3617 41055
rect 3651 41052 3663 41055
rect 4154 41052 4160 41064
rect 3651 41024 4160 41052
rect 3651 41021 3663 41024
rect 3605 41015 3663 41021
rect 4154 41012 4160 41024
rect 4212 41012 4218 41064
rect 5810 41052 5816 41064
rect 5771 41024 5816 41052
rect 5810 41012 5816 41024
rect 5868 41012 5874 41064
rect 8478 41012 8484 41064
rect 8536 41052 8542 41064
rect 8573 41055 8631 41061
rect 8573 41052 8585 41055
rect 8536 41024 8585 41052
rect 8536 41012 8542 41024
rect 8573 41021 8585 41024
rect 8619 41021 8631 41055
rect 8573 41015 8631 41021
rect 4522 40984 4528 40996
rect 4264 40956 4528 40984
rect 4264 40916 4292 40956
rect 4522 40944 4528 40956
rect 4580 40984 4586 40996
rect 4580 40956 4948 40984
rect 4580 40944 4586 40956
rect 4430 40916 4436 40928
rect 3252 40888 4292 40916
rect 4391 40888 4436 40916
rect 4430 40876 4436 40888
rect 4488 40876 4494 40928
rect 4920 40916 4948 40956
rect 5166 40916 5172 40928
rect 4920 40888 5172 40916
rect 5166 40876 5172 40888
rect 5224 40876 5230 40928
rect 16758 40916 16764 40928
rect 16719 40888 16764 40916
rect 16758 40876 16764 40888
rect 16816 40876 16822 40928
rect 29914 40916 29920 40928
rect 29875 40888 29920 40916
rect 29914 40876 29920 40888
rect 29972 40876 29978 40928
rect 1104 40826 30820 40848
rect 1104 40774 5915 40826
rect 5967 40774 5979 40826
rect 6031 40774 6043 40826
rect 6095 40774 6107 40826
rect 6159 40774 6171 40826
rect 6223 40774 15846 40826
rect 15898 40774 15910 40826
rect 15962 40774 15974 40826
rect 16026 40774 16038 40826
rect 16090 40774 16102 40826
rect 16154 40774 25776 40826
rect 25828 40774 25840 40826
rect 25892 40774 25904 40826
rect 25956 40774 25968 40826
rect 26020 40774 26032 40826
rect 26084 40774 30820 40826
rect 1104 40752 30820 40774
rect 2406 40672 2412 40724
rect 2464 40712 2470 40724
rect 2501 40715 2559 40721
rect 2501 40712 2513 40715
rect 2464 40684 2513 40712
rect 2464 40672 2470 40684
rect 2501 40681 2513 40684
rect 2547 40681 2559 40715
rect 2501 40675 2559 40681
rect 2685 40715 2743 40721
rect 2685 40681 2697 40715
rect 2731 40712 2743 40715
rect 2866 40712 2872 40724
rect 2731 40684 2872 40712
rect 2731 40681 2743 40684
rect 2685 40675 2743 40681
rect 2866 40672 2872 40684
rect 2924 40672 2930 40724
rect 4338 40712 4344 40724
rect 4299 40684 4344 40712
rect 4338 40672 4344 40684
rect 4396 40672 4402 40724
rect 2133 40647 2191 40653
rect 2133 40613 2145 40647
rect 2179 40644 2191 40647
rect 2222 40644 2228 40656
rect 2179 40616 2228 40644
rect 2179 40613 2191 40616
rect 2133 40607 2191 40613
rect 2222 40604 2228 40616
rect 2280 40604 2286 40656
rect 3694 40604 3700 40656
rect 3752 40644 3758 40656
rect 8018 40644 8024 40656
rect 3752 40616 8024 40644
rect 3752 40604 3758 40616
rect 8018 40604 8024 40616
rect 8076 40604 8082 40656
rect 14476 40616 15240 40644
rect 4798 40536 4804 40588
rect 4856 40576 4862 40588
rect 4856 40548 4901 40576
rect 4856 40536 4862 40548
rect 5626 40536 5632 40588
rect 5684 40576 5690 40588
rect 7190 40576 7196 40588
rect 5684 40548 6408 40576
rect 7151 40548 7196 40576
rect 5684 40536 5690 40548
rect 1673 40511 1731 40517
rect 1673 40477 1685 40511
rect 1719 40508 1731 40511
rect 1762 40508 1768 40520
rect 1719 40480 1768 40508
rect 1719 40477 1731 40480
rect 1673 40471 1731 40477
rect 1762 40468 1768 40480
rect 1820 40468 1826 40520
rect 4430 40508 4436 40520
rect 2516 40480 4436 40508
rect 2516 40449 2544 40480
rect 4430 40468 4436 40480
rect 4488 40508 4494 40520
rect 4525 40511 4583 40517
rect 4525 40508 4537 40511
rect 4488 40480 4537 40508
rect 4488 40468 4494 40480
rect 4525 40477 4537 40480
rect 4571 40477 4583 40511
rect 4525 40471 4583 40477
rect 4706 40468 4712 40520
rect 4764 40508 4770 40520
rect 4893 40511 4951 40517
rect 4764 40480 4809 40508
rect 4764 40468 4770 40480
rect 4893 40477 4905 40511
rect 4939 40477 4951 40511
rect 4893 40471 4951 40477
rect 5077 40511 5135 40517
rect 5077 40477 5089 40511
rect 5123 40508 5135 40511
rect 5166 40508 5172 40520
rect 5123 40480 5172 40508
rect 5123 40477 5135 40480
rect 5077 40471 5135 40477
rect 2501 40443 2559 40449
rect 2501 40409 2513 40443
rect 2547 40409 2559 40443
rect 4908 40440 4936 40471
rect 5166 40468 5172 40480
rect 5224 40468 5230 40520
rect 5350 40468 5356 40520
rect 5408 40508 5414 40520
rect 6089 40511 6147 40517
rect 6089 40508 6101 40511
rect 5408 40480 6101 40508
rect 5408 40468 5414 40480
rect 6089 40477 6101 40480
rect 6135 40508 6147 40511
rect 6270 40508 6276 40520
rect 6135 40480 6276 40508
rect 6135 40477 6147 40480
rect 6089 40471 6147 40477
rect 6270 40468 6276 40480
rect 6328 40468 6334 40520
rect 6380 40517 6408 40548
rect 7190 40536 7196 40548
rect 7248 40536 7254 40588
rect 14476 40520 14504 40616
rect 15102 40576 15108 40588
rect 15063 40548 15108 40576
rect 15102 40536 15108 40548
rect 15160 40536 15166 40588
rect 15212 40576 15240 40616
rect 15381 40579 15439 40585
rect 15381 40576 15393 40579
rect 15212 40548 15393 40576
rect 15381 40545 15393 40548
rect 15427 40545 15439 40579
rect 15381 40539 15439 40545
rect 15657 40579 15715 40585
rect 15657 40545 15669 40579
rect 15703 40576 15715 40579
rect 16298 40576 16304 40588
rect 15703 40548 16304 40576
rect 15703 40545 15715 40548
rect 15657 40539 15715 40545
rect 16298 40536 16304 40548
rect 16356 40536 16362 40588
rect 6365 40511 6423 40517
rect 6365 40477 6377 40511
rect 6411 40508 6423 40511
rect 6546 40508 6552 40520
rect 6411 40480 6552 40508
rect 6411 40477 6423 40480
rect 6365 40471 6423 40477
rect 6546 40468 6552 40480
rect 6604 40468 6610 40520
rect 6917 40511 6975 40517
rect 6917 40477 6929 40511
rect 6963 40508 6975 40511
rect 7006 40508 7012 40520
rect 6963 40480 7012 40508
rect 6963 40477 6975 40480
rect 6917 40471 6975 40477
rect 7006 40468 7012 40480
rect 7064 40468 7070 40520
rect 8294 40468 8300 40520
rect 8352 40508 8358 40520
rect 9122 40508 9128 40520
rect 8352 40480 9128 40508
rect 8352 40468 8358 40480
rect 9122 40468 9128 40480
rect 9180 40468 9186 40520
rect 9582 40508 9588 40520
rect 9543 40480 9588 40508
rect 9582 40468 9588 40480
rect 9640 40468 9646 40520
rect 12158 40468 12164 40520
rect 12216 40508 12222 40520
rect 12345 40511 12403 40517
rect 12345 40508 12357 40511
rect 12216 40480 12357 40508
rect 12216 40468 12222 40480
rect 12345 40477 12357 40480
rect 12391 40477 12403 40511
rect 12986 40508 12992 40520
rect 12947 40480 12992 40508
rect 12345 40471 12403 40477
rect 12986 40468 12992 40480
rect 13044 40468 13050 40520
rect 14458 40508 14464 40520
rect 14419 40480 14464 40508
rect 14458 40468 14464 40480
rect 14516 40468 14522 40520
rect 14642 40508 14648 40520
rect 14603 40480 14648 40508
rect 14642 40468 14648 40480
rect 14700 40468 14706 40520
rect 15470 40468 15476 40520
rect 15528 40517 15534 40520
rect 15528 40511 15556 40517
rect 15544 40477 15556 40511
rect 16945 40511 17003 40517
rect 16945 40508 16957 40511
rect 15528 40471 15556 40477
rect 16224 40480 16957 40508
rect 15528 40468 15534 40471
rect 9030 40440 9036 40452
rect 4908 40412 9036 40440
rect 2501 40403 2559 40409
rect 9030 40400 9036 40412
rect 9088 40400 9094 40452
rect 1486 40372 1492 40384
rect 1447 40344 1492 40372
rect 1486 40332 1492 40344
rect 1544 40332 1550 40384
rect 8938 40372 8944 40384
rect 8899 40344 8944 40372
rect 8938 40332 8944 40344
rect 8996 40332 9002 40384
rect 9769 40375 9827 40381
rect 9769 40341 9781 40375
rect 9815 40372 9827 40375
rect 10410 40372 10416 40384
rect 9815 40344 10416 40372
rect 9815 40341 9827 40344
rect 9769 40335 9827 40341
rect 10410 40332 10416 40344
rect 10468 40332 10474 40384
rect 12526 40372 12532 40384
rect 12487 40344 12532 40372
rect 12526 40332 12532 40344
rect 12584 40332 12590 40384
rect 13173 40375 13231 40381
rect 13173 40341 13185 40375
rect 13219 40372 13231 40375
rect 13538 40372 13544 40384
rect 13219 40344 13544 40372
rect 13219 40341 13231 40344
rect 13173 40335 13231 40341
rect 13538 40332 13544 40344
rect 13596 40332 13602 40384
rect 15194 40332 15200 40384
rect 15252 40372 15258 40384
rect 15746 40372 15752 40384
rect 15252 40344 15752 40372
rect 15252 40332 15258 40344
rect 15746 40332 15752 40344
rect 15804 40372 15810 40384
rect 16224 40372 16252 40480
rect 16945 40477 16957 40480
rect 16991 40477 17003 40511
rect 16945 40471 17003 40477
rect 17402 40468 17408 40520
rect 17460 40508 17466 40520
rect 17681 40511 17739 40517
rect 17681 40508 17693 40511
rect 17460 40480 17693 40508
rect 17460 40468 17466 40480
rect 17681 40477 17693 40480
rect 17727 40477 17739 40511
rect 17681 40471 17739 40477
rect 16574 40400 16580 40452
rect 16632 40440 16638 40452
rect 16761 40443 16819 40449
rect 16761 40440 16773 40443
rect 16632 40412 16773 40440
rect 16632 40400 16638 40412
rect 16761 40409 16773 40412
rect 16807 40409 16819 40443
rect 17586 40440 17592 40452
rect 17547 40412 17592 40440
rect 16761 40403 16819 40409
rect 17586 40400 17592 40412
rect 17644 40400 17650 40452
rect 15804 40344 16252 40372
rect 16301 40375 16359 40381
rect 15804 40332 15810 40344
rect 16301 40341 16313 40375
rect 16347 40372 16359 40375
rect 17034 40372 17040 40384
rect 16347 40344 17040 40372
rect 16347 40341 16359 40344
rect 16301 40335 16359 40341
rect 17034 40332 17040 40344
rect 17092 40332 17098 40384
rect 17126 40332 17132 40384
rect 17184 40372 17190 40384
rect 17184 40344 17229 40372
rect 17184 40332 17190 40344
rect 1104 40282 30820 40304
rect 1104 40230 10880 40282
rect 10932 40230 10944 40282
rect 10996 40230 11008 40282
rect 11060 40230 11072 40282
rect 11124 40230 11136 40282
rect 11188 40230 20811 40282
rect 20863 40230 20875 40282
rect 20927 40230 20939 40282
rect 20991 40230 21003 40282
rect 21055 40230 21067 40282
rect 21119 40230 30820 40282
rect 1104 40208 30820 40230
rect 3418 40168 3424 40180
rect 1688 40140 3424 40168
rect 1688 40041 1716 40140
rect 3418 40128 3424 40140
rect 3476 40128 3482 40180
rect 3970 40128 3976 40180
rect 4028 40168 4034 40180
rect 4525 40171 4583 40177
rect 4525 40168 4537 40171
rect 4028 40140 4537 40168
rect 4028 40128 4034 40140
rect 4525 40137 4537 40140
rect 4571 40137 4583 40171
rect 4525 40131 4583 40137
rect 5169 40171 5227 40177
rect 5169 40137 5181 40171
rect 5215 40168 5227 40171
rect 5810 40168 5816 40180
rect 5215 40140 5816 40168
rect 5215 40137 5227 40140
rect 5169 40131 5227 40137
rect 5810 40128 5816 40140
rect 5868 40128 5874 40180
rect 7929 40171 7987 40177
rect 6564 40140 7052 40168
rect 4890 40060 4896 40112
rect 4948 40100 4954 40112
rect 4948 40072 5028 40100
rect 4948 40060 4954 40072
rect 1673 40035 1731 40041
rect 1673 40001 1685 40035
rect 1719 40001 1731 40035
rect 1673 39995 1731 40001
rect 2501 40035 2559 40041
rect 2501 40001 2513 40035
rect 2547 40032 2559 40035
rect 3050 40032 3056 40044
rect 2547 40004 3056 40032
rect 2547 40001 2559 40004
rect 2501 39995 2559 40001
rect 3050 39992 3056 40004
rect 3108 39992 3114 40044
rect 3412 40035 3470 40041
rect 3412 40001 3424 40035
rect 3458 40032 3470 40035
rect 3786 40032 3792 40044
rect 3458 40004 3792 40032
rect 3458 40001 3470 40004
rect 3412 39995 3470 40001
rect 3786 39992 3792 40004
rect 3844 39992 3850 40044
rect 5000 40041 5028 40072
rect 4985 40035 5043 40041
rect 4985 40001 4997 40035
rect 5031 40001 5043 40035
rect 5626 40032 5632 40044
rect 5587 40004 5632 40032
rect 4985 39995 5043 40001
rect 5626 39992 5632 40004
rect 5684 39992 5690 40044
rect 6365 40035 6423 40041
rect 6365 40001 6377 40035
rect 6411 40032 6423 40035
rect 6454 40032 6460 40044
rect 6411 40004 6460 40032
rect 6411 40001 6423 40004
rect 6365 39995 6423 40001
rect 6454 39992 6460 40004
rect 6512 39992 6518 40044
rect 6564 40041 6592 40140
rect 6730 40060 6736 40112
rect 6788 40100 6794 40112
rect 7024 40100 7052 40140
rect 7929 40137 7941 40171
rect 7975 40168 7987 40171
rect 9582 40168 9588 40180
rect 7975 40140 9588 40168
rect 7975 40137 7987 40140
rect 7929 40131 7987 40137
rect 9582 40128 9588 40140
rect 9640 40128 9646 40180
rect 12158 40168 12164 40180
rect 12119 40140 12164 40168
rect 12158 40128 12164 40140
rect 12216 40128 12222 40180
rect 13170 40128 13176 40180
rect 13228 40168 13234 40180
rect 15194 40168 15200 40180
rect 13228 40140 15200 40168
rect 13228 40128 13234 40140
rect 15194 40128 15200 40140
rect 15252 40128 15258 40180
rect 15657 40171 15715 40177
rect 15657 40137 15669 40171
rect 15703 40168 15715 40171
rect 17862 40168 17868 40180
rect 15703 40140 17868 40168
rect 15703 40137 15715 40140
rect 15657 40131 15715 40137
rect 17862 40128 17868 40140
rect 17920 40128 17926 40180
rect 8294 40100 8300 40112
rect 6788 40072 6960 40100
rect 7024 40072 7696 40100
rect 6788 40060 6794 40072
rect 6932 40041 6960 40072
rect 6549 40035 6607 40041
rect 6549 40001 6561 40035
rect 6595 40001 6607 40035
rect 6549 39995 6607 40001
rect 6917 40035 6975 40041
rect 6917 40001 6929 40035
rect 6963 40001 6975 40035
rect 7098 40032 7104 40044
rect 7059 40004 7104 40032
rect 6917 39995 6975 40001
rect 7098 39992 7104 40004
rect 7156 39992 7162 40044
rect 3145 39967 3203 39973
rect 3145 39933 3157 39967
rect 3191 39933 3203 39967
rect 6638 39964 6644 39976
rect 6599 39936 6644 39964
rect 3145 39927 3203 39933
rect 1394 39788 1400 39840
rect 1452 39828 1458 39840
rect 1489 39831 1547 39837
rect 1489 39828 1501 39831
rect 1452 39800 1501 39828
rect 1452 39788 1458 39800
rect 1489 39797 1501 39800
rect 1535 39797 1547 39831
rect 1489 39791 1547 39797
rect 2685 39831 2743 39837
rect 2685 39797 2697 39831
rect 2731 39828 2743 39831
rect 3160 39828 3188 39927
rect 6638 39924 6644 39936
rect 6696 39924 6702 39976
rect 6733 39967 6791 39973
rect 6733 39933 6745 39967
rect 6779 39964 6791 39967
rect 7006 39964 7012 39976
rect 6779 39936 7012 39964
rect 6779 39933 6791 39936
rect 6733 39927 6791 39933
rect 7006 39924 7012 39936
rect 7064 39924 7070 39976
rect 7668 39964 7696 40072
rect 7760 40072 8300 40100
rect 7760 40041 7788 40072
rect 8294 40060 8300 40072
rect 8352 40060 8358 40112
rect 8938 40100 8944 40112
rect 8404 40072 8944 40100
rect 8404 40041 8432 40072
rect 8938 40060 8944 40072
rect 8996 40060 9002 40112
rect 9030 40060 9036 40112
rect 9088 40100 9094 40112
rect 9490 40100 9496 40112
rect 9088 40072 9496 40100
rect 9088 40060 9094 40072
rect 9490 40060 9496 40072
rect 9548 40100 9554 40112
rect 9858 40100 9864 40112
rect 9548 40072 9864 40100
rect 9548 40060 9554 40072
rect 9858 40060 9864 40072
rect 9916 40060 9922 40112
rect 15289 40103 15347 40109
rect 11992 40072 12848 40100
rect 7745 40035 7803 40041
rect 7745 40001 7757 40035
rect 7791 40001 7803 40035
rect 7745 39995 7803 40001
rect 8389 40035 8447 40041
rect 8389 40001 8401 40035
rect 8435 40001 8447 40035
rect 8389 39995 8447 40001
rect 9674 39992 9680 40044
rect 9732 40032 9738 40044
rect 10146 40035 10204 40041
rect 10146 40032 10158 40035
rect 9732 40004 10158 40032
rect 9732 39992 9738 40004
rect 10146 40001 10158 40004
rect 10192 40001 10204 40035
rect 10410 40032 10416 40044
rect 10371 40004 10416 40032
rect 10146 39995 10204 40001
rect 10410 39992 10416 40004
rect 10468 39992 10474 40044
rect 11992 40041 12020 40072
rect 11977 40035 12035 40041
rect 11977 40001 11989 40035
rect 12023 40001 12035 40035
rect 11977 39995 12035 40001
rect 12526 39992 12532 40044
rect 12584 40032 12590 40044
rect 12621 40035 12679 40041
rect 12621 40032 12633 40035
rect 12584 40004 12633 40032
rect 12584 39992 12590 40004
rect 12621 40001 12633 40004
rect 12667 40001 12679 40035
rect 12820 40032 12848 40072
rect 15289 40069 15301 40103
rect 15335 40069 15347 40103
rect 15289 40063 15347 40069
rect 14461 40035 14519 40041
rect 12820 40004 12940 40032
rect 12621 39995 12679 40001
rect 8754 39964 8760 39976
rect 7668 39936 8760 39964
rect 8754 39924 8760 39936
rect 8812 39924 8818 39976
rect 12805 39967 12863 39973
rect 12805 39964 12817 39967
rect 12636 39936 12817 39964
rect 12636 39908 12664 39936
rect 12805 39933 12817 39936
rect 12851 39933 12863 39967
rect 12912 39964 12940 40004
rect 14461 40001 14473 40035
rect 14507 40032 14519 40035
rect 15304 40032 15332 40063
rect 14507 40004 15332 40032
rect 16669 40035 16727 40041
rect 14507 40001 14519 40004
rect 14461 39995 14519 40001
rect 16669 40001 16681 40035
rect 16715 40032 16727 40035
rect 16758 40032 16764 40044
rect 16715 40004 16764 40032
rect 16715 40001 16727 40004
rect 16669 39995 16727 40001
rect 16758 39992 16764 40004
rect 16816 39992 16822 40044
rect 16850 39992 16856 40044
rect 16908 40032 16914 40044
rect 16908 40004 16953 40032
rect 16908 39992 16914 40004
rect 17586 39992 17592 40044
rect 17644 40032 17650 40044
rect 19153 40035 19211 40041
rect 17644 40004 17689 40032
rect 17644 39992 17650 40004
rect 19153 40001 19165 40035
rect 19199 40032 19211 40035
rect 19334 40032 19340 40044
rect 19199 40004 19340 40032
rect 19199 40001 19211 40004
rect 19153 39995 19211 40001
rect 19334 39992 19340 40004
rect 19392 39992 19398 40044
rect 22094 39992 22100 40044
rect 22152 40032 22158 40044
rect 22281 40035 22339 40041
rect 22281 40032 22293 40035
rect 22152 40004 22293 40032
rect 22152 39992 22158 40004
rect 22281 40001 22293 40004
rect 22327 40001 22339 40035
rect 22281 39995 22339 40001
rect 13541 39967 13599 39973
rect 13541 39964 13553 39967
rect 12912 39936 13553 39964
rect 12805 39927 12863 39933
rect 4338 39856 4344 39908
rect 4396 39896 4402 39908
rect 7650 39896 7656 39908
rect 4396 39868 7656 39896
rect 4396 39856 4402 39868
rect 7650 39856 7656 39868
rect 7708 39856 7714 39908
rect 12618 39856 12624 39908
rect 12676 39856 12682 39908
rect 13262 39896 13268 39908
rect 13223 39868 13268 39896
rect 13262 39856 13268 39868
rect 13320 39856 13326 39908
rect 13372 39840 13400 39936
rect 13541 39933 13553 39936
rect 13587 39933 13599 39967
rect 13541 39927 13599 39933
rect 13630 39924 13636 39976
rect 13688 39973 13694 39976
rect 13688 39967 13716 39973
rect 13704 39933 13716 39967
rect 13814 39964 13820 39976
rect 13775 39936 13820 39964
rect 13688 39927 13716 39933
rect 13688 39924 13694 39927
rect 13814 39924 13820 39936
rect 13872 39924 13878 39976
rect 15013 39967 15071 39973
rect 15013 39933 15025 39967
rect 15059 39933 15071 39967
rect 15194 39964 15200 39976
rect 15155 39936 15200 39964
rect 15013 39927 15071 39933
rect 15028 39896 15056 39927
rect 15194 39924 15200 39936
rect 15252 39924 15258 39976
rect 16298 39924 16304 39976
rect 16356 39964 16362 39976
rect 17313 39967 17371 39973
rect 17313 39964 17325 39967
rect 16356 39936 17325 39964
rect 16356 39924 16362 39936
rect 17313 39933 17325 39936
rect 17359 39933 17371 39967
rect 17313 39927 17371 39933
rect 17402 39924 17408 39976
rect 17460 39964 17466 39976
rect 17706 39967 17764 39973
rect 17706 39964 17718 39967
rect 17460 39936 17718 39964
rect 17460 39924 17466 39936
rect 17706 39933 17718 39936
rect 17752 39933 17764 39967
rect 17706 39927 17764 39933
rect 17865 39967 17923 39973
rect 17865 39933 17877 39967
rect 17911 39964 17923 39967
rect 18046 39964 18052 39976
rect 17911 39936 18052 39964
rect 17911 39933 17923 39936
rect 17865 39927 17923 39933
rect 18046 39924 18052 39936
rect 18104 39924 18110 39976
rect 21818 39964 21824 39976
rect 21779 39936 21824 39964
rect 21818 39924 21824 39936
rect 21876 39924 21882 39976
rect 22373 39967 22431 39973
rect 22373 39933 22385 39967
rect 22419 39964 22431 39967
rect 29914 39964 29920 39976
rect 22419 39936 29920 39964
rect 22419 39933 22431 39936
rect 22373 39927 22431 39933
rect 29914 39924 29920 39936
rect 29972 39924 29978 39976
rect 16850 39896 16856 39908
rect 15028 39868 16856 39896
rect 16850 39856 16856 39868
rect 16908 39856 16914 39908
rect 5810 39828 5816 39840
rect 2731 39800 3188 39828
rect 5771 39800 5816 39828
rect 2731 39797 2743 39800
rect 2685 39791 2743 39797
rect 5810 39788 5816 39800
rect 5868 39788 5874 39840
rect 8570 39828 8576 39840
rect 8531 39800 8576 39828
rect 8570 39788 8576 39800
rect 8628 39788 8634 39840
rect 9033 39831 9091 39837
rect 9033 39797 9045 39831
rect 9079 39828 9091 39831
rect 9490 39828 9496 39840
rect 9079 39800 9496 39828
rect 9079 39797 9091 39800
rect 9033 39791 9091 39797
rect 9490 39788 9496 39800
rect 9548 39788 9554 39840
rect 13354 39828 13360 39840
rect 13267 39800 13360 39828
rect 13354 39788 13360 39800
rect 13412 39828 13418 39840
rect 15470 39828 15476 39840
rect 13412 39800 15476 39828
rect 13412 39788 13418 39800
rect 15470 39788 15476 39800
rect 15528 39788 15534 39840
rect 17770 39788 17776 39840
rect 17828 39828 17834 39840
rect 18509 39831 18567 39837
rect 18509 39828 18521 39831
rect 17828 39800 18521 39828
rect 17828 39788 17834 39800
rect 18509 39797 18521 39800
rect 18555 39797 18567 39831
rect 18966 39828 18972 39840
rect 18927 39800 18972 39828
rect 18509 39791 18567 39797
rect 18966 39788 18972 39800
rect 19024 39788 19030 39840
rect 1104 39738 30820 39760
rect 1104 39686 5915 39738
rect 5967 39686 5979 39738
rect 6031 39686 6043 39738
rect 6095 39686 6107 39738
rect 6159 39686 6171 39738
rect 6223 39686 15846 39738
rect 15898 39686 15910 39738
rect 15962 39686 15974 39738
rect 16026 39686 16038 39738
rect 16090 39686 16102 39738
rect 16154 39686 25776 39738
rect 25828 39686 25840 39738
rect 25892 39686 25904 39738
rect 25956 39686 25968 39738
rect 26020 39686 26032 39738
rect 26084 39686 30820 39738
rect 1104 39664 30820 39686
rect 2317 39627 2375 39633
rect 2317 39593 2329 39627
rect 2363 39593 2375 39627
rect 2317 39587 2375 39593
rect 1949 39559 2007 39565
rect 1949 39525 1961 39559
rect 1995 39556 2007 39559
rect 2130 39556 2136 39568
rect 1995 39528 2136 39556
rect 1995 39525 2007 39528
rect 1949 39519 2007 39525
rect 2130 39516 2136 39528
rect 2188 39516 2194 39568
rect 2332 39556 2360 39587
rect 2406 39584 2412 39636
rect 2464 39624 2470 39636
rect 2501 39627 2559 39633
rect 2501 39624 2513 39627
rect 2464 39596 2513 39624
rect 2464 39584 2470 39596
rect 2501 39593 2513 39596
rect 2547 39593 2559 39627
rect 3050 39624 3056 39636
rect 3011 39596 3056 39624
rect 2501 39587 2559 39593
rect 3050 39584 3056 39596
rect 3108 39584 3114 39636
rect 3786 39624 3792 39636
rect 3747 39596 3792 39624
rect 3786 39584 3792 39596
rect 3844 39584 3850 39636
rect 5626 39584 5632 39636
rect 5684 39624 5690 39636
rect 5721 39627 5779 39633
rect 5721 39624 5733 39627
rect 5684 39596 5733 39624
rect 5684 39584 5690 39596
rect 5721 39593 5733 39596
rect 5767 39593 5779 39627
rect 9030 39624 9036 39636
rect 5721 39587 5779 39593
rect 6564 39596 9036 39624
rect 4985 39559 5043 39565
rect 4985 39556 4997 39559
rect 2332 39528 4997 39556
rect 2424 39500 2452 39528
rect 4985 39525 4997 39528
rect 5031 39525 5043 39559
rect 4985 39519 5043 39525
rect 2406 39448 2412 39500
rect 2464 39448 2470 39500
rect 4154 39488 4160 39500
rect 4067 39460 4160 39488
rect 4154 39448 4160 39460
rect 4212 39488 4218 39500
rect 4706 39488 4712 39500
rect 4212 39460 4712 39488
rect 4212 39448 4218 39460
rect 4706 39448 4712 39460
rect 4764 39448 4770 39500
rect 3234 39420 3240 39432
rect 3195 39392 3240 39420
rect 3234 39380 3240 39392
rect 3292 39380 3298 39432
rect 3970 39420 3976 39432
rect 3931 39392 3976 39420
rect 3970 39380 3976 39392
rect 4028 39380 4034 39432
rect 4246 39420 4252 39432
rect 4207 39392 4252 39420
rect 4246 39380 4252 39392
rect 4304 39380 4310 39432
rect 4338 39380 4344 39432
rect 4396 39420 4402 39432
rect 4396 39392 4441 39420
rect 4396 39380 4402 39392
rect 4522 39380 4528 39432
rect 4580 39420 4586 39432
rect 4580 39392 4625 39420
rect 4580 39380 4586 39392
rect 5074 39380 5080 39432
rect 5132 39420 5138 39432
rect 5169 39423 5227 39429
rect 5169 39420 5181 39423
rect 5132 39392 5181 39420
rect 5132 39380 5138 39392
rect 5169 39389 5181 39392
rect 5215 39389 5227 39423
rect 5169 39383 5227 39389
rect 5718 39380 5724 39432
rect 5776 39420 5782 39432
rect 6564 39429 6592 39596
rect 9030 39584 9036 39596
rect 9088 39584 9094 39636
rect 12986 39624 12992 39636
rect 12947 39596 12992 39624
rect 12986 39584 12992 39596
rect 13044 39584 13050 39636
rect 15654 39624 15660 39636
rect 15120 39596 15660 39624
rect 12161 39559 12219 39565
rect 12161 39525 12173 39559
rect 12207 39556 12219 39559
rect 12207 39528 12434 39556
rect 12207 39525 12219 39528
rect 12161 39519 12219 39525
rect 6733 39491 6791 39497
rect 6733 39457 6745 39491
rect 6779 39488 6791 39491
rect 7006 39488 7012 39500
rect 6779 39460 7012 39488
rect 6779 39457 6791 39460
rect 6733 39451 6791 39457
rect 7006 39448 7012 39460
rect 7064 39488 7070 39500
rect 7653 39491 7711 39497
rect 7653 39488 7665 39491
rect 7064 39460 7665 39488
rect 7064 39448 7070 39460
rect 7653 39457 7665 39460
rect 7699 39457 7711 39491
rect 7653 39451 7711 39457
rect 8570 39448 8576 39500
rect 8628 39488 8634 39500
rect 9033 39491 9091 39497
rect 9033 39488 9045 39491
rect 8628 39460 9045 39488
rect 8628 39448 8634 39460
rect 9033 39457 9045 39460
rect 9079 39457 9091 39491
rect 12406 39488 12434 39528
rect 13262 39516 13268 39568
rect 13320 39556 13326 39568
rect 15120 39565 15148 39596
rect 15654 39584 15660 39596
rect 15712 39584 15718 39636
rect 16850 39584 16856 39636
rect 16908 39624 16914 39636
rect 18046 39624 18052 39636
rect 16908 39596 18052 39624
rect 16908 39584 16914 39596
rect 18046 39584 18052 39596
rect 18104 39584 18110 39636
rect 15105 39559 15163 39565
rect 15105 39556 15117 39559
rect 13320 39528 15117 39556
rect 13320 39516 13326 39528
rect 15105 39525 15117 39528
rect 15151 39525 15163 39559
rect 15105 39519 15163 39525
rect 17497 39559 17555 39565
rect 17497 39525 17509 39559
rect 17543 39556 17555 39559
rect 18782 39556 18788 39568
rect 17543 39528 18788 39556
rect 17543 39525 17555 39528
rect 17497 39519 17555 39525
rect 18782 39516 18788 39528
rect 18840 39516 18846 39568
rect 14642 39488 14648 39500
rect 12406 39460 14648 39488
rect 9033 39451 9091 39457
rect 14642 39448 14648 39460
rect 14700 39448 14706 39500
rect 15381 39491 15439 39497
rect 15381 39488 15393 39491
rect 14844 39460 15393 39488
rect 5905 39423 5963 39429
rect 5905 39420 5917 39423
rect 5776 39392 5917 39420
rect 5776 39380 5782 39392
rect 5905 39389 5917 39392
rect 5951 39389 5963 39423
rect 5905 39383 5963 39389
rect 6365 39423 6423 39429
rect 6365 39389 6377 39423
rect 6411 39389 6423 39423
rect 6365 39383 6423 39389
rect 6549 39423 6607 39429
rect 6549 39389 6561 39423
rect 6595 39389 6607 39423
rect 6549 39383 6607 39389
rect 2317 39355 2375 39361
rect 2317 39321 2329 39355
rect 2363 39352 2375 39355
rect 3988 39352 4016 39380
rect 6380 39352 6408 39383
rect 6638 39380 6644 39432
rect 6696 39420 6702 39432
rect 6914 39420 6920 39432
rect 6696 39392 6741 39420
rect 6875 39392 6920 39420
rect 6696 39380 6702 39392
rect 6914 39380 6920 39392
rect 6972 39380 6978 39432
rect 7745 39423 7803 39429
rect 7745 39389 7757 39423
rect 7791 39389 7803 39423
rect 7745 39383 7803 39389
rect 6454 39352 6460 39364
rect 2363 39324 4016 39352
rect 6367 39324 6460 39352
rect 2363 39321 2375 39324
rect 2317 39315 2375 39321
rect 6454 39312 6460 39324
rect 6512 39352 6518 39364
rect 6822 39352 6828 39364
rect 6512 39324 6828 39352
rect 6512 39312 6518 39324
rect 6822 39312 6828 39324
rect 6880 39312 6886 39364
rect 7760 39352 7788 39383
rect 8110 39380 8116 39432
rect 8168 39420 8174 39432
rect 8389 39423 8447 39429
rect 8389 39420 8401 39423
rect 8168 39392 8401 39420
rect 8168 39380 8174 39392
rect 8389 39389 8401 39392
rect 8435 39389 8447 39423
rect 8389 39383 8447 39389
rect 11977 39423 12035 39429
rect 11977 39389 11989 39423
rect 12023 39420 12035 39423
rect 13722 39420 13728 39432
rect 12023 39392 13728 39420
rect 12023 39389 12035 39392
rect 11977 39383 12035 39389
rect 13722 39380 13728 39392
rect 13780 39380 13786 39432
rect 14458 39420 14464 39432
rect 14419 39392 14464 39420
rect 14458 39380 14464 39392
rect 14516 39420 14522 39432
rect 14844 39420 14872 39460
rect 15381 39457 15393 39460
rect 15427 39457 15439 39491
rect 15381 39451 15439 39457
rect 15470 39448 15476 39500
rect 15528 39497 15534 39500
rect 15528 39491 15556 39497
rect 15544 39457 15556 39491
rect 15528 39451 15556 39457
rect 15657 39491 15715 39497
rect 15657 39457 15669 39491
rect 15703 39488 15715 39491
rect 16298 39488 16304 39500
rect 15703 39460 16304 39488
rect 15703 39457 15715 39460
rect 15657 39451 15715 39457
rect 15528 39448 15534 39451
rect 16298 39448 16304 39460
rect 16356 39448 16362 39500
rect 16850 39488 16856 39500
rect 16811 39460 16856 39488
rect 16850 39448 16856 39460
rect 16908 39448 16914 39500
rect 17034 39488 17040 39500
rect 16995 39460 17040 39488
rect 17034 39448 17040 39460
rect 17092 39448 17098 39500
rect 18138 39420 18144 39432
rect 14516 39392 14872 39420
rect 18099 39392 18144 39420
rect 14516 39380 14522 39392
rect 18138 39380 18144 39392
rect 18196 39380 18202 39432
rect 19426 39380 19432 39432
rect 19484 39420 19490 39432
rect 19797 39423 19855 39429
rect 19797 39420 19809 39423
rect 19484 39392 19809 39420
rect 19484 39380 19490 39392
rect 19797 39389 19809 39392
rect 19843 39389 19855 39423
rect 30098 39420 30104 39432
rect 30059 39392 30104 39420
rect 19797 39383 19855 39389
rect 30098 39380 30104 39392
rect 30156 39380 30162 39432
rect 8478 39352 8484 39364
rect 6932 39324 8484 39352
rect 6638 39244 6644 39296
rect 6696 39284 6702 39296
rect 6932 39284 6960 39324
rect 8478 39312 8484 39324
rect 8536 39312 8542 39364
rect 9306 39361 9312 39364
rect 9300 39315 9312 39361
rect 9364 39352 9370 39364
rect 12618 39352 12624 39364
rect 9364 39324 9400 39352
rect 12579 39324 12624 39352
rect 9306 39312 9312 39315
rect 9364 39312 9370 39324
rect 12618 39312 12624 39324
rect 12676 39312 12682 39364
rect 12805 39355 12863 39361
rect 12805 39321 12817 39355
rect 12851 39321 12863 39355
rect 12805 39315 12863 39321
rect 16301 39355 16359 39361
rect 16301 39321 16313 39355
rect 16347 39352 16359 39355
rect 17129 39355 17187 39361
rect 17129 39352 17141 39355
rect 16347 39324 17141 39352
rect 16347 39321 16359 39324
rect 16301 39315 16359 39321
rect 17129 39321 17141 39324
rect 17175 39321 17187 39355
rect 17129 39315 17187 39321
rect 7098 39284 7104 39296
rect 6696 39256 6960 39284
rect 7059 39256 7104 39284
rect 6696 39244 6702 39256
rect 7098 39244 7104 39256
rect 7156 39244 7162 39296
rect 8202 39284 8208 39296
rect 8163 39256 8208 39284
rect 8202 39244 8208 39256
rect 8260 39244 8266 39296
rect 9122 39244 9128 39296
rect 9180 39284 9186 39296
rect 10413 39287 10471 39293
rect 10413 39284 10425 39287
rect 9180 39256 10425 39284
rect 9180 39244 9186 39256
rect 10413 39253 10425 39256
rect 10459 39253 10471 39287
rect 12820 39284 12848 39315
rect 17862 39312 17868 39364
rect 17920 39352 17926 39364
rect 19610 39352 19616 39364
rect 17920 39324 19616 39352
rect 17920 39312 17926 39324
rect 19610 39312 19616 39324
rect 19668 39312 19674 39364
rect 14826 39284 14832 39296
rect 12820 39256 14832 39284
rect 10413 39247 10471 39253
rect 14826 39244 14832 39256
rect 14884 39244 14890 39296
rect 17678 39244 17684 39296
rect 17736 39284 17742 39296
rect 17957 39287 18015 39293
rect 17957 39284 17969 39287
rect 17736 39256 17969 39284
rect 17736 39244 17742 39256
rect 17957 39253 17969 39256
rect 18003 39253 18015 39287
rect 17957 39247 18015 39253
rect 19981 39287 20039 39293
rect 19981 39253 19993 39287
rect 20027 39284 20039 39287
rect 20254 39284 20260 39296
rect 20027 39256 20260 39284
rect 20027 39253 20039 39256
rect 19981 39247 20039 39253
rect 20254 39244 20260 39256
rect 20312 39244 20318 39296
rect 29914 39284 29920 39296
rect 29875 39256 29920 39284
rect 29914 39244 29920 39256
rect 29972 39244 29978 39296
rect 1104 39194 30820 39216
rect 1104 39142 10880 39194
rect 10932 39142 10944 39194
rect 10996 39142 11008 39194
rect 11060 39142 11072 39194
rect 11124 39142 11136 39194
rect 11188 39142 20811 39194
rect 20863 39142 20875 39194
rect 20927 39142 20939 39194
rect 20991 39142 21003 39194
rect 21055 39142 21067 39194
rect 21119 39142 30820 39194
rect 1104 39120 30820 39142
rect 2593 39083 2651 39089
rect 2593 39049 2605 39083
rect 2639 39080 2651 39083
rect 3602 39080 3608 39092
rect 2639 39052 3608 39080
rect 2639 39049 2651 39052
rect 2593 39043 2651 39049
rect 3602 39040 3608 39052
rect 3660 39040 3666 39092
rect 5169 39083 5227 39089
rect 5169 39049 5181 39083
rect 5215 39080 5227 39083
rect 5718 39080 5724 39092
rect 5215 39052 5724 39080
rect 5215 39049 5227 39052
rect 5169 39043 5227 39049
rect 5718 39040 5724 39052
rect 5776 39040 5782 39092
rect 6914 39040 6920 39092
rect 6972 39080 6978 39092
rect 7929 39083 7987 39089
rect 7929 39080 7941 39083
rect 6972 39052 7941 39080
rect 6972 39040 6978 39052
rect 7929 39049 7941 39052
rect 7975 39049 7987 39083
rect 9306 39080 9312 39092
rect 9267 39052 9312 39080
rect 7929 39043 7987 39049
rect 9306 39040 9312 39052
rect 9364 39040 9370 39092
rect 14369 39083 14427 39089
rect 14369 39049 14381 39083
rect 14415 39080 14427 39083
rect 15194 39080 15200 39092
rect 14415 39052 15200 39080
rect 14415 39049 14427 39052
rect 14369 39043 14427 39049
rect 15194 39040 15200 39052
rect 15252 39040 15258 39092
rect 16117 39083 16175 39089
rect 16117 39049 16129 39083
rect 16163 39080 16175 39083
rect 16206 39080 16212 39092
rect 16163 39052 16212 39080
rect 16163 39049 16175 39052
rect 16117 39043 16175 39049
rect 16206 39040 16212 39052
rect 16264 39040 16270 39092
rect 16853 39083 16911 39089
rect 16853 39049 16865 39083
rect 16899 39080 16911 39083
rect 17402 39080 17408 39092
rect 16899 39052 17408 39080
rect 16899 39049 16911 39052
rect 16853 39043 16911 39049
rect 17402 39040 17408 39052
rect 17460 39040 17466 39092
rect 17678 39080 17684 39092
rect 17639 39052 17684 39080
rect 17678 39040 17684 39052
rect 17736 39040 17742 39092
rect 17770 39040 17776 39092
rect 17828 39080 17834 39092
rect 18782 39080 18788 39092
rect 17828 39052 17873 39080
rect 18743 39052 18788 39080
rect 17828 39040 17834 39052
rect 18782 39040 18788 39052
rect 18840 39040 18846 39092
rect 18877 39083 18935 39089
rect 18877 39049 18889 39083
rect 18923 39080 18935 39083
rect 18966 39080 18972 39092
rect 18923 39052 18972 39080
rect 18923 39049 18935 39052
rect 18877 39043 18935 39049
rect 18966 39040 18972 39052
rect 19024 39040 19030 39092
rect 19610 39040 19616 39092
rect 19668 39080 19674 39092
rect 19981 39083 20039 39089
rect 19981 39080 19993 39083
rect 19668 39052 19993 39080
rect 19668 39040 19674 39052
rect 19981 39049 19993 39052
rect 20027 39049 20039 39083
rect 21910 39080 21916 39092
rect 21871 39052 21916 39080
rect 19981 39043 20039 39049
rect 21910 39040 21916 39052
rect 21968 39040 21974 39092
rect 2409 39015 2467 39021
rect 2409 38981 2421 39015
rect 2455 39012 2467 39015
rect 2498 39012 2504 39024
rect 2455 38984 2504 39012
rect 2455 38981 2467 38984
rect 2409 38975 2467 38981
rect 2498 38972 2504 38984
rect 2556 38972 2562 39024
rect 8018 39012 8024 39024
rect 5000 38984 8024 39012
rect 1397 38947 1455 38953
rect 1397 38913 1409 38947
rect 1443 38944 1455 38947
rect 1854 38944 1860 38956
rect 1443 38916 1860 38944
rect 1443 38913 1455 38916
rect 1397 38907 1455 38913
rect 1854 38904 1860 38916
rect 1912 38904 1918 38956
rect 2041 38947 2099 38953
rect 2041 38913 2053 38947
rect 2087 38944 2099 38947
rect 2130 38944 2136 38956
rect 2087 38916 2136 38944
rect 2087 38913 2099 38916
rect 2041 38907 2099 38913
rect 2130 38904 2136 38916
rect 2188 38904 2194 38956
rect 2774 38904 2780 38956
rect 2832 38944 2838 38956
rect 3050 38944 3056 38956
rect 2832 38916 3056 38944
rect 2832 38904 2838 38916
rect 3050 38904 3056 38916
rect 3108 38904 3114 38956
rect 3237 38947 3295 38953
rect 3237 38913 3249 38947
rect 3283 38944 3295 38947
rect 3510 38944 3516 38956
rect 3283 38916 3516 38944
rect 3283 38913 3295 38916
rect 3237 38907 3295 38913
rect 3510 38904 3516 38916
rect 3568 38904 3574 38956
rect 3970 38944 3976 38956
rect 3931 38916 3976 38944
rect 3970 38904 3976 38916
rect 4028 38904 4034 38956
rect 5000 38953 5028 38984
rect 8018 38972 8024 38984
rect 8076 38972 8082 39024
rect 15749 39015 15807 39021
rect 15749 39012 15761 39015
rect 15212 38984 15761 39012
rect 4985 38947 5043 38953
rect 4985 38913 4997 38947
rect 5031 38913 5043 38947
rect 5626 38944 5632 38956
rect 5587 38916 5632 38944
rect 4985 38907 5043 38913
rect 5626 38904 5632 38916
rect 5684 38904 5690 38956
rect 5810 38904 5816 38956
rect 5868 38944 5874 38956
rect 6549 38947 6607 38953
rect 6549 38944 6561 38947
rect 5868 38916 6561 38944
rect 5868 38904 5874 38916
rect 6549 38913 6561 38916
rect 6595 38913 6607 38947
rect 6549 38907 6607 38913
rect 6816 38947 6874 38953
rect 6816 38913 6828 38947
rect 6862 38944 6874 38947
rect 7098 38944 7104 38956
rect 6862 38916 7104 38944
rect 6862 38913 6874 38916
rect 6816 38907 6874 38913
rect 7098 38904 7104 38916
rect 7156 38904 7162 38956
rect 8570 38944 8576 38956
rect 8531 38916 8576 38944
rect 8570 38904 8576 38916
rect 8628 38904 8634 38956
rect 8754 38944 8760 38956
rect 8715 38916 8760 38944
rect 8754 38904 8760 38916
rect 8812 38904 8818 38956
rect 9122 38944 9128 38956
rect 9083 38916 9128 38944
rect 9122 38904 9128 38916
rect 9180 38904 9186 38956
rect 10321 38947 10379 38953
rect 10321 38913 10333 38947
rect 10367 38944 10379 38947
rect 11422 38944 11428 38956
rect 10367 38916 11428 38944
rect 10367 38913 10379 38916
rect 10321 38907 10379 38913
rect 11422 38904 11428 38916
rect 11480 38904 11486 38956
rect 12526 38944 12532 38956
rect 12487 38916 12532 38944
rect 12526 38904 12532 38916
rect 12584 38904 12590 38956
rect 13446 38904 13452 38956
rect 13504 38944 13510 38956
rect 13504 38916 13549 38944
rect 13504 38904 13510 38916
rect 14826 38904 14832 38956
rect 14884 38944 14890 38956
rect 15212 38953 15240 38984
rect 15749 38981 15761 38984
rect 15795 39012 15807 39015
rect 16574 39012 16580 39024
rect 15795 38984 16580 39012
rect 15795 38981 15807 38984
rect 15749 38975 15807 38981
rect 16574 38972 16580 38984
rect 16632 38972 16638 39024
rect 15105 38947 15163 38953
rect 15105 38944 15117 38947
rect 14884 38916 15117 38944
rect 14884 38904 14890 38916
rect 15105 38913 15117 38916
rect 15151 38913 15163 38947
rect 15105 38907 15163 38913
rect 15197 38947 15255 38953
rect 15197 38913 15209 38947
rect 15243 38913 15255 38947
rect 15197 38907 15255 38913
rect 15654 38904 15660 38956
rect 15712 38944 15718 38956
rect 15933 38947 15991 38953
rect 15933 38944 15945 38947
rect 15712 38916 15945 38944
rect 15712 38904 15718 38916
rect 15933 38913 15945 38916
rect 15979 38913 15991 38947
rect 15933 38907 15991 38913
rect 16669 38947 16727 38953
rect 16669 38913 16681 38947
rect 16715 38944 16727 38947
rect 17126 38944 17132 38956
rect 16715 38916 17132 38944
rect 16715 38913 16727 38916
rect 16669 38907 16727 38913
rect 17126 38904 17132 38916
rect 17184 38904 17190 38956
rect 20070 38944 20076 38956
rect 20031 38916 20076 38944
rect 20070 38904 20076 38916
rect 20128 38904 20134 38956
rect 22094 38944 22100 38956
rect 22055 38916 22100 38944
rect 22094 38904 22100 38916
rect 22152 38904 22158 38956
rect 8849 38879 8907 38885
rect 8849 38845 8861 38879
rect 8895 38845 8907 38879
rect 8849 38839 8907 38845
rect 8941 38879 8999 38885
rect 8941 38845 8953 38879
rect 8987 38876 8999 38879
rect 9306 38876 9312 38888
rect 8987 38848 9312 38876
rect 8987 38845 8999 38848
rect 8941 38839 8999 38845
rect 2774 38808 2780 38820
rect 2148 38780 2780 38808
rect 1581 38743 1639 38749
rect 1581 38709 1593 38743
rect 1627 38740 1639 38743
rect 2148 38740 2176 38780
rect 2774 38768 2780 38780
rect 2832 38768 2838 38820
rect 2406 38740 2412 38752
rect 1627 38712 2176 38740
rect 2367 38712 2412 38740
rect 1627 38709 1639 38712
rect 1581 38703 1639 38709
rect 2406 38700 2412 38712
rect 2464 38700 2470 38752
rect 2866 38700 2872 38752
rect 2924 38740 2930 38752
rect 3053 38743 3111 38749
rect 3053 38740 3065 38743
rect 2924 38712 3065 38740
rect 2924 38700 2930 38712
rect 3053 38709 3065 38712
rect 3099 38709 3111 38743
rect 4154 38740 4160 38752
rect 4115 38712 4160 38740
rect 3053 38703 3111 38709
rect 4154 38700 4160 38712
rect 4212 38700 4218 38752
rect 5721 38743 5779 38749
rect 5721 38709 5733 38743
rect 5767 38740 5779 38743
rect 6730 38740 6736 38752
rect 5767 38712 6736 38740
rect 5767 38709 5779 38712
rect 5721 38703 5779 38709
rect 6730 38700 6736 38712
rect 6788 38740 6794 38752
rect 8864 38740 8892 38839
rect 9306 38836 9312 38848
rect 9364 38836 9370 38888
rect 12618 38836 12624 38888
rect 12676 38876 12682 38888
rect 12713 38879 12771 38885
rect 12713 38876 12725 38879
rect 12676 38848 12725 38876
rect 12676 38836 12682 38848
rect 12713 38845 12725 38848
rect 12759 38876 12771 38879
rect 13262 38876 13268 38888
rect 12759 38848 13268 38876
rect 12759 38845 12771 38848
rect 12713 38839 12771 38845
rect 13262 38836 13268 38848
rect 13320 38836 13326 38888
rect 13538 38836 13544 38888
rect 13596 38885 13602 38888
rect 13596 38879 13624 38885
rect 13612 38845 13624 38879
rect 13596 38839 13624 38845
rect 13725 38879 13783 38885
rect 13725 38845 13737 38879
rect 13771 38876 13783 38879
rect 13906 38876 13912 38888
rect 13771 38848 13912 38876
rect 13771 38845 13783 38848
rect 13725 38839 13783 38845
rect 13596 38836 13602 38839
rect 13906 38836 13912 38848
rect 13964 38876 13970 38888
rect 16298 38876 16304 38888
rect 13964 38848 16304 38876
rect 13964 38836 13970 38848
rect 16298 38836 16304 38848
rect 16356 38836 16362 38888
rect 17954 38876 17960 38888
rect 17915 38848 17960 38876
rect 17954 38836 17960 38848
rect 18012 38876 18018 38888
rect 18601 38879 18659 38885
rect 18601 38876 18613 38879
rect 18012 38848 18613 38876
rect 18012 38836 18018 38848
rect 18601 38845 18613 38848
rect 18647 38876 18659 38879
rect 19797 38879 19855 38885
rect 19797 38876 19809 38879
rect 18647 38848 19809 38876
rect 18647 38845 18659 38848
rect 18601 38839 18659 38845
rect 19797 38845 19809 38848
rect 19843 38845 19855 38879
rect 19797 38839 19855 38845
rect 22281 38879 22339 38885
rect 22281 38845 22293 38879
rect 22327 38876 22339 38879
rect 29914 38876 29920 38888
rect 22327 38848 29920 38876
rect 22327 38845 22339 38848
rect 22281 38839 22339 38845
rect 29914 38836 29920 38848
rect 29972 38836 29978 38888
rect 13170 38808 13176 38820
rect 13131 38780 13176 38808
rect 13170 38768 13176 38780
rect 13228 38768 13234 38820
rect 9214 38740 9220 38752
rect 6788 38712 9220 38740
rect 6788 38700 6794 38712
rect 9214 38700 9220 38712
rect 9272 38700 9278 38752
rect 10505 38743 10563 38749
rect 10505 38709 10517 38743
rect 10551 38740 10563 38743
rect 10594 38740 10600 38752
rect 10551 38712 10600 38740
rect 10551 38709 10563 38712
rect 10505 38703 10563 38709
rect 10594 38700 10600 38712
rect 10652 38700 10658 38752
rect 16758 38700 16764 38752
rect 16816 38740 16822 38752
rect 17313 38743 17371 38749
rect 17313 38740 17325 38743
rect 16816 38712 17325 38740
rect 16816 38700 16822 38712
rect 17313 38709 17325 38712
rect 17359 38709 17371 38743
rect 17313 38703 17371 38709
rect 19150 38700 19156 38752
rect 19208 38740 19214 38752
rect 19245 38743 19303 38749
rect 19245 38740 19257 38743
rect 19208 38712 19257 38740
rect 19208 38700 19214 38712
rect 19245 38709 19257 38712
rect 19291 38709 19303 38743
rect 19245 38703 19303 38709
rect 20441 38743 20499 38749
rect 20441 38709 20453 38743
rect 20487 38740 20499 38743
rect 21358 38740 21364 38752
rect 20487 38712 21364 38740
rect 20487 38709 20499 38712
rect 20441 38703 20499 38709
rect 21358 38700 21364 38712
rect 21416 38700 21422 38752
rect 1104 38650 30820 38672
rect 1104 38598 5915 38650
rect 5967 38598 5979 38650
rect 6031 38598 6043 38650
rect 6095 38598 6107 38650
rect 6159 38598 6171 38650
rect 6223 38598 15846 38650
rect 15898 38598 15910 38650
rect 15962 38598 15974 38650
rect 16026 38598 16038 38650
rect 16090 38598 16102 38650
rect 16154 38598 25776 38650
rect 25828 38598 25840 38650
rect 25892 38598 25904 38650
rect 25956 38598 25968 38650
rect 26020 38598 26032 38650
rect 26084 38598 30820 38650
rect 1104 38576 30820 38598
rect 2317 38539 2375 38545
rect 2317 38505 2329 38539
rect 2363 38536 2375 38539
rect 2406 38536 2412 38548
rect 2363 38508 2412 38536
rect 2363 38505 2375 38508
rect 2317 38499 2375 38505
rect 2406 38496 2412 38508
rect 2464 38496 2470 38548
rect 2501 38539 2559 38545
rect 2501 38505 2513 38539
rect 2547 38536 2559 38539
rect 2590 38536 2596 38548
rect 2547 38508 2596 38536
rect 2547 38505 2559 38508
rect 2501 38499 2559 38505
rect 2590 38496 2596 38508
rect 2648 38496 2654 38548
rect 4246 38496 4252 38548
rect 4304 38536 4310 38548
rect 6963 38539 7021 38545
rect 6963 38536 6975 38539
rect 4304 38508 6975 38536
rect 4304 38496 4310 38508
rect 6963 38505 6975 38508
rect 7009 38505 7021 38539
rect 6963 38499 7021 38505
rect 8294 38496 8300 38548
rect 8352 38536 8358 38548
rect 8389 38539 8447 38545
rect 8389 38536 8401 38539
rect 8352 38508 8401 38536
rect 8352 38496 8358 38508
rect 8389 38505 8401 38508
rect 8435 38505 8447 38539
rect 9674 38536 9680 38548
rect 9635 38508 9680 38536
rect 8389 38499 8447 38505
rect 9674 38496 9680 38508
rect 9732 38496 9738 38548
rect 13722 38496 13728 38548
rect 13780 38536 13786 38548
rect 14093 38539 14151 38545
rect 14093 38536 14105 38539
rect 13780 38508 14105 38536
rect 13780 38496 13786 38508
rect 14093 38505 14105 38508
rect 14139 38505 14151 38539
rect 14093 38499 14151 38505
rect 18138 38496 18144 38548
rect 18196 38536 18202 38548
rect 18233 38539 18291 38545
rect 18233 38536 18245 38539
rect 18196 38508 18245 38536
rect 18196 38496 18202 38508
rect 18233 38505 18245 38508
rect 18279 38505 18291 38539
rect 18233 38499 18291 38505
rect 19334 38496 19340 38548
rect 19392 38536 19398 38548
rect 19613 38539 19671 38545
rect 19613 38536 19625 38539
rect 19392 38508 19625 38536
rect 19392 38496 19398 38508
rect 19613 38505 19625 38508
rect 19659 38505 19671 38539
rect 20070 38536 20076 38548
rect 20031 38508 20076 38536
rect 19613 38499 19671 38505
rect 20070 38496 20076 38508
rect 20128 38496 20134 38548
rect 1949 38471 2007 38477
rect 1949 38437 1961 38471
rect 1995 38468 2007 38471
rect 2130 38468 2136 38480
rect 1995 38440 2136 38468
rect 1995 38437 2007 38440
rect 1949 38431 2007 38437
rect 2130 38428 2136 38440
rect 2188 38428 2194 38480
rect 9122 38468 9128 38480
rect 2332 38440 9128 38468
rect 2332 38273 2360 38440
rect 9122 38428 9128 38440
rect 9180 38428 9186 38480
rect 12345 38471 12403 38477
rect 12345 38437 12357 38471
rect 12391 38468 12403 38471
rect 13262 38468 13268 38480
rect 12391 38440 13268 38468
rect 12391 38437 12403 38440
rect 12345 38431 12403 38437
rect 13262 38428 13268 38440
rect 13320 38428 13326 38480
rect 13354 38428 13360 38480
rect 13412 38428 13418 38480
rect 2498 38360 2504 38412
rect 2556 38400 2562 38412
rect 4157 38403 4215 38409
rect 2556 38372 4016 38400
rect 2556 38360 2562 38372
rect 2958 38332 2964 38344
rect 2919 38304 2964 38332
rect 2958 38292 2964 38304
rect 3016 38292 3022 38344
rect 3988 38341 4016 38372
rect 4157 38369 4169 38403
rect 4203 38400 4215 38403
rect 4706 38400 4712 38412
rect 4203 38372 4712 38400
rect 4203 38369 4215 38372
rect 4157 38363 4215 38369
rect 4706 38360 4712 38372
rect 4764 38400 4770 38412
rect 5721 38403 5779 38409
rect 5721 38400 5733 38403
rect 4764 38372 5733 38400
rect 4764 38360 4770 38372
rect 5721 38369 5733 38372
rect 5767 38369 5779 38403
rect 6730 38400 6736 38412
rect 6691 38372 6736 38400
rect 5721 38363 5779 38369
rect 6730 38360 6736 38372
rect 6788 38360 6794 38412
rect 9214 38400 9220 38412
rect 9175 38372 9220 38400
rect 9214 38360 9220 38372
rect 9272 38360 9278 38412
rect 13081 38403 13139 38409
rect 13081 38369 13093 38403
rect 13127 38400 13139 38403
rect 13372 38400 13400 38428
rect 13127 38372 13400 38400
rect 13449 38403 13507 38409
rect 13127 38369 13139 38372
rect 13081 38363 13139 38369
rect 13449 38369 13461 38403
rect 13495 38400 13507 38403
rect 14366 38400 14372 38412
rect 13495 38372 14372 38400
rect 13495 38369 13507 38372
rect 13449 38363 13507 38369
rect 14366 38360 14372 38372
rect 14424 38400 14430 38412
rect 15013 38403 15071 38409
rect 15013 38400 15025 38403
rect 14424 38372 15025 38400
rect 14424 38360 14430 38372
rect 15013 38369 15025 38372
rect 15059 38369 15071 38403
rect 15013 38363 15071 38369
rect 3973 38335 4031 38341
rect 3973 38301 3985 38335
rect 4019 38301 4031 38335
rect 4246 38332 4252 38344
rect 4207 38304 4252 38332
rect 3973 38295 4031 38301
rect 4246 38292 4252 38304
rect 4304 38292 4310 38344
rect 4341 38335 4399 38341
rect 4341 38301 4353 38335
rect 4387 38301 4399 38335
rect 4341 38295 4399 38301
rect 4525 38335 4583 38341
rect 4525 38301 4537 38335
rect 4571 38332 4583 38335
rect 4614 38332 4620 38344
rect 4571 38304 4620 38332
rect 4571 38301 4583 38304
rect 4525 38295 4583 38301
rect 2317 38267 2375 38273
rect 2317 38233 2329 38267
rect 2363 38233 2375 38267
rect 2317 38227 2375 38233
rect 3142 38196 3148 38208
rect 3103 38168 3148 38196
rect 3142 38156 3148 38168
rect 3200 38156 3206 38208
rect 3786 38196 3792 38208
rect 3747 38168 3792 38196
rect 3786 38156 3792 38168
rect 3844 38156 3850 38208
rect 4264 38196 4292 38292
rect 4356 38264 4384 38295
rect 4614 38292 4620 38304
rect 4672 38292 4678 38344
rect 5445 38335 5503 38341
rect 5445 38301 5457 38335
rect 5491 38301 5503 38335
rect 5445 38295 5503 38301
rect 4890 38264 4896 38276
rect 4356 38236 4896 38264
rect 4890 38224 4896 38236
rect 4948 38224 4954 38276
rect 5460 38264 5488 38295
rect 8018 38292 8024 38344
rect 8076 38332 8082 38344
rect 8205 38335 8263 38341
rect 8205 38332 8217 38335
rect 8076 38304 8217 38332
rect 8076 38292 8082 38304
rect 8205 38301 8217 38304
rect 8251 38301 8263 38335
rect 8205 38295 8263 38301
rect 8570 38292 8576 38344
rect 8628 38332 8634 38344
rect 8941 38335 8999 38341
rect 8941 38332 8953 38335
rect 8628 38304 8953 38332
rect 8628 38292 8634 38304
rect 8941 38301 8953 38304
rect 8987 38301 8999 38335
rect 8941 38295 8999 38301
rect 5626 38264 5632 38276
rect 5460 38236 5632 38264
rect 5626 38224 5632 38236
rect 5684 38264 5690 38276
rect 8956 38264 8984 38295
rect 9030 38292 9036 38344
rect 9088 38332 9094 38344
rect 9125 38335 9183 38341
rect 9125 38332 9137 38335
rect 9088 38304 9137 38332
rect 9088 38292 9094 38304
rect 9125 38301 9137 38304
rect 9171 38301 9183 38335
rect 9306 38332 9312 38344
rect 9267 38304 9312 38332
rect 9125 38295 9183 38301
rect 9306 38292 9312 38304
rect 9364 38292 9370 38344
rect 9490 38332 9496 38344
rect 9451 38304 9496 38332
rect 9490 38292 9496 38304
rect 9548 38292 9554 38344
rect 10410 38332 10416 38344
rect 10371 38304 10416 38332
rect 10410 38292 10416 38304
rect 10468 38292 10474 38344
rect 11057 38335 11115 38341
rect 11057 38332 11069 38335
rect 10612 38304 11069 38332
rect 9674 38264 9680 38276
rect 5684 38236 8340 38264
rect 8956 38236 9680 38264
rect 5684 38224 5690 38236
rect 4522 38196 4528 38208
rect 4264 38168 4528 38196
rect 4522 38156 4528 38168
rect 4580 38156 4586 38208
rect 4908 38196 4936 38224
rect 7558 38196 7564 38208
rect 4908 38168 7564 38196
rect 7558 38156 7564 38168
rect 7616 38156 7622 38208
rect 8312 38196 8340 38236
rect 9674 38224 9680 38236
rect 9732 38224 9738 38276
rect 9306 38196 9312 38208
rect 8312 38168 9312 38196
rect 9306 38156 9312 38168
rect 9364 38156 9370 38208
rect 10612 38205 10640 38304
rect 11057 38301 11069 38304
rect 11103 38301 11115 38335
rect 11057 38295 11115 38301
rect 12161 38335 12219 38341
rect 12161 38301 12173 38335
rect 12207 38332 12219 38335
rect 12710 38332 12716 38344
rect 12207 38304 12716 38332
rect 12207 38301 12219 38304
rect 12161 38295 12219 38301
rect 12710 38292 12716 38304
rect 12768 38292 12774 38344
rect 13354 38332 13360 38344
rect 13315 38304 13360 38332
rect 13354 38292 13360 38304
rect 13412 38292 13418 38344
rect 14274 38332 14280 38344
rect 14235 38304 14280 38332
rect 14274 38292 14280 38304
rect 14332 38292 14338 38344
rect 14461 38335 14519 38341
rect 14461 38301 14473 38335
rect 14507 38301 14519 38335
rect 14918 38332 14924 38344
rect 14879 38304 14924 38332
rect 14461 38295 14519 38301
rect 12805 38267 12863 38273
rect 12805 38233 12817 38267
rect 12851 38264 12863 38267
rect 13538 38264 13544 38276
rect 12851 38236 13544 38264
rect 12851 38233 12863 38236
rect 12805 38227 12863 38233
rect 13538 38224 13544 38236
rect 13596 38224 13602 38276
rect 10597 38199 10655 38205
rect 10597 38165 10609 38199
rect 10643 38165 10655 38199
rect 10597 38159 10655 38165
rect 11241 38199 11299 38205
rect 11241 38165 11253 38199
rect 11287 38196 11299 38199
rect 11514 38196 11520 38208
rect 11287 38168 11520 38196
rect 11287 38165 11299 38168
rect 11241 38159 11299 38165
rect 11514 38156 11520 38168
rect 11572 38156 11578 38208
rect 13262 38156 13268 38208
rect 13320 38196 13326 38208
rect 14476 38196 14504 38295
rect 14918 38292 14924 38304
rect 14976 38292 14982 38344
rect 15102 38332 15108 38344
rect 15063 38304 15108 38332
rect 15102 38292 15108 38304
rect 15160 38292 15166 38344
rect 17770 38292 17776 38344
rect 17828 38332 17834 38344
rect 17865 38335 17923 38341
rect 17865 38332 17877 38335
rect 17828 38304 17877 38332
rect 17828 38292 17834 38304
rect 17865 38301 17877 38304
rect 17911 38301 17923 38335
rect 17865 38295 17923 38301
rect 18782 38292 18788 38344
rect 18840 38332 18846 38344
rect 19245 38335 19303 38341
rect 19245 38332 19257 38335
rect 18840 38304 19257 38332
rect 18840 38292 18846 38304
rect 19245 38301 19257 38304
rect 19291 38301 19303 38335
rect 20254 38332 20260 38344
rect 20215 38304 20260 38332
rect 19245 38295 19303 38301
rect 20254 38292 20260 38304
rect 20312 38292 20318 38344
rect 18049 38267 18107 38273
rect 18049 38233 18061 38267
rect 18095 38264 18107 38267
rect 19426 38264 19432 38276
rect 18095 38236 19432 38264
rect 18095 38233 18107 38236
rect 18049 38227 18107 38233
rect 19426 38224 19432 38236
rect 19484 38224 19490 38276
rect 13320 38168 14504 38196
rect 13320 38156 13326 38168
rect 1104 38106 30820 38128
rect 1104 38054 10880 38106
rect 10932 38054 10944 38106
rect 10996 38054 11008 38106
rect 11060 38054 11072 38106
rect 11124 38054 11136 38106
rect 11188 38054 20811 38106
rect 20863 38054 20875 38106
rect 20927 38054 20939 38106
rect 20991 38054 21003 38106
rect 21055 38054 21067 38106
rect 21119 38054 30820 38106
rect 1104 38032 30820 38054
rect 2317 37995 2375 38001
rect 2317 37961 2329 37995
rect 2363 37992 2375 37995
rect 2498 37992 2504 38004
rect 2363 37964 2504 37992
rect 2363 37961 2375 37964
rect 2317 37955 2375 37961
rect 2498 37952 2504 37964
rect 2556 37952 2562 38004
rect 7561 37995 7619 38001
rect 7561 37992 7573 37995
rect 2746 37964 7573 37992
rect 1673 37859 1731 37865
rect 1673 37825 1685 37859
rect 1719 37856 1731 37859
rect 2746 37856 2774 37964
rect 7561 37961 7573 37964
rect 7607 37961 7619 37995
rect 13357 37995 13415 38001
rect 7561 37955 7619 37961
rect 8036 37964 12434 37992
rect 3452 37927 3510 37933
rect 3452 37893 3464 37927
rect 3498 37924 3510 37927
rect 3786 37924 3792 37936
rect 3498 37896 3792 37924
rect 3498 37893 3510 37896
rect 3452 37887 3510 37893
rect 3786 37884 3792 37896
rect 3844 37884 3850 37936
rect 7006 37924 7012 37936
rect 6748 37896 7012 37924
rect 4154 37856 4160 37868
rect 1719 37828 2774 37856
rect 4115 37828 4160 37856
rect 1719 37825 1731 37828
rect 1673 37819 1731 37825
rect 4154 37816 4160 37828
rect 4212 37816 4218 37868
rect 4430 37865 4436 37868
rect 4424 37819 4436 37865
rect 4488 37856 4494 37868
rect 4488 37828 4524 37856
rect 4430 37816 4436 37819
rect 4488 37816 4494 37828
rect 6362 37816 6368 37868
rect 6420 37856 6426 37868
rect 6748 37865 6776 37896
rect 7006 37884 7012 37896
rect 7064 37884 7070 37936
rect 6549 37859 6607 37865
rect 6549 37856 6561 37859
rect 6420 37828 6561 37856
rect 6420 37816 6426 37828
rect 6549 37825 6561 37828
rect 6595 37825 6607 37859
rect 6549 37819 6607 37825
rect 6733 37859 6791 37865
rect 6733 37825 6745 37859
rect 6779 37825 6791 37859
rect 6733 37819 6791 37825
rect 6917 37859 6975 37865
rect 6917 37825 6929 37859
rect 6963 37825 6975 37859
rect 6917 37819 6975 37825
rect 3694 37788 3700 37800
rect 3655 37760 3700 37788
rect 3694 37748 3700 37760
rect 3752 37748 3758 37800
rect 6638 37748 6644 37800
rect 6696 37788 6702 37800
rect 6825 37791 6883 37797
rect 6825 37788 6837 37791
rect 6696 37760 6837 37788
rect 6696 37748 6702 37760
rect 6825 37757 6837 37760
rect 6871 37757 6883 37791
rect 6932 37788 6960 37819
rect 7098 37816 7104 37868
rect 7156 37856 7162 37868
rect 7742 37856 7748 37868
rect 7156 37828 7201 37856
rect 7703 37828 7748 37856
rect 7156 37816 7162 37828
rect 7742 37816 7748 37828
rect 7800 37816 7806 37868
rect 7926 37788 7932 37800
rect 6932 37760 7932 37788
rect 6825 37751 6883 37757
rect 5626 37680 5632 37732
rect 5684 37720 5690 37732
rect 6840 37720 6868 37751
rect 7926 37748 7932 37760
rect 7984 37748 7990 37800
rect 8036 37720 8064 37964
rect 10318 37924 10324 37936
rect 10244 37896 10324 37924
rect 8202 37856 8208 37868
rect 8163 37828 8208 37856
rect 8202 37816 8208 37828
rect 8260 37816 8266 37868
rect 8472 37859 8530 37865
rect 8472 37825 8484 37859
rect 8518 37856 8530 37859
rect 8938 37856 8944 37868
rect 8518 37828 8944 37856
rect 8518 37825 8530 37828
rect 8472 37819 8530 37825
rect 8938 37816 8944 37828
rect 8996 37816 9002 37868
rect 10045 37859 10103 37865
rect 10045 37825 10057 37859
rect 10091 37856 10103 37859
rect 10134 37856 10140 37868
rect 10091 37828 10140 37856
rect 10091 37825 10103 37828
rect 10045 37819 10103 37825
rect 10134 37816 10140 37828
rect 10192 37816 10198 37868
rect 10244 37865 10272 37896
rect 10318 37884 10324 37896
rect 10376 37884 10382 37936
rect 11238 37884 11244 37936
rect 11296 37924 11302 37936
rect 11762 37927 11820 37933
rect 11762 37924 11774 37927
rect 11296 37896 11774 37924
rect 11296 37884 11302 37896
rect 11762 37893 11774 37896
rect 11808 37893 11820 37927
rect 11762 37887 11820 37893
rect 10229 37859 10287 37865
rect 10229 37825 10241 37859
rect 10275 37825 10287 37859
rect 10229 37819 10287 37825
rect 10597 37859 10655 37865
rect 10597 37825 10609 37859
rect 10643 37825 10655 37859
rect 11514 37856 11520 37868
rect 11475 37828 11520 37856
rect 10597 37819 10655 37825
rect 9766 37748 9772 37800
rect 9824 37788 9830 37800
rect 10321 37791 10379 37797
rect 10321 37788 10333 37791
rect 9824 37760 10333 37788
rect 9824 37748 9830 37760
rect 10321 37757 10333 37760
rect 10367 37757 10379 37791
rect 10321 37751 10379 37757
rect 10413 37791 10471 37797
rect 10413 37757 10425 37791
rect 10459 37788 10471 37791
rect 10502 37788 10508 37800
rect 10459 37760 10508 37788
rect 10459 37757 10471 37760
rect 10413 37751 10471 37757
rect 10502 37748 10508 37760
rect 10560 37748 10566 37800
rect 5684 37692 6500 37720
rect 6840 37692 8064 37720
rect 9140 37692 9720 37720
rect 5684 37680 5690 37692
rect 1486 37652 1492 37664
rect 1447 37624 1492 37652
rect 1486 37612 1492 37624
rect 1544 37612 1550 37664
rect 5534 37652 5540 37664
rect 5495 37624 5540 37652
rect 5534 37612 5540 37624
rect 5592 37612 5598 37664
rect 6362 37652 6368 37664
rect 6323 37624 6368 37652
rect 6362 37612 6368 37624
rect 6420 37612 6426 37664
rect 6472 37652 6500 37692
rect 9140 37652 9168 37692
rect 9582 37652 9588 37664
rect 6472 37624 9168 37652
rect 9543 37624 9588 37652
rect 9582 37612 9588 37624
rect 9640 37612 9646 37664
rect 9692 37652 9720 37692
rect 10042 37680 10048 37732
rect 10100 37720 10106 37732
rect 10612 37720 10640 37819
rect 11514 37816 11520 37828
rect 11572 37816 11578 37868
rect 12406 37856 12434 37964
rect 13357 37961 13369 37995
rect 13403 37992 13415 37995
rect 14274 37992 14280 38004
rect 13403 37964 14280 37992
rect 13403 37961 13415 37964
rect 13357 37955 13415 37961
rect 14274 37952 14280 37964
rect 14332 37952 14338 38004
rect 14458 37952 14464 38004
rect 14516 37992 14522 38004
rect 14553 37995 14611 38001
rect 14553 37992 14565 37995
rect 14516 37964 14565 37992
rect 14516 37952 14522 37964
rect 14553 37961 14565 37964
rect 14599 37992 14611 37995
rect 16206 37992 16212 38004
rect 14599 37964 16212 37992
rect 14599 37961 14611 37964
rect 14553 37955 14611 37961
rect 16206 37952 16212 37964
rect 16264 37952 16270 38004
rect 17865 37927 17923 37933
rect 13832 37896 15056 37924
rect 13832 37868 13860 37896
rect 13633 37859 13691 37865
rect 12406 37828 13584 37856
rect 12986 37748 12992 37800
rect 13044 37788 13050 37800
rect 13354 37788 13360 37800
rect 13044 37760 13360 37788
rect 13044 37748 13050 37760
rect 13354 37748 13360 37760
rect 13412 37748 13418 37800
rect 13556 37788 13584 37828
rect 13633 37825 13645 37859
rect 13679 37856 13691 37859
rect 13814 37856 13820 37868
rect 13679 37828 13820 37856
rect 13679 37825 13691 37828
rect 13633 37819 13691 37825
rect 13814 37816 13820 37828
rect 13872 37816 13878 37868
rect 14093 37859 14151 37865
rect 14093 37825 14105 37859
rect 14139 37856 14151 37859
rect 14182 37856 14188 37868
rect 14139 37828 14188 37856
rect 14139 37825 14151 37828
rect 14093 37819 14151 37825
rect 14182 37816 14188 37828
rect 14240 37816 14246 37868
rect 14366 37856 14372 37868
rect 14327 37828 14372 37856
rect 14366 37816 14372 37828
rect 14424 37816 14430 37868
rect 15028 37865 15056 37896
rect 17865 37893 17877 37927
rect 17911 37924 17923 37927
rect 19426 37924 19432 37936
rect 17911 37896 19432 37924
rect 17911 37893 17923 37896
rect 17865 37887 17923 37893
rect 19426 37884 19432 37896
rect 19484 37884 19490 37936
rect 15013 37859 15071 37865
rect 15013 37825 15025 37859
rect 15059 37825 15071 37859
rect 17678 37856 17684 37868
rect 17639 37828 17684 37856
rect 15013 37819 15071 37825
rect 17678 37816 17684 37828
rect 17736 37816 17742 37868
rect 18049 37859 18107 37865
rect 18049 37825 18061 37859
rect 18095 37856 18107 37859
rect 18693 37859 18751 37865
rect 18693 37856 18705 37859
rect 18095 37828 18705 37856
rect 18095 37825 18107 37828
rect 18049 37819 18107 37825
rect 18693 37825 18705 37828
rect 18739 37825 18751 37859
rect 18693 37819 18751 37825
rect 13998 37788 14004 37800
rect 13556 37760 14004 37788
rect 13998 37748 14004 37760
rect 14056 37748 14062 37800
rect 14200 37788 14228 37816
rect 15102 37788 15108 37800
rect 14200 37760 15108 37788
rect 15102 37748 15108 37760
rect 15160 37748 15166 37800
rect 14185 37723 14243 37729
rect 10100 37692 10640 37720
rect 10704 37692 11008 37720
rect 10100 37680 10106 37692
rect 10704 37652 10732 37692
rect 9692 37624 10732 37652
rect 10781 37655 10839 37661
rect 10781 37621 10793 37655
rect 10827 37652 10839 37655
rect 10870 37652 10876 37664
rect 10827 37624 10876 37652
rect 10827 37621 10839 37624
rect 10781 37615 10839 37621
rect 10870 37612 10876 37624
rect 10928 37612 10934 37664
rect 10980 37652 11008 37692
rect 14185 37689 14197 37723
rect 14231 37720 14243 37723
rect 14918 37720 14924 37732
rect 14231 37692 14924 37720
rect 14231 37689 14243 37692
rect 14185 37683 14243 37689
rect 14918 37680 14924 37692
rect 14976 37680 14982 37732
rect 12434 37652 12440 37664
rect 10980 37624 12440 37652
rect 12434 37612 12440 37624
rect 12492 37612 12498 37664
rect 12894 37652 12900 37664
rect 12855 37624 12900 37652
rect 12894 37612 12900 37624
rect 12952 37612 12958 37664
rect 13541 37655 13599 37661
rect 13541 37621 13553 37655
rect 13587 37652 13599 37655
rect 13722 37652 13728 37664
rect 13587 37624 13728 37652
rect 13587 37621 13599 37624
rect 13541 37615 13599 37621
rect 13722 37612 13728 37624
rect 13780 37612 13786 37664
rect 18506 37652 18512 37664
rect 18467 37624 18512 37652
rect 18506 37612 18512 37624
rect 18564 37612 18570 37664
rect 1104 37562 30820 37584
rect 1104 37510 5915 37562
rect 5967 37510 5979 37562
rect 6031 37510 6043 37562
rect 6095 37510 6107 37562
rect 6159 37510 6171 37562
rect 6223 37510 15846 37562
rect 15898 37510 15910 37562
rect 15962 37510 15974 37562
rect 16026 37510 16038 37562
rect 16090 37510 16102 37562
rect 16154 37510 25776 37562
rect 25828 37510 25840 37562
rect 25892 37510 25904 37562
rect 25956 37510 25968 37562
rect 26020 37510 26032 37562
rect 26084 37510 30820 37562
rect 1104 37488 30820 37510
rect 2317 37451 2375 37457
rect 2317 37417 2329 37451
rect 2363 37448 2375 37451
rect 2406 37448 2412 37460
rect 2363 37420 2412 37448
rect 2363 37417 2375 37420
rect 2317 37411 2375 37417
rect 2406 37408 2412 37420
rect 2464 37408 2470 37460
rect 6454 37408 6460 37460
rect 6512 37448 6518 37460
rect 7469 37451 7527 37457
rect 7469 37448 7481 37451
rect 6512 37420 7481 37448
rect 6512 37408 6518 37420
rect 7469 37417 7481 37420
rect 7515 37417 7527 37451
rect 8938 37448 8944 37460
rect 8899 37420 8944 37448
rect 7469 37411 7527 37417
rect 8938 37408 8944 37420
rect 8996 37408 9002 37460
rect 12710 37448 12716 37460
rect 12671 37420 12716 37448
rect 12710 37408 12716 37420
rect 12768 37408 12774 37460
rect 13081 37451 13139 37457
rect 13081 37417 13093 37451
rect 13127 37448 13139 37451
rect 13814 37448 13820 37460
rect 13127 37420 13820 37448
rect 13127 37417 13139 37420
rect 13081 37411 13139 37417
rect 13814 37408 13820 37420
rect 13872 37408 13878 37460
rect 13998 37408 14004 37460
rect 14056 37448 14062 37460
rect 20346 37448 20352 37460
rect 14056 37420 20352 37448
rect 14056 37408 14062 37420
rect 20346 37408 20352 37420
rect 20404 37408 20410 37460
rect 2501 37383 2559 37389
rect 2501 37349 2513 37383
rect 2547 37349 2559 37383
rect 9582 37380 9588 37392
rect 2501 37343 2559 37349
rect 9140 37352 9588 37380
rect 2516 37312 2544 37343
rect 2516 37284 4099 37312
rect 1946 37244 1952 37256
rect 1907 37216 1952 37244
rect 1946 37204 1952 37216
rect 2004 37204 2010 37256
rect 2961 37247 3019 37253
rect 2961 37213 2973 37247
rect 3007 37213 3019 37247
rect 2961 37207 3019 37213
rect 2317 37179 2375 37185
rect 2317 37145 2329 37179
rect 2363 37176 2375 37179
rect 2976 37176 3004 37207
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 3786 37244 3792 37256
rect 3292 37216 3792 37244
rect 3292 37204 3298 37216
rect 3786 37204 3792 37216
rect 3844 37244 3850 37256
rect 3973 37247 4031 37253
rect 3973 37244 3985 37247
rect 3844 37216 3985 37244
rect 3844 37204 3850 37216
rect 3973 37213 3985 37216
rect 4019 37213 4031 37247
rect 3973 37207 4031 37213
rect 3326 37176 3332 37188
rect 2363 37148 2774 37176
rect 2976 37148 3332 37176
rect 2363 37145 2375 37148
rect 2317 37139 2375 37145
rect 2746 37108 2774 37148
rect 3326 37136 3332 37148
rect 3384 37136 3390 37188
rect 4071 37176 4099 37284
rect 4614 37272 4620 37324
rect 4672 37312 4678 37324
rect 4798 37312 4804 37324
rect 4672 37284 4804 37312
rect 4672 37272 4678 37284
rect 4798 37272 4804 37284
rect 4856 37312 4862 37324
rect 5353 37315 5411 37321
rect 5353 37312 5365 37315
rect 4856 37284 5365 37312
rect 4856 37272 4862 37284
rect 5353 37281 5365 37284
rect 5399 37281 5411 37315
rect 5626 37312 5632 37324
rect 5587 37284 5632 37312
rect 5353 37275 5411 37281
rect 5626 37272 5632 37284
rect 5684 37312 5690 37324
rect 5810 37312 5816 37324
rect 5684 37284 5816 37312
rect 5684 37272 5690 37284
rect 5810 37272 5816 37284
rect 5868 37272 5874 37324
rect 9140 37256 9168 37352
rect 9582 37340 9588 37352
rect 9640 37340 9646 37392
rect 15194 37340 15200 37392
rect 15252 37380 15258 37392
rect 15252 37352 15884 37380
rect 15252 37340 15258 37352
rect 9214 37272 9220 37324
rect 9272 37312 9278 37324
rect 9401 37315 9459 37321
rect 9401 37312 9413 37315
rect 9272 37284 9413 37312
rect 9272 37272 9278 37284
rect 9401 37281 9413 37284
rect 9447 37281 9459 37315
rect 9401 37275 9459 37281
rect 15378 37272 15384 37324
rect 15436 37312 15442 37324
rect 15654 37312 15660 37324
rect 15436 37284 15660 37312
rect 15436 37272 15442 37284
rect 15654 37272 15660 37284
rect 15712 37312 15718 37324
rect 15749 37315 15807 37321
rect 15749 37312 15761 37315
rect 15712 37284 15761 37312
rect 15712 37272 15718 37284
rect 15749 37281 15761 37284
rect 15795 37281 15807 37315
rect 15856 37312 15884 37352
rect 16025 37315 16083 37321
rect 16025 37312 16037 37315
rect 15856 37284 16037 37312
rect 15749 37275 15807 37281
rect 16025 37281 16037 37284
rect 16071 37281 16083 37315
rect 16025 37275 16083 37281
rect 16114 37272 16120 37324
rect 16172 37321 16178 37324
rect 16172 37315 16200 37321
rect 16188 37281 16200 37315
rect 16298 37312 16304 37324
rect 16259 37284 16304 37312
rect 16172 37275 16200 37281
rect 16172 37272 16178 37275
rect 16298 37272 16304 37284
rect 16356 37312 16362 37324
rect 17954 37312 17960 37324
rect 16356 37284 17960 37312
rect 16356 37272 16362 37284
rect 17954 37272 17960 37284
rect 18012 37272 18018 37324
rect 5718 37204 5724 37256
rect 5776 37244 5782 37256
rect 6362 37253 6368 37256
rect 6089 37247 6147 37253
rect 6089 37244 6101 37247
rect 5776 37216 6101 37244
rect 5776 37204 5782 37216
rect 6089 37213 6101 37216
rect 6135 37213 6147 37247
rect 6356 37244 6368 37253
rect 6323 37216 6368 37244
rect 6089 37207 6147 37213
rect 6356 37207 6368 37216
rect 6362 37204 6368 37207
rect 6420 37204 6426 37256
rect 8294 37204 8300 37256
rect 8352 37244 8358 37256
rect 8389 37247 8447 37253
rect 8389 37244 8401 37247
rect 8352 37216 8401 37244
rect 8352 37204 8358 37216
rect 8389 37213 8401 37216
rect 8435 37213 8447 37247
rect 9122 37244 9128 37256
rect 9083 37216 9128 37244
rect 8389 37207 8447 37213
rect 9122 37204 9128 37216
rect 9180 37204 9186 37256
rect 9306 37244 9312 37256
rect 9267 37216 9312 37244
rect 9306 37204 9312 37216
rect 9364 37204 9370 37256
rect 9493 37247 9551 37253
rect 9493 37213 9505 37247
rect 9539 37213 9551 37247
rect 9493 37207 9551 37213
rect 7742 37176 7748 37188
rect 4071 37148 7748 37176
rect 7742 37136 7748 37148
rect 7800 37136 7806 37188
rect 7926 37136 7932 37188
rect 7984 37176 7990 37188
rect 9508 37176 9536 37207
rect 9674 37204 9680 37256
rect 9732 37244 9738 37256
rect 10594 37244 10600 37256
rect 9732 37216 9825 37244
rect 10555 37216 10600 37244
rect 9732 37204 9738 37216
rect 10594 37204 10600 37216
rect 10652 37204 10658 37256
rect 10870 37253 10876 37256
rect 10864 37244 10876 37253
rect 10831 37216 10876 37244
rect 10864 37207 10876 37216
rect 10870 37204 10876 37207
rect 10928 37204 10934 37256
rect 12986 37244 12992 37256
rect 12947 37216 12992 37244
rect 12986 37204 12992 37216
rect 13044 37204 13050 37256
rect 13078 37204 13084 37256
rect 13136 37244 13142 37256
rect 14090 37244 14096 37256
rect 13136 37216 13181 37244
rect 14051 37216 14096 37244
rect 13136 37204 13142 37216
rect 14090 37204 14096 37216
rect 14148 37204 14154 37256
rect 14277 37247 14335 37253
rect 14277 37213 14289 37247
rect 14323 37213 14335 37247
rect 14277 37207 14335 37213
rect 14645 37247 14703 37253
rect 14645 37213 14657 37247
rect 14691 37244 14703 37247
rect 14918 37244 14924 37256
rect 14691 37216 14924 37244
rect 14691 37213 14703 37216
rect 14645 37207 14703 37213
rect 7984 37148 9536 37176
rect 9692 37176 9720 37204
rect 11330 37176 11336 37188
rect 9692 37148 11336 37176
rect 7984 37136 7990 37148
rect 8312 37120 8340 37148
rect 11330 37136 11336 37148
rect 11388 37136 11394 37188
rect 13722 37136 13728 37188
rect 13780 37176 13786 37188
rect 14292 37176 14320 37207
rect 14918 37204 14924 37216
rect 14976 37204 14982 37256
rect 15105 37247 15163 37253
rect 15105 37213 15117 37247
rect 15151 37213 15163 37247
rect 15286 37244 15292 37256
rect 15247 37216 15292 37244
rect 15105 37207 15163 37213
rect 13780 37148 14320 37176
rect 14553 37179 14611 37185
rect 13780 37136 13786 37148
rect 14553 37145 14565 37179
rect 14599 37176 14611 37179
rect 15120 37176 15148 37207
rect 15286 37204 15292 37216
rect 15344 37204 15350 37256
rect 17678 37204 17684 37256
rect 17736 37244 17742 37256
rect 18049 37247 18107 37253
rect 18049 37244 18061 37247
rect 17736 37216 18061 37244
rect 17736 37204 17742 37216
rect 18049 37213 18061 37216
rect 18095 37213 18107 37247
rect 18049 37207 18107 37213
rect 18141 37247 18199 37253
rect 18141 37213 18153 37247
rect 18187 37244 18199 37247
rect 18506 37244 18512 37256
rect 18187 37216 18512 37244
rect 18187 37213 18199 37216
rect 18141 37207 18199 37213
rect 18506 37204 18512 37216
rect 18564 37204 18570 37256
rect 18782 37204 18788 37256
rect 18840 37244 18846 37256
rect 19429 37247 19487 37253
rect 19429 37244 19441 37247
rect 18840 37216 19441 37244
rect 18840 37204 18846 37216
rect 19429 37213 19441 37216
rect 19475 37213 19487 37247
rect 30098 37244 30104 37256
rect 30059 37216 30104 37244
rect 19429 37207 19487 37213
rect 30098 37204 30104 37216
rect 30156 37204 30162 37256
rect 15194 37176 15200 37188
rect 14599 37148 15200 37176
rect 14599 37145 14611 37148
rect 14553 37139 14611 37145
rect 15194 37136 15200 37148
rect 15252 37136 15258 37188
rect 2958 37108 2964 37120
rect 2746 37080 2964 37108
rect 2958 37068 2964 37080
rect 3016 37068 3022 37120
rect 3142 37108 3148 37120
rect 3103 37080 3148 37108
rect 3142 37068 3148 37080
rect 3200 37068 3206 37120
rect 3418 37068 3424 37120
rect 3476 37108 3482 37120
rect 3789 37111 3847 37117
rect 3789 37108 3801 37111
rect 3476 37080 3801 37108
rect 3476 37068 3482 37080
rect 3789 37077 3801 37080
rect 3835 37077 3847 37111
rect 3789 37071 3847 37077
rect 4614 37068 4620 37120
rect 4672 37108 4678 37120
rect 4982 37108 4988 37120
rect 4672 37080 4988 37108
rect 4672 37068 4678 37080
rect 4982 37068 4988 37080
rect 5040 37108 5046 37120
rect 7282 37108 7288 37120
rect 5040 37080 7288 37108
rect 5040 37068 5046 37080
rect 7282 37068 7288 37080
rect 7340 37068 7346 37120
rect 8110 37068 8116 37120
rect 8168 37108 8174 37120
rect 8205 37111 8263 37117
rect 8205 37108 8217 37111
rect 8168 37080 8217 37108
rect 8168 37068 8174 37080
rect 8205 37077 8217 37080
rect 8251 37077 8263 37111
rect 8205 37071 8263 37077
rect 8294 37068 8300 37120
rect 8352 37068 8358 37120
rect 10042 37068 10048 37120
rect 10100 37108 10106 37120
rect 11977 37111 12035 37117
rect 11977 37108 11989 37111
rect 10100 37080 11989 37108
rect 10100 37068 10106 37080
rect 11977 37077 11989 37080
rect 12023 37077 12035 37111
rect 11977 37071 12035 37077
rect 14090 37068 14096 37120
rect 14148 37108 14154 37120
rect 14826 37108 14832 37120
rect 14148 37080 14832 37108
rect 14148 37068 14154 37080
rect 14826 37068 14832 37080
rect 14884 37068 14890 37120
rect 16942 37108 16948 37120
rect 16903 37080 16948 37108
rect 16942 37068 16948 37080
rect 17000 37068 17006 37120
rect 18138 37068 18144 37120
rect 18196 37108 18202 37120
rect 18509 37111 18567 37117
rect 18509 37108 18521 37111
rect 18196 37080 18521 37108
rect 18196 37068 18202 37080
rect 18509 37077 18521 37080
rect 18555 37077 18567 37111
rect 19242 37108 19248 37120
rect 19203 37080 19248 37108
rect 18509 37071 18567 37077
rect 19242 37068 19248 37080
rect 19300 37068 19306 37120
rect 29914 37108 29920 37120
rect 29875 37080 29920 37108
rect 29914 37068 29920 37080
rect 29972 37068 29978 37120
rect 1104 37018 30820 37040
rect 1104 36966 10880 37018
rect 10932 36966 10944 37018
rect 10996 36966 11008 37018
rect 11060 36966 11072 37018
rect 11124 36966 11136 37018
rect 11188 36966 20811 37018
rect 20863 36966 20875 37018
rect 20927 36966 20939 37018
rect 20991 36966 21003 37018
rect 21055 36966 21067 37018
rect 21119 36966 30820 37018
rect 1104 36944 30820 36966
rect 1581 36907 1639 36913
rect 1581 36873 1593 36907
rect 1627 36904 1639 36907
rect 1946 36904 1952 36916
rect 1627 36876 1952 36904
rect 1627 36873 1639 36876
rect 1581 36867 1639 36873
rect 1946 36864 1952 36876
rect 2004 36864 2010 36916
rect 2593 36907 2651 36913
rect 2593 36873 2605 36907
rect 2639 36904 2651 36907
rect 3050 36904 3056 36916
rect 2639 36876 3056 36904
rect 2639 36873 2651 36876
rect 2593 36867 2651 36873
rect 3050 36864 3056 36876
rect 3108 36864 3114 36916
rect 3605 36907 3663 36913
rect 3605 36873 3617 36907
rect 3651 36904 3663 36907
rect 3694 36904 3700 36916
rect 3651 36876 3700 36904
rect 3651 36873 3663 36876
rect 3605 36867 3663 36873
rect 3694 36864 3700 36876
rect 3752 36864 3758 36916
rect 3786 36864 3792 36916
rect 3844 36904 3850 36916
rect 5445 36907 5503 36913
rect 5445 36904 5457 36907
rect 3844 36876 5457 36904
rect 3844 36864 3850 36876
rect 5445 36873 5457 36876
rect 5491 36873 5503 36907
rect 5445 36867 5503 36873
rect 10873 36907 10931 36913
rect 10873 36873 10885 36907
rect 10919 36904 10931 36907
rect 11238 36904 11244 36916
rect 10919 36876 11244 36904
rect 10919 36873 10931 36876
rect 10873 36867 10931 36873
rect 11238 36864 11244 36876
rect 11296 36864 11302 36916
rect 11422 36864 11428 36916
rect 11480 36904 11486 36916
rect 11517 36907 11575 36913
rect 11517 36904 11529 36907
rect 11480 36876 11529 36904
rect 11480 36864 11486 36876
rect 11517 36873 11529 36876
rect 11563 36873 11575 36907
rect 14918 36904 14924 36916
rect 14879 36876 14924 36904
rect 11517 36867 11575 36873
rect 14918 36864 14924 36876
rect 14976 36864 14982 36916
rect 16942 36864 16948 36916
rect 17000 36904 17006 36916
rect 17221 36907 17279 36913
rect 17221 36904 17233 36907
rect 17000 36876 17233 36904
rect 17000 36864 17006 36876
rect 17221 36873 17233 36876
rect 17267 36873 17279 36907
rect 17221 36867 17279 36873
rect 17589 36907 17647 36913
rect 17589 36873 17601 36907
rect 17635 36904 17647 36907
rect 17678 36904 17684 36916
rect 17635 36876 17684 36904
rect 17635 36873 17647 36876
rect 17589 36867 17647 36873
rect 17678 36864 17684 36876
rect 17736 36864 17742 36916
rect 18782 36904 18788 36916
rect 18743 36876 18788 36904
rect 18782 36864 18788 36876
rect 18840 36864 18846 36916
rect 2409 36839 2467 36845
rect 2409 36805 2421 36839
rect 2455 36836 2467 36839
rect 4065 36839 4123 36845
rect 2455 36808 4016 36836
rect 2455 36805 2467 36808
rect 2409 36799 2467 36805
rect 1397 36771 1455 36777
rect 1397 36737 1409 36771
rect 1443 36768 1455 36771
rect 1762 36768 1768 36780
rect 1443 36740 1768 36768
rect 1443 36737 1455 36740
rect 1397 36731 1455 36737
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 2041 36771 2099 36777
rect 2041 36737 2053 36771
rect 2087 36768 2099 36771
rect 2130 36768 2136 36780
rect 2087 36740 2136 36768
rect 2087 36737 2099 36740
rect 2041 36731 2099 36737
rect 2130 36728 2136 36740
rect 2188 36728 2194 36780
rect 3418 36768 3424 36780
rect 3379 36740 3424 36768
rect 3418 36728 3424 36740
rect 3476 36728 3482 36780
rect 3988 36768 4016 36808
rect 4065 36805 4077 36839
rect 4111 36836 4123 36839
rect 4430 36836 4436 36848
rect 4111 36808 4436 36836
rect 4111 36805 4123 36808
rect 4065 36799 4123 36805
rect 4430 36796 4436 36808
rect 4488 36796 4494 36848
rect 5534 36836 5540 36848
rect 4540 36808 5540 36836
rect 4249 36771 4307 36777
rect 4249 36768 4261 36771
rect 3988 36740 4261 36768
rect 4249 36737 4261 36740
rect 4295 36768 4307 36771
rect 4540 36768 4568 36808
rect 5534 36796 5540 36808
rect 5592 36796 5598 36848
rect 12894 36836 12900 36848
rect 7392 36808 12900 36836
rect 4295 36740 4568 36768
rect 4295 36737 4307 36740
rect 4249 36731 4307 36737
rect 4614 36728 4620 36780
rect 4672 36768 4678 36780
rect 4672 36740 4717 36768
rect 4672 36728 4678 36740
rect 4798 36728 4804 36780
rect 4856 36768 4862 36780
rect 5626 36768 5632 36780
rect 4856 36740 4901 36768
rect 5587 36740 5632 36768
rect 4856 36728 4862 36740
rect 5626 36728 5632 36740
rect 5684 36728 5690 36780
rect 7392 36777 7420 36808
rect 7377 36771 7435 36777
rect 7377 36737 7389 36771
rect 7423 36737 7435 36771
rect 7377 36731 7435 36737
rect 7466 36728 7472 36780
rect 7524 36768 7530 36780
rect 8021 36771 8079 36777
rect 8021 36768 8033 36771
rect 7524 36740 8033 36768
rect 7524 36728 7530 36740
rect 8021 36737 8033 36740
rect 8067 36737 8079 36771
rect 8021 36731 8079 36737
rect 8110 36728 8116 36780
rect 8168 36768 8174 36780
rect 9033 36771 9091 36777
rect 9033 36768 9045 36771
rect 8168 36740 9045 36768
rect 8168 36728 8174 36740
rect 9033 36737 9045 36740
rect 9079 36737 9091 36771
rect 10134 36768 10140 36780
rect 10095 36740 10140 36768
rect 9033 36731 9091 36737
rect 10134 36728 10140 36740
rect 10192 36728 10198 36780
rect 10318 36768 10324 36780
rect 10279 36740 10324 36768
rect 10318 36728 10324 36740
rect 10376 36728 10382 36780
rect 10502 36768 10508 36780
rect 10463 36740 10508 36768
rect 10502 36728 10508 36740
rect 10560 36728 10566 36780
rect 10704 36777 10732 36808
rect 12894 36796 12900 36808
rect 12952 36796 12958 36848
rect 19334 36836 19340 36848
rect 13740 36808 14872 36836
rect 13740 36780 13768 36808
rect 10689 36771 10747 36777
rect 10689 36737 10701 36771
rect 10735 36737 10747 36771
rect 10689 36731 10747 36737
rect 10778 36728 10784 36780
rect 10836 36768 10842 36780
rect 11701 36771 11759 36777
rect 11701 36768 11713 36771
rect 10836 36740 11713 36768
rect 10836 36728 10842 36740
rect 11701 36737 11713 36740
rect 11747 36737 11759 36771
rect 11701 36731 11759 36737
rect 12434 36728 12440 36780
rect 12492 36768 12498 36780
rect 12492 36740 12537 36768
rect 12492 36728 12498 36740
rect 13078 36728 13084 36780
rect 13136 36768 13142 36780
rect 13173 36771 13231 36777
rect 13173 36768 13185 36771
rect 13136 36740 13185 36768
rect 13136 36728 13142 36740
rect 13173 36737 13185 36740
rect 13219 36768 13231 36771
rect 13722 36768 13728 36780
rect 13219 36740 13728 36768
rect 13219 36737 13231 36740
rect 13173 36731 13231 36737
rect 13722 36728 13728 36740
rect 13780 36728 13786 36780
rect 13814 36728 13820 36780
rect 13872 36768 13878 36780
rect 14093 36771 14151 36777
rect 13872 36740 13917 36768
rect 13872 36728 13878 36740
rect 14093 36737 14105 36771
rect 14139 36737 14151 36771
rect 14093 36731 14151 36737
rect 4433 36703 4491 36709
rect 4433 36669 4445 36703
rect 4479 36669 4491 36703
rect 4433 36663 4491 36669
rect 4448 36632 4476 36663
rect 4522 36660 4528 36712
rect 4580 36700 4586 36712
rect 9490 36700 9496 36712
rect 4580 36672 4625 36700
rect 6840 36672 9496 36700
rect 4580 36660 4586 36672
rect 4706 36632 4712 36644
rect 4448 36604 4712 36632
rect 4706 36592 4712 36604
rect 4764 36592 4770 36644
rect 2406 36564 2412 36576
rect 2367 36536 2412 36564
rect 2406 36524 2412 36536
rect 2464 36524 2470 36576
rect 2958 36524 2964 36576
rect 3016 36564 3022 36576
rect 6840 36564 6868 36672
rect 9490 36660 9496 36672
rect 9548 36660 9554 36712
rect 9766 36660 9772 36712
rect 9824 36700 9830 36712
rect 10413 36703 10471 36709
rect 10413 36700 10425 36703
rect 9824 36672 10425 36700
rect 9824 36660 9830 36672
rect 10413 36669 10425 36672
rect 10459 36669 10471 36703
rect 10413 36663 10471 36669
rect 11882 36660 11888 36712
rect 11940 36700 11946 36712
rect 13265 36703 13323 36709
rect 13265 36700 13277 36703
rect 11940 36672 13277 36700
rect 11940 36660 11946 36672
rect 13265 36669 13277 36672
rect 13311 36700 13323 36703
rect 14108 36700 14136 36731
rect 14182 36728 14188 36780
rect 14240 36768 14246 36780
rect 14844 36777 14872 36808
rect 18616 36808 19340 36836
rect 14829 36771 14887 36777
rect 14240 36740 14285 36768
rect 14240 36728 14246 36740
rect 14829 36737 14841 36771
rect 14875 36737 14887 36771
rect 14829 36731 14887 36737
rect 14918 36728 14924 36780
rect 14976 36768 14982 36780
rect 18616 36777 18644 36808
rect 19334 36796 19340 36808
rect 19392 36836 19398 36848
rect 20162 36836 20168 36848
rect 19392 36808 20168 36836
rect 19392 36796 19398 36808
rect 20162 36796 20168 36808
rect 20220 36796 20226 36848
rect 15013 36771 15071 36777
rect 15013 36768 15025 36771
rect 14976 36740 15025 36768
rect 14976 36728 14982 36740
rect 15013 36737 15025 36740
rect 15059 36737 15071 36771
rect 15013 36731 15071 36737
rect 18601 36771 18659 36777
rect 18601 36737 18613 36771
rect 18647 36737 18659 36771
rect 19242 36768 19248 36780
rect 19203 36740 19248 36768
rect 18601 36731 18659 36737
rect 13311 36672 14136 36700
rect 14369 36703 14427 36709
rect 13311 36669 13323 36672
rect 13265 36663 13323 36669
rect 14369 36669 14381 36703
rect 14415 36700 14427 36703
rect 15286 36700 15292 36712
rect 14415 36672 15292 36700
rect 14415 36669 14427 36672
rect 14369 36663 14427 36669
rect 15286 36660 15292 36672
rect 15344 36660 15350 36712
rect 16574 36660 16580 36712
rect 16632 36700 16638 36712
rect 16850 36700 16856 36712
rect 16632 36672 16856 36700
rect 16632 36660 16638 36672
rect 16850 36660 16856 36672
rect 16908 36700 16914 36712
rect 16945 36703 17003 36709
rect 16945 36700 16957 36703
rect 16908 36672 16957 36700
rect 16908 36660 16914 36672
rect 16945 36669 16957 36672
rect 16991 36669 17003 36703
rect 17126 36700 17132 36712
rect 17087 36672 17132 36700
rect 16945 36663 17003 36669
rect 17126 36660 17132 36672
rect 17184 36660 17190 36712
rect 6917 36635 6975 36641
rect 6917 36601 6929 36635
rect 6963 36632 6975 36635
rect 7558 36632 7564 36644
rect 6963 36604 7564 36632
rect 6963 36601 6975 36604
rect 6917 36595 6975 36601
rect 7558 36592 7564 36604
rect 7616 36592 7622 36644
rect 8018 36592 8024 36644
rect 8076 36632 8082 36644
rect 18616 36632 18644 36731
rect 19242 36728 19248 36740
rect 19300 36728 19306 36780
rect 19518 36777 19524 36780
rect 19512 36731 19524 36777
rect 19576 36768 19582 36780
rect 22094 36768 22100 36780
rect 19576 36740 19612 36768
rect 22055 36740 22100 36768
rect 19518 36728 19524 36731
rect 19576 36728 19582 36740
rect 22094 36728 22100 36740
rect 22152 36728 22158 36780
rect 22281 36703 22339 36709
rect 22281 36669 22293 36703
rect 22327 36700 22339 36703
rect 29914 36700 29920 36712
rect 22327 36672 29920 36700
rect 22327 36669 22339 36672
rect 22281 36663 22339 36669
rect 29914 36660 29920 36672
rect 29972 36660 29978 36712
rect 8076 36604 18644 36632
rect 8076 36592 8082 36604
rect 7190 36564 7196 36576
rect 3016 36536 6868 36564
rect 7151 36536 7196 36564
rect 3016 36524 3022 36536
rect 7190 36524 7196 36536
rect 7248 36524 7254 36576
rect 7742 36524 7748 36576
rect 7800 36564 7806 36576
rect 7837 36567 7895 36573
rect 7837 36564 7849 36567
rect 7800 36536 7849 36564
rect 7800 36524 7806 36536
rect 7837 36533 7849 36536
rect 7883 36533 7895 36567
rect 7837 36527 7895 36533
rect 9217 36567 9275 36573
rect 9217 36533 9229 36567
rect 9263 36564 9275 36567
rect 10410 36564 10416 36576
rect 9263 36536 10416 36564
rect 9263 36533 9275 36536
rect 9217 36527 9275 36533
rect 10410 36524 10416 36536
rect 10468 36564 10474 36576
rect 10778 36564 10784 36576
rect 10468 36536 10784 36564
rect 10468 36524 10474 36536
rect 10778 36524 10784 36536
rect 10836 36524 10842 36576
rect 11330 36524 11336 36576
rect 11388 36564 11394 36576
rect 12621 36567 12679 36573
rect 12621 36564 12633 36567
rect 11388 36536 12633 36564
rect 11388 36524 11394 36536
rect 12621 36533 12633 36536
rect 12667 36564 12679 36567
rect 13538 36564 13544 36576
rect 12667 36536 13544 36564
rect 12667 36533 12679 36536
rect 12621 36527 12679 36533
rect 13538 36524 13544 36536
rect 13596 36524 13602 36576
rect 13722 36524 13728 36576
rect 13780 36564 13786 36576
rect 13909 36567 13967 36573
rect 13909 36564 13921 36567
rect 13780 36536 13921 36564
rect 13780 36524 13786 36536
rect 13909 36533 13921 36536
rect 13955 36533 13967 36567
rect 20622 36564 20628 36576
rect 20583 36536 20628 36564
rect 13909 36527 13967 36533
rect 20622 36524 20628 36536
rect 20680 36524 20686 36576
rect 21266 36524 21272 36576
rect 21324 36564 21330 36576
rect 21913 36567 21971 36573
rect 21913 36564 21925 36567
rect 21324 36536 21925 36564
rect 21324 36524 21330 36536
rect 21913 36533 21925 36536
rect 21959 36533 21971 36567
rect 21913 36527 21971 36533
rect 1104 36474 30820 36496
rect 1104 36422 5915 36474
rect 5967 36422 5979 36474
rect 6031 36422 6043 36474
rect 6095 36422 6107 36474
rect 6159 36422 6171 36474
rect 6223 36422 15846 36474
rect 15898 36422 15910 36474
rect 15962 36422 15974 36474
rect 16026 36422 16038 36474
rect 16090 36422 16102 36474
rect 16154 36422 25776 36474
rect 25828 36422 25840 36474
rect 25892 36422 25904 36474
rect 25956 36422 25968 36474
rect 26020 36422 26032 36474
rect 26084 36422 30820 36474
rect 1104 36400 30820 36422
rect 3970 36360 3976 36372
rect 3931 36332 3976 36360
rect 3970 36320 3976 36332
rect 4028 36320 4034 36372
rect 5261 36363 5319 36369
rect 5261 36329 5273 36363
rect 5307 36360 5319 36363
rect 5718 36360 5724 36372
rect 5307 36332 5724 36360
rect 5307 36329 5319 36332
rect 5261 36323 5319 36329
rect 5718 36320 5724 36332
rect 5776 36320 5782 36372
rect 7190 36360 7196 36372
rect 7103 36332 7196 36360
rect 7190 36320 7196 36332
rect 7248 36320 7254 36372
rect 9306 36320 9312 36372
rect 9364 36360 9370 36372
rect 16945 36363 17003 36369
rect 9364 36332 12434 36360
rect 9364 36320 9370 36332
rect 1762 36252 1768 36304
rect 1820 36292 1826 36304
rect 2314 36292 2320 36304
rect 1820 36264 2320 36292
rect 1820 36252 1826 36264
rect 2314 36252 2320 36264
rect 2372 36292 2378 36304
rect 7208 36292 7236 36320
rect 9674 36292 9680 36304
rect 2372 36264 7236 36292
rect 7300 36264 9680 36292
rect 2372 36252 2378 36264
rect 2866 36224 2872 36236
rect 1688 36196 2872 36224
rect 1688 36165 1716 36196
rect 2866 36184 2872 36196
rect 2924 36184 2930 36236
rect 6012 36233 6040 36264
rect 5997 36227 6055 36233
rect 5997 36193 6009 36227
rect 6043 36193 6055 36227
rect 5997 36187 6055 36193
rect 1673 36159 1731 36165
rect 1673 36125 1685 36159
rect 1719 36125 1731 36159
rect 1673 36119 1731 36125
rect 2409 36159 2467 36165
rect 2409 36125 2421 36159
rect 2455 36156 2467 36159
rect 2455 36128 2774 36156
rect 2455 36125 2467 36128
rect 2409 36119 2467 36125
rect 2746 36088 2774 36128
rect 2958 36116 2964 36168
rect 3016 36156 3022 36168
rect 3053 36159 3111 36165
rect 3053 36156 3065 36159
rect 3016 36128 3065 36156
rect 3016 36116 3022 36128
rect 3053 36125 3065 36128
rect 3099 36125 3111 36159
rect 3786 36156 3792 36168
rect 3747 36128 3792 36156
rect 3053 36119 3111 36125
rect 3786 36116 3792 36128
rect 3844 36116 3850 36168
rect 3970 36116 3976 36168
rect 4028 36156 4034 36168
rect 4617 36159 4675 36165
rect 4617 36156 4629 36159
rect 4028 36128 4629 36156
rect 4028 36116 4034 36128
rect 4617 36125 4629 36128
rect 4663 36125 4675 36159
rect 4617 36119 4675 36125
rect 5077 36159 5135 36165
rect 5077 36125 5089 36159
rect 5123 36156 5135 36159
rect 5534 36156 5540 36168
rect 5123 36128 5540 36156
rect 5123 36125 5135 36128
rect 5077 36119 5135 36125
rect 5534 36116 5540 36128
rect 5592 36116 5598 36168
rect 5721 36159 5779 36165
rect 5721 36125 5733 36159
rect 5767 36156 5779 36159
rect 6546 36156 6552 36168
rect 5767 36128 6552 36156
rect 5767 36125 5779 36128
rect 5721 36119 5779 36125
rect 6546 36116 6552 36128
rect 6604 36156 6610 36168
rect 7300 36156 7328 36264
rect 9674 36252 9680 36264
rect 9732 36252 9738 36304
rect 9769 36295 9827 36301
rect 9769 36261 9781 36295
rect 9815 36292 9827 36295
rect 12406 36292 12434 36332
rect 15120 36332 16712 36360
rect 15120 36292 15148 36332
rect 9815 36264 10272 36292
rect 12406 36264 15148 36292
rect 9815 36261 9827 36264
rect 9769 36255 9827 36261
rect 10042 36224 10048 36236
rect 7484 36196 10048 36224
rect 7484 36165 7512 36196
rect 10042 36184 10048 36196
rect 10100 36184 10106 36236
rect 10244 36233 10272 36264
rect 15194 36252 15200 36304
rect 15252 36292 15258 36304
rect 16684 36292 16712 36332
rect 16945 36329 16957 36363
rect 16991 36360 17003 36363
rect 17126 36360 17132 36372
rect 16991 36332 17132 36360
rect 16991 36329 17003 36332
rect 16945 36323 17003 36329
rect 17126 36320 17132 36332
rect 17184 36320 17190 36372
rect 21542 36292 21548 36304
rect 15252 36264 15884 36292
rect 16684 36264 21548 36292
rect 15252 36252 15258 36264
rect 10229 36227 10287 36233
rect 10229 36193 10241 36227
rect 10275 36193 10287 36227
rect 10229 36187 10287 36193
rect 12894 36184 12900 36236
rect 12952 36224 12958 36236
rect 15286 36224 15292 36236
rect 12952 36196 13216 36224
rect 15247 36196 15292 36224
rect 12952 36184 12958 36196
rect 6604 36128 7328 36156
rect 7469 36159 7527 36165
rect 6604 36116 6610 36128
rect 7469 36125 7481 36159
rect 7515 36125 7527 36159
rect 8110 36156 8116 36168
rect 8071 36128 8116 36156
rect 7469 36119 7527 36125
rect 8110 36116 8116 36128
rect 8168 36116 8174 36168
rect 8478 36116 8484 36168
rect 8536 36156 8542 36168
rect 9125 36159 9183 36165
rect 9125 36156 9137 36159
rect 8536 36128 9137 36156
rect 8536 36116 8542 36128
rect 9125 36125 9137 36128
rect 9171 36125 9183 36159
rect 9125 36119 9183 36125
rect 9585 36159 9643 36165
rect 9585 36125 9597 36159
rect 9631 36156 9643 36159
rect 10318 36156 10324 36168
rect 9631 36128 10324 36156
rect 9631 36125 9643 36128
rect 9585 36119 9643 36125
rect 10318 36116 10324 36128
rect 10376 36116 10382 36168
rect 12800 36159 12858 36165
rect 12800 36125 12812 36159
rect 12846 36156 12858 36159
rect 13078 36156 13084 36168
rect 12846 36128 13084 36156
rect 12846 36125 12858 36128
rect 12800 36119 12858 36125
rect 13078 36116 13084 36128
rect 13136 36116 13142 36168
rect 13188 36165 13216 36196
rect 15286 36184 15292 36196
rect 15344 36184 15350 36236
rect 15746 36224 15752 36236
rect 15707 36196 15752 36224
rect 15746 36184 15752 36196
rect 15804 36184 15810 36236
rect 15856 36224 15884 36264
rect 21542 36252 21548 36264
rect 21600 36252 21606 36304
rect 16025 36227 16083 36233
rect 16025 36224 16037 36227
rect 15856 36196 16037 36224
rect 16025 36193 16037 36196
rect 16071 36193 16083 36227
rect 16025 36187 16083 36193
rect 16114 36184 16120 36236
rect 16172 36233 16178 36236
rect 16172 36227 16200 36233
rect 16188 36193 16200 36227
rect 19334 36224 19340 36236
rect 16172 36187 16200 36193
rect 17604 36196 19340 36224
rect 16172 36184 16178 36187
rect 13172 36159 13230 36165
rect 13172 36125 13184 36159
rect 13218 36125 13230 36159
rect 13172 36119 13230 36125
rect 13262 36116 13268 36168
rect 13320 36156 13326 36168
rect 15105 36159 15163 36165
rect 13320 36128 13365 36156
rect 13320 36116 13326 36128
rect 15105 36125 15117 36159
rect 15151 36156 15163 36159
rect 15194 36156 15200 36168
rect 15151 36128 15200 36156
rect 15151 36125 15163 36128
rect 15105 36119 15163 36125
rect 15194 36116 15200 36128
rect 15252 36116 15258 36168
rect 16298 36156 16304 36168
rect 16259 36128 16304 36156
rect 16298 36116 16304 36128
rect 16356 36116 16362 36168
rect 17604 36165 17632 36196
rect 19334 36184 19340 36196
rect 19392 36184 19398 36236
rect 19794 36184 19800 36236
rect 19852 36224 19858 36236
rect 20254 36224 20260 36236
rect 19852 36196 20260 36224
rect 19852 36184 19858 36196
rect 20254 36184 20260 36196
rect 20312 36184 20318 36236
rect 17589 36159 17647 36165
rect 17589 36125 17601 36159
rect 17635 36125 17647 36159
rect 18417 36159 18475 36165
rect 18417 36156 18429 36159
rect 17589 36119 17647 36125
rect 17788 36128 18429 36156
rect 10496 36091 10554 36097
rect 2746 36060 8984 36088
rect 1486 36020 1492 36032
rect 1447 35992 1492 36020
rect 1486 35980 1492 35992
rect 1544 35980 1550 36032
rect 2222 36020 2228 36032
rect 2183 35992 2228 36020
rect 2222 35980 2228 35992
rect 2280 35980 2286 36032
rect 2866 36020 2872 36032
rect 2827 35992 2872 36020
rect 2866 35980 2872 35992
rect 2924 35980 2930 36032
rect 3142 35980 3148 36032
rect 3200 36020 3206 36032
rect 4433 36023 4491 36029
rect 4433 36020 4445 36023
rect 3200 35992 4445 36020
rect 3200 35980 3206 35992
rect 4433 35989 4445 35992
rect 4479 35989 4491 36023
rect 4433 35983 4491 35989
rect 7009 36023 7067 36029
rect 7009 35989 7021 36023
rect 7055 36020 7067 36023
rect 7190 36020 7196 36032
rect 7055 35992 7196 36020
rect 7055 35989 7067 35992
rect 7009 35983 7067 35989
rect 7190 35980 7196 35992
rect 7248 35980 7254 36032
rect 7926 36020 7932 36032
rect 7887 35992 7932 36020
rect 7926 35980 7932 35992
rect 7984 35980 7990 36032
rect 8956 36029 8984 36060
rect 10496 36057 10508 36091
rect 10542 36088 10554 36091
rect 10686 36088 10692 36100
rect 10542 36060 10692 36088
rect 10542 36057 10554 36060
rect 10496 36051 10554 36057
rect 10686 36048 10692 36060
rect 10744 36048 10750 36100
rect 12897 36091 12955 36097
rect 12897 36057 12909 36091
rect 12943 36057 12955 36091
rect 12897 36051 12955 36057
rect 12989 36091 13047 36097
rect 12989 36057 13001 36091
rect 13035 36088 13047 36091
rect 13354 36088 13360 36100
rect 13035 36060 13360 36088
rect 13035 36057 13047 36060
rect 12989 36051 13047 36057
rect 8941 36023 8999 36029
rect 8941 35989 8953 36023
rect 8987 35989 8999 36023
rect 8941 35983 8999 35989
rect 10594 35980 10600 36032
rect 10652 36020 10658 36032
rect 11609 36023 11667 36029
rect 11609 36020 11621 36023
rect 10652 35992 11621 36020
rect 10652 35980 10658 35992
rect 11609 35989 11621 35992
rect 11655 35989 11667 36023
rect 12618 36020 12624 36032
rect 12579 35992 12624 36020
rect 11609 35983 11667 35989
rect 12618 35980 12624 35992
rect 12676 35980 12682 36032
rect 12912 36020 12940 36051
rect 13354 36048 13360 36060
rect 13412 36048 13418 36100
rect 13170 36020 13176 36032
rect 12912 35992 13176 36020
rect 13170 35980 13176 35992
rect 13228 35980 13234 36032
rect 13372 36020 13400 36048
rect 16574 36020 16580 36032
rect 13372 35992 16580 36020
rect 16574 35980 16580 35992
rect 16632 35980 16638 36032
rect 17788 36029 17816 36128
rect 18417 36125 18429 36128
rect 18463 36125 18475 36159
rect 18417 36119 18475 36125
rect 20622 36116 20628 36168
rect 20680 36156 20686 36168
rect 20809 36159 20867 36165
rect 20809 36156 20821 36159
rect 20680 36128 20821 36156
rect 20680 36116 20686 36128
rect 20809 36125 20821 36128
rect 20855 36125 20867 36159
rect 20809 36119 20867 36125
rect 21085 36159 21143 36165
rect 21085 36125 21097 36159
rect 21131 36156 21143 36159
rect 21174 36156 21180 36168
rect 21131 36128 21180 36156
rect 21131 36125 21143 36128
rect 21085 36119 21143 36125
rect 21174 36116 21180 36128
rect 21232 36116 21238 36168
rect 18506 36048 18512 36100
rect 18564 36088 18570 36100
rect 19426 36088 19432 36100
rect 18564 36060 19432 36088
rect 18564 36048 18570 36060
rect 19426 36048 19432 36060
rect 19484 36088 19490 36100
rect 19981 36091 20039 36097
rect 19981 36088 19993 36091
rect 19484 36060 19993 36088
rect 19484 36048 19490 36060
rect 19981 36057 19993 36060
rect 20027 36057 20039 36091
rect 19981 36051 20039 36057
rect 20073 36091 20131 36097
rect 20073 36057 20085 36091
rect 20119 36088 20131 36091
rect 21269 36091 21327 36097
rect 21269 36088 21281 36091
rect 20119 36060 21281 36088
rect 20119 36057 20131 36060
rect 20073 36051 20131 36057
rect 21269 36057 21281 36060
rect 21315 36057 21327 36091
rect 21269 36051 21327 36057
rect 17773 36023 17831 36029
rect 17773 35989 17785 36023
rect 17819 35989 17831 36023
rect 18230 36020 18236 36032
rect 18191 35992 18236 36020
rect 17773 35983 17831 35989
rect 18230 35980 18236 35992
rect 18288 35980 18294 36032
rect 19610 36020 19616 36032
rect 19571 35992 19616 36020
rect 19610 35980 19616 35992
rect 19668 35980 19674 36032
rect 20254 35980 20260 36032
rect 20312 36020 20318 36032
rect 20901 36023 20959 36029
rect 20901 36020 20913 36023
rect 20312 35992 20913 36020
rect 20312 35980 20318 35992
rect 20901 35989 20913 35992
rect 20947 35989 20959 36023
rect 20901 35983 20959 35989
rect 1104 35930 30820 35952
rect 1104 35878 10880 35930
rect 10932 35878 10944 35930
rect 10996 35878 11008 35930
rect 11060 35878 11072 35930
rect 11124 35878 11136 35930
rect 11188 35878 20811 35930
rect 20863 35878 20875 35930
rect 20927 35878 20939 35930
rect 20991 35878 21003 35930
rect 21055 35878 21067 35930
rect 21119 35878 30820 35930
rect 1104 35856 30820 35878
rect 2225 35819 2283 35825
rect 2225 35785 2237 35819
rect 2271 35816 2283 35819
rect 5534 35816 5540 35828
rect 2271 35788 5396 35816
rect 5495 35788 5540 35816
rect 2271 35785 2283 35788
rect 2225 35779 2283 35785
rect 3234 35748 3240 35760
rect 2884 35720 3240 35748
rect 1857 35683 1915 35689
rect 1857 35649 1869 35683
rect 1903 35680 1915 35683
rect 1946 35680 1952 35692
rect 1903 35652 1952 35680
rect 1903 35649 1915 35652
rect 1857 35643 1915 35649
rect 1946 35640 1952 35652
rect 2004 35640 2010 35692
rect 2884 35689 2912 35720
rect 3234 35708 3240 35720
rect 3292 35748 3298 35760
rect 5368 35748 5396 35788
rect 5534 35776 5540 35788
rect 5592 35776 5598 35828
rect 6825 35819 6883 35825
rect 6825 35785 6837 35819
rect 6871 35816 6883 35819
rect 7466 35816 7472 35828
rect 6871 35788 7472 35816
rect 6871 35785 6883 35788
rect 6825 35779 6883 35785
rect 7466 35776 7472 35788
rect 7524 35776 7530 35828
rect 7745 35819 7803 35825
rect 7745 35785 7757 35819
rect 7791 35816 7803 35819
rect 8202 35816 8208 35828
rect 7791 35788 8208 35816
rect 7791 35785 7803 35788
rect 7745 35779 7803 35785
rect 8202 35776 8208 35788
rect 8260 35816 8266 35828
rect 9217 35819 9275 35825
rect 9217 35816 9229 35819
rect 8260 35788 9229 35816
rect 8260 35776 8266 35788
rect 9217 35785 9229 35788
rect 9263 35785 9275 35819
rect 9217 35779 9275 35785
rect 9398 35776 9404 35828
rect 9456 35816 9462 35828
rect 10686 35816 10692 35828
rect 9456 35788 10548 35816
rect 10647 35788 10692 35816
rect 9456 35776 9462 35788
rect 9122 35748 9128 35760
rect 3292 35720 4936 35748
rect 5368 35720 9128 35748
rect 3292 35708 3298 35720
rect 4908 35689 4936 35720
rect 9122 35708 9128 35720
rect 9180 35708 9186 35760
rect 10410 35748 10416 35760
rect 10152 35720 10416 35748
rect 2869 35683 2927 35689
rect 2869 35649 2881 35683
rect 2915 35649 2927 35683
rect 3513 35683 3571 35689
rect 3513 35680 3525 35683
rect 2869 35643 2927 35649
rect 3068 35652 3525 35680
rect 3068 35553 3096 35652
rect 3513 35649 3525 35652
rect 3559 35649 3571 35683
rect 3513 35643 3571 35649
rect 4893 35683 4951 35689
rect 4893 35649 4905 35683
rect 4939 35680 4951 35683
rect 5534 35680 5540 35692
rect 4939 35652 5540 35680
rect 4939 35649 4951 35652
rect 4893 35643 4951 35649
rect 5534 35640 5540 35652
rect 5592 35680 5598 35692
rect 5721 35683 5779 35689
rect 5721 35680 5733 35683
rect 5592 35652 5733 35680
rect 5592 35640 5598 35652
rect 5721 35649 5733 35652
rect 5767 35649 5779 35683
rect 5721 35643 5779 35649
rect 6365 35683 6423 35689
rect 6365 35649 6377 35683
rect 6411 35680 6423 35683
rect 7745 35683 7803 35689
rect 7745 35680 7757 35683
rect 6411 35652 7757 35680
rect 6411 35649 6423 35652
rect 6365 35643 6423 35649
rect 7745 35649 7757 35652
rect 7791 35649 7803 35683
rect 7745 35643 7803 35649
rect 7837 35683 7895 35689
rect 7837 35649 7849 35683
rect 7883 35680 7895 35683
rect 7926 35680 7932 35692
rect 7883 35652 7932 35680
rect 7883 35649 7895 35652
rect 7837 35643 7895 35649
rect 7926 35640 7932 35652
rect 7984 35640 7990 35692
rect 8104 35683 8162 35689
rect 8104 35649 8116 35683
rect 8150 35680 8162 35683
rect 8386 35680 8392 35692
rect 8150 35652 8392 35680
rect 8150 35649 8162 35652
rect 8104 35643 8162 35649
rect 8386 35640 8392 35652
rect 8444 35640 8450 35692
rect 9953 35683 10011 35689
rect 9953 35649 9965 35683
rect 9999 35680 10011 35683
rect 10042 35680 10048 35692
rect 9999 35652 10048 35680
rect 9999 35649 10011 35652
rect 9953 35643 10011 35649
rect 10042 35640 10048 35652
rect 10100 35640 10106 35692
rect 10152 35689 10180 35720
rect 10410 35708 10416 35720
rect 10468 35708 10474 35760
rect 10520 35748 10548 35788
rect 10686 35776 10692 35788
rect 10744 35776 10750 35828
rect 13262 35816 13268 35828
rect 12636 35788 13268 35816
rect 10594 35748 10600 35760
rect 10520 35720 10600 35748
rect 10137 35683 10195 35689
rect 10137 35649 10149 35683
rect 10183 35649 10195 35683
rect 10137 35643 10195 35649
rect 10226 35640 10232 35692
rect 10284 35680 10290 35692
rect 10520 35689 10548 35720
rect 10594 35708 10600 35720
rect 10652 35708 10658 35760
rect 10505 35683 10563 35689
rect 10284 35652 10329 35680
rect 10284 35640 10290 35652
rect 10505 35649 10517 35683
rect 10551 35649 10563 35683
rect 10505 35643 10563 35649
rect 11793 35683 11851 35689
rect 11793 35649 11805 35683
rect 11839 35680 11851 35683
rect 11974 35680 11980 35692
rect 11839 35652 11980 35680
rect 11839 35649 11851 35652
rect 11793 35643 11851 35649
rect 11974 35640 11980 35652
rect 12032 35640 12038 35692
rect 12636 35689 12664 35788
rect 13262 35776 13268 35788
rect 13320 35776 13326 35828
rect 19426 35776 19432 35828
rect 19484 35816 19490 35828
rect 19521 35819 19579 35825
rect 19521 35816 19533 35819
rect 19484 35788 19533 35816
rect 19484 35776 19490 35788
rect 19521 35785 19533 35788
rect 19567 35816 19579 35819
rect 20254 35816 20260 35828
rect 19567 35788 20260 35816
rect 19567 35785 19579 35788
rect 19521 35779 19579 35785
rect 20254 35776 20260 35788
rect 20312 35776 20318 35828
rect 20349 35819 20407 35825
rect 20349 35785 20361 35819
rect 20395 35816 20407 35819
rect 20714 35816 20720 35828
rect 20395 35788 20720 35816
rect 20395 35785 20407 35788
rect 20349 35779 20407 35785
rect 20714 35776 20720 35788
rect 20772 35816 20778 35828
rect 21174 35816 21180 35828
rect 20772 35788 21180 35816
rect 20772 35776 20778 35788
rect 21174 35776 21180 35788
rect 21232 35776 21238 35828
rect 12897 35751 12955 35757
rect 12897 35717 12909 35751
rect 12943 35748 12955 35751
rect 15746 35748 15752 35760
rect 12943 35720 15752 35748
rect 12943 35717 12955 35720
rect 12897 35711 12955 35717
rect 15746 35708 15752 35720
rect 15804 35708 15810 35760
rect 12802 35689 12808 35692
rect 12621 35683 12679 35689
rect 12621 35649 12633 35683
rect 12667 35649 12679 35683
rect 12621 35643 12679 35649
rect 12769 35683 12808 35689
rect 12769 35649 12781 35683
rect 12769 35643 12808 35649
rect 12802 35640 12808 35643
rect 12860 35640 12866 35692
rect 12989 35683 13047 35689
rect 12989 35649 13001 35683
rect 13035 35649 13047 35683
rect 12989 35643 13047 35649
rect 10321 35615 10379 35621
rect 10321 35581 10333 35615
rect 10367 35581 10379 35615
rect 10321 35575 10379 35581
rect 3053 35547 3111 35553
rect 3053 35513 3065 35547
rect 3099 35513 3111 35547
rect 10336 35544 10364 35575
rect 10502 35544 10508 35556
rect 3053 35507 3111 35513
rect 3620 35516 6592 35544
rect 10336 35516 10508 35544
rect 2222 35476 2228 35488
rect 2183 35448 2228 35476
rect 2222 35436 2228 35448
rect 2280 35436 2286 35488
rect 2409 35479 2467 35485
rect 2409 35445 2421 35479
rect 2455 35476 2467 35479
rect 3620 35476 3648 35516
rect 2455 35448 3648 35476
rect 3697 35479 3755 35485
rect 2455 35445 2467 35448
rect 2409 35439 2467 35445
rect 3697 35445 3709 35479
rect 3743 35476 3755 35479
rect 3786 35476 3792 35488
rect 3743 35448 3792 35476
rect 3743 35445 3755 35448
rect 3697 35439 3755 35445
rect 3786 35436 3792 35448
rect 3844 35436 3850 35488
rect 4709 35479 4767 35485
rect 4709 35445 4721 35479
rect 4755 35476 4767 35479
rect 4890 35476 4896 35488
rect 4755 35448 4896 35476
rect 4755 35445 4767 35448
rect 4709 35439 4767 35445
rect 4890 35436 4896 35448
rect 4948 35436 4954 35488
rect 6270 35436 6276 35488
rect 6328 35476 6334 35488
rect 6457 35479 6515 35485
rect 6457 35476 6469 35479
rect 6328 35448 6469 35476
rect 6328 35436 6334 35448
rect 6457 35445 6469 35448
rect 6503 35445 6515 35479
rect 6564 35476 6592 35516
rect 10502 35504 10508 35516
rect 10560 35504 10566 35556
rect 12894 35544 12900 35556
rect 12406 35516 12900 35544
rect 8478 35476 8484 35488
rect 6564 35448 8484 35476
rect 6457 35439 6515 35445
rect 8478 35436 8484 35448
rect 8536 35436 8542 35488
rect 10134 35436 10140 35488
rect 10192 35476 10198 35488
rect 11885 35479 11943 35485
rect 11885 35476 11897 35479
rect 10192 35448 11897 35476
rect 10192 35436 10198 35448
rect 11885 35445 11897 35448
rect 11931 35476 11943 35479
rect 12406 35476 12434 35516
rect 12894 35504 12900 35516
rect 12952 35504 12958 35556
rect 11931 35448 12434 35476
rect 11931 35445 11943 35448
rect 11885 35439 11943 35445
rect 12710 35436 12716 35488
rect 12768 35476 12774 35488
rect 13004 35476 13032 35643
rect 13078 35640 13084 35692
rect 13136 35689 13142 35692
rect 13136 35680 13144 35689
rect 13136 35652 13181 35680
rect 13136 35643 13144 35652
rect 13136 35640 13142 35643
rect 16574 35640 16580 35692
rect 16632 35680 16638 35692
rect 17037 35683 17095 35689
rect 17037 35680 17049 35683
rect 16632 35652 17049 35680
rect 16632 35640 16638 35652
rect 17037 35649 17049 35652
rect 17083 35649 17095 35683
rect 17037 35643 17095 35649
rect 18141 35683 18199 35689
rect 18141 35649 18153 35683
rect 18187 35680 18199 35683
rect 18230 35680 18236 35692
rect 18187 35652 18236 35680
rect 18187 35649 18199 35652
rect 18141 35643 18199 35649
rect 18230 35640 18236 35652
rect 18288 35640 18294 35692
rect 18414 35689 18420 35692
rect 18408 35643 18420 35689
rect 18472 35680 18478 35692
rect 20254 35680 20260 35692
rect 18472 35652 18508 35680
rect 20215 35652 20260 35680
rect 18414 35640 18420 35643
rect 18472 35640 18478 35652
rect 20254 35640 20260 35652
rect 20312 35640 20318 35692
rect 20441 35683 20499 35689
rect 20441 35649 20453 35683
rect 20487 35680 20499 35683
rect 20622 35680 20628 35692
rect 20487 35652 20628 35680
rect 20487 35649 20499 35652
rect 20441 35643 20499 35649
rect 20622 35640 20628 35652
rect 20680 35640 20686 35692
rect 16666 35572 16672 35624
rect 16724 35612 16730 35624
rect 16761 35615 16819 35621
rect 16761 35612 16773 35615
rect 16724 35584 16773 35612
rect 16724 35572 16730 35584
rect 16761 35581 16773 35584
rect 16807 35581 16819 35615
rect 16942 35612 16948 35624
rect 16903 35584 16948 35612
rect 16761 35575 16819 35581
rect 16942 35572 16948 35584
rect 17000 35572 17006 35624
rect 12768 35448 13032 35476
rect 13265 35479 13323 35485
rect 12768 35436 12774 35448
rect 13265 35445 13277 35479
rect 13311 35476 13323 35479
rect 14366 35476 14372 35488
rect 13311 35448 14372 35476
rect 13311 35445 13323 35448
rect 13265 35439 13323 35445
rect 14366 35436 14372 35448
rect 14424 35436 14430 35488
rect 17310 35436 17316 35488
rect 17368 35476 17374 35488
rect 17405 35479 17463 35485
rect 17405 35476 17417 35479
rect 17368 35448 17417 35476
rect 17368 35436 17374 35448
rect 17405 35445 17417 35448
rect 17451 35445 17463 35479
rect 17405 35439 17463 35445
rect 1104 35386 30820 35408
rect 1104 35334 5915 35386
rect 5967 35334 5979 35386
rect 6031 35334 6043 35386
rect 6095 35334 6107 35386
rect 6159 35334 6171 35386
rect 6223 35334 15846 35386
rect 15898 35334 15910 35386
rect 15962 35334 15974 35386
rect 16026 35334 16038 35386
rect 16090 35334 16102 35386
rect 16154 35334 25776 35386
rect 25828 35334 25840 35386
rect 25892 35334 25904 35386
rect 25956 35334 25968 35386
rect 26020 35334 26032 35386
rect 26084 35334 30820 35386
rect 1104 35312 30820 35334
rect 2222 35272 2228 35284
rect 2183 35244 2228 35272
rect 2222 35232 2228 35244
rect 2280 35232 2286 35284
rect 2409 35275 2467 35281
rect 2409 35241 2421 35275
rect 2455 35272 2467 35275
rect 3510 35272 3516 35284
rect 2455 35244 3516 35272
rect 2455 35241 2467 35244
rect 2409 35235 2467 35241
rect 3510 35232 3516 35244
rect 3568 35232 3574 35284
rect 5626 35232 5632 35284
rect 5684 35272 5690 35284
rect 5813 35275 5871 35281
rect 5813 35272 5825 35275
rect 5684 35244 5825 35272
rect 5684 35232 5690 35244
rect 5813 35241 5825 35244
rect 5859 35272 5871 35275
rect 8018 35272 8024 35284
rect 5859 35244 8024 35272
rect 5859 35241 5871 35244
rect 5813 35235 5871 35241
rect 8018 35232 8024 35244
rect 8076 35232 8082 35284
rect 8386 35272 8392 35284
rect 8347 35244 8392 35272
rect 8386 35232 8392 35244
rect 8444 35232 8450 35284
rect 10318 35232 10324 35284
rect 10376 35272 10382 35284
rect 10597 35275 10655 35281
rect 10597 35272 10609 35275
rect 10376 35244 10609 35272
rect 10376 35232 10382 35244
rect 10597 35241 10609 35244
rect 10643 35241 10655 35275
rect 10597 35235 10655 35241
rect 12894 35232 12900 35284
rect 12952 35272 12958 35284
rect 16574 35272 16580 35284
rect 12952 35244 16436 35272
rect 16535 35244 16580 35272
rect 12952 35232 12958 35244
rect 1857 35207 1915 35213
rect 1857 35173 1869 35207
rect 1903 35204 1915 35207
rect 1946 35204 1952 35216
rect 1903 35176 1952 35204
rect 1903 35173 1915 35176
rect 1857 35167 1915 35173
rect 1946 35164 1952 35176
rect 2004 35164 2010 35216
rect 8294 35204 8300 35216
rect 7944 35176 8300 35204
rect 3786 35136 3792 35148
rect 3747 35108 3792 35136
rect 3786 35096 3792 35108
rect 3844 35096 3850 35148
rect 7944 35145 7972 35176
rect 8294 35164 8300 35176
rect 8352 35204 8358 35216
rect 8846 35204 8852 35216
rect 8352 35176 8852 35204
rect 8352 35164 8358 35176
rect 8846 35164 8852 35176
rect 8904 35164 8910 35216
rect 15194 35164 15200 35216
rect 15252 35204 15258 35216
rect 16408 35204 16436 35244
rect 16574 35232 16580 35244
rect 16632 35232 16638 35284
rect 20441 35275 20499 35281
rect 20441 35241 20453 35275
rect 20487 35272 20499 35275
rect 20714 35272 20720 35284
rect 20487 35244 20720 35272
rect 20487 35241 20499 35244
rect 20441 35235 20499 35241
rect 20714 35232 20720 35244
rect 20772 35232 20778 35284
rect 17218 35204 17224 35216
rect 15252 35176 15516 35204
rect 16408 35176 17224 35204
rect 15252 35164 15258 35176
rect 7929 35139 7987 35145
rect 7929 35105 7941 35139
rect 7975 35105 7987 35139
rect 9585 35139 9643 35145
rect 7929 35099 7987 35105
rect 8128 35108 8800 35136
rect 2774 35028 2780 35080
rect 2832 35068 2838 35080
rect 2869 35071 2927 35077
rect 2869 35068 2881 35071
rect 2832 35040 2881 35068
rect 2832 35028 2838 35040
rect 2869 35037 2881 35040
rect 2915 35037 2927 35071
rect 4430 35068 4436 35080
rect 2869 35031 2927 35037
rect 3988 35040 4436 35068
rect 2225 35003 2283 35009
rect 2225 34969 2237 35003
rect 2271 35000 2283 35003
rect 3988 35000 4016 35040
rect 4430 35028 4436 35040
rect 4488 35028 4494 35080
rect 5997 35071 6055 35077
rect 5997 35037 6009 35071
rect 6043 35068 6055 35071
rect 6549 35071 6607 35077
rect 6549 35068 6561 35071
rect 6043 35040 6561 35068
rect 6043 35037 6055 35040
rect 5997 35031 6055 35037
rect 6549 35037 6561 35040
rect 6595 35037 6607 35071
rect 6549 35031 6607 35037
rect 6638 35028 6644 35080
rect 6696 35068 6702 35080
rect 7650 35068 7656 35080
rect 6696 35040 6741 35068
rect 7611 35040 7656 35068
rect 6696 35028 6702 35040
rect 7650 35028 7656 35040
rect 7708 35028 7714 35080
rect 8128 35078 8156 35108
rect 8772 35080 8800 35108
rect 9585 35105 9597 35139
rect 9631 35136 9643 35139
rect 9950 35136 9956 35148
rect 9631 35108 9956 35136
rect 9631 35105 9643 35108
rect 9585 35099 9643 35105
rect 9950 35096 9956 35108
rect 10008 35136 10014 35148
rect 10502 35136 10508 35148
rect 10008 35108 10508 35136
rect 10008 35096 10014 35108
rect 10502 35096 10508 35108
rect 10560 35096 10566 35148
rect 15378 35136 15384 35148
rect 15339 35108 15384 35136
rect 15378 35096 15384 35108
rect 15436 35096 15442 35148
rect 15488 35136 15516 35176
rect 17218 35164 17224 35176
rect 17276 35164 17282 35216
rect 15774 35139 15832 35145
rect 15774 35136 15786 35139
rect 15488 35108 15786 35136
rect 15774 35105 15786 35108
rect 15820 35105 15832 35139
rect 16298 35136 16304 35148
rect 15774 35099 15832 35105
rect 15948 35108 16304 35136
rect 15948 35080 15976 35108
rect 16298 35096 16304 35108
rect 16356 35136 16362 35148
rect 17129 35139 17187 35145
rect 17129 35136 17141 35139
rect 16356 35108 17141 35136
rect 16356 35096 16362 35108
rect 17129 35105 17141 35108
rect 17175 35105 17187 35139
rect 17310 35136 17316 35148
rect 17271 35108 17316 35136
rect 17129 35099 17187 35105
rect 17310 35096 17316 35108
rect 17368 35136 17374 35148
rect 20732 35136 20760 35232
rect 17368 35108 18276 35136
rect 20732 35108 21220 35136
rect 17368 35096 17374 35108
rect 8036 35077 8156 35078
rect 8202 35077 8208 35080
rect 8021 35071 8156 35077
rect 7837 35065 7895 35071
rect 7837 35031 7849 35065
rect 7883 35031 7895 35065
rect 8021 35037 8033 35071
rect 8067 35050 8156 35071
rect 8067 35037 8079 35050
rect 8021 35031 8079 35037
rect 7837 35025 7895 35031
rect 4062 35009 4068 35012
rect 2271 34972 4016 35000
rect 2271 34969 2283 34972
rect 2225 34963 2283 34969
rect 4056 34963 4068 35009
rect 4120 35000 4126 35012
rect 4120 34972 4156 35000
rect 4062 34960 4068 34963
rect 4120 34960 4126 34972
rect 3050 34932 3056 34944
rect 3011 34904 3056 34932
rect 3050 34892 3056 34904
rect 3108 34892 3114 34944
rect 3786 34892 3792 34944
rect 3844 34932 3850 34944
rect 5169 34935 5227 34941
rect 5169 34932 5181 34935
rect 3844 34904 5181 34932
rect 3844 34892 3850 34904
rect 5169 34901 5181 34904
rect 5215 34901 5227 34935
rect 7852 34932 7880 35025
rect 7926 34960 7932 35012
rect 7984 35000 7990 35012
rect 8128 35000 8156 35050
rect 8188 35071 8208 35077
rect 8188 35037 8200 35071
rect 8188 35031 8208 35037
rect 8202 35028 8208 35031
rect 8260 35028 8266 35080
rect 8754 35028 8760 35080
rect 8812 35068 8818 35080
rect 9309 35071 9367 35077
rect 9309 35068 9321 35071
rect 8812 35040 9321 35068
rect 8812 35028 8818 35040
rect 9309 35037 9321 35040
rect 9355 35037 9367 35071
rect 10778 35068 10784 35080
rect 10739 35040 10784 35068
rect 9309 35031 9367 35037
rect 10778 35028 10784 35040
rect 10836 35028 10842 35080
rect 11606 35028 11612 35080
rect 11664 35068 11670 35080
rect 11701 35071 11759 35077
rect 11701 35068 11713 35071
rect 11664 35040 11713 35068
rect 11664 35028 11670 35040
rect 11701 35037 11713 35040
rect 11747 35037 11759 35071
rect 11701 35031 11759 35037
rect 14642 35028 14648 35080
rect 14700 35068 14706 35080
rect 14737 35071 14795 35077
rect 14737 35068 14749 35071
rect 14700 35040 14749 35068
rect 14700 35028 14706 35040
rect 14737 35037 14749 35040
rect 14783 35037 14795 35071
rect 14737 35031 14795 35037
rect 14921 35071 14979 35077
rect 14921 35037 14933 35071
rect 14967 35037 14979 35071
rect 14921 35031 14979 35037
rect 7984 34972 8156 35000
rect 11968 35003 12026 35009
rect 7984 34960 7990 34972
rect 11968 34969 11980 35003
rect 12014 35000 12026 35003
rect 12066 35000 12072 35012
rect 12014 34972 12072 35000
rect 12014 34969 12026 34972
rect 11968 34963 12026 34969
rect 12066 34960 12072 34972
rect 12124 34960 12130 35012
rect 13722 35000 13728 35012
rect 13096 34972 13728 35000
rect 8662 34932 8668 34944
rect 7852 34904 8668 34932
rect 5169 34895 5227 34901
rect 8662 34892 8668 34904
rect 8720 34892 8726 34944
rect 13096 34941 13124 34972
rect 13722 34960 13728 34972
rect 13780 35000 13786 35012
rect 14458 35000 14464 35012
rect 13780 34972 14464 35000
rect 13780 34960 13786 34972
rect 14458 34960 14464 34972
rect 14516 35000 14522 35012
rect 14936 35000 14964 35031
rect 15654 35028 15660 35080
rect 15712 35068 15718 35080
rect 15930 35068 15936 35080
rect 15712 35040 15757 35068
rect 15891 35040 15936 35068
rect 15712 35028 15718 35040
rect 15930 35028 15936 35040
rect 15988 35028 15994 35080
rect 18248 35077 18276 35108
rect 18233 35071 18291 35077
rect 18233 35037 18245 35071
rect 18279 35037 18291 35071
rect 18233 35031 18291 35037
rect 20257 35071 20315 35077
rect 20257 35037 20269 35071
rect 20303 35037 20315 35071
rect 20257 35031 20315 35037
rect 14516 34972 14964 35000
rect 18417 35003 18475 35009
rect 14516 34960 14522 34972
rect 18417 34969 18429 35003
rect 18463 35000 18475 35003
rect 18506 35000 18512 35012
rect 18463 34972 18512 35000
rect 18463 34969 18475 34972
rect 18417 34963 18475 34969
rect 18506 34960 18512 34972
rect 18564 34960 18570 35012
rect 20272 35000 20300 35031
rect 20438 35028 20444 35080
rect 20496 35068 20502 35080
rect 21192 35077 21220 35108
rect 20533 35071 20591 35077
rect 20533 35068 20545 35071
rect 20496 35040 20545 35068
rect 20496 35028 20502 35040
rect 20533 35037 20545 35040
rect 20579 35068 20591 35071
rect 20993 35071 21051 35077
rect 20993 35068 21005 35071
rect 20579 35040 21005 35068
rect 20579 35037 20591 35040
rect 20533 35031 20591 35037
rect 20993 35037 21005 35040
rect 21039 35037 21051 35071
rect 20993 35031 21051 35037
rect 21177 35071 21235 35077
rect 21177 35037 21189 35071
rect 21223 35037 21235 35071
rect 21177 35031 21235 35037
rect 22097 35071 22155 35077
rect 22097 35037 22109 35071
rect 22143 35068 22155 35071
rect 22186 35068 22192 35080
rect 22143 35040 22192 35068
rect 22143 35037 22155 35040
rect 22097 35031 22155 35037
rect 22186 35028 22192 35040
rect 22244 35028 22250 35080
rect 22281 35071 22339 35077
rect 22281 35037 22293 35071
rect 22327 35068 22339 35071
rect 30098 35068 30104 35080
rect 22327 35040 26234 35068
rect 30059 35040 30104 35068
rect 22327 35037 22339 35040
rect 22281 35031 22339 35037
rect 20622 35000 20628 35012
rect 20272 34972 20628 35000
rect 20622 34960 20628 34972
rect 20680 35000 20686 35012
rect 21085 35003 21143 35009
rect 21085 35000 21097 35003
rect 20680 34972 21097 35000
rect 20680 34960 20686 34972
rect 21085 34969 21097 34972
rect 21131 34969 21143 35003
rect 21085 34963 21143 34969
rect 13081 34935 13139 34941
rect 13081 34901 13093 34935
rect 13127 34901 13139 34935
rect 13081 34895 13139 34901
rect 14642 34892 14648 34944
rect 14700 34932 14706 34944
rect 14918 34932 14924 34944
rect 14700 34904 14924 34932
rect 14700 34892 14706 34904
rect 14918 34892 14924 34904
rect 14976 34932 14982 34944
rect 15654 34932 15660 34944
rect 14976 34904 15660 34932
rect 14976 34892 14982 34904
rect 15654 34892 15660 34904
rect 15712 34892 15718 34944
rect 17402 34892 17408 34944
rect 17460 34932 17466 34944
rect 17773 34935 17831 34941
rect 17460 34904 17505 34932
rect 17460 34892 17466 34904
rect 17773 34901 17785 34935
rect 17819 34932 17831 34935
rect 18322 34932 18328 34944
rect 17819 34904 18328 34932
rect 17819 34901 17831 34904
rect 17773 34895 17831 34901
rect 18322 34892 18328 34904
rect 18380 34892 18386 34944
rect 18598 34932 18604 34944
rect 18559 34904 18604 34932
rect 18598 34892 18604 34904
rect 18656 34892 18662 34944
rect 19978 34892 19984 34944
rect 20036 34932 20042 34944
rect 20073 34935 20131 34941
rect 20073 34932 20085 34935
rect 20036 34904 20085 34932
rect 20036 34892 20042 34904
rect 20073 34901 20085 34904
rect 20119 34901 20131 34935
rect 21910 34932 21916 34944
rect 21871 34904 21916 34932
rect 20073 34895 20131 34901
rect 21910 34892 21916 34904
rect 21968 34892 21974 34944
rect 26206 34932 26234 35040
rect 30098 35028 30104 35040
rect 30156 35028 30162 35080
rect 29917 34935 29975 34941
rect 29917 34932 29929 34935
rect 26206 34904 29929 34932
rect 29917 34901 29929 34904
rect 29963 34901 29975 34935
rect 29917 34895 29975 34901
rect 1104 34842 30820 34864
rect 1104 34790 10880 34842
rect 10932 34790 10944 34842
rect 10996 34790 11008 34842
rect 11060 34790 11072 34842
rect 11124 34790 11136 34842
rect 11188 34790 20811 34842
rect 20863 34790 20875 34842
rect 20927 34790 20939 34842
rect 20991 34790 21003 34842
rect 21055 34790 21067 34842
rect 21119 34790 30820 34842
rect 1104 34768 30820 34790
rect 1854 34688 1860 34740
rect 1912 34728 1918 34740
rect 2409 34731 2467 34737
rect 2409 34728 2421 34731
rect 1912 34700 2421 34728
rect 1912 34688 1918 34700
rect 2409 34697 2421 34700
rect 2455 34697 2467 34731
rect 2409 34691 2467 34697
rect 3973 34731 4031 34737
rect 3973 34697 3985 34731
rect 4019 34728 4031 34731
rect 4062 34728 4068 34740
rect 4019 34700 4068 34728
rect 4019 34697 4031 34700
rect 3973 34691 4031 34697
rect 4062 34688 4068 34700
rect 4120 34688 4126 34740
rect 4430 34728 4436 34740
rect 4391 34700 4436 34728
rect 4430 34688 4436 34700
rect 4488 34728 4494 34740
rect 5810 34728 5816 34740
rect 4488 34700 5816 34728
rect 4488 34688 4494 34700
rect 5810 34688 5816 34700
rect 5868 34688 5874 34740
rect 6365 34731 6423 34737
rect 6365 34697 6377 34731
rect 6411 34728 6423 34731
rect 6822 34728 6828 34740
rect 6411 34700 6828 34728
rect 6411 34697 6423 34700
rect 6365 34691 6423 34697
rect 6822 34688 6828 34700
rect 6880 34688 6886 34740
rect 7009 34731 7067 34737
rect 7009 34697 7021 34731
rect 7055 34728 7067 34731
rect 7834 34728 7840 34740
rect 7055 34700 7840 34728
rect 7055 34697 7067 34700
rect 7009 34691 7067 34697
rect 2225 34663 2283 34669
rect 2225 34629 2237 34663
rect 2271 34660 2283 34663
rect 2271 34632 3843 34660
rect 2271 34629 2283 34632
rect 2225 34623 2283 34629
rect 3815 34604 3843 34632
rect 4706 34620 4712 34672
rect 4764 34660 4770 34672
rect 4764 34632 5856 34660
rect 4764 34620 4770 34632
rect 1857 34595 1915 34601
rect 1857 34561 1869 34595
rect 1903 34592 1915 34595
rect 1946 34592 1952 34604
rect 1903 34564 1952 34592
rect 1903 34561 1915 34564
rect 1857 34555 1915 34561
rect 1946 34552 1952 34564
rect 2004 34552 2010 34604
rect 3237 34595 3295 34601
rect 3237 34561 3249 34595
rect 3283 34561 3295 34595
rect 3418 34592 3424 34604
rect 3379 34564 3424 34592
rect 3237 34555 3295 34561
rect 3252 34524 3280 34555
rect 3418 34552 3424 34564
rect 3476 34552 3482 34604
rect 3510 34552 3516 34604
rect 3568 34592 3574 34604
rect 3568 34564 3613 34592
rect 3568 34552 3574 34564
rect 3786 34552 3792 34604
rect 3844 34592 3850 34604
rect 5557 34595 5615 34601
rect 3844 34564 3889 34592
rect 3844 34552 3850 34564
rect 5557 34561 5569 34595
rect 5603 34592 5615 34595
rect 5718 34592 5724 34604
rect 5603 34564 5724 34592
rect 5603 34561 5615 34564
rect 5557 34555 5615 34561
rect 5718 34552 5724 34564
rect 5776 34552 5782 34604
rect 5828 34601 5856 34632
rect 5813 34595 5871 34601
rect 5813 34561 5825 34595
rect 5859 34561 5871 34595
rect 5813 34555 5871 34561
rect 6270 34552 6276 34604
rect 6328 34592 6334 34604
rect 6549 34595 6607 34601
rect 6549 34592 6561 34595
rect 6328 34564 6561 34592
rect 6328 34552 6334 34564
rect 6549 34561 6561 34564
rect 6595 34592 6607 34595
rect 7024 34592 7052 34691
rect 7834 34688 7840 34700
rect 7892 34688 7898 34740
rect 8754 34728 8760 34740
rect 8715 34700 8760 34728
rect 8754 34688 8760 34700
rect 8812 34688 8818 34740
rect 13354 34688 13360 34740
rect 13412 34728 13418 34740
rect 13725 34731 13783 34737
rect 13725 34728 13737 34731
rect 13412 34700 13737 34728
rect 13412 34688 13418 34700
rect 13725 34697 13737 34700
rect 13771 34697 13783 34731
rect 13725 34691 13783 34697
rect 16117 34731 16175 34737
rect 16117 34697 16129 34731
rect 16163 34728 16175 34731
rect 16942 34728 16948 34740
rect 16163 34700 16948 34728
rect 16163 34697 16175 34700
rect 16117 34691 16175 34697
rect 16942 34688 16948 34700
rect 17000 34688 17006 34740
rect 17037 34731 17095 34737
rect 17037 34697 17049 34731
rect 17083 34728 17095 34731
rect 17402 34728 17408 34740
rect 17083 34700 17408 34728
rect 17083 34697 17095 34700
rect 17037 34691 17095 34697
rect 17402 34688 17408 34700
rect 17460 34688 17466 34740
rect 18877 34731 18935 34737
rect 18877 34697 18889 34731
rect 18923 34697 18935 34731
rect 18877 34691 18935 34697
rect 12618 34669 12624 34672
rect 11609 34663 11667 34669
rect 11609 34660 11621 34663
rect 7208 34632 11621 34660
rect 7208 34601 7236 34632
rect 11609 34629 11621 34632
rect 11655 34629 11667 34663
rect 12612 34660 12624 34669
rect 12579 34632 12624 34660
rect 11609 34623 11667 34629
rect 12612 34623 12624 34632
rect 12618 34620 12624 34623
rect 12676 34620 12682 34672
rect 18598 34660 18604 34672
rect 16868 34632 18604 34660
rect 6595 34564 7052 34592
rect 7193 34595 7251 34601
rect 6595 34561 6607 34564
rect 6549 34555 6607 34561
rect 7193 34561 7205 34595
rect 7239 34561 7251 34595
rect 7193 34555 7251 34561
rect 7837 34595 7895 34601
rect 7837 34561 7849 34595
rect 7883 34592 7895 34595
rect 8018 34592 8024 34604
rect 7883 34564 8024 34592
rect 7883 34561 7895 34564
rect 7837 34555 7895 34561
rect 8018 34552 8024 34564
rect 8076 34552 8082 34604
rect 8662 34592 8668 34604
rect 8623 34564 8668 34592
rect 8662 34552 8668 34564
rect 8720 34592 8726 34604
rect 8720 34564 8800 34592
rect 8720 34552 8726 34564
rect 3602 34524 3608 34536
rect 3252 34496 3464 34524
rect 3563 34496 3608 34524
rect 3436 34456 3464 34496
rect 3602 34484 3608 34496
rect 3660 34484 3666 34536
rect 4522 34524 4528 34536
rect 3712 34496 4528 34524
rect 3712 34456 3740 34496
rect 4522 34484 4528 34496
rect 4580 34484 4586 34536
rect 7650 34484 7656 34536
rect 7708 34524 7714 34536
rect 8478 34524 8484 34536
rect 7708 34496 8484 34524
rect 7708 34484 7714 34496
rect 8478 34484 8484 34496
rect 8536 34484 8542 34536
rect 3436 34428 3740 34456
rect 8772 34456 8800 34564
rect 8938 34552 8944 34604
rect 8996 34592 9002 34604
rect 11517 34595 11575 34601
rect 11517 34592 11529 34595
rect 8996 34564 11529 34592
rect 8996 34552 9002 34564
rect 11517 34561 11529 34564
rect 11563 34561 11575 34595
rect 11517 34555 11575 34561
rect 11698 34552 11704 34604
rect 11756 34592 11762 34604
rect 13078 34592 13084 34604
rect 11756 34564 13084 34592
rect 11756 34552 11762 34564
rect 13078 34552 13084 34564
rect 13136 34552 13142 34604
rect 14458 34592 14464 34604
rect 14419 34564 14464 34592
rect 14458 34552 14464 34564
rect 14516 34552 14522 34604
rect 15286 34552 15292 34604
rect 15344 34601 15350 34604
rect 16868 34601 16896 34632
rect 18598 34620 18604 34632
rect 18656 34620 18662 34672
rect 18892 34660 18920 34691
rect 19150 34688 19156 34740
rect 19208 34728 19214 34740
rect 19521 34731 19579 34737
rect 19521 34728 19533 34731
rect 19208 34700 19533 34728
rect 19208 34688 19214 34700
rect 19521 34697 19533 34700
rect 19567 34697 19579 34731
rect 19521 34691 19579 34697
rect 20346 34688 20352 34740
rect 20404 34728 20410 34740
rect 20533 34731 20591 34737
rect 20533 34728 20545 34731
rect 20404 34700 20545 34728
rect 20404 34688 20410 34700
rect 20533 34697 20545 34700
rect 20579 34697 20591 34731
rect 20714 34728 20720 34740
rect 20675 34700 20720 34728
rect 20533 34691 20591 34697
rect 20714 34688 20720 34700
rect 20772 34688 20778 34740
rect 20809 34731 20867 34737
rect 20809 34697 20821 34731
rect 20855 34728 20867 34731
rect 21174 34728 21180 34740
rect 20855 34700 21180 34728
rect 20855 34697 20867 34700
rect 20809 34691 20867 34697
rect 21174 34688 21180 34700
rect 21232 34688 21238 34740
rect 20438 34660 20444 34672
rect 18892 34632 20444 34660
rect 20438 34620 20444 34632
rect 20496 34620 20502 34672
rect 20622 34660 20628 34672
rect 20583 34632 20628 34660
rect 20622 34620 20628 34632
rect 20680 34620 20686 34672
rect 15344 34595 15372 34601
rect 15360 34561 15372 34595
rect 15344 34555 15372 34561
rect 16853 34595 16911 34601
rect 16853 34561 16865 34595
rect 16899 34561 16911 34595
rect 16853 34555 16911 34561
rect 17764 34595 17822 34601
rect 17764 34561 17776 34595
rect 17810 34592 17822 34595
rect 18046 34592 18052 34604
rect 17810 34564 18052 34592
rect 17810 34561 17822 34564
rect 17764 34555 17822 34561
rect 15344 34552 15350 34555
rect 18046 34552 18052 34564
rect 18104 34552 18110 34604
rect 19518 34595 19576 34601
rect 19518 34561 19530 34595
rect 19564 34592 19576 34595
rect 19610 34592 19616 34604
rect 19564 34564 19616 34592
rect 19564 34561 19576 34564
rect 19518 34555 19576 34561
rect 19610 34552 19616 34564
rect 19668 34552 19674 34604
rect 20990 34592 20996 34604
rect 20951 34564 20996 34592
rect 20990 34552 20996 34564
rect 21048 34552 21054 34604
rect 9858 34524 9864 34536
rect 9819 34496 9864 34524
rect 9858 34484 9864 34496
rect 9916 34484 9922 34536
rect 10134 34524 10140 34536
rect 10047 34496 10140 34524
rect 10134 34484 10140 34496
rect 10192 34524 10198 34536
rect 10410 34524 10416 34536
rect 10192 34496 10416 34524
rect 10192 34484 10198 34496
rect 10410 34484 10416 34496
rect 10468 34484 10474 34536
rect 11606 34484 11612 34536
rect 11664 34524 11670 34536
rect 12345 34527 12403 34533
rect 12345 34524 12357 34527
rect 11664 34496 12357 34524
rect 11664 34484 11670 34496
rect 12345 34493 12357 34496
rect 12391 34493 12403 34527
rect 12345 34487 12403 34493
rect 14182 34484 14188 34536
rect 14240 34524 14246 34536
rect 14277 34527 14335 34533
rect 14277 34524 14289 34527
rect 14240 34496 14289 34524
rect 14240 34484 14246 34496
rect 14277 34493 14289 34496
rect 14323 34524 14335 34527
rect 14642 34524 14648 34536
rect 14323 34496 14648 34524
rect 14323 34493 14335 34496
rect 14277 34487 14335 34493
rect 14642 34484 14648 34496
rect 14700 34524 14706 34536
rect 15197 34527 15255 34533
rect 15197 34524 15209 34527
rect 14700 34496 15209 34524
rect 14700 34484 14706 34496
rect 15197 34493 15209 34496
rect 15243 34493 15255 34527
rect 15197 34487 15255 34493
rect 15473 34527 15531 34533
rect 15473 34493 15485 34527
rect 15519 34524 15531 34527
rect 15654 34524 15660 34536
rect 15519 34496 15660 34524
rect 15519 34493 15531 34496
rect 15473 34487 15531 34493
rect 15654 34484 15660 34496
rect 15712 34524 15718 34536
rect 15838 34524 15844 34536
rect 15712 34496 15844 34524
rect 15712 34484 15718 34496
rect 15838 34484 15844 34496
rect 15896 34484 15902 34536
rect 17494 34524 17500 34536
rect 17455 34496 17500 34524
rect 17494 34484 17500 34496
rect 17552 34484 17558 34536
rect 19981 34527 20039 34533
rect 19981 34493 19993 34527
rect 20027 34524 20039 34527
rect 20070 34524 20076 34536
rect 20027 34496 20076 34524
rect 20027 34493 20039 34496
rect 19981 34487 20039 34493
rect 20070 34484 20076 34496
rect 20128 34484 20134 34536
rect 9876 34456 9904 34484
rect 14921 34459 14979 34465
rect 8772 34428 9904 34456
rect 13648 34428 13860 34456
rect 2222 34388 2228 34400
rect 2183 34360 2228 34388
rect 2222 34348 2228 34360
rect 2280 34348 2286 34400
rect 7650 34388 7656 34400
rect 7611 34360 7656 34388
rect 7650 34348 7656 34360
rect 7708 34348 7714 34400
rect 9030 34348 9036 34400
rect 9088 34388 9094 34400
rect 13648 34388 13676 34428
rect 9088 34360 13676 34388
rect 13832 34388 13860 34428
rect 14921 34425 14933 34459
rect 14967 34456 14979 34459
rect 15010 34456 15016 34468
rect 14967 34428 15016 34456
rect 14967 34425 14979 34428
rect 14921 34419 14979 34425
rect 15010 34416 15016 34428
rect 15068 34416 15074 34468
rect 18432 34428 20024 34456
rect 18432 34388 18460 34428
rect 19334 34388 19340 34400
rect 13832 34360 18460 34388
rect 19295 34360 19340 34388
rect 9088 34348 9094 34360
rect 19334 34348 19340 34360
rect 19392 34348 19398 34400
rect 19886 34388 19892 34400
rect 19847 34360 19892 34388
rect 19886 34348 19892 34360
rect 19944 34348 19950 34400
rect 19996 34388 20024 34428
rect 21910 34388 21916 34400
rect 19996 34360 21916 34388
rect 21910 34348 21916 34360
rect 21968 34348 21974 34400
rect 1104 34298 30820 34320
rect 1104 34246 5915 34298
rect 5967 34246 5979 34298
rect 6031 34246 6043 34298
rect 6095 34246 6107 34298
rect 6159 34246 6171 34298
rect 6223 34246 15846 34298
rect 15898 34246 15910 34298
rect 15962 34246 15974 34298
rect 16026 34246 16038 34298
rect 16090 34246 16102 34298
rect 16154 34246 25776 34298
rect 25828 34246 25840 34298
rect 25892 34246 25904 34298
rect 25956 34246 25968 34298
rect 26020 34246 26032 34298
rect 26084 34246 30820 34298
rect 1104 34224 30820 34246
rect 2222 34184 2228 34196
rect 2183 34156 2228 34184
rect 2222 34144 2228 34156
rect 2280 34144 2286 34196
rect 2409 34187 2467 34193
rect 2409 34153 2421 34187
rect 2455 34184 2467 34187
rect 3970 34184 3976 34196
rect 2455 34156 3976 34184
rect 2455 34153 2467 34156
rect 2409 34147 2467 34153
rect 3970 34144 3976 34156
rect 4028 34144 4034 34196
rect 5629 34187 5687 34193
rect 5629 34153 5641 34187
rect 5675 34184 5687 34187
rect 5718 34184 5724 34196
rect 5675 34156 5724 34184
rect 5675 34153 5687 34156
rect 5629 34147 5687 34153
rect 5718 34144 5724 34156
rect 5776 34144 5782 34196
rect 7193 34187 7251 34193
rect 7193 34153 7205 34187
rect 7239 34184 7251 34187
rect 8110 34184 8116 34196
rect 7239 34156 8116 34184
rect 7239 34153 7251 34156
rect 7193 34147 7251 34153
rect 8110 34144 8116 34156
rect 8168 34144 8174 34196
rect 8938 34184 8944 34196
rect 8220 34156 8944 34184
rect 1857 34119 1915 34125
rect 1857 34085 1869 34119
rect 1903 34116 1915 34119
rect 1946 34116 1952 34128
rect 1903 34088 1952 34116
rect 1903 34085 1915 34088
rect 1857 34079 1915 34085
rect 1946 34076 1952 34088
rect 2004 34076 2010 34128
rect 6089 34051 6147 34057
rect 6089 34048 6101 34051
rect 4816 34020 6101 34048
rect 3142 33980 3148 33992
rect 3103 33952 3148 33980
rect 3142 33940 3148 33952
rect 3200 33940 3206 33992
rect 3786 33980 3792 33992
rect 3747 33952 3792 33980
rect 3786 33940 3792 33952
rect 3844 33940 3850 33992
rect 4430 33940 4436 33992
rect 4488 33980 4494 33992
rect 4816 33980 4844 34020
rect 6089 34017 6101 34020
rect 6135 34017 6147 34051
rect 6089 34011 6147 34017
rect 7926 34008 7932 34060
rect 7984 34048 7990 34060
rect 8021 34051 8079 34057
rect 8021 34048 8033 34051
rect 7984 34020 8033 34048
rect 7984 34008 7990 34020
rect 8021 34017 8033 34020
rect 8067 34017 8079 34051
rect 8021 34011 8079 34017
rect 5810 33980 5816 33992
rect 4488 33952 4844 33980
rect 5771 33952 5816 33980
rect 4488 33940 4494 33952
rect 5810 33940 5816 33952
rect 5868 33940 5874 33992
rect 5997 33983 6055 33989
rect 5997 33949 6009 33983
rect 6043 33949 6055 33983
rect 5997 33943 6055 33949
rect 2225 33915 2283 33921
rect 2225 33881 2237 33915
rect 2271 33912 2283 33915
rect 2271 33884 3648 33912
rect 2271 33881 2283 33884
rect 2225 33875 2283 33881
rect 2958 33844 2964 33856
rect 2919 33816 2964 33844
rect 2958 33804 2964 33816
rect 3016 33804 3022 33856
rect 3620 33844 3648 33884
rect 3878 33872 3884 33924
rect 3936 33912 3942 33924
rect 4034 33915 4092 33921
rect 4034 33912 4046 33915
rect 3936 33884 4046 33912
rect 3936 33872 3942 33884
rect 4034 33881 4046 33884
rect 4080 33881 4092 33915
rect 4034 33875 4092 33881
rect 4154 33872 4160 33924
rect 4212 33912 4218 33924
rect 6012 33912 6040 33943
rect 6178 33940 6184 33992
rect 6236 33980 6242 33992
rect 6362 33980 6368 33992
rect 6236 33952 6281 33980
rect 6323 33952 6368 33980
rect 6236 33940 6242 33952
rect 6362 33940 6368 33952
rect 6420 33980 6426 33992
rect 6730 33980 6736 33992
rect 6420 33952 6736 33980
rect 6420 33940 6426 33952
rect 6730 33940 6736 33952
rect 6788 33940 6794 33992
rect 7006 33980 7012 33992
rect 6967 33952 7012 33980
rect 7006 33940 7012 33952
rect 7064 33940 7070 33992
rect 7837 33983 7895 33989
rect 7837 33949 7849 33983
rect 7883 33949 7895 33983
rect 8110 33980 8116 33992
rect 8071 33952 8116 33980
rect 7837 33943 7895 33949
rect 4212 33884 6040 33912
rect 7852 33912 7880 33943
rect 8110 33940 8116 33952
rect 8168 33940 8174 33992
rect 8220 33989 8248 34156
rect 8938 34144 8944 34156
rect 8996 34144 9002 34196
rect 9858 34144 9864 34196
rect 9916 34184 9922 34196
rect 18046 34184 18052 34196
rect 9916 34156 16620 34184
rect 18007 34156 18052 34184
rect 9916 34144 9922 34156
rect 8294 34076 8300 34128
rect 8352 34116 8358 34128
rect 9766 34116 9772 34128
rect 8352 34088 9772 34116
rect 8352 34076 8358 34088
rect 9766 34076 9772 34088
rect 9824 34076 9830 34128
rect 8938 34008 8944 34060
rect 8996 34048 9002 34060
rect 9876 34048 9904 34144
rect 15194 34076 15200 34128
rect 15252 34116 15258 34128
rect 15473 34119 15531 34125
rect 15473 34116 15485 34119
rect 15252 34088 15485 34116
rect 15252 34076 15258 34088
rect 15473 34085 15485 34088
rect 15519 34116 15531 34119
rect 15746 34116 15752 34128
rect 15519 34088 15752 34116
rect 15519 34085 15531 34088
rect 15473 34079 15531 34085
rect 15746 34076 15752 34088
rect 15804 34076 15810 34128
rect 16592 34116 16620 34156
rect 18046 34144 18052 34156
rect 18104 34144 18110 34196
rect 18601 34187 18659 34193
rect 18601 34153 18613 34187
rect 18647 34184 18659 34187
rect 20070 34184 20076 34196
rect 18647 34156 20076 34184
rect 18647 34153 18659 34156
rect 18601 34147 18659 34153
rect 20070 34144 20076 34156
rect 20128 34144 20134 34196
rect 20717 34119 20775 34125
rect 20717 34116 20729 34119
rect 16592 34088 20729 34116
rect 20717 34085 20729 34088
rect 20763 34085 20775 34119
rect 20717 34079 20775 34085
rect 20806 34076 20812 34128
rect 20864 34116 20870 34128
rect 22002 34116 22008 34128
rect 20864 34088 22008 34116
rect 20864 34076 20870 34088
rect 22002 34076 22008 34088
rect 22060 34076 22066 34128
rect 12069 34051 12127 34057
rect 12069 34048 12081 34051
rect 8996 34020 9904 34048
rect 11256 34020 12081 34048
rect 8996 34008 9002 34020
rect 8205 33983 8263 33989
rect 8205 33949 8217 33983
rect 8251 33949 8263 33983
rect 8205 33943 8263 33949
rect 8389 33983 8447 33989
rect 8389 33949 8401 33983
rect 8435 33976 8447 33983
rect 8478 33976 8484 33992
rect 8435 33949 8484 33976
rect 8389 33948 8484 33949
rect 8389 33943 8447 33948
rect 8478 33940 8484 33948
rect 8536 33940 8542 33992
rect 9306 33980 9312 33992
rect 9267 33952 9312 33980
rect 9306 33940 9312 33952
rect 9364 33940 9370 33992
rect 11256 33980 11284 34020
rect 12069 34017 12081 34020
rect 12115 34017 12127 34051
rect 19978 34048 19984 34060
rect 19939 34020 19984 34048
rect 12069 34011 12127 34017
rect 19978 34008 19984 34020
rect 20036 34008 20042 34060
rect 20073 34051 20131 34057
rect 20073 34017 20085 34051
rect 20119 34017 20131 34051
rect 20073 34011 20131 34017
rect 10428 33952 11284 33980
rect 11333 33983 11391 33989
rect 8294 33912 8300 33924
rect 7852 33884 8300 33912
rect 4212 33872 4218 33884
rect 8294 33872 8300 33884
rect 8352 33872 8358 33924
rect 8496 33912 8524 33940
rect 10428 33924 10456 33952
rect 11333 33949 11345 33983
rect 11379 33980 11391 33983
rect 11514 33980 11520 33992
rect 11379 33952 11520 33980
rect 11379 33949 11391 33952
rect 11333 33943 11391 33949
rect 11514 33940 11520 33952
rect 11572 33940 11578 33992
rect 11793 33983 11851 33989
rect 11793 33949 11805 33983
rect 11839 33980 11851 33983
rect 11974 33980 11980 33992
rect 11839 33952 11980 33980
rect 11839 33949 11851 33952
rect 11793 33943 11851 33949
rect 11974 33940 11980 33952
rect 12032 33940 12038 33992
rect 14093 33983 14151 33989
rect 14093 33949 14105 33983
rect 14139 33980 14151 33983
rect 17865 33983 17923 33989
rect 14139 33952 14596 33980
rect 14139 33949 14151 33952
rect 14093 33943 14151 33949
rect 14568 33924 14596 33952
rect 17865 33949 17877 33983
rect 17911 33949 17923 33983
rect 17865 33943 17923 33949
rect 18049 33983 18107 33989
rect 18049 33949 18061 33983
rect 18095 33980 18107 33983
rect 18598 33980 18604 33992
rect 18095 33952 18604 33980
rect 18095 33949 18107 33952
rect 18049 33943 18107 33949
rect 9582 33912 9588 33924
rect 8496 33884 9588 33912
rect 9582 33872 9588 33884
rect 9640 33912 9646 33924
rect 10410 33912 10416 33924
rect 9640 33884 10416 33912
rect 9640 33872 9646 33884
rect 10410 33872 10416 33884
rect 10468 33872 10474 33924
rect 11088 33915 11146 33921
rect 11088 33881 11100 33915
rect 11134 33912 11146 33915
rect 11238 33912 11244 33924
rect 11134 33884 11244 33912
rect 11134 33881 11146 33884
rect 11088 33875 11146 33881
rect 11238 33872 11244 33884
rect 11296 33872 11302 33924
rect 11422 33872 11428 33924
rect 11480 33912 11486 33924
rect 13998 33912 14004 33924
rect 11480 33884 14004 33912
rect 11480 33872 11486 33884
rect 13998 33872 14004 33884
rect 14056 33872 14062 33924
rect 14366 33921 14372 33924
rect 14360 33912 14372 33921
rect 14327 33884 14372 33912
rect 14360 33875 14372 33884
rect 14366 33872 14372 33875
rect 14424 33872 14430 33924
rect 14550 33872 14556 33924
rect 14608 33872 14614 33924
rect 17880 33912 17908 33943
rect 18598 33940 18604 33952
rect 18656 33940 18662 33992
rect 18693 33983 18751 33989
rect 18693 33949 18705 33983
rect 18739 33980 18751 33983
rect 19426 33980 19432 33992
rect 18739 33952 19432 33980
rect 18739 33949 18751 33952
rect 18693 33943 18751 33949
rect 19426 33940 19432 33952
rect 19484 33980 19490 33992
rect 19610 33980 19616 33992
rect 19484 33952 19616 33980
rect 19484 33940 19490 33952
rect 19610 33940 19616 33952
rect 19668 33940 19674 33992
rect 19794 33940 19800 33992
rect 19852 33980 19858 33992
rect 20088 33980 20116 34011
rect 20162 34008 20168 34060
rect 20220 34048 20226 34060
rect 20220 34020 22416 34048
rect 20220 34008 20226 34020
rect 20346 33980 20352 33992
rect 19852 33952 20352 33980
rect 19852 33940 19858 33952
rect 20346 33940 20352 33952
rect 20404 33940 20410 33992
rect 20806 33980 20812 33992
rect 20640 33952 20812 33980
rect 18230 33912 18236 33924
rect 17880 33884 18236 33912
rect 18230 33872 18236 33884
rect 18288 33872 18294 33924
rect 5166 33844 5172 33856
rect 3620 33816 5172 33844
rect 5166 33804 5172 33816
rect 5224 33804 5230 33856
rect 7282 33804 7288 33856
rect 7340 33844 7346 33856
rect 7653 33847 7711 33853
rect 7653 33844 7665 33847
rect 7340 33816 7665 33844
rect 7340 33804 7346 33816
rect 7653 33813 7665 33816
rect 7699 33813 7711 33847
rect 7653 33807 7711 33813
rect 8110 33804 8116 33856
rect 8168 33844 8174 33856
rect 9030 33844 9036 33856
rect 8168 33816 9036 33844
rect 8168 33804 8174 33816
rect 9030 33804 9036 33816
rect 9088 33804 9094 33856
rect 9490 33844 9496 33856
rect 9451 33816 9496 33844
rect 9490 33804 9496 33816
rect 9548 33804 9554 33856
rect 9953 33847 10011 33853
rect 9953 33813 9965 33847
rect 9999 33844 10011 33847
rect 10318 33844 10324 33856
rect 9999 33816 10324 33844
rect 9999 33813 10011 33816
rect 9953 33807 10011 33813
rect 10318 33804 10324 33816
rect 10376 33804 10382 33856
rect 10778 33804 10784 33856
rect 10836 33844 10842 33856
rect 15378 33844 15384 33856
rect 10836 33816 15384 33844
rect 10836 33804 10842 33816
rect 15378 33804 15384 33816
rect 15436 33804 15442 33856
rect 19058 33804 19064 33856
rect 19116 33844 19122 33856
rect 19521 33847 19579 33853
rect 19521 33844 19533 33847
rect 19116 33816 19533 33844
rect 19116 33804 19122 33816
rect 19521 33813 19533 33816
rect 19567 33813 19579 33847
rect 19521 33807 19579 33813
rect 19889 33847 19947 33853
rect 19889 33813 19901 33847
rect 19935 33844 19947 33847
rect 20070 33844 20076 33856
rect 19935 33816 20076 33844
rect 19935 33813 19947 33816
rect 19889 33807 19947 33813
rect 20070 33804 20076 33816
rect 20128 33804 20134 33856
rect 20640 33844 20668 33952
rect 20806 33940 20812 33952
rect 20864 33940 20870 33992
rect 20990 33940 20996 33992
rect 21048 33980 21054 33992
rect 21269 33983 21327 33989
rect 21269 33980 21281 33983
rect 21048 33952 21281 33980
rect 21048 33940 21054 33952
rect 21269 33949 21281 33952
rect 21315 33949 21327 33983
rect 21726 33980 21732 33992
rect 21687 33952 21732 33980
rect 21269 33943 21327 33949
rect 20714 33872 20720 33924
rect 20772 33912 20778 33924
rect 20901 33915 20959 33921
rect 20901 33912 20913 33915
rect 20772 33884 20913 33912
rect 20772 33872 20778 33884
rect 20901 33881 20913 33884
rect 20947 33881 20959 33915
rect 21284 33912 21312 33943
rect 21726 33940 21732 33952
rect 21784 33940 21790 33992
rect 22388 33989 22416 34020
rect 22373 33983 22431 33989
rect 22373 33949 22385 33983
rect 22419 33949 22431 33983
rect 22373 33943 22431 33949
rect 21821 33915 21879 33921
rect 21821 33912 21833 33915
rect 21284 33884 21833 33912
rect 20901 33875 20959 33881
rect 21821 33881 21833 33884
rect 21867 33881 21879 33915
rect 21821 33875 21879 33881
rect 20993 33847 21051 33853
rect 20993 33844 21005 33847
rect 20640 33816 21005 33844
rect 20993 33813 21005 33816
rect 21039 33813 21051 33847
rect 20993 33807 21051 33813
rect 21085 33847 21143 33853
rect 21085 33813 21097 33847
rect 21131 33844 21143 33847
rect 21174 33844 21180 33856
rect 21131 33816 21180 33844
rect 21131 33813 21143 33816
rect 21085 33807 21143 33813
rect 21174 33804 21180 33816
rect 21232 33804 21238 33856
rect 22370 33804 22376 33856
rect 22428 33844 22434 33856
rect 22557 33847 22615 33853
rect 22557 33844 22569 33847
rect 22428 33816 22569 33844
rect 22428 33804 22434 33816
rect 22557 33813 22569 33816
rect 22603 33813 22615 33847
rect 22557 33807 22615 33813
rect 1104 33754 30820 33776
rect 1104 33702 10880 33754
rect 10932 33702 10944 33754
rect 10996 33702 11008 33754
rect 11060 33702 11072 33754
rect 11124 33702 11136 33754
rect 11188 33702 20811 33754
rect 20863 33702 20875 33754
rect 20927 33702 20939 33754
rect 20991 33702 21003 33754
rect 21055 33702 21067 33754
rect 21119 33702 30820 33754
rect 1104 33680 30820 33702
rect 2593 33643 2651 33649
rect 2593 33609 2605 33643
rect 2639 33640 2651 33643
rect 3786 33640 3792 33652
rect 2639 33612 3792 33640
rect 2639 33609 2651 33612
rect 2593 33603 2651 33609
rect 3786 33600 3792 33612
rect 3844 33600 3850 33652
rect 5534 33640 5540 33652
rect 5495 33612 5540 33640
rect 5534 33600 5540 33612
rect 5592 33600 5598 33652
rect 8386 33600 8392 33652
rect 8444 33640 8450 33652
rect 10965 33643 11023 33649
rect 8444 33612 10916 33640
rect 8444 33600 8450 33612
rect 2866 33572 2872 33584
rect 1688 33544 2872 33572
rect 1688 33513 1716 33544
rect 2866 33532 2872 33544
rect 2924 33532 2930 33584
rect 5166 33572 5172 33584
rect 3988 33544 5172 33572
rect 1673 33507 1731 33513
rect 1673 33473 1685 33507
rect 1719 33473 1731 33507
rect 1673 33467 1731 33473
rect 2409 33507 2467 33513
rect 2409 33473 2421 33507
rect 2455 33504 2467 33507
rect 3234 33504 3240 33516
rect 2455 33476 2774 33504
rect 3195 33476 3240 33504
rect 2455 33473 2467 33476
rect 2409 33467 2467 33473
rect 2746 33368 2774 33476
rect 3234 33464 3240 33476
rect 3292 33464 3298 33516
rect 3789 33507 3847 33513
rect 3789 33473 3801 33507
rect 3835 33504 3847 33507
rect 3878 33504 3884 33516
rect 3835 33476 3884 33504
rect 3835 33473 3847 33476
rect 3789 33467 3847 33473
rect 3878 33464 3884 33476
rect 3936 33464 3942 33516
rect 3988 33513 4016 33544
rect 5166 33532 5172 33544
rect 5224 33532 5230 33584
rect 7006 33572 7012 33584
rect 6472 33544 7012 33572
rect 3973 33507 4031 33513
rect 3973 33473 3985 33507
rect 4019 33473 4031 33507
rect 4338 33504 4344 33516
rect 4299 33476 4344 33504
rect 3973 33467 4031 33473
rect 4338 33464 4344 33476
rect 4396 33464 4402 33516
rect 4522 33504 4528 33516
rect 4483 33476 4528 33504
rect 4522 33464 4528 33476
rect 4580 33464 4586 33516
rect 5721 33507 5779 33513
rect 5721 33473 5733 33507
rect 5767 33504 5779 33507
rect 6270 33504 6276 33516
rect 5767 33476 6276 33504
rect 5767 33473 5779 33476
rect 5721 33467 5779 33473
rect 6270 33464 6276 33476
rect 6328 33464 6334 33516
rect 6472 33513 6500 33544
rect 7006 33532 7012 33544
rect 7064 33572 7070 33584
rect 7650 33572 7656 33584
rect 7064 33544 7656 33572
rect 7064 33532 7070 33544
rect 7300 33513 7328 33544
rect 7650 33532 7656 33544
rect 7708 33572 7714 33584
rect 9306 33572 9312 33584
rect 7708 33544 9312 33572
rect 7708 33532 7714 33544
rect 9306 33532 9312 33544
rect 9364 33532 9370 33584
rect 9490 33532 9496 33584
rect 9548 33572 9554 33584
rect 10888 33572 10916 33612
rect 10965 33609 10977 33643
rect 11011 33640 11023 33643
rect 11514 33640 11520 33652
rect 11011 33612 11520 33640
rect 11011 33609 11023 33612
rect 10965 33603 11023 33609
rect 11514 33600 11520 33612
rect 11572 33600 11578 33652
rect 12066 33640 12072 33652
rect 12027 33612 12072 33640
rect 12066 33600 12072 33612
rect 12124 33600 12130 33652
rect 15657 33643 15715 33649
rect 15657 33609 15669 33643
rect 15703 33609 15715 33643
rect 15657 33603 15715 33609
rect 18325 33643 18383 33649
rect 18325 33609 18337 33643
rect 18371 33640 18383 33643
rect 18414 33640 18420 33652
rect 18371 33612 18420 33640
rect 18371 33609 18383 33612
rect 18325 33603 18383 33609
rect 11422 33572 11428 33584
rect 9548 33544 10824 33572
rect 10888 33544 11428 33572
rect 9548 33532 9554 33544
rect 6457 33507 6515 33513
rect 6457 33473 6469 33507
rect 6503 33473 6515 33507
rect 6457 33467 6515 33473
rect 7285 33507 7343 33513
rect 7285 33473 7297 33507
rect 7331 33473 7343 33507
rect 7285 33467 7343 33473
rect 8113 33507 8171 33513
rect 8113 33473 8125 33507
rect 8159 33473 8171 33507
rect 8113 33467 8171 33473
rect 3602 33396 3608 33448
rect 3660 33436 3666 33448
rect 4154 33436 4160 33448
rect 3660 33408 4160 33436
rect 3660 33396 3666 33408
rect 4154 33396 4160 33408
rect 4212 33396 4218 33448
rect 4249 33439 4307 33445
rect 4249 33405 4261 33439
rect 4295 33405 4307 33439
rect 4249 33399 4307 33405
rect 3053 33371 3111 33377
rect 3053 33368 3065 33371
rect 2746 33340 3065 33368
rect 3053 33337 3065 33340
rect 3099 33337 3111 33371
rect 3053 33331 3111 33337
rect 3510 33328 3516 33380
rect 3568 33368 3574 33380
rect 4264 33368 4292 33399
rect 4338 33368 4344 33380
rect 3568 33340 4344 33368
rect 3568 33328 3574 33340
rect 4338 33328 4344 33340
rect 4396 33328 4402 33380
rect 8128 33368 8156 33467
rect 8202 33464 8208 33516
rect 8260 33504 8266 33516
rect 8297 33507 8355 33513
rect 8297 33504 8309 33507
rect 8260 33476 8309 33504
rect 8260 33464 8266 33476
rect 8297 33473 8309 33476
rect 8343 33473 8355 33507
rect 8297 33467 8355 33473
rect 8481 33507 8539 33513
rect 8481 33473 8493 33507
rect 8527 33473 8539 33507
rect 8481 33467 8539 33473
rect 8386 33436 8392 33448
rect 8347 33408 8392 33436
rect 8386 33396 8392 33408
rect 8444 33396 8450 33448
rect 8496 33436 8524 33467
rect 8570 33464 8576 33516
rect 8628 33504 8634 33516
rect 8665 33507 8723 33513
rect 8665 33504 8677 33507
rect 8628 33476 8677 33504
rect 8628 33464 8634 33476
rect 8665 33473 8677 33476
rect 8711 33473 8723 33507
rect 9766 33504 9772 33516
rect 9727 33476 9772 33504
rect 8665 33467 8723 33473
rect 9766 33464 9772 33476
rect 9824 33464 9830 33516
rect 9950 33504 9956 33516
rect 9911 33476 9956 33504
rect 9950 33464 9956 33476
rect 10008 33464 10014 33516
rect 10134 33504 10140 33516
rect 10095 33476 10140 33504
rect 10134 33464 10140 33476
rect 10192 33464 10198 33516
rect 10321 33507 10379 33513
rect 10321 33473 10333 33507
rect 10367 33504 10379 33507
rect 10410 33504 10416 33516
rect 10367 33476 10416 33504
rect 10367 33473 10379 33476
rect 10321 33467 10379 33473
rect 10410 33464 10416 33476
rect 10468 33464 10474 33516
rect 10796 33513 10824 33544
rect 11422 33532 11428 33544
rect 11480 33532 11486 33584
rect 11532 33544 12434 33572
rect 11532 33513 11560 33544
rect 10781 33507 10839 33513
rect 10781 33473 10793 33507
rect 10827 33473 10839 33507
rect 10781 33467 10839 33473
rect 11517 33507 11575 33513
rect 11517 33473 11529 33507
rect 11563 33473 11575 33507
rect 11517 33467 11575 33473
rect 11698 33464 11704 33516
rect 11756 33504 11762 33516
rect 11793 33507 11851 33513
rect 11793 33504 11805 33507
rect 11756 33476 11805 33504
rect 11756 33464 11762 33476
rect 11793 33473 11805 33476
rect 11839 33473 11851 33507
rect 11793 33467 11851 33473
rect 11882 33464 11888 33516
rect 11940 33504 11946 33516
rect 11940 33476 11985 33504
rect 11940 33464 11946 33476
rect 12066 33464 12072 33516
rect 12124 33504 12130 33516
rect 12124 33476 12169 33504
rect 12124 33464 12130 33476
rect 8938 33436 8944 33448
rect 8496 33408 8944 33436
rect 8938 33396 8944 33408
rect 8996 33396 9002 33448
rect 10042 33436 10048 33448
rect 10003 33408 10048 33436
rect 10042 33396 10048 33408
rect 10100 33396 10106 33448
rect 12406 33436 12434 33544
rect 13998 33532 14004 33584
rect 14056 33572 14062 33584
rect 14056 33544 14688 33572
rect 14056 33532 14062 33544
rect 14274 33504 14280 33516
rect 14332 33513 14338 33516
rect 14244 33476 14280 33504
rect 14274 33464 14280 33476
rect 14332 33467 14344 33513
rect 14550 33504 14556 33516
rect 14511 33476 14556 33504
rect 14332 33464 14338 33467
rect 14550 33464 14556 33476
rect 14608 33464 14614 33516
rect 12802 33436 12808 33448
rect 12406 33408 12808 33436
rect 12802 33396 12808 33408
rect 12860 33396 12866 33448
rect 8754 33368 8760 33380
rect 8128 33340 8760 33368
rect 8754 33328 8760 33340
rect 8812 33328 8818 33380
rect 14660 33368 14688 33544
rect 15378 33464 15384 33516
rect 15436 33504 15442 33516
rect 15473 33507 15531 33513
rect 15473 33504 15485 33507
rect 15436 33476 15485 33504
rect 15436 33464 15442 33476
rect 15473 33473 15485 33476
rect 15519 33473 15531 33507
rect 15672 33504 15700 33603
rect 18414 33600 18420 33612
rect 18472 33600 18478 33652
rect 18598 33600 18604 33652
rect 18656 33640 18662 33652
rect 18877 33643 18935 33649
rect 18877 33640 18889 33643
rect 18656 33612 18889 33640
rect 18656 33600 18662 33612
rect 18877 33609 18889 33612
rect 18923 33609 18935 33643
rect 18877 33603 18935 33609
rect 19061 33643 19119 33649
rect 19061 33609 19073 33643
rect 19107 33640 19119 33643
rect 19150 33640 19156 33652
rect 19107 33612 19156 33640
rect 19107 33609 19119 33612
rect 19061 33603 19119 33609
rect 19150 33600 19156 33612
rect 19208 33600 19214 33652
rect 21269 33643 21327 33649
rect 21269 33609 21281 33643
rect 21315 33640 21327 33643
rect 21726 33640 21732 33652
rect 21315 33612 21732 33640
rect 21315 33609 21327 33612
rect 21269 33603 21327 33609
rect 21726 33600 21732 33612
rect 21784 33600 21790 33652
rect 19334 33572 19340 33584
rect 18432 33544 19340 33572
rect 16669 33507 16727 33513
rect 16669 33504 16681 33507
rect 15672 33476 16681 33504
rect 15473 33467 15531 33473
rect 16669 33473 16681 33476
rect 16715 33473 16727 33507
rect 18230 33504 18236 33516
rect 18191 33476 18236 33504
rect 16669 33467 16727 33473
rect 18230 33464 18236 33476
rect 18288 33464 18294 33516
rect 18432 33513 18460 33544
rect 19334 33532 19340 33544
rect 19392 33532 19398 33584
rect 19702 33532 19708 33584
rect 19760 33572 19766 33584
rect 20901 33575 20959 33581
rect 20901 33572 20913 33575
rect 19760 33544 20913 33572
rect 19760 33532 19766 33544
rect 20901 33541 20913 33544
rect 20947 33541 20959 33575
rect 20901 33535 20959 33541
rect 18417 33507 18475 33513
rect 18417 33473 18429 33507
rect 18463 33473 18475 33507
rect 19058 33504 19064 33516
rect 19019 33476 19064 33504
rect 18417 33467 18475 33473
rect 19058 33464 19064 33476
rect 19116 33464 19122 33516
rect 19426 33504 19432 33516
rect 19339 33476 19432 33504
rect 19426 33464 19432 33476
rect 19484 33504 19490 33516
rect 19886 33504 19892 33516
rect 19484 33476 19892 33504
rect 19484 33464 19490 33476
rect 19886 33464 19892 33476
rect 19944 33464 19950 33516
rect 20346 33464 20352 33516
rect 20404 33504 20410 33516
rect 22370 33504 22376 33516
rect 20404 33476 20668 33504
rect 22331 33476 22376 33504
rect 20404 33464 20410 33476
rect 19521 33439 19579 33445
rect 19521 33405 19533 33439
rect 19567 33436 19579 33439
rect 20530 33436 20536 33448
rect 19567 33408 20536 33436
rect 19567 33405 19579 33408
rect 19521 33399 19579 33405
rect 20530 33396 20536 33408
rect 20588 33396 20594 33448
rect 20640 33445 20668 33476
rect 22370 33464 22376 33476
rect 22428 33464 22434 33516
rect 30098 33504 30104 33516
rect 30059 33476 30104 33504
rect 30098 33464 30104 33476
rect 30156 33464 30162 33516
rect 20625 33439 20683 33445
rect 20625 33405 20637 33439
rect 20671 33405 20683 33439
rect 20806 33436 20812 33448
rect 20767 33408 20812 33436
rect 20625 33399 20683 33405
rect 20806 33396 20812 33408
rect 20864 33436 20870 33448
rect 21174 33436 21180 33448
rect 20864 33408 21180 33436
rect 20864 33396 20870 33408
rect 21174 33396 21180 33408
rect 21232 33396 21238 33448
rect 21266 33368 21272 33380
rect 14660 33340 21272 33368
rect 21266 33328 21272 33340
rect 21324 33328 21330 33380
rect 1486 33300 1492 33312
rect 1447 33272 1492 33300
rect 1486 33260 1492 33272
rect 1544 33260 1550 33312
rect 6641 33303 6699 33309
rect 6641 33269 6653 33303
rect 6687 33300 6699 33303
rect 6730 33300 6736 33312
rect 6687 33272 6736 33300
rect 6687 33269 6699 33272
rect 6641 33263 6699 33269
rect 6730 33260 6736 33272
rect 6788 33260 6794 33312
rect 7098 33300 7104 33312
rect 7059 33272 7104 33300
rect 7098 33260 7104 33272
rect 7156 33260 7162 33312
rect 7926 33300 7932 33312
rect 7887 33272 7932 33300
rect 7926 33260 7932 33272
rect 7984 33260 7990 33312
rect 9585 33303 9643 33309
rect 9585 33269 9597 33303
rect 9631 33300 9643 33303
rect 10686 33300 10692 33312
rect 9631 33272 10692 33300
rect 9631 33269 9643 33272
rect 9585 33263 9643 33269
rect 10686 33260 10692 33272
rect 10744 33260 10750 33312
rect 11330 33260 11336 33312
rect 11388 33300 11394 33312
rect 11609 33303 11667 33309
rect 11609 33300 11621 33303
rect 11388 33272 11621 33300
rect 11388 33260 11394 33272
rect 11609 33269 11621 33272
rect 11655 33269 11667 33303
rect 11609 33263 11667 33269
rect 13173 33303 13231 33309
rect 13173 33269 13185 33303
rect 13219 33300 13231 33303
rect 13814 33300 13820 33312
rect 13219 33272 13820 33300
rect 13219 33269 13231 33272
rect 13173 33263 13231 33269
rect 13814 33260 13820 33272
rect 13872 33300 13878 33312
rect 14366 33300 14372 33312
rect 13872 33272 14372 33300
rect 13872 33260 13878 33272
rect 14366 33260 14372 33272
rect 14424 33260 14430 33312
rect 16850 33300 16856 33312
rect 16811 33272 16856 33300
rect 16850 33260 16856 33272
rect 16908 33260 16914 33312
rect 16942 33260 16948 33312
rect 17000 33300 17006 33312
rect 21818 33300 21824 33312
rect 17000 33272 21824 33300
rect 17000 33260 17006 33272
rect 21818 33260 21824 33272
rect 21876 33260 21882 33312
rect 22554 33300 22560 33312
rect 22515 33272 22560 33300
rect 22554 33260 22560 33272
rect 22612 33260 22618 33312
rect 29914 33300 29920 33312
rect 29875 33272 29920 33300
rect 29914 33260 29920 33272
rect 29972 33260 29978 33312
rect 1104 33210 30820 33232
rect 1104 33158 5915 33210
rect 5967 33158 5979 33210
rect 6031 33158 6043 33210
rect 6095 33158 6107 33210
rect 6159 33158 6171 33210
rect 6223 33158 15846 33210
rect 15898 33158 15910 33210
rect 15962 33158 15974 33210
rect 16026 33158 16038 33210
rect 16090 33158 16102 33210
rect 16154 33158 25776 33210
rect 25828 33158 25840 33210
rect 25892 33158 25904 33210
rect 25956 33158 25968 33210
rect 26020 33158 26032 33210
rect 26084 33158 30820 33210
rect 1104 33136 30820 33158
rect 4706 33096 4712 33108
rect 4667 33068 4712 33096
rect 4706 33056 4712 33068
rect 4764 33056 4770 33108
rect 5644 33068 8248 33096
rect 4614 32988 4620 33040
rect 4672 33028 4678 33040
rect 5644 33028 5672 33068
rect 4672 33000 5672 33028
rect 5721 33031 5779 33037
rect 4672 32988 4678 33000
rect 5721 32997 5733 33031
rect 5767 33028 5779 33031
rect 6362 33028 6368 33040
rect 5767 33000 6368 33028
rect 5767 32997 5779 33000
rect 5721 32991 5779 32997
rect 6362 32988 6368 33000
rect 6420 32988 6426 33040
rect 8220 33028 8248 33068
rect 8294 33056 8300 33108
rect 8352 33096 8358 33108
rect 8389 33099 8447 33105
rect 8389 33096 8401 33099
rect 8352 33068 8401 33096
rect 8352 33056 8358 33068
rect 8389 33065 8401 33068
rect 8435 33065 8447 33099
rect 10042 33096 10048 33108
rect 8389 33059 8447 33065
rect 9646 33068 10048 33096
rect 9646 33028 9674 33068
rect 10042 33056 10048 33068
rect 10100 33056 10106 33108
rect 10505 33099 10563 33105
rect 10505 33065 10517 33099
rect 10551 33096 10563 33099
rect 11238 33096 11244 33108
rect 10551 33068 11244 33096
rect 10551 33065 10563 33068
rect 10505 33059 10563 33065
rect 11238 33056 11244 33068
rect 11296 33056 11302 33108
rect 15378 33096 15384 33108
rect 15120 33068 15384 33096
rect 8220 33000 9674 33028
rect 9950 32988 9956 33040
rect 10008 33028 10014 33040
rect 10008 33000 10180 33028
rect 10008 32988 10014 33000
rect 6822 32960 6828 32972
rect 4080 32932 6828 32960
rect 4080 32904 4108 32932
rect 6822 32920 6828 32932
rect 6880 32920 6886 32972
rect 9674 32920 9680 32972
rect 9732 32960 9738 32972
rect 10152 32969 10180 33000
rect 15120 32969 15148 33068
rect 15378 33056 15384 33068
rect 15436 33056 15442 33108
rect 15470 33056 15476 33108
rect 15528 33096 15534 33108
rect 16485 33099 16543 33105
rect 16485 33096 16497 33099
rect 15528 33068 16497 33096
rect 15528 33056 15534 33068
rect 16485 33065 16497 33068
rect 16531 33065 16543 33099
rect 16485 33059 16543 33065
rect 19610 33056 19616 33108
rect 19668 33096 19674 33108
rect 20346 33096 20352 33108
rect 19668 33068 20352 33096
rect 19668 33056 19674 33068
rect 20346 33056 20352 33068
rect 20404 33056 20410 33108
rect 20714 33096 20720 33108
rect 20675 33068 20720 33096
rect 20714 33056 20720 33068
rect 20772 33056 20778 33108
rect 10045 32963 10103 32969
rect 10045 32960 10057 32963
rect 9732 32932 10057 32960
rect 9732 32920 9738 32932
rect 10045 32929 10057 32932
rect 10091 32929 10103 32963
rect 10045 32923 10103 32929
rect 10137 32963 10195 32969
rect 10137 32929 10149 32963
rect 10183 32929 10195 32963
rect 10137 32923 10195 32929
rect 15105 32963 15163 32969
rect 15105 32929 15117 32963
rect 15151 32929 15163 32963
rect 15105 32923 15163 32929
rect 16850 32920 16856 32972
rect 16908 32960 16914 32972
rect 17037 32963 17095 32969
rect 17037 32960 17049 32963
rect 16908 32932 17049 32960
rect 16908 32920 16914 32932
rect 17037 32929 17049 32932
rect 17083 32929 17095 32963
rect 20438 32960 20444 32972
rect 20399 32932 20444 32960
rect 17037 32923 17095 32929
rect 20438 32920 20444 32932
rect 20496 32920 20502 32972
rect 1394 32892 1400 32904
rect 1355 32864 1400 32892
rect 1394 32852 1400 32864
rect 1452 32852 1458 32904
rect 2314 32892 2320 32904
rect 2275 32864 2320 32892
rect 2314 32852 2320 32864
rect 2372 32852 2378 32904
rect 3145 32895 3203 32901
rect 3145 32861 3157 32895
rect 3191 32892 3203 32895
rect 3234 32892 3240 32904
rect 3191 32864 3240 32892
rect 3191 32861 3203 32864
rect 3145 32855 3203 32861
rect 3234 32852 3240 32864
rect 3292 32852 3298 32904
rect 4062 32892 4068 32904
rect 3975 32864 4068 32892
rect 4062 32852 4068 32864
rect 4120 32852 4126 32904
rect 4890 32892 4896 32904
rect 4851 32864 4896 32892
rect 4890 32852 4896 32864
rect 4948 32852 4954 32904
rect 6365 32895 6423 32901
rect 6365 32861 6377 32895
rect 6411 32861 6423 32895
rect 6365 32855 6423 32861
rect 5537 32827 5595 32833
rect 5537 32793 5549 32827
rect 5583 32824 5595 32827
rect 5718 32824 5724 32836
rect 5583 32796 5724 32824
rect 5583 32793 5595 32796
rect 5537 32787 5595 32793
rect 5718 32784 5724 32796
rect 5776 32784 5782 32836
rect 6380 32824 6408 32855
rect 6914 32852 6920 32904
rect 6972 32892 6978 32904
rect 7282 32901 7288 32904
rect 7009 32895 7067 32901
rect 7009 32892 7021 32895
rect 6972 32864 7021 32892
rect 6972 32852 6978 32864
rect 7009 32861 7021 32864
rect 7055 32861 7067 32895
rect 7276 32892 7288 32901
rect 7243 32864 7288 32892
rect 7009 32855 7067 32861
rect 7276 32855 7288 32864
rect 7282 32852 7288 32855
rect 7340 32852 7346 32904
rect 9033 32895 9091 32901
rect 9033 32861 9045 32895
rect 9079 32892 9091 32895
rect 9306 32892 9312 32904
rect 9079 32864 9312 32892
rect 9079 32861 9091 32864
rect 9033 32855 9091 32861
rect 9306 32852 9312 32864
rect 9364 32852 9370 32904
rect 9582 32852 9588 32904
rect 9640 32892 9646 32904
rect 9769 32895 9827 32901
rect 9769 32892 9781 32895
rect 9640 32864 9781 32892
rect 9640 32852 9646 32864
rect 9769 32861 9781 32864
rect 9815 32861 9827 32895
rect 9950 32892 9956 32904
rect 9911 32864 9956 32892
rect 9769 32855 9827 32861
rect 9950 32852 9956 32864
rect 10008 32852 10014 32904
rect 10318 32892 10324 32904
rect 10279 32864 10324 32892
rect 10318 32852 10324 32864
rect 10376 32852 10382 32904
rect 11149 32895 11207 32901
rect 11149 32861 11161 32895
rect 11195 32861 11207 32895
rect 11606 32892 11612 32904
rect 11567 32864 11612 32892
rect 11149 32855 11207 32861
rect 7098 32824 7104 32836
rect 6380 32796 7104 32824
rect 7098 32784 7104 32796
rect 7156 32784 7162 32836
rect 11164 32824 11192 32855
rect 11606 32852 11612 32864
rect 11664 32852 11670 32904
rect 18874 32852 18880 32904
rect 18932 32892 18938 32904
rect 19705 32895 19763 32901
rect 19705 32892 19717 32895
rect 18932 32864 19717 32892
rect 18932 32852 18938 32864
rect 19705 32861 19717 32864
rect 19751 32892 19763 32895
rect 19794 32892 19800 32904
rect 19751 32864 19800 32892
rect 19751 32861 19763 32864
rect 19705 32855 19763 32861
rect 19794 32852 19800 32864
rect 19852 32852 19858 32904
rect 20349 32895 20407 32901
rect 20349 32892 20361 32895
rect 19904 32864 20361 32892
rect 9232 32796 11192 32824
rect 11876 32827 11934 32833
rect 1578 32756 1584 32768
rect 1539 32728 1584 32756
rect 1578 32716 1584 32728
rect 1636 32716 1642 32768
rect 2130 32756 2136 32768
rect 2091 32728 2136 32756
rect 2130 32716 2136 32728
rect 2188 32716 2194 32768
rect 2590 32716 2596 32768
rect 2648 32756 2654 32768
rect 2961 32759 3019 32765
rect 2961 32756 2973 32759
rect 2648 32728 2973 32756
rect 2648 32716 2654 32728
rect 2961 32725 2973 32728
rect 3007 32725 3019 32759
rect 4246 32756 4252 32768
rect 4207 32728 4252 32756
rect 2961 32719 3019 32725
rect 4246 32716 4252 32728
rect 4304 32716 4310 32768
rect 6549 32759 6607 32765
rect 6549 32725 6561 32759
rect 6595 32756 6607 32759
rect 7374 32756 7380 32768
rect 6595 32728 7380 32756
rect 6595 32725 6607 32728
rect 6549 32719 6607 32725
rect 7374 32716 7380 32728
rect 7432 32716 7438 32768
rect 9232 32765 9260 32796
rect 11876 32793 11888 32827
rect 11922 32824 11934 32827
rect 11974 32824 11980 32836
rect 11922 32796 11980 32824
rect 11922 32793 11934 32796
rect 11876 32787 11934 32793
rect 11974 32784 11980 32796
rect 12032 32784 12038 32836
rect 15372 32827 15430 32833
rect 15372 32793 15384 32827
rect 15418 32824 15430 32827
rect 15746 32824 15752 32836
rect 15418 32796 15752 32824
rect 15418 32793 15430 32796
rect 15372 32787 15430 32793
rect 15746 32784 15752 32796
rect 15804 32784 15810 32836
rect 17304 32827 17362 32833
rect 17304 32793 17316 32827
rect 17350 32824 17362 32827
rect 17954 32824 17960 32836
rect 17350 32796 17960 32824
rect 17350 32793 17362 32796
rect 17304 32787 17362 32793
rect 17954 32784 17960 32796
rect 18012 32784 18018 32836
rect 19904 32768 19932 32864
rect 20349 32861 20361 32864
rect 20395 32861 20407 32895
rect 22278 32892 22284 32904
rect 22239 32864 22284 32892
rect 20349 32855 20407 32861
rect 22278 32852 22284 32864
rect 22336 32852 22342 32904
rect 22465 32895 22523 32901
rect 22465 32861 22477 32895
rect 22511 32892 22523 32895
rect 29914 32892 29920 32904
rect 22511 32864 29920 32892
rect 22511 32861 22523 32864
rect 22465 32855 22523 32861
rect 29914 32852 29920 32864
rect 29972 32852 29978 32904
rect 9217 32759 9275 32765
rect 9217 32725 9229 32759
rect 9263 32725 9275 32759
rect 9217 32719 9275 32725
rect 10778 32716 10784 32768
rect 10836 32756 10842 32768
rect 10965 32759 11023 32765
rect 10965 32756 10977 32759
rect 10836 32728 10977 32756
rect 10836 32716 10842 32728
rect 10965 32725 10977 32728
rect 11011 32725 11023 32759
rect 10965 32719 11023 32725
rect 12894 32716 12900 32768
rect 12952 32756 12958 32768
rect 12989 32759 13047 32765
rect 12989 32756 13001 32759
rect 12952 32728 13001 32756
rect 12952 32716 12958 32728
rect 12989 32725 13001 32728
rect 13035 32725 13047 32759
rect 18414 32756 18420 32768
rect 18375 32728 18420 32756
rect 12989 32719 13047 32725
rect 18414 32716 18420 32728
rect 18472 32716 18478 32768
rect 19797 32759 19855 32765
rect 19797 32725 19809 32759
rect 19843 32756 19855 32759
rect 19886 32756 19892 32768
rect 19843 32728 19892 32756
rect 19843 32725 19855 32728
rect 19797 32719 19855 32725
rect 19886 32716 19892 32728
rect 19944 32716 19950 32768
rect 22094 32756 22100 32768
rect 22055 32728 22100 32756
rect 22094 32716 22100 32728
rect 22152 32716 22158 32768
rect 1104 32666 30820 32688
rect 1104 32614 10880 32666
rect 10932 32614 10944 32666
rect 10996 32614 11008 32666
rect 11060 32614 11072 32666
rect 11124 32614 11136 32666
rect 11188 32614 20811 32666
rect 20863 32614 20875 32666
rect 20927 32614 20939 32666
rect 20991 32614 21003 32666
rect 21055 32614 21067 32666
rect 21119 32614 30820 32666
rect 1104 32592 30820 32614
rect 2225 32555 2283 32561
rect 2225 32521 2237 32555
rect 2271 32552 2283 32555
rect 3970 32552 3976 32564
rect 2271 32524 3976 32552
rect 2271 32521 2283 32524
rect 2225 32515 2283 32521
rect 3970 32512 3976 32524
rect 4028 32552 4034 32564
rect 4249 32555 4307 32561
rect 4249 32552 4261 32555
rect 4028 32524 4261 32552
rect 4028 32512 4034 32524
rect 4249 32521 4261 32524
rect 4295 32521 4307 32555
rect 6914 32552 6920 32564
rect 6875 32524 6920 32552
rect 4249 32515 4307 32521
rect 6914 32512 6920 32524
rect 6972 32512 6978 32564
rect 8754 32552 8760 32564
rect 8715 32524 8760 32552
rect 8754 32512 8760 32524
rect 8812 32512 8818 32564
rect 9585 32555 9643 32561
rect 9585 32521 9597 32555
rect 9631 32552 9643 32555
rect 9766 32552 9772 32564
rect 9631 32524 9772 32552
rect 9631 32521 9643 32524
rect 9585 32515 9643 32521
rect 9766 32512 9772 32524
rect 9824 32512 9830 32564
rect 10778 32512 10784 32564
rect 10836 32512 10842 32564
rect 12986 32512 12992 32564
rect 13044 32552 13050 32564
rect 13262 32552 13268 32564
rect 13044 32524 13268 32552
rect 13044 32512 13050 32524
rect 13262 32512 13268 32524
rect 13320 32552 13326 32564
rect 14642 32552 14648 32564
rect 13320 32524 14648 32552
rect 13320 32512 13326 32524
rect 14642 32512 14648 32524
rect 14700 32512 14706 32564
rect 15746 32552 15752 32564
rect 15707 32524 15752 32552
rect 15746 32512 15752 32524
rect 15804 32512 15810 32564
rect 17954 32552 17960 32564
rect 17915 32524 17960 32552
rect 17954 32512 17960 32524
rect 18012 32512 18018 32564
rect 18414 32552 18420 32564
rect 18156 32524 18420 32552
rect 7644 32487 7702 32493
rect 7644 32453 7656 32487
rect 7690 32484 7702 32487
rect 7926 32484 7932 32496
rect 7690 32456 7932 32484
rect 7690 32453 7702 32456
rect 7644 32447 7702 32453
rect 7926 32444 7932 32456
rect 7984 32444 7990 32496
rect 10686 32484 10692 32496
rect 10744 32493 10750 32496
rect 10656 32456 10692 32484
rect 10686 32444 10692 32456
rect 10744 32447 10756 32493
rect 10744 32444 10750 32447
rect 1857 32419 1915 32425
rect 1857 32385 1869 32419
rect 1903 32416 1915 32419
rect 2130 32416 2136 32428
rect 1903 32388 2136 32416
rect 1903 32385 1915 32388
rect 1857 32379 1915 32385
rect 2130 32376 2136 32388
rect 2188 32376 2194 32428
rect 3136 32419 3194 32425
rect 3136 32385 3148 32419
rect 3182 32416 3194 32419
rect 3694 32416 3700 32428
rect 3182 32388 3700 32416
rect 3182 32385 3194 32388
rect 3136 32379 3194 32385
rect 3694 32376 3700 32388
rect 3752 32376 3758 32428
rect 4522 32376 4528 32428
rect 4580 32416 4586 32428
rect 5353 32419 5411 32425
rect 5353 32416 5365 32419
rect 4580 32388 5365 32416
rect 4580 32376 4586 32388
rect 5353 32385 5365 32388
rect 5399 32385 5411 32419
rect 6730 32416 6736 32428
rect 6691 32388 6736 32416
rect 5353 32379 5411 32385
rect 6730 32376 6736 32388
rect 6788 32376 6794 32428
rect 7374 32416 7380 32428
rect 7335 32388 7380 32416
rect 7374 32376 7380 32388
rect 7432 32376 7438 32428
rect 10796 32416 10824 32512
rect 15470 32484 15476 32496
rect 15431 32456 15476 32484
rect 15470 32444 15476 32456
rect 15528 32444 15534 32496
rect 18046 32484 18052 32496
rect 17512 32456 18052 32484
rect 10965 32419 11023 32425
rect 10965 32416 10977 32419
rect 10796 32388 10977 32416
rect 10965 32385 10977 32388
rect 11011 32385 11023 32419
rect 10965 32379 11023 32385
rect 11876 32419 11934 32425
rect 11876 32385 11888 32419
rect 11922 32416 11934 32419
rect 12250 32416 12256 32428
rect 11922 32388 12256 32416
rect 11922 32385 11934 32388
rect 11876 32379 11934 32385
rect 12250 32376 12256 32388
rect 12308 32376 12314 32428
rect 14642 32376 14648 32428
rect 14700 32416 14706 32428
rect 15105 32419 15163 32425
rect 15105 32416 15117 32419
rect 14700 32388 15117 32416
rect 14700 32376 14706 32388
rect 15105 32385 15117 32388
rect 15151 32385 15163 32419
rect 15105 32379 15163 32385
rect 15253 32419 15311 32425
rect 15253 32385 15265 32419
rect 15299 32416 15311 32419
rect 15299 32385 15332 32416
rect 15253 32379 15332 32385
rect 2774 32308 2780 32360
rect 2832 32348 2838 32360
rect 2869 32351 2927 32357
rect 2869 32348 2881 32351
rect 2832 32320 2881 32348
rect 2832 32308 2838 32320
rect 2869 32317 2881 32320
rect 2915 32317 2927 32351
rect 2869 32311 2927 32317
rect 5629 32351 5687 32357
rect 5629 32317 5641 32351
rect 5675 32348 5687 32351
rect 11606 32348 11612 32360
rect 5675 32320 5764 32348
rect 11567 32320 11612 32348
rect 5675 32317 5687 32320
rect 5629 32311 5687 32317
rect 5736 32224 5764 32320
rect 11606 32308 11612 32320
rect 11664 32308 11670 32360
rect 15304 32348 15332 32379
rect 15378 32376 15384 32428
rect 15436 32416 15442 32428
rect 15611 32419 15669 32425
rect 15436 32388 15481 32416
rect 15436 32376 15442 32388
rect 15611 32385 15623 32419
rect 15657 32416 15669 32419
rect 15746 32416 15752 32428
rect 15657 32388 15752 32416
rect 15657 32385 15669 32388
rect 15611 32379 15669 32385
rect 15746 32376 15752 32388
rect 15804 32376 15810 32428
rect 16574 32376 16580 32428
rect 16632 32416 16638 32428
rect 17218 32416 17224 32428
rect 16632 32388 17224 32416
rect 16632 32376 16638 32388
rect 17218 32376 17224 32388
rect 17276 32376 17282 32428
rect 17512 32425 17540 32456
rect 18046 32444 18052 32456
rect 18104 32444 18110 32496
rect 17405 32419 17463 32425
rect 17405 32385 17417 32419
rect 17451 32385 17463 32419
rect 17405 32379 17463 32385
rect 17497 32419 17555 32425
rect 17497 32385 17509 32419
rect 17543 32385 17555 32419
rect 17497 32379 17555 32385
rect 17773 32419 17831 32425
rect 17773 32385 17785 32419
rect 17819 32416 17831 32419
rect 18156 32416 18184 32524
rect 18414 32512 18420 32524
rect 18472 32552 18478 32564
rect 18601 32555 18659 32561
rect 18601 32552 18613 32555
rect 18472 32524 18613 32552
rect 18472 32512 18478 32524
rect 18601 32521 18613 32524
rect 18647 32521 18659 32555
rect 18601 32515 18659 32521
rect 20530 32512 20536 32564
rect 20588 32561 20594 32564
rect 20588 32555 20607 32561
rect 20595 32521 20607 32555
rect 20588 32515 20607 32521
rect 20588 32512 20594 32515
rect 18782 32484 18788 32496
rect 17819 32388 18184 32416
rect 18340 32456 18788 32484
rect 17819 32385 17831 32388
rect 17773 32379 17831 32385
rect 17126 32348 17132 32360
rect 15304 32320 17132 32348
rect 17126 32308 17132 32320
rect 17184 32308 17190 32360
rect 17420 32292 17448 32379
rect 17589 32351 17647 32357
rect 17589 32317 17601 32351
rect 17635 32348 17647 32351
rect 17862 32348 17868 32360
rect 17635 32320 17868 32348
rect 17635 32317 17647 32320
rect 17589 32311 17647 32317
rect 17862 32308 17868 32320
rect 17920 32308 17926 32360
rect 18046 32308 18052 32360
rect 18104 32348 18110 32360
rect 18340 32348 18368 32456
rect 18782 32444 18788 32456
rect 18840 32484 18846 32496
rect 20346 32484 20352 32496
rect 18840 32456 19656 32484
rect 20307 32456 20352 32484
rect 18840 32444 18846 32456
rect 18509 32419 18567 32425
rect 18509 32385 18521 32419
rect 18555 32416 18567 32419
rect 18874 32416 18880 32428
rect 18555 32388 18880 32416
rect 18555 32385 18567 32388
rect 18509 32379 18567 32385
rect 18874 32376 18880 32388
rect 18932 32376 18938 32428
rect 19628 32425 19656 32456
rect 20346 32444 20352 32456
rect 20404 32444 20410 32496
rect 19613 32419 19671 32425
rect 19613 32385 19625 32419
rect 19659 32385 19671 32419
rect 19613 32379 19671 32385
rect 19794 32376 19800 32428
rect 19852 32416 19858 32428
rect 19978 32416 19984 32428
rect 19852 32388 19984 32416
rect 19852 32376 19858 32388
rect 19978 32376 19984 32388
rect 20036 32416 20042 32428
rect 20622 32416 20628 32428
rect 20036 32388 20628 32416
rect 20036 32376 20042 32388
rect 20622 32376 20628 32388
rect 20680 32376 20686 32428
rect 18104 32320 18368 32348
rect 18693 32351 18751 32357
rect 18104 32308 18110 32320
rect 18693 32317 18705 32351
rect 18739 32348 18751 32351
rect 29822 32348 29828 32360
rect 18739 32320 29828 32348
rect 18739 32317 18751 32320
rect 18693 32311 18751 32317
rect 14182 32280 14188 32292
rect 13004 32252 14188 32280
rect 2222 32212 2228 32224
rect 2183 32184 2228 32212
rect 2222 32172 2228 32184
rect 2280 32172 2286 32224
rect 2409 32215 2467 32221
rect 2409 32181 2421 32215
rect 2455 32212 2467 32215
rect 3050 32212 3056 32224
rect 2455 32184 3056 32212
rect 2455 32181 2467 32184
rect 2409 32175 2467 32181
rect 3050 32172 3056 32184
rect 3108 32172 3114 32224
rect 5718 32172 5724 32224
rect 5776 32212 5782 32224
rect 10042 32212 10048 32224
rect 5776 32184 10048 32212
rect 5776 32172 5782 32184
rect 10042 32172 10048 32184
rect 10100 32172 10106 32224
rect 12710 32172 12716 32224
rect 12768 32212 12774 32224
rect 13004 32221 13032 32252
rect 14182 32240 14188 32252
rect 14240 32240 14246 32292
rect 17402 32280 17408 32292
rect 17315 32252 17408 32280
rect 17402 32240 17408 32252
rect 17460 32280 17466 32292
rect 18708 32280 18736 32311
rect 29822 32308 29828 32320
rect 29880 32308 29886 32360
rect 20254 32280 20260 32292
rect 17460 32252 18736 32280
rect 18800 32252 20260 32280
rect 17460 32240 17466 32252
rect 12989 32215 13047 32221
rect 12989 32212 13001 32215
rect 12768 32184 13001 32212
rect 12768 32172 12774 32184
rect 12989 32181 13001 32184
rect 13035 32181 13047 32215
rect 12989 32175 13047 32181
rect 13814 32172 13820 32224
rect 13872 32212 13878 32224
rect 15102 32212 15108 32224
rect 13872 32184 15108 32212
rect 13872 32172 13878 32184
rect 15102 32172 15108 32184
rect 15160 32172 15166 32224
rect 17862 32172 17868 32224
rect 17920 32212 17926 32224
rect 18800 32212 18828 32252
rect 20254 32240 20260 32252
rect 20312 32240 20318 32292
rect 19058 32212 19064 32224
rect 17920 32184 18828 32212
rect 19019 32184 19064 32212
rect 17920 32172 17926 32184
rect 19058 32172 19064 32184
rect 19116 32172 19122 32224
rect 19610 32212 19616 32224
rect 19571 32184 19616 32212
rect 19610 32172 19616 32184
rect 19668 32172 19674 32224
rect 20533 32215 20591 32221
rect 20533 32181 20545 32215
rect 20579 32212 20591 32215
rect 20622 32212 20628 32224
rect 20579 32184 20628 32212
rect 20579 32181 20591 32184
rect 20533 32175 20591 32181
rect 20622 32172 20628 32184
rect 20680 32172 20686 32224
rect 20717 32215 20775 32221
rect 20717 32181 20729 32215
rect 20763 32212 20775 32215
rect 21634 32212 21640 32224
rect 20763 32184 21640 32212
rect 20763 32181 20775 32184
rect 20717 32175 20775 32181
rect 21634 32172 21640 32184
rect 21692 32172 21698 32224
rect 1104 32122 30820 32144
rect 1104 32070 5915 32122
rect 5967 32070 5979 32122
rect 6031 32070 6043 32122
rect 6095 32070 6107 32122
rect 6159 32070 6171 32122
rect 6223 32070 15846 32122
rect 15898 32070 15910 32122
rect 15962 32070 15974 32122
rect 16026 32070 16038 32122
rect 16090 32070 16102 32122
rect 16154 32070 25776 32122
rect 25828 32070 25840 32122
rect 25892 32070 25904 32122
rect 25956 32070 25968 32122
rect 26020 32070 26032 32122
rect 26084 32070 30820 32122
rect 1104 32048 30820 32070
rect 2774 31968 2780 32020
rect 2832 32008 2838 32020
rect 2832 31980 2877 32008
rect 2832 31968 2838 31980
rect 3694 31968 3700 32020
rect 3752 32008 3758 32020
rect 3789 32011 3847 32017
rect 3789 32008 3801 32011
rect 3752 31980 3801 32008
rect 3752 31968 3758 31980
rect 3789 31977 3801 31980
rect 3835 31977 3847 32011
rect 3789 31971 3847 31977
rect 4246 31968 4252 32020
rect 4304 32008 4310 32020
rect 9769 32011 9827 32017
rect 4304 31980 7696 32008
rect 4304 31968 4310 31980
rect 7101 31943 7159 31949
rect 7101 31909 7113 31943
rect 7147 31909 7159 31943
rect 7101 31903 7159 31909
rect 3050 31872 3056 31884
rect 1688 31844 3056 31872
rect 1688 31813 1716 31844
rect 3050 31832 3056 31844
rect 3108 31832 3114 31884
rect 4154 31872 4160 31884
rect 4115 31844 4160 31872
rect 4154 31832 4160 31844
rect 4212 31872 4218 31884
rect 5537 31875 5595 31881
rect 5537 31872 5549 31875
rect 4212 31844 5549 31872
rect 4212 31832 4218 31844
rect 5537 31841 5549 31844
rect 5583 31841 5595 31875
rect 5537 31835 5595 31841
rect 1673 31807 1731 31813
rect 1673 31773 1685 31807
rect 1719 31773 1731 31807
rect 2590 31804 2596 31816
rect 2551 31776 2596 31804
rect 1673 31767 1731 31773
rect 2590 31764 2596 31776
rect 2648 31764 2654 31816
rect 3970 31804 3976 31816
rect 3931 31776 3976 31804
rect 3970 31764 3976 31776
rect 4028 31764 4034 31816
rect 4246 31804 4252 31816
rect 4207 31776 4252 31804
rect 4246 31764 4252 31776
rect 4304 31764 4310 31816
rect 4341 31807 4399 31813
rect 4341 31773 4353 31807
rect 4387 31804 4399 31807
rect 4522 31804 4528 31816
rect 4387 31776 4421 31804
rect 4483 31776 4528 31804
rect 4387 31773 4399 31776
rect 4341 31767 4399 31773
rect 4356 31736 4384 31767
rect 4522 31764 4528 31776
rect 4580 31764 4586 31816
rect 4614 31764 4620 31816
rect 4672 31764 4678 31816
rect 5813 31807 5871 31813
rect 5813 31773 5825 31807
rect 5859 31804 5871 31807
rect 6454 31804 6460 31816
rect 5859 31776 6460 31804
rect 5859 31773 5871 31776
rect 5813 31767 5871 31773
rect 6454 31764 6460 31776
rect 6512 31764 6518 31816
rect 6822 31764 6828 31816
rect 6880 31804 6886 31816
rect 6917 31807 6975 31813
rect 6917 31804 6929 31807
rect 6880 31776 6929 31804
rect 6880 31764 6886 31776
rect 6917 31773 6929 31776
rect 6963 31773 6975 31807
rect 7116 31804 7144 31903
rect 7561 31807 7619 31813
rect 7561 31804 7573 31807
rect 7116 31776 7573 31804
rect 6917 31767 6975 31773
rect 7561 31773 7573 31776
rect 7607 31773 7619 31807
rect 7668 31804 7696 31980
rect 9769 31977 9781 32011
rect 9815 32008 9827 32011
rect 9858 32008 9864 32020
rect 9815 31980 9864 32008
rect 9815 31977 9827 31980
rect 9769 31971 9827 31977
rect 9858 31968 9864 31980
rect 9916 31968 9922 32020
rect 14458 32008 14464 32020
rect 10520 31980 12434 32008
rect 8389 31943 8447 31949
rect 8389 31909 8401 31943
rect 8435 31940 8447 31943
rect 10520 31940 10548 31980
rect 8435 31912 10548 31940
rect 10597 31943 10655 31949
rect 8435 31909 8447 31912
rect 8389 31903 8447 31909
rect 10597 31909 10609 31943
rect 10643 31909 10655 31943
rect 12406 31940 12434 31980
rect 14108 31980 14464 32008
rect 12406 31912 13952 31940
rect 10597 31903 10655 31909
rect 9401 31875 9459 31881
rect 9401 31841 9413 31875
rect 9447 31872 9459 31875
rect 9674 31872 9680 31884
rect 9447 31844 9680 31872
rect 9447 31841 9459 31844
rect 9401 31835 9459 31841
rect 9674 31832 9680 31844
rect 9732 31832 9738 31884
rect 10226 31832 10232 31884
rect 10284 31872 10290 31884
rect 10612 31872 10640 31903
rect 11238 31872 11244 31884
rect 10284 31844 10640 31872
rect 11151 31844 11244 31872
rect 10284 31832 10290 31844
rect 11238 31832 11244 31844
rect 11296 31872 11302 31884
rect 13722 31872 13728 31884
rect 11296 31844 13728 31872
rect 11296 31832 11302 31844
rect 13722 31832 13728 31844
rect 13780 31832 13786 31884
rect 13814 31832 13820 31884
rect 13872 31832 13878 31884
rect 8205 31807 8263 31813
rect 8205 31804 8217 31807
rect 7668 31776 8217 31804
rect 7561 31767 7619 31773
rect 8205 31773 8217 31776
rect 8251 31773 8263 31807
rect 8205 31767 8263 31773
rect 9766 31764 9772 31816
rect 9824 31804 9830 31816
rect 9861 31807 9919 31813
rect 9861 31804 9873 31807
rect 9824 31776 9873 31804
rect 9824 31764 9830 31776
rect 9861 31773 9873 31776
rect 9907 31773 9919 31807
rect 9861 31767 9919 31773
rect 10042 31764 10048 31816
rect 10100 31804 10106 31816
rect 10413 31807 10471 31813
rect 10413 31804 10425 31807
rect 10100 31776 10425 31804
rect 10100 31764 10106 31776
rect 10413 31773 10425 31776
rect 10459 31804 10471 31807
rect 10502 31804 10508 31816
rect 10459 31776 10508 31804
rect 10459 31773 10471 31776
rect 10413 31767 10471 31773
rect 10502 31764 10508 31776
rect 10560 31764 10566 31816
rect 11514 31804 11520 31816
rect 11475 31776 11520 31804
rect 11514 31764 11520 31776
rect 11572 31804 11578 31816
rect 12066 31804 12072 31816
rect 11572 31776 12072 31804
rect 11572 31764 11578 31776
rect 12066 31764 12072 31776
rect 12124 31764 12130 31816
rect 13832 31804 13860 31832
rect 13740 31776 13860 31804
rect 13924 31804 13952 31912
rect 14108 31884 14136 31980
rect 14458 31968 14464 31980
rect 14516 31968 14522 32020
rect 15746 31968 15752 32020
rect 15804 32008 15810 32020
rect 16025 32011 16083 32017
rect 16025 32008 16037 32011
rect 15804 31980 16037 32008
rect 15804 31968 15810 31980
rect 16025 31977 16037 31980
rect 16071 31977 16083 32011
rect 16025 31971 16083 31977
rect 17126 31968 17132 32020
rect 17184 32008 17190 32020
rect 17221 32011 17279 32017
rect 17221 32008 17233 32011
rect 17184 31980 17233 32008
rect 17184 31968 17190 31980
rect 17221 31977 17233 31980
rect 17267 31977 17279 32011
rect 17221 31971 17279 31977
rect 19150 31968 19156 32020
rect 19208 32008 19214 32020
rect 19245 32011 19303 32017
rect 19245 32008 19257 32011
rect 19208 31980 19257 32008
rect 19208 31968 19214 31980
rect 19245 31977 19257 31980
rect 19291 31977 19303 32011
rect 19245 31971 19303 31977
rect 19613 32011 19671 32017
rect 19613 31977 19625 32011
rect 19659 31977 19671 32011
rect 19794 32008 19800 32020
rect 19707 31980 19800 32008
rect 19613 31971 19671 31977
rect 15102 31900 15108 31952
rect 15160 31940 15166 31952
rect 18690 31940 18696 31952
rect 15160 31912 18696 31940
rect 15160 31900 15166 31912
rect 18690 31900 18696 31912
rect 18748 31900 18754 31952
rect 14090 31872 14096 31884
rect 14003 31844 14096 31872
rect 14090 31832 14096 31844
rect 14148 31832 14154 31884
rect 17494 31872 17500 31884
rect 15120 31844 17500 31872
rect 15120 31804 15148 31844
rect 17494 31832 17500 31844
rect 17552 31832 17558 31884
rect 13924 31776 15148 31804
rect 4632 31736 4660 31764
rect 4356 31708 4660 31736
rect 4982 31696 4988 31748
rect 5040 31736 5046 31748
rect 9490 31736 9496 31748
rect 5040 31708 9496 31736
rect 5040 31696 5046 31708
rect 9490 31696 9496 31708
rect 9548 31696 9554 31748
rect 13740 31736 13768 31776
rect 15378 31764 15384 31816
rect 15436 31804 15442 31816
rect 15933 31807 15991 31813
rect 15933 31804 15945 31807
rect 15436 31776 15945 31804
rect 15436 31764 15442 31776
rect 15933 31773 15945 31776
rect 15979 31773 15991 31807
rect 17402 31804 17408 31816
rect 17363 31776 17408 31804
rect 15933 31767 15991 31773
rect 17402 31764 17408 31776
rect 17460 31764 17466 31816
rect 18506 31804 18512 31816
rect 18467 31776 18512 31804
rect 18506 31764 18512 31776
rect 18564 31764 18570 31816
rect 18601 31807 18659 31813
rect 18601 31773 18613 31807
rect 18647 31804 18659 31807
rect 19426 31804 19432 31816
rect 18647 31776 19432 31804
rect 18647 31773 18659 31776
rect 18601 31767 18659 31773
rect 19426 31764 19432 31776
rect 19484 31804 19490 31816
rect 19521 31807 19579 31813
rect 19521 31804 19533 31807
rect 19484 31776 19533 31804
rect 19484 31764 19490 31776
rect 19521 31773 19533 31776
rect 19567 31773 19579 31807
rect 19521 31767 19579 31773
rect 12406 31708 13768 31736
rect 1486 31668 1492 31680
rect 1447 31640 1492 31668
rect 1486 31628 1492 31640
rect 1544 31628 1550 31680
rect 6362 31668 6368 31680
rect 6323 31640 6368 31668
rect 6362 31628 6368 31640
rect 6420 31628 6426 31680
rect 7742 31668 7748 31680
rect 7703 31640 7748 31668
rect 7742 31628 7748 31640
rect 7800 31628 7806 31680
rect 8846 31628 8852 31680
rect 8904 31668 8910 31680
rect 12406 31668 12434 31708
rect 13814 31696 13820 31748
rect 13872 31736 13878 31748
rect 14338 31739 14396 31745
rect 14338 31736 14350 31739
rect 13872 31708 14350 31736
rect 13872 31696 13878 31708
rect 14338 31705 14350 31708
rect 14384 31705 14396 31739
rect 17586 31736 17592 31748
rect 14338 31699 14396 31705
rect 14476 31708 15608 31736
rect 17547 31708 17592 31736
rect 8904 31640 12434 31668
rect 8904 31628 8910 31640
rect 13906 31628 13912 31680
rect 13964 31668 13970 31680
rect 14476 31668 14504 31708
rect 15470 31668 15476 31680
rect 13964 31640 14504 31668
rect 15431 31640 15476 31668
rect 13964 31628 13970 31640
rect 15470 31628 15476 31640
rect 15528 31628 15534 31680
rect 15580 31668 15608 31708
rect 17586 31696 17592 31708
rect 17644 31696 17650 31748
rect 18966 31696 18972 31748
rect 19024 31736 19030 31748
rect 19628 31736 19656 31971
rect 19794 31968 19800 31980
rect 19852 32008 19858 32020
rect 20346 32008 20352 32020
rect 19852 31980 20352 32008
rect 19852 31968 19858 31980
rect 20346 31968 20352 31980
rect 20404 31968 20410 32020
rect 19705 31943 19763 31949
rect 19705 31909 19717 31943
rect 19751 31940 19763 31943
rect 19978 31940 19984 31952
rect 19751 31912 19984 31940
rect 19751 31909 19763 31912
rect 19705 31903 19763 31909
rect 19978 31900 19984 31912
rect 20036 31900 20042 31952
rect 20254 31900 20260 31952
rect 20312 31940 20318 31952
rect 20625 31943 20683 31949
rect 20625 31940 20637 31943
rect 20312 31912 20637 31940
rect 20312 31900 20318 31912
rect 20625 31909 20637 31912
rect 20671 31909 20683 31943
rect 20625 31903 20683 31909
rect 22002 31872 22008 31884
rect 21963 31844 22008 31872
rect 22002 31832 22008 31844
rect 22060 31832 22066 31884
rect 19981 31807 20039 31813
rect 19981 31773 19993 31807
rect 20027 31804 20039 31807
rect 20346 31804 20352 31816
rect 20027 31776 20352 31804
rect 20027 31773 20039 31776
rect 19981 31767 20039 31773
rect 20346 31764 20352 31776
rect 20404 31764 20410 31816
rect 20441 31807 20499 31813
rect 20441 31773 20453 31807
rect 20487 31804 20499 31807
rect 21174 31804 21180 31816
rect 20487 31776 21180 31804
rect 20487 31773 20499 31776
rect 20441 31767 20499 31773
rect 21174 31764 21180 31776
rect 21232 31804 21238 31816
rect 21729 31807 21787 31813
rect 21729 31804 21741 31807
rect 21232 31776 21741 31804
rect 21232 31764 21238 31776
rect 21729 31773 21741 31776
rect 21775 31773 21787 31807
rect 21729 31767 21787 31773
rect 19024 31708 19656 31736
rect 19024 31696 19030 31708
rect 21450 31668 21456 31680
rect 15580 31640 21456 31668
rect 21450 31628 21456 31640
rect 21508 31628 21514 31680
rect 1104 31578 30820 31600
rect 1104 31526 10880 31578
rect 10932 31526 10944 31578
rect 10996 31526 11008 31578
rect 11060 31526 11072 31578
rect 11124 31526 11136 31578
rect 11188 31526 20811 31578
rect 20863 31526 20875 31578
rect 20927 31526 20939 31578
rect 20991 31526 21003 31578
rect 21055 31526 21067 31578
rect 21119 31526 30820 31578
rect 1104 31504 30820 31526
rect 1394 31464 1400 31476
rect 1355 31436 1400 31464
rect 1394 31424 1400 31436
rect 1452 31424 1458 31476
rect 2222 31424 2228 31476
rect 2280 31464 2286 31476
rect 3053 31467 3111 31473
rect 3053 31464 3065 31467
rect 2280 31436 3065 31464
rect 2280 31424 2286 31436
rect 3053 31433 3065 31436
rect 3099 31433 3111 31467
rect 3053 31427 3111 31433
rect 3234 31424 3240 31476
rect 3292 31464 3298 31476
rect 3878 31464 3884 31476
rect 3292 31436 3884 31464
rect 3292 31424 3298 31436
rect 3878 31424 3884 31436
rect 3936 31464 3942 31476
rect 5074 31464 5080 31476
rect 3936 31436 5080 31464
rect 3936 31424 3942 31436
rect 5074 31424 5080 31436
rect 5132 31424 5138 31476
rect 9674 31424 9680 31476
rect 9732 31464 9738 31476
rect 10781 31467 10839 31473
rect 10781 31464 10793 31467
rect 9732 31436 10793 31464
rect 9732 31424 9738 31436
rect 10781 31433 10793 31436
rect 10827 31464 10839 31467
rect 11606 31464 11612 31476
rect 10827 31436 11612 31464
rect 10827 31433 10839 31436
rect 10781 31427 10839 31433
rect 11606 31424 11612 31436
rect 11664 31424 11670 31476
rect 12250 31464 12256 31476
rect 12211 31436 12256 31464
rect 12250 31424 12256 31436
rect 12308 31424 12314 31476
rect 12897 31467 12955 31473
rect 12897 31433 12909 31467
rect 12943 31464 12955 31467
rect 13633 31467 13691 31473
rect 12943 31436 13400 31464
rect 12943 31433 12955 31436
rect 12897 31427 12955 31433
rect 2409 31399 2467 31405
rect 2409 31365 2421 31399
rect 2455 31396 2467 31399
rect 4154 31396 4160 31408
rect 2455 31368 3924 31396
rect 2455 31365 2467 31368
rect 2409 31359 2467 31365
rect 1581 31331 1639 31337
rect 1581 31297 1593 31331
rect 1627 31328 1639 31331
rect 3234 31328 3240 31340
rect 1627 31300 2636 31328
rect 3195 31300 3240 31328
rect 1627 31297 1639 31300
rect 1581 31291 1639 31297
rect 2041 31263 2099 31269
rect 2041 31229 2053 31263
rect 2087 31260 2099 31263
rect 2130 31260 2136 31272
rect 2087 31232 2136 31260
rect 2087 31229 2099 31232
rect 2041 31223 2099 31229
rect 2130 31220 2136 31232
rect 2188 31220 2194 31272
rect 2608 31201 2636 31300
rect 3234 31288 3240 31300
rect 3292 31288 3298 31340
rect 3896 31337 3924 31368
rect 4080 31368 4160 31396
rect 4080 31337 4108 31368
rect 4154 31356 4160 31368
rect 4212 31356 4218 31408
rect 4982 31396 4988 31408
rect 4264 31368 4988 31396
rect 4264 31337 4292 31368
rect 4982 31356 4988 31368
rect 5040 31356 5046 31408
rect 5258 31356 5264 31408
rect 5316 31396 5322 31408
rect 8570 31396 8576 31408
rect 5316 31368 8576 31396
rect 5316 31356 5322 31368
rect 8570 31356 8576 31368
rect 8628 31356 8634 31408
rect 12802 31396 12808 31408
rect 11716 31368 12808 31396
rect 3881 31331 3939 31337
rect 3881 31297 3893 31331
rect 3927 31328 3939 31331
rect 4065 31331 4123 31337
rect 3927 31300 4016 31328
rect 3927 31297 3939 31300
rect 3881 31291 3939 31297
rect 2593 31195 2651 31201
rect 2593 31161 2605 31195
rect 2639 31161 2651 31195
rect 3988 31192 4016 31300
rect 4065 31297 4077 31331
rect 4111 31297 4123 31331
rect 4065 31291 4123 31297
rect 4249 31331 4307 31337
rect 4249 31297 4261 31331
rect 4295 31297 4307 31331
rect 4249 31291 4307 31297
rect 4433 31331 4491 31337
rect 4433 31297 4445 31331
rect 4479 31328 4491 31331
rect 4522 31328 4528 31340
rect 4479 31300 4528 31328
rect 4479 31297 4491 31300
rect 4433 31291 4491 31297
rect 4522 31288 4528 31300
rect 4580 31328 4586 31340
rect 5350 31328 5356 31340
rect 4580 31300 5356 31328
rect 4580 31288 4586 31300
rect 5350 31288 5356 31300
rect 5408 31288 5414 31340
rect 6270 31288 6276 31340
rect 6328 31328 6334 31340
rect 7478 31331 7536 31337
rect 7478 31328 7490 31331
rect 6328 31300 7490 31328
rect 6328 31288 6334 31300
rect 7478 31297 7490 31300
rect 7524 31297 7536 31331
rect 7742 31328 7748 31340
rect 7703 31300 7748 31328
rect 7478 31291 7536 31297
rect 7742 31288 7748 31300
rect 7800 31288 7806 31340
rect 8297 31331 8355 31337
rect 8297 31297 8309 31331
rect 8343 31328 8355 31331
rect 9398 31328 9404 31340
rect 8343 31300 9404 31328
rect 8343 31297 8355 31300
rect 8297 31291 8355 31297
rect 9398 31288 9404 31300
rect 9456 31288 9462 31340
rect 9493 31331 9551 31337
rect 9493 31297 9505 31331
rect 9539 31328 9551 31331
rect 10318 31328 10324 31340
rect 9539 31300 10324 31328
rect 9539 31297 9551 31300
rect 9493 31291 9551 31297
rect 10318 31288 10324 31300
rect 10376 31288 10382 31340
rect 10870 31328 10876 31340
rect 10831 31300 10876 31328
rect 10870 31288 10876 31300
rect 10928 31288 10934 31340
rect 11514 31328 11520 31340
rect 11475 31300 11520 31328
rect 11514 31288 11520 31300
rect 11572 31288 11578 31340
rect 11716 31337 11744 31368
rect 12802 31356 12808 31368
rect 12860 31396 12866 31408
rect 13372 31405 13400 31436
rect 13633 31433 13645 31467
rect 13679 31464 13691 31467
rect 13814 31464 13820 31476
rect 13679 31436 13820 31464
rect 13679 31433 13691 31436
rect 13633 31427 13691 31433
rect 13814 31424 13820 31436
rect 13872 31424 13878 31476
rect 14550 31464 14556 31476
rect 14292 31436 14556 31464
rect 13357 31399 13415 31405
rect 12860 31368 13124 31396
rect 12860 31356 12866 31368
rect 13096 31340 13124 31368
rect 13357 31365 13369 31399
rect 13403 31365 13415 31399
rect 13357 31359 13415 31365
rect 11701 31331 11759 31337
rect 11701 31297 11713 31331
rect 11747 31297 11759 31331
rect 11701 31291 11759 31297
rect 12069 31331 12127 31337
rect 12069 31297 12081 31331
rect 12115 31328 12127 31331
rect 12710 31328 12716 31340
rect 12115 31300 12716 31328
rect 12115 31297 12127 31300
rect 12069 31291 12127 31297
rect 12710 31288 12716 31300
rect 12768 31288 12774 31340
rect 12986 31328 12992 31340
rect 12947 31300 12992 31328
rect 12986 31288 12992 31300
rect 13044 31288 13050 31340
rect 13078 31288 13084 31340
rect 13136 31328 13142 31340
rect 13265 31331 13323 31337
rect 13136 31300 13181 31328
rect 13136 31288 13142 31300
rect 13265 31297 13277 31331
rect 13311 31297 13323 31331
rect 13265 31291 13323 31297
rect 13495 31331 13553 31337
rect 13495 31297 13507 31331
rect 13541 31328 13553 31331
rect 13541 31300 13768 31328
rect 13541 31297 13553 31300
rect 13495 31291 13553 31297
rect 4157 31263 4215 31269
rect 4157 31229 4169 31263
rect 4203 31260 4215 31263
rect 4338 31260 4344 31272
rect 4203 31232 4344 31260
rect 4203 31229 4215 31232
rect 4157 31223 4215 31229
rect 4338 31220 4344 31232
rect 4396 31260 4402 31272
rect 5445 31263 5503 31269
rect 5445 31260 5457 31263
rect 4396 31232 5457 31260
rect 4396 31220 4402 31232
rect 5445 31229 5457 31232
rect 5491 31229 5503 31263
rect 5445 31223 5503 31229
rect 5721 31263 5779 31269
rect 5721 31229 5733 31263
rect 5767 31260 5779 31263
rect 6362 31260 6368 31272
rect 5767 31232 6368 31260
rect 5767 31229 5779 31232
rect 5721 31223 5779 31229
rect 6362 31220 6368 31232
rect 6420 31220 6426 31272
rect 9306 31220 9312 31272
rect 9364 31260 9370 31272
rect 11790 31260 11796 31272
rect 9364 31232 10824 31260
rect 11751 31232 11796 31260
rect 9364 31220 9370 31232
rect 4614 31192 4620 31204
rect 3988 31164 4620 31192
rect 2593 31155 2651 31161
rect 4614 31152 4620 31164
rect 4672 31152 4678 31204
rect 8757 31195 8815 31201
rect 8757 31161 8769 31195
rect 8803 31192 8815 31195
rect 10042 31192 10048 31204
rect 8803 31164 10048 31192
rect 8803 31161 8815 31164
rect 8757 31155 8815 31161
rect 10042 31152 10048 31164
rect 10100 31152 10106 31204
rect 2314 31084 2320 31136
rect 2372 31124 2378 31136
rect 2409 31127 2467 31133
rect 2409 31124 2421 31127
rect 2372 31096 2421 31124
rect 2372 31084 2378 31096
rect 2409 31093 2421 31096
rect 2455 31093 2467 31127
rect 3694 31124 3700 31136
rect 3655 31096 3700 31124
rect 2409 31087 2467 31093
rect 3694 31084 3700 31096
rect 3752 31084 3758 31136
rect 5810 31084 5816 31136
rect 5868 31124 5874 31136
rect 6365 31127 6423 31133
rect 6365 31124 6377 31127
rect 5868 31096 6377 31124
rect 5868 31084 5874 31096
rect 6365 31093 6377 31096
rect 6411 31093 6423 31127
rect 6365 31087 6423 31093
rect 7006 31084 7012 31136
rect 7064 31124 7070 31136
rect 8110 31124 8116 31136
rect 7064 31096 8116 31124
rect 7064 31084 7070 31096
rect 8110 31084 8116 31096
rect 8168 31084 8174 31136
rect 8570 31124 8576 31136
rect 8483 31096 8576 31124
rect 8570 31084 8576 31096
rect 8628 31124 8634 31136
rect 9769 31127 9827 31133
rect 9769 31124 9781 31127
rect 8628 31096 9781 31124
rect 8628 31084 8634 31096
rect 9769 31093 9781 31096
rect 9815 31124 9827 31127
rect 9858 31124 9864 31136
rect 9815 31096 9864 31124
rect 9815 31093 9827 31096
rect 9769 31087 9827 31093
rect 9858 31084 9864 31096
rect 9916 31084 9922 31136
rect 9953 31127 10011 31133
rect 9953 31093 9965 31127
rect 9999 31124 10011 31127
rect 10686 31124 10692 31136
rect 9999 31096 10692 31124
rect 9999 31093 10011 31096
rect 9953 31087 10011 31093
rect 10686 31084 10692 31096
rect 10744 31084 10750 31136
rect 10796 31124 10824 31232
rect 11790 31220 11796 31232
rect 11848 31220 11854 31272
rect 11885 31263 11943 31269
rect 11885 31229 11897 31263
rect 11931 31229 11943 31263
rect 11885 31223 11943 31229
rect 11698 31152 11704 31204
rect 11756 31192 11762 31204
rect 11900 31192 11928 31223
rect 12897 31195 12955 31201
rect 12897 31192 12909 31195
rect 11756 31164 11928 31192
rect 12406 31164 12909 31192
rect 11756 31152 11762 31164
rect 12406 31124 12434 31164
rect 12897 31161 12909 31164
rect 12943 31161 12955 31195
rect 13280 31192 13308 31291
rect 13740 31272 13768 31300
rect 13998 31288 14004 31340
rect 14056 31328 14062 31340
rect 14292 31337 14320 31436
rect 14550 31424 14556 31436
rect 14608 31424 14614 31476
rect 15378 31464 15384 31476
rect 15339 31436 15384 31464
rect 15378 31424 15384 31436
rect 15436 31424 15442 31476
rect 17862 31464 17868 31476
rect 17823 31436 17868 31464
rect 17862 31424 17868 31436
rect 17920 31424 17926 31476
rect 19058 31424 19064 31476
rect 19116 31464 19122 31476
rect 19429 31467 19487 31473
rect 19116 31436 19380 31464
rect 19116 31424 19122 31436
rect 14369 31399 14427 31405
rect 14369 31365 14381 31399
rect 14415 31396 14427 31399
rect 15562 31396 15568 31408
rect 14415 31368 15568 31396
rect 14415 31365 14427 31368
rect 14369 31359 14427 31365
rect 15562 31356 15568 31368
rect 15620 31356 15626 31408
rect 17773 31399 17831 31405
rect 17773 31396 17785 31399
rect 16316 31368 17785 31396
rect 16316 31340 16344 31368
rect 17773 31365 17785 31368
rect 17819 31365 17831 31399
rect 17773 31359 17831 31365
rect 18506 31356 18512 31408
rect 18564 31396 18570 31408
rect 19352 31396 19380 31436
rect 19429 31433 19441 31467
rect 19475 31464 19487 31467
rect 19518 31464 19524 31476
rect 19475 31436 19524 31464
rect 19475 31433 19487 31436
rect 19429 31427 19487 31433
rect 19518 31424 19524 31436
rect 19576 31424 19582 31476
rect 18564 31368 19288 31396
rect 19352 31368 20668 31396
rect 18564 31356 18570 31368
rect 14093 31331 14151 31337
rect 14093 31328 14105 31331
rect 14056 31300 14105 31328
rect 14056 31288 14062 31300
rect 14093 31297 14105 31300
rect 14139 31297 14151 31331
rect 14093 31291 14151 31297
rect 14241 31331 14320 31337
rect 14241 31297 14253 31331
rect 14287 31300 14320 31331
rect 14458 31328 14464 31340
rect 14419 31300 14464 31328
rect 14287 31297 14299 31300
rect 14241 31291 14299 31297
rect 14458 31288 14464 31300
rect 14516 31288 14522 31340
rect 14558 31331 14616 31337
rect 14558 31297 14570 31331
rect 14604 31297 14616 31331
rect 14558 31291 14616 31297
rect 13722 31220 13728 31272
rect 13780 31260 13786 31272
rect 14568 31260 14596 31291
rect 15194 31288 15200 31340
rect 15252 31328 15258 31340
rect 15749 31331 15807 31337
rect 15749 31328 15761 31331
rect 15252 31300 15761 31328
rect 15252 31288 15258 31300
rect 15749 31297 15761 31300
rect 15795 31297 15807 31331
rect 15749 31291 15807 31297
rect 15841 31331 15899 31337
rect 15841 31297 15853 31331
rect 15887 31328 15899 31331
rect 16298 31328 16304 31340
rect 15887 31300 16304 31328
rect 15887 31297 15899 31300
rect 15841 31291 15899 31297
rect 16298 31288 16304 31300
rect 16356 31288 16362 31340
rect 16666 31328 16672 31340
rect 16627 31300 16672 31328
rect 16666 31288 16672 31300
rect 16724 31288 16730 31340
rect 18690 31328 18696 31340
rect 18651 31300 18696 31328
rect 18690 31288 18696 31300
rect 18748 31288 18754 31340
rect 18874 31328 18880 31340
rect 18835 31300 18880 31328
rect 18874 31288 18880 31300
rect 18932 31288 18938 31340
rect 18969 31331 19027 31337
rect 18969 31297 18981 31331
rect 19015 31328 19027 31331
rect 19150 31328 19156 31340
rect 19015 31300 19156 31328
rect 19015 31297 19027 31300
rect 18969 31291 19027 31297
rect 19150 31288 19156 31300
rect 19208 31288 19214 31340
rect 19260 31337 19288 31368
rect 19245 31331 19303 31337
rect 19245 31297 19257 31331
rect 19291 31297 19303 31331
rect 19245 31291 19303 31297
rect 19889 31331 19947 31337
rect 19889 31297 19901 31331
rect 19935 31328 19947 31331
rect 20346 31328 20352 31340
rect 19935 31300 20352 31328
rect 19935 31297 19947 31300
rect 19889 31291 19947 31297
rect 20346 31288 20352 31300
rect 20404 31288 20410 31340
rect 20640 31328 20668 31368
rect 21450 31356 21456 31408
rect 21508 31396 21514 31408
rect 22094 31396 22100 31408
rect 21508 31368 22100 31396
rect 21508 31356 21514 31368
rect 22094 31356 22100 31368
rect 22152 31356 22158 31408
rect 20714 31328 20720 31340
rect 20627 31300 20720 31328
rect 20714 31288 20720 31300
rect 20772 31288 20778 31340
rect 21103 31331 21161 31337
rect 21103 31297 21115 31331
rect 21149 31328 21161 31331
rect 21269 31331 21327 31337
rect 21149 31300 21220 31328
rect 21149 31297 21161 31300
rect 21103 31291 21161 31297
rect 13780 31232 14596 31260
rect 16025 31263 16083 31269
rect 13780 31220 13786 31232
rect 16025 31229 16037 31263
rect 16071 31260 16083 31263
rect 17589 31263 17647 31269
rect 17589 31260 17601 31263
rect 16071 31232 17601 31260
rect 16071 31229 16083 31232
rect 16025 31223 16083 31229
rect 17589 31229 17601 31232
rect 17635 31260 17647 31263
rect 19061 31263 19119 31269
rect 17635 31232 19012 31260
rect 17635 31229 17647 31232
rect 17589 31223 17647 31229
rect 15470 31192 15476 31204
rect 13280 31164 15476 31192
rect 12897 31155 12955 31161
rect 15470 31152 15476 31164
rect 15528 31152 15534 31204
rect 10796 31096 12434 31124
rect 13814 31084 13820 31136
rect 13872 31124 13878 31136
rect 14458 31124 14464 31136
rect 13872 31096 14464 31124
rect 13872 31084 13878 31096
rect 14458 31084 14464 31096
rect 14516 31084 14522 31136
rect 14734 31124 14740 31136
rect 14695 31096 14740 31124
rect 14734 31084 14740 31096
rect 14792 31084 14798 31136
rect 16761 31127 16819 31133
rect 16761 31093 16773 31127
rect 16807 31124 16819 31127
rect 17218 31124 17224 31136
rect 16807 31096 17224 31124
rect 16807 31093 16819 31096
rect 16761 31087 16819 31093
rect 17218 31084 17224 31096
rect 17276 31084 17282 31136
rect 18233 31127 18291 31133
rect 18233 31093 18245 31127
rect 18279 31124 18291 31127
rect 18414 31124 18420 31136
rect 18279 31096 18420 31124
rect 18279 31093 18291 31096
rect 18233 31087 18291 31093
rect 18414 31084 18420 31096
rect 18472 31084 18478 31136
rect 18984 31124 19012 31232
rect 19061 31229 19073 31263
rect 19107 31260 19119 31263
rect 19610 31260 19616 31272
rect 19107 31232 19616 31260
rect 19107 31229 19119 31232
rect 19061 31223 19119 31229
rect 19610 31220 19616 31232
rect 19668 31220 19674 31272
rect 20806 31220 20812 31272
rect 20864 31260 20870 31272
rect 20901 31263 20959 31269
rect 20901 31260 20913 31263
rect 20864 31232 20913 31260
rect 20864 31220 20870 31232
rect 20901 31229 20913 31232
rect 20947 31229 20959 31263
rect 20901 31223 20959 31229
rect 20990 31220 20996 31272
rect 21048 31260 21054 31272
rect 21192 31260 21220 31300
rect 21269 31297 21281 31331
rect 21315 31328 21327 31331
rect 22002 31328 22008 31340
rect 21315 31300 22008 31328
rect 21315 31297 21327 31300
rect 21269 31291 21327 31297
rect 22002 31288 22008 31300
rect 22060 31288 22066 31340
rect 29822 31328 29828 31340
rect 29783 31300 29828 31328
rect 29822 31288 29828 31300
rect 29880 31288 29886 31340
rect 21726 31260 21732 31272
rect 21048 31232 21093 31260
rect 21192 31232 21732 31260
rect 21048 31220 21054 31232
rect 21726 31220 21732 31232
rect 21784 31220 21790 31272
rect 21821 31263 21879 31269
rect 21821 31229 21833 31263
rect 21867 31229 21879 31263
rect 21821 31223 21879 31229
rect 22097 31263 22155 31269
rect 22097 31229 22109 31263
rect 22143 31260 22155 31263
rect 22278 31260 22284 31272
rect 22143 31232 22284 31260
rect 22143 31229 22155 31232
rect 22097 31223 22155 31229
rect 19150 31152 19156 31204
rect 19208 31192 19214 31204
rect 20533 31195 20591 31201
rect 20533 31192 20545 31195
rect 19208 31164 20545 31192
rect 19208 31152 19214 31164
rect 20533 31161 20545 31164
rect 20579 31161 20591 31195
rect 20533 31155 20591 31161
rect 21174 31152 21180 31204
rect 21232 31192 21238 31204
rect 21450 31192 21456 31204
rect 21232 31164 21456 31192
rect 21232 31152 21238 31164
rect 21450 31152 21456 31164
rect 21508 31192 21514 31204
rect 21836 31192 21864 31223
rect 22278 31220 22284 31232
rect 22336 31220 22342 31272
rect 30098 31260 30104 31272
rect 30059 31232 30104 31260
rect 30098 31220 30104 31232
rect 30156 31220 30162 31272
rect 21508 31164 21864 31192
rect 21508 31152 21514 31164
rect 19610 31124 19616 31136
rect 18984 31096 19616 31124
rect 19610 31084 19616 31096
rect 19668 31084 19674 31136
rect 19978 31124 19984 31136
rect 19939 31096 19984 31124
rect 19978 31084 19984 31096
rect 20036 31084 20042 31136
rect 1104 31034 30820 31056
rect 1104 30982 5915 31034
rect 5967 30982 5979 31034
rect 6031 30982 6043 31034
rect 6095 30982 6107 31034
rect 6159 30982 6171 31034
rect 6223 30982 15846 31034
rect 15898 30982 15910 31034
rect 15962 30982 15974 31034
rect 16026 30982 16038 31034
rect 16090 30982 16102 31034
rect 16154 30982 25776 31034
rect 25828 30982 25840 31034
rect 25892 30982 25904 31034
rect 25956 30982 25968 31034
rect 26020 30982 26032 31034
rect 26084 30982 30820 31034
rect 1104 30960 30820 30982
rect 1412 30892 2268 30920
rect 1412 30725 1440 30892
rect 1581 30855 1639 30861
rect 1581 30821 1593 30855
rect 1627 30821 1639 30855
rect 1581 30815 1639 30821
rect 2041 30855 2099 30861
rect 2041 30821 2053 30855
rect 2087 30852 2099 30855
rect 2130 30852 2136 30864
rect 2087 30824 2136 30852
rect 2087 30821 2099 30824
rect 2041 30815 2099 30821
rect 1596 30784 1624 30815
rect 2130 30812 2136 30824
rect 2188 30812 2194 30864
rect 2240 30852 2268 30892
rect 2314 30880 2320 30932
rect 2372 30920 2378 30932
rect 2409 30923 2467 30929
rect 2409 30920 2421 30923
rect 2372 30892 2421 30920
rect 2372 30880 2378 30892
rect 2409 30889 2421 30892
rect 2455 30889 2467 30923
rect 3050 30920 3056 30932
rect 3011 30892 3056 30920
rect 2409 30883 2467 30889
rect 3050 30880 3056 30892
rect 3108 30880 3114 30932
rect 5905 30923 5963 30929
rect 5905 30889 5917 30923
rect 5951 30920 5963 30923
rect 6270 30920 6276 30932
rect 5951 30892 6276 30920
rect 5951 30889 5963 30892
rect 5905 30883 5963 30889
rect 6270 30880 6276 30892
rect 6328 30880 6334 30932
rect 9309 30923 9367 30929
rect 9309 30889 9321 30923
rect 9355 30920 9367 30923
rect 9858 30920 9864 30932
rect 9355 30892 9864 30920
rect 9355 30889 9367 30892
rect 9309 30883 9367 30889
rect 9858 30880 9864 30892
rect 9916 30880 9922 30932
rect 10870 30880 10876 30932
rect 10928 30920 10934 30932
rect 15381 30923 15439 30929
rect 15381 30920 15393 30923
rect 10928 30892 15393 30920
rect 10928 30880 10934 30892
rect 15381 30889 15393 30892
rect 15427 30889 15439 30923
rect 18506 30920 18512 30932
rect 18467 30892 18512 30920
rect 15381 30883 15439 30889
rect 2593 30855 2651 30861
rect 2593 30852 2605 30855
rect 2240 30824 2605 30852
rect 2593 30821 2605 30824
rect 2639 30821 2651 30855
rect 6454 30852 6460 30864
rect 2593 30815 2651 30821
rect 5092 30824 6460 30852
rect 5092 30793 5120 30824
rect 6454 30812 6460 30824
rect 6512 30812 6518 30864
rect 7098 30852 7104 30864
rect 7059 30824 7104 30852
rect 7098 30812 7104 30824
rect 7156 30812 7162 30864
rect 8846 30852 8852 30864
rect 7668 30824 8852 30852
rect 5077 30787 5135 30793
rect 1596 30756 3832 30784
rect 1397 30719 1455 30725
rect 1397 30685 1409 30719
rect 1443 30685 1455 30719
rect 1397 30679 1455 30685
rect 2958 30676 2964 30728
rect 3016 30716 3022 30728
rect 3804 30725 3832 30756
rect 5077 30753 5089 30787
rect 5123 30753 5135 30787
rect 5077 30747 5135 30753
rect 5169 30787 5227 30793
rect 5169 30753 5181 30787
rect 5215 30784 5227 30787
rect 6362 30784 6368 30796
rect 5215 30756 6368 30784
rect 5215 30753 5227 30756
rect 5169 30747 5227 30753
rect 6362 30744 6368 30756
rect 6420 30784 6426 30796
rect 7561 30787 7619 30793
rect 7561 30784 7573 30787
rect 6420 30756 7573 30784
rect 6420 30744 6426 30756
rect 7561 30753 7573 30756
rect 7607 30753 7619 30787
rect 7561 30747 7619 30753
rect 3237 30719 3295 30725
rect 3237 30716 3249 30719
rect 3016 30688 3249 30716
rect 3016 30676 3022 30688
rect 3237 30685 3249 30688
rect 3283 30685 3295 30719
rect 3237 30679 3295 30685
rect 3789 30719 3847 30725
rect 3789 30685 3801 30719
rect 3835 30685 3847 30719
rect 4890 30716 4896 30728
rect 4851 30688 4896 30716
rect 3789 30679 3847 30685
rect 4890 30676 4896 30688
rect 4948 30676 4954 30728
rect 5258 30716 5264 30728
rect 5219 30688 5264 30716
rect 5258 30676 5264 30688
rect 5316 30676 5322 30728
rect 5350 30676 5356 30728
rect 5408 30716 5414 30728
rect 5445 30719 5503 30725
rect 5445 30716 5457 30719
rect 5408 30688 5457 30716
rect 5408 30676 5414 30688
rect 5445 30685 5457 30688
rect 5491 30685 5503 30719
rect 5445 30679 5503 30685
rect 6089 30719 6147 30725
rect 6089 30685 6101 30719
rect 6135 30685 6147 30719
rect 6089 30679 6147 30685
rect 6273 30719 6331 30725
rect 6273 30685 6285 30719
rect 6319 30716 6331 30719
rect 6457 30719 6515 30725
rect 6319 30688 6408 30716
rect 6319 30685 6331 30688
rect 6273 30679 6331 30685
rect 5810 30648 5816 30660
rect 2746 30620 5816 30648
rect 2409 30583 2467 30589
rect 2409 30549 2421 30583
rect 2455 30580 2467 30583
rect 2746 30580 2774 30620
rect 5810 30608 5816 30620
rect 5868 30648 5874 30660
rect 6104 30648 6132 30679
rect 5868 30620 6132 30648
rect 5868 30608 5874 30620
rect 3970 30580 3976 30592
rect 2455 30552 2774 30580
rect 3931 30552 3976 30580
rect 2455 30549 2467 30552
rect 2409 30543 2467 30549
rect 3970 30540 3976 30552
rect 4028 30540 4034 30592
rect 4706 30580 4712 30592
rect 4667 30552 4712 30580
rect 4706 30540 4712 30552
rect 4764 30540 4770 30592
rect 6380 30580 6408 30688
rect 6457 30685 6469 30719
rect 6503 30685 6515 30719
rect 6457 30679 6515 30685
rect 6641 30719 6699 30725
rect 6641 30685 6653 30719
rect 6687 30716 6699 30719
rect 7285 30719 7343 30725
rect 6687 30688 7236 30716
rect 6687 30685 6699 30688
rect 6641 30679 6699 30685
rect 6472 30648 6500 30679
rect 7006 30648 7012 30660
rect 6472 30620 7012 30648
rect 7006 30608 7012 30620
rect 7064 30608 7070 30660
rect 7208 30648 7236 30688
rect 7285 30685 7297 30719
rect 7331 30716 7343 30719
rect 7374 30716 7380 30728
rect 7331 30688 7380 30716
rect 7331 30685 7343 30688
rect 7285 30679 7343 30685
rect 7374 30676 7380 30688
rect 7432 30676 7438 30728
rect 7466 30676 7472 30728
rect 7524 30716 7530 30728
rect 7668 30725 7696 30824
rect 8846 30812 8852 30824
rect 8904 30812 8910 30864
rect 11238 30812 11244 30864
rect 11296 30812 11302 30864
rect 11974 30852 11980 30864
rect 11935 30824 11980 30852
rect 11974 30812 11980 30824
rect 12032 30812 12038 30864
rect 12434 30812 12440 30864
rect 12492 30852 12498 30864
rect 14093 30855 14151 30861
rect 12492 30824 13492 30852
rect 12492 30812 12498 30824
rect 11256 30784 11284 30812
rect 7944 30756 11284 30784
rect 11517 30787 11575 30793
rect 7653 30719 7711 30725
rect 7524 30688 7569 30716
rect 7524 30676 7530 30688
rect 7653 30685 7665 30719
rect 7699 30685 7711 30719
rect 7837 30719 7895 30725
rect 7837 30718 7849 30719
rect 7653 30679 7711 30685
rect 7760 30690 7849 30718
rect 7760 30648 7788 30690
rect 7837 30685 7849 30690
rect 7883 30718 7895 30719
rect 7944 30718 7972 30756
rect 11517 30753 11529 30787
rect 11563 30784 11575 30787
rect 11882 30784 11888 30796
rect 11563 30756 11888 30784
rect 11563 30753 11575 30756
rect 11517 30747 11575 30753
rect 11882 30744 11888 30756
rect 11940 30744 11946 30796
rect 12066 30744 12072 30796
rect 12124 30784 12130 30796
rect 13464 30784 13492 30824
rect 14093 30821 14105 30855
rect 14139 30852 14151 30855
rect 14274 30852 14280 30864
rect 14139 30824 14280 30852
rect 14139 30821 14151 30824
rect 14093 30815 14151 30821
rect 14274 30812 14280 30824
rect 14332 30812 14338 30864
rect 12124 30756 13400 30784
rect 13464 30756 15332 30784
rect 12124 30744 12130 30756
rect 7883 30690 7972 30718
rect 7883 30685 7895 30690
rect 7837 30679 7895 30685
rect 8294 30676 8300 30728
rect 8352 30716 8358 30728
rect 9401 30719 9459 30725
rect 9401 30716 9413 30719
rect 8352 30688 9413 30716
rect 8352 30676 8358 30688
rect 9401 30685 9413 30688
rect 9447 30685 9459 30719
rect 9401 30679 9459 30685
rect 9950 30676 9956 30728
rect 10008 30716 10014 30728
rect 10045 30719 10103 30725
rect 10045 30716 10057 30719
rect 10008 30688 10057 30716
rect 10008 30676 10014 30688
rect 10045 30685 10057 30688
rect 10091 30716 10103 30719
rect 10134 30716 10140 30728
rect 10091 30688 10140 30716
rect 10091 30685 10103 30688
rect 10045 30679 10103 30685
rect 10134 30676 10140 30688
rect 10192 30676 10198 30728
rect 10686 30716 10692 30728
rect 10647 30688 10692 30716
rect 10686 30676 10692 30688
rect 10744 30676 10750 30728
rect 11241 30719 11299 30725
rect 11241 30685 11253 30719
rect 11287 30685 11299 30719
rect 11422 30716 11428 30728
rect 11383 30688 11428 30716
rect 11241 30679 11299 30685
rect 11256 30648 11284 30679
rect 11422 30676 11428 30688
rect 11480 30676 11486 30728
rect 11609 30719 11667 30725
rect 11609 30685 11621 30719
rect 11655 30716 11667 30719
rect 11698 30716 11704 30728
rect 11655 30688 11704 30716
rect 11655 30685 11667 30688
rect 11609 30679 11667 30685
rect 11698 30676 11704 30688
rect 11756 30676 11762 30728
rect 11793 30719 11851 30725
rect 11793 30685 11805 30719
rect 11839 30716 11851 30719
rect 12894 30716 12900 30728
rect 11839 30688 12900 30716
rect 11839 30685 11851 30688
rect 11793 30679 11851 30685
rect 12894 30676 12900 30688
rect 12952 30676 12958 30728
rect 12989 30719 13047 30725
rect 12989 30685 13001 30719
rect 13035 30716 13047 30719
rect 13078 30716 13084 30728
rect 13035 30688 13084 30716
rect 13035 30685 13047 30688
rect 12989 30679 13047 30685
rect 13078 30676 13084 30688
rect 13136 30676 13142 30728
rect 13262 30716 13268 30728
rect 13223 30688 13268 30716
rect 13262 30676 13268 30688
rect 13320 30676 13326 30728
rect 11514 30648 11520 30660
rect 7208 30620 7788 30648
rect 7852 30620 10640 30648
rect 11256 30620 11520 30648
rect 6454 30580 6460 30592
rect 6367 30552 6460 30580
rect 6454 30540 6460 30552
rect 6512 30580 6518 30592
rect 7466 30580 7472 30592
rect 6512 30552 7472 30580
rect 6512 30540 6518 30552
rect 7466 30540 7472 30552
rect 7524 30580 7530 30592
rect 7852 30580 7880 30620
rect 8938 30580 8944 30592
rect 7524 30552 7880 30580
rect 8899 30552 8944 30580
rect 7524 30540 7530 30552
rect 8938 30540 8944 30552
rect 8996 30540 9002 30592
rect 9398 30540 9404 30592
rect 9456 30580 9462 30592
rect 10505 30583 10563 30589
rect 10505 30580 10517 30583
rect 9456 30552 10517 30580
rect 9456 30540 9462 30552
rect 10505 30549 10517 30552
rect 10551 30549 10563 30583
rect 10612 30580 10640 30620
rect 11514 30608 11520 30620
rect 11572 30648 11578 30660
rect 12250 30648 12256 30660
rect 11572 30620 12256 30648
rect 11572 30608 11578 30620
rect 12250 30608 12256 30620
rect 12308 30608 12314 30660
rect 13372 30648 13400 30756
rect 13722 30676 13728 30728
rect 13780 30716 13786 30728
rect 14231 30719 14289 30725
rect 14231 30716 14243 30719
rect 13780 30688 14243 30716
rect 13780 30676 13786 30688
rect 14231 30685 14243 30688
rect 14277 30685 14289 30719
rect 14458 30716 14464 30728
rect 14419 30688 14464 30716
rect 14231 30679 14289 30685
rect 14458 30676 14464 30688
rect 14516 30676 14522 30728
rect 14550 30676 14556 30728
rect 14608 30725 14614 30728
rect 14608 30719 14647 30725
rect 14635 30685 14647 30719
rect 14608 30679 14647 30685
rect 14737 30719 14795 30725
rect 14737 30685 14749 30719
rect 14783 30716 14795 30719
rect 15102 30716 15108 30728
rect 14783 30688 15108 30716
rect 14783 30685 14795 30688
rect 14737 30679 14795 30685
rect 14608 30676 14614 30679
rect 15102 30676 15108 30688
rect 15160 30676 15166 30728
rect 15304 30725 15332 30756
rect 15289 30719 15347 30725
rect 15289 30685 15301 30719
rect 15335 30685 15347 30719
rect 15396 30716 15424 30883
rect 18506 30880 18512 30892
rect 18564 30880 18570 30932
rect 19794 30880 19800 30932
rect 19852 30920 19858 30932
rect 19981 30923 20039 30929
rect 19981 30920 19993 30923
rect 19852 30892 19993 30920
rect 19852 30880 19858 30892
rect 19981 30889 19993 30892
rect 20027 30889 20039 30923
rect 19981 30883 20039 30889
rect 20165 30923 20223 30929
rect 20165 30889 20177 30923
rect 20211 30920 20223 30923
rect 20990 30920 20996 30932
rect 20211 30892 20996 30920
rect 20211 30889 20223 30892
rect 20165 30883 20223 30889
rect 20990 30880 20996 30892
rect 21048 30880 21054 30932
rect 17405 30855 17463 30861
rect 17405 30821 17417 30855
rect 17451 30852 17463 30855
rect 17586 30852 17592 30864
rect 17451 30824 17592 30852
rect 17451 30821 17463 30824
rect 17405 30815 17463 30821
rect 17586 30812 17592 30824
rect 17644 30852 17650 30864
rect 18601 30855 18659 30861
rect 17644 30824 18552 30852
rect 17644 30812 17650 30824
rect 18414 30784 18420 30796
rect 16500 30756 17356 30784
rect 18375 30756 18420 30784
rect 16025 30719 16083 30725
rect 16025 30716 16037 30719
rect 15396 30688 16037 30716
rect 15289 30679 15347 30685
rect 16025 30685 16037 30688
rect 16071 30685 16083 30719
rect 16025 30679 16083 30685
rect 14369 30651 14427 30657
rect 14369 30648 14381 30651
rect 13372 30620 14381 30648
rect 14369 30617 14381 30620
rect 14415 30617 14427 30651
rect 16206 30648 16212 30660
rect 16167 30620 16212 30648
rect 14369 30611 14427 30617
rect 16206 30608 16212 30620
rect 16264 30608 16270 30660
rect 16500 30580 16528 30756
rect 17126 30716 17132 30728
rect 17087 30688 17132 30716
rect 17126 30676 17132 30688
rect 17184 30676 17190 30728
rect 17221 30719 17279 30725
rect 17221 30685 17233 30719
rect 17267 30685 17279 30719
rect 17221 30679 17279 30685
rect 17034 30608 17040 30660
rect 17092 30648 17098 30660
rect 17236 30648 17264 30679
rect 17092 30620 17264 30648
rect 17328 30648 17356 30756
rect 18414 30744 18420 30756
rect 18472 30744 18478 30796
rect 18524 30784 18552 30824
rect 18601 30821 18613 30855
rect 18647 30852 18659 30855
rect 20806 30852 20812 30864
rect 18647 30824 20812 30852
rect 18647 30821 18659 30824
rect 18601 30815 18659 30821
rect 20806 30812 20812 30824
rect 20864 30812 20870 30864
rect 20901 30855 20959 30861
rect 20901 30821 20913 30855
rect 20947 30852 20959 30855
rect 21542 30852 21548 30864
rect 20947 30824 21548 30852
rect 20947 30821 20959 30824
rect 20901 30815 20959 30821
rect 21542 30812 21548 30824
rect 21600 30812 21606 30864
rect 18782 30784 18788 30796
rect 18524 30756 18788 30784
rect 18782 30744 18788 30756
rect 18840 30744 18846 30796
rect 20714 30744 20720 30796
rect 20772 30784 20778 30796
rect 21177 30787 21235 30793
rect 21177 30784 21189 30787
rect 20772 30756 21189 30784
rect 20772 30744 20778 30756
rect 21177 30753 21189 30756
rect 21223 30753 21235 30787
rect 23293 30787 23351 30793
rect 23293 30784 23305 30787
rect 21177 30747 21235 30753
rect 22066 30756 23305 30784
rect 22066 30728 22094 30756
rect 23293 30753 23305 30756
rect 23339 30753 23351 30787
rect 23293 30747 23351 30753
rect 17494 30716 17500 30728
rect 17455 30688 17500 30716
rect 17494 30676 17500 30688
rect 17552 30676 17558 30728
rect 18693 30719 18751 30725
rect 18693 30685 18705 30719
rect 18739 30716 18751 30719
rect 19058 30716 19064 30728
rect 18739 30688 19064 30716
rect 18739 30685 18751 30688
rect 18693 30679 18751 30685
rect 19058 30676 19064 30688
rect 19116 30676 19122 30728
rect 21266 30716 21272 30728
rect 21227 30688 21272 30716
rect 21266 30676 21272 30688
rect 21324 30676 21330 30728
rect 21634 30676 21640 30728
rect 21692 30716 21698 30728
rect 21692 30688 21737 30716
rect 21692 30676 21698 30688
rect 21818 30676 21824 30728
rect 21876 30716 21882 30728
rect 22002 30716 22008 30728
rect 21876 30688 21921 30716
rect 21963 30688 22008 30716
rect 21876 30676 21882 30688
rect 22002 30676 22008 30688
rect 22060 30688 22094 30728
rect 22060 30676 22066 30688
rect 22370 30676 22376 30728
rect 22428 30716 22434 30728
rect 23201 30719 23259 30725
rect 23201 30716 23213 30719
rect 22428 30688 23213 30716
rect 22428 30676 22434 30688
rect 23201 30685 23213 30688
rect 23247 30685 23259 30719
rect 23201 30679 23259 30685
rect 19150 30648 19156 30660
rect 17328 30620 19156 30648
rect 17092 30608 17098 30620
rect 19150 30608 19156 30620
rect 19208 30608 19214 30660
rect 19797 30651 19855 30657
rect 19797 30617 19809 30651
rect 19843 30617 19855 30651
rect 19797 30611 19855 30617
rect 10612 30552 16528 30580
rect 16945 30583 17003 30589
rect 10505 30543 10563 30549
rect 16945 30549 16957 30583
rect 16991 30580 17003 30583
rect 18046 30580 18052 30592
rect 16991 30552 18052 30580
rect 16991 30549 17003 30552
rect 16945 30543 17003 30549
rect 18046 30540 18052 30552
rect 18104 30540 18110 30592
rect 19812 30580 19840 30611
rect 19886 30608 19892 30660
rect 19944 30648 19950 30660
rect 19997 30651 20055 30657
rect 19997 30648 20009 30651
rect 19944 30620 20009 30648
rect 19944 30608 19950 30620
rect 19997 30617 20009 30620
rect 20043 30617 20055 30651
rect 21284 30648 21312 30676
rect 22465 30651 22523 30657
rect 22465 30648 22477 30651
rect 21284 30620 22477 30648
rect 19997 30611 20055 30617
rect 22465 30617 22477 30620
rect 22511 30617 22523 30651
rect 22646 30648 22652 30660
rect 22607 30620 22652 30648
rect 22465 30611 22523 30617
rect 22646 30608 22652 30620
rect 22704 30608 22710 30660
rect 20530 30580 20536 30592
rect 19812 30552 20536 30580
rect 20530 30540 20536 30552
rect 20588 30540 20594 30592
rect 1104 30490 30820 30512
rect 1104 30438 10880 30490
rect 10932 30438 10944 30490
rect 10996 30438 11008 30490
rect 11060 30438 11072 30490
rect 11124 30438 11136 30490
rect 11188 30438 20811 30490
rect 20863 30438 20875 30490
rect 20927 30438 20939 30490
rect 20991 30438 21003 30490
rect 21055 30438 21067 30490
rect 21119 30438 30820 30490
rect 1104 30416 30820 30438
rect 2317 30379 2375 30385
rect 2317 30345 2329 30379
rect 2363 30376 2375 30379
rect 4614 30376 4620 30388
rect 2363 30348 4476 30376
rect 4575 30348 4620 30376
rect 2363 30345 2375 30348
rect 2317 30339 2375 30345
rect 3504 30311 3562 30317
rect 3504 30277 3516 30311
rect 3550 30308 3562 30311
rect 3694 30308 3700 30320
rect 3550 30280 3700 30308
rect 3550 30277 3562 30280
rect 3504 30271 3562 30277
rect 3694 30268 3700 30280
rect 3752 30268 3758 30320
rect 4448 30308 4476 30348
rect 4614 30336 4620 30348
rect 4672 30336 4678 30388
rect 7374 30376 7380 30388
rect 4724 30348 7380 30376
rect 4724 30308 4752 30348
rect 7374 30336 7380 30348
rect 7432 30376 7438 30388
rect 7745 30379 7803 30385
rect 7745 30376 7757 30379
rect 7432 30348 7757 30376
rect 7432 30336 7438 30348
rect 7745 30345 7757 30348
rect 7791 30345 7803 30379
rect 7745 30339 7803 30345
rect 10778 30336 10784 30388
rect 10836 30376 10842 30388
rect 12066 30376 12072 30388
rect 10836 30348 12072 30376
rect 10836 30336 10842 30348
rect 12066 30336 12072 30348
rect 12124 30336 12130 30388
rect 12802 30336 12808 30388
rect 12860 30376 12866 30388
rect 14550 30376 14556 30388
rect 12860 30348 14556 30376
rect 12860 30336 12866 30348
rect 14550 30336 14556 30348
rect 14608 30336 14614 30388
rect 16206 30376 16212 30388
rect 15120 30348 16212 30376
rect 4448 30280 4752 30308
rect 6632 30311 6690 30317
rect 6632 30277 6644 30311
rect 6678 30308 6690 30311
rect 7098 30308 7104 30320
rect 6678 30280 7104 30308
rect 6678 30277 6690 30280
rect 6632 30271 6690 30277
rect 7098 30268 7104 30280
rect 7156 30268 7162 30320
rect 15120 30308 15148 30348
rect 16206 30336 16212 30348
rect 16264 30336 16270 30388
rect 16666 30376 16672 30388
rect 16627 30348 16672 30376
rect 16666 30336 16672 30348
rect 16724 30336 16730 30388
rect 17494 30336 17500 30388
rect 17552 30376 17558 30388
rect 17865 30379 17923 30385
rect 17865 30376 17877 30379
rect 17552 30348 17877 30376
rect 17552 30336 17558 30348
rect 17865 30345 17877 30348
rect 17911 30345 17923 30379
rect 21266 30376 21272 30388
rect 17865 30339 17923 30345
rect 19168 30348 21272 30376
rect 18322 30308 18328 30320
rect 14200 30280 15148 30308
rect 18283 30280 18328 30308
rect 1949 30243 2007 30249
rect 1949 30209 1961 30243
rect 1995 30240 2007 30243
rect 2130 30240 2136 30252
rect 1995 30212 2136 30240
rect 1995 30209 2007 30212
rect 1949 30203 2007 30209
rect 2130 30200 2136 30212
rect 2188 30200 2194 30252
rect 5629 30243 5687 30249
rect 5629 30209 5641 30243
rect 5675 30240 5687 30243
rect 7190 30240 7196 30252
rect 5675 30212 7196 30240
rect 5675 30209 5687 30212
rect 5629 30203 5687 30209
rect 7190 30200 7196 30212
rect 7248 30200 7254 30252
rect 8665 30243 8723 30249
rect 8665 30209 8677 30243
rect 8711 30240 8723 30243
rect 8754 30240 8760 30252
rect 8711 30212 8760 30240
rect 8711 30209 8723 30212
rect 8665 30203 8723 30209
rect 8754 30200 8760 30212
rect 8812 30200 8818 30252
rect 9585 30243 9643 30249
rect 9585 30209 9597 30243
rect 9631 30240 9643 30243
rect 9674 30240 9680 30252
rect 9631 30212 9680 30240
rect 9631 30209 9643 30212
rect 9585 30203 9643 30209
rect 9674 30200 9680 30212
rect 9732 30200 9738 30252
rect 9858 30249 9864 30252
rect 9852 30203 9864 30249
rect 9916 30240 9922 30252
rect 11793 30243 11851 30249
rect 9916 30212 9952 30240
rect 9858 30200 9864 30203
rect 9916 30200 9922 30212
rect 11793 30209 11805 30243
rect 11839 30240 11851 30243
rect 12066 30240 12072 30252
rect 11839 30212 12072 30240
rect 11839 30209 11851 30212
rect 11793 30203 11851 30209
rect 12066 30200 12072 30212
rect 12124 30240 12130 30252
rect 12345 30243 12403 30249
rect 12345 30240 12357 30243
rect 12124 30212 12357 30240
rect 12124 30200 12130 30212
rect 12345 30209 12357 30212
rect 12391 30209 12403 30243
rect 12345 30203 12403 30209
rect 12621 30243 12679 30249
rect 12621 30209 12633 30243
rect 12667 30240 12679 30243
rect 12710 30240 12716 30252
rect 12667 30212 12716 30240
rect 12667 30209 12679 30212
rect 12621 30203 12679 30209
rect 12710 30200 12716 30212
rect 12768 30240 12774 30252
rect 13722 30240 13728 30252
rect 12768 30212 13728 30240
rect 12768 30200 12774 30212
rect 13722 30200 13728 30212
rect 13780 30200 13786 30252
rect 14090 30200 14096 30252
rect 14148 30240 14154 30252
rect 14200 30249 14228 30280
rect 18322 30268 18328 30280
rect 18380 30268 18386 30320
rect 14185 30243 14243 30249
rect 14185 30240 14197 30243
rect 14148 30212 14197 30240
rect 14148 30200 14154 30212
rect 14185 30209 14197 30212
rect 14231 30209 14243 30243
rect 14185 30203 14243 30209
rect 14452 30243 14510 30249
rect 14452 30209 14464 30243
rect 14498 30240 14510 30243
rect 14734 30240 14740 30252
rect 14498 30212 14740 30240
rect 14498 30209 14510 30212
rect 14452 30203 14510 30209
rect 14734 30200 14740 30212
rect 14792 30200 14798 30252
rect 17037 30243 17095 30249
rect 17037 30209 17049 30243
rect 17083 30240 17095 30243
rect 17310 30240 17316 30252
rect 17083 30212 17316 30240
rect 17083 30209 17095 30212
rect 17037 30203 17095 30209
rect 17310 30200 17316 30212
rect 17368 30200 17374 30252
rect 17402 30200 17408 30252
rect 17460 30240 17466 30252
rect 18233 30243 18291 30249
rect 18233 30240 18245 30243
rect 17460 30212 18245 30240
rect 17460 30200 17466 30212
rect 18233 30209 18245 30212
rect 18279 30209 18291 30243
rect 18233 30203 18291 30209
rect 18690 30200 18696 30252
rect 18748 30240 18754 30252
rect 18966 30240 18972 30252
rect 18748 30212 18972 30240
rect 18748 30200 18754 30212
rect 18966 30200 18972 30212
rect 19024 30240 19030 30252
rect 19168 30249 19196 30348
rect 21266 30336 21272 30348
rect 21324 30336 21330 30388
rect 21836 30348 22094 30376
rect 20714 30268 20720 30320
rect 20772 30308 20778 30320
rect 21836 30317 21864 30348
rect 21821 30311 21879 30317
rect 21821 30308 21833 30311
rect 20772 30280 21833 30308
rect 20772 30268 20778 30280
rect 21821 30277 21833 30280
rect 21867 30277 21879 30311
rect 22066 30308 22094 30348
rect 22066 30280 22508 30308
rect 21821 30271 21879 30277
rect 19153 30243 19211 30249
rect 19153 30240 19165 30243
rect 19024 30212 19165 30240
rect 19024 30200 19030 30212
rect 19153 30209 19165 30212
rect 19199 30209 19211 30243
rect 19978 30240 19984 30252
rect 19939 30212 19984 30240
rect 19153 30203 19211 30209
rect 19978 30200 19984 30212
rect 20036 30200 20042 30252
rect 20257 30243 20315 30249
rect 20257 30209 20269 30243
rect 20303 30240 20315 30243
rect 20530 30240 20536 30252
rect 20303 30212 20536 30240
rect 20303 30209 20315 30212
rect 20257 30203 20315 30209
rect 20530 30200 20536 30212
rect 20588 30200 20594 30252
rect 22005 30243 22063 30249
rect 22005 30240 22017 30243
rect 21836 30212 22017 30240
rect 21836 30184 21864 30212
rect 22005 30209 22017 30212
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 22189 30243 22247 30249
rect 22189 30209 22201 30243
rect 22235 30240 22247 30243
rect 22370 30240 22376 30252
rect 22235 30212 22376 30240
rect 22235 30209 22247 30212
rect 22189 30203 22247 30209
rect 22370 30200 22376 30212
rect 22428 30200 22434 30252
rect 22480 30240 22508 30280
rect 22646 30249 22652 30252
rect 22641 30240 22652 30249
rect 22480 30212 22652 30240
rect 22641 30203 22652 30212
rect 22646 30200 22652 30203
rect 22704 30200 22710 30252
rect 3234 30172 3240 30184
rect 3195 30144 3240 30172
rect 3234 30132 3240 30144
rect 3292 30132 3298 30184
rect 6362 30172 6368 30184
rect 6323 30144 6368 30172
rect 6362 30132 6368 30144
rect 6420 30132 6426 30184
rect 17129 30175 17187 30181
rect 17129 30141 17141 30175
rect 17175 30141 17187 30175
rect 17129 30135 17187 30141
rect 17221 30175 17279 30181
rect 17221 30141 17233 30175
rect 17267 30172 17279 30175
rect 18322 30172 18328 30184
rect 17267 30144 18328 30172
rect 17267 30141 17279 30144
rect 17221 30135 17279 30141
rect 10686 30064 10692 30116
rect 10744 30104 10750 30116
rect 10965 30107 11023 30113
rect 10965 30104 10977 30107
rect 10744 30076 10977 30104
rect 10744 30064 10750 30076
rect 10965 30073 10977 30076
rect 11011 30104 11023 30107
rect 13170 30104 13176 30116
rect 11011 30076 13176 30104
rect 11011 30073 11023 30076
rect 10965 30067 11023 30073
rect 13170 30064 13176 30076
rect 13228 30064 13234 30116
rect 15562 30104 15568 30116
rect 15523 30076 15568 30104
rect 15562 30064 15568 30076
rect 15620 30104 15626 30116
rect 17144 30104 17172 30135
rect 18322 30132 18328 30144
rect 18380 30172 18386 30184
rect 18417 30175 18475 30181
rect 18417 30172 18429 30175
rect 18380 30144 18429 30172
rect 18380 30132 18386 30144
rect 18417 30141 18429 30144
rect 18463 30141 18475 30175
rect 18417 30135 18475 30141
rect 21818 30132 21824 30184
rect 21876 30132 21882 30184
rect 15620 30076 17172 30104
rect 15620 30064 15626 30076
rect 17770 30064 17776 30116
rect 17828 30104 17834 30116
rect 18874 30104 18880 30116
rect 17828 30076 18880 30104
rect 17828 30064 17834 30076
rect 18874 30064 18880 30076
rect 18932 30104 18938 30116
rect 19337 30107 19395 30113
rect 19337 30104 19349 30107
rect 18932 30076 19349 30104
rect 18932 30064 18938 30076
rect 19337 30073 19349 30076
rect 19383 30073 19395 30107
rect 19337 30067 19395 30073
rect 2314 30036 2320 30048
rect 2275 30008 2320 30036
rect 2314 29996 2320 30008
rect 2372 29996 2378 30048
rect 2498 30036 2504 30048
rect 2459 30008 2504 30036
rect 2498 29996 2504 30008
rect 2556 29996 2562 30048
rect 5810 30036 5816 30048
rect 5771 30008 5816 30036
rect 5810 29996 5816 30008
rect 5868 29996 5874 30048
rect 8202 30036 8208 30048
rect 8163 30008 8208 30036
rect 8202 29996 8208 30008
rect 8260 29996 8266 30048
rect 8570 30036 8576 30048
rect 8531 30008 8576 30036
rect 8570 29996 8576 30008
rect 8628 29996 8634 30048
rect 11606 29996 11612 30048
rect 11664 30036 11670 30048
rect 11701 30039 11759 30045
rect 11701 30036 11713 30039
rect 11664 30008 11713 30036
rect 11664 29996 11670 30008
rect 11701 30005 11713 30008
rect 11747 30036 11759 30039
rect 13078 30036 13084 30048
rect 11747 30008 13084 30036
rect 11747 30005 11759 30008
rect 11701 29999 11759 30005
rect 13078 29996 13084 30008
rect 13136 29996 13142 30048
rect 22002 29996 22008 30048
rect 22060 30036 22066 30048
rect 22186 30036 22192 30048
rect 22060 30008 22192 30036
rect 22060 29996 22066 30008
rect 22186 29996 22192 30008
rect 22244 30036 22250 30048
rect 22741 30039 22799 30045
rect 22741 30036 22753 30039
rect 22244 30008 22753 30036
rect 22244 29996 22250 30008
rect 22741 30005 22753 30008
rect 22787 30005 22799 30039
rect 22741 29999 22799 30005
rect 1104 29946 30820 29968
rect 1104 29894 5915 29946
rect 5967 29894 5979 29946
rect 6031 29894 6043 29946
rect 6095 29894 6107 29946
rect 6159 29894 6171 29946
rect 6223 29894 15846 29946
rect 15898 29894 15910 29946
rect 15962 29894 15974 29946
rect 16026 29894 16038 29946
rect 16090 29894 16102 29946
rect 16154 29894 25776 29946
rect 25828 29894 25840 29946
rect 25892 29894 25904 29946
rect 25956 29894 25968 29946
rect 26020 29894 26032 29946
rect 26084 29894 30820 29946
rect 1104 29872 30820 29894
rect 2314 29792 2320 29844
rect 2372 29832 2378 29844
rect 2409 29835 2467 29841
rect 2409 29832 2421 29835
rect 2372 29804 2421 29832
rect 2372 29792 2378 29804
rect 2409 29801 2421 29804
rect 2455 29801 2467 29835
rect 2409 29795 2467 29801
rect 2593 29835 2651 29841
rect 2593 29801 2605 29835
rect 2639 29832 2651 29835
rect 2958 29832 2964 29844
rect 2639 29804 2964 29832
rect 2639 29801 2651 29804
rect 2593 29795 2651 29801
rect 2041 29767 2099 29773
rect 2041 29733 2053 29767
rect 2087 29764 2099 29767
rect 2130 29764 2136 29776
rect 2087 29736 2136 29764
rect 2087 29733 2099 29736
rect 2041 29727 2099 29733
rect 2130 29724 2136 29736
rect 2188 29724 2194 29776
rect 2424 29764 2452 29795
rect 2958 29792 2964 29804
rect 3016 29792 3022 29844
rect 6181 29835 6239 29841
rect 6181 29801 6193 29835
rect 6227 29832 6239 29835
rect 6362 29832 6368 29844
rect 6227 29804 6368 29832
rect 6227 29801 6239 29804
rect 6181 29795 6239 29801
rect 6362 29792 6368 29804
rect 6420 29792 6426 29844
rect 6638 29792 6644 29844
rect 6696 29832 6702 29844
rect 7377 29835 7435 29841
rect 7377 29832 7389 29835
rect 6696 29804 7389 29832
rect 6696 29792 6702 29804
rect 7377 29801 7389 29804
rect 7423 29832 7435 29835
rect 8846 29832 8852 29844
rect 7423 29804 8852 29832
rect 7423 29801 7435 29804
rect 7377 29795 7435 29801
rect 8846 29792 8852 29804
rect 8904 29792 8910 29844
rect 10689 29835 10747 29841
rect 10689 29801 10701 29835
rect 10735 29832 10747 29835
rect 10778 29832 10784 29844
rect 10735 29804 10784 29832
rect 10735 29801 10747 29804
rect 10689 29795 10747 29801
rect 10778 29792 10784 29804
rect 10836 29792 10842 29844
rect 11057 29835 11115 29841
rect 11057 29801 11069 29835
rect 11103 29832 11115 29835
rect 11330 29832 11336 29844
rect 11103 29804 11336 29832
rect 11103 29801 11115 29804
rect 11057 29795 11115 29801
rect 11330 29792 11336 29804
rect 11388 29792 11394 29844
rect 17126 29792 17132 29844
rect 17184 29832 17190 29844
rect 17497 29835 17555 29841
rect 17497 29832 17509 29835
rect 17184 29804 17509 29832
rect 17184 29792 17190 29804
rect 17497 29801 17509 29804
rect 17543 29801 17555 29835
rect 17497 29795 17555 29801
rect 18414 29792 18420 29844
rect 18472 29832 18478 29844
rect 18472 29804 21404 29832
rect 18472 29792 18478 29804
rect 2866 29764 2872 29776
rect 2424 29736 2872 29764
rect 2866 29724 2872 29736
rect 2924 29724 2930 29776
rect 15102 29724 15108 29776
rect 15160 29764 15166 29776
rect 15160 29736 18000 29764
rect 15160 29724 15166 29736
rect 2498 29696 2504 29708
rect 1412 29668 2504 29696
rect 1412 29637 1440 29668
rect 2498 29656 2504 29668
rect 2556 29656 2562 29708
rect 10597 29699 10655 29705
rect 10597 29665 10609 29699
rect 10643 29696 10655 29699
rect 11422 29696 11428 29708
rect 10643 29668 11428 29696
rect 10643 29665 10655 29668
rect 10597 29659 10655 29665
rect 11422 29656 11428 29668
rect 11480 29696 11486 29708
rect 11606 29696 11612 29708
rect 11480 29668 11612 29696
rect 11480 29656 11486 29668
rect 11606 29656 11612 29668
rect 11664 29656 11670 29708
rect 14090 29696 14096 29708
rect 14051 29668 14096 29696
rect 14090 29656 14096 29668
rect 14148 29656 14154 29708
rect 16945 29699 17003 29705
rect 16945 29665 16957 29699
rect 16991 29696 17003 29699
rect 16991 29668 17724 29696
rect 16991 29665 17003 29668
rect 16945 29659 17003 29665
rect 1397 29631 1455 29637
rect 1397 29597 1409 29631
rect 1443 29597 1455 29631
rect 1397 29591 1455 29597
rect 3053 29631 3111 29637
rect 3053 29597 3065 29631
rect 3099 29628 3111 29631
rect 3970 29628 3976 29640
rect 3099 29600 3976 29628
rect 3099 29597 3111 29600
rect 3053 29591 3111 29597
rect 3970 29588 3976 29600
rect 4028 29588 4034 29640
rect 4154 29628 4160 29640
rect 4115 29600 4160 29628
rect 4154 29588 4160 29600
rect 4212 29588 4218 29640
rect 4424 29631 4482 29637
rect 4424 29597 4436 29631
rect 4470 29628 4482 29631
rect 4706 29628 4712 29640
rect 4470 29600 4712 29628
rect 4470 29597 4482 29600
rect 4424 29591 4482 29597
rect 4706 29588 4712 29600
rect 4764 29588 4770 29640
rect 5258 29588 5264 29640
rect 5316 29628 5322 29640
rect 5997 29631 6055 29637
rect 5997 29628 6009 29631
rect 5316 29600 6009 29628
rect 5316 29588 5322 29600
rect 5997 29597 6009 29600
rect 6043 29597 6055 29631
rect 5997 29591 6055 29597
rect 8205 29631 8263 29637
rect 8205 29597 8217 29631
rect 8251 29628 8263 29631
rect 8938 29628 8944 29640
rect 8251 29600 8944 29628
rect 8251 29597 8263 29600
rect 8205 29591 8263 29597
rect 8938 29588 8944 29600
rect 8996 29588 9002 29640
rect 9677 29631 9735 29637
rect 9677 29597 9689 29631
rect 9723 29628 9735 29631
rect 9766 29628 9772 29640
rect 9723 29600 9772 29628
rect 9723 29597 9735 29600
rect 9677 29591 9735 29597
rect 9766 29588 9772 29600
rect 9824 29588 9830 29640
rect 9950 29588 9956 29640
rect 10008 29628 10014 29640
rect 10873 29631 10931 29637
rect 10873 29628 10885 29631
rect 10008 29600 10885 29628
rect 10008 29588 10014 29600
rect 10873 29597 10885 29600
rect 10919 29597 10931 29631
rect 10873 29591 10931 29597
rect 12526 29588 12532 29640
rect 12584 29628 12590 29640
rect 12621 29631 12679 29637
rect 12621 29628 12633 29631
rect 12584 29600 12633 29628
rect 12584 29588 12590 29600
rect 12621 29597 12633 29600
rect 12667 29597 12679 29631
rect 12621 29591 12679 29597
rect 12802 29588 12808 29640
rect 12860 29628 12866 29640
rect 12897 29631 12955 29637
rect 12897 29628 12909 29631
rect 12860 29600 12909 29628
rect 12860 29588 12866 29600
rect 12897 29597 12909 29600
rect 12943 29597 12955 29631
rect 12897 29591 12955 29597
rect 16301 29631 16359 29637
rect 16301 29597 16313 29631
rect 16347 29628 16359 29631
rect 17310 29628 17316 29640
rect 16347 29600 17316 29628
rect 16347 29597 16359 29600
rect 16301 29591 16359 29597
rect 17310 29588 17316 29600
rect 17368 29588 17374 29640
rect 2409 29563 2467 29569
rect 2409 29529 2421 29563
rect 2455 29560 2467 29563
rect 4890 29560 4896 29572
rect 2455 29532 4896 29560
rect 2455 29529 2467 29532
rect 2409 29523 2467 29529
rect 4890 29520 4896 29532
rect 4948 29560 4954 29572
rect 4948 29532 5580 29560
rect 4948 29520 4954 29532
rect 1581 29495 1639 29501
rect 1581 29461 1593 29495
rect 1627 29492 1639 29495
rect 2130 29492 2136 29504
rect 1627 29464 2136 29492
rect 1627 29461 1639 29464
rect 1581 29455 1639 29461
rect 2130 29452 2136 29464
rect 2188 29452 2194 29504
rect 3237 29495 3295 29501
rect 3237 29461 3249 29495
rect 3283 29492 3295 29495
rect 3602 29492 3608 29504
rect 3283 29464 3608 29492
rect 3283 29461 3295 29464
rect 3237 29455 3295 29461
rect 3602 29452 3608 29464
rect 3660 29452 3666 29504
rect 5552 29501 5580 29532
rect 6546 29520 6552 29572
rect 6604 29560 6610 29572
rect 7285 29563 7343 29569
rect 7285 29560 7297 29563
rect 6604 29532 7297 29560
rect 6604 29520 6610 29532
rect 7285 29529 7297 29532
rect 7331 29529 7343 29563
rect 12066 29560 12072 29572
rect 12027 29532 12072 29560
rect 7285 29523 7343 29529
rect 12066 29520 12072 29532
rect 12124 29520 12130 29572
rect 13170 29520 13176 29572
rect 13228 29560 13234 29572
rect 14338 29563 14396 29569
rect 14338 29560 14350 29563
rect 13228 29532 14350 29560
rect 13228 29520 13234 29532
rect 14338 29529 14350 29532
rect 14384 29529 14396 29563
rect 14338 29523 14396 29529
rect 16209 29563 16267 29569
rect 16209 29529 16221 29563
rect 16255 29560 16267 29563
rect 17696 29560 17724 29668
rect 17972 29637 18000 29736
rect 18322 29724 18328 29776
rect 18380 29764 18386 29776
rect 20530 29764 20536 29776
rect 18380 29736 20536 29764
rect 18380 29724 18386 29736
rect 20530 29724 20536 29736
rect 20588 29724 20594 29776
rect 20622 29724 20628 29776
rect 20680 29764 20686 29776
rect 21376 29773 21404 29804
rect 21542 29792 21548 29844
rect 21600 29832 21606 29844
rect 21600 29804 22094 29832
rect 21600 29792 21606 29804
rect 21361 29767 21419 29773
rect 20680 29736 21220 29764
rect 20680 29724 20686 29736
rect 19886 29656 19892 29708
rect 19944 29696 19950 29708
rect 19944 29668 21128 29696
rect 19944 29656 19950 29668
rect 17957 29631 18015 29637
rect 17957 29597 17969 29631
rect 18003 29628 18015 29631
rect 19334 29628 19340 29640
rect 18003 29600 19340 29628
rect 18003 29597 18015 29600
rect 17957 29591 18015 29597
rect 19334 29588 19340 29600
rect 19392 29588 19398 29640
rect 19978 29628 19984 29640
rect 19939 29600 19984 29628
rect 19978 29588 19984 29600
rect 20036 29588 20042 29640
rect 20349 29631 20407 29637
rect 20349 29597 20361 29631
rect 20395 29628 20407 29631
rect 20714 29628 20720 29640
rect 20395 29600 20720 29628
rect 20395 29597 20407 29600
rect 20349 29591 20407 29597
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 18322 29560 18328 29572
rect 16255 29532 17172 29560
rect 17696 29532 18328 29560
rect 16255 29529 16267 29532
rect 16209 29523 16267 29529
rect 5537 29495 5595 29501
rect 5537 29461 5549 29495
rect 5583 29461 5595 29495
rect 5537 29455 5595 29461
rect 7650 29452 7656 29504
rect 7708 29492 7714 29504
rect 8021 29495 8079 29501
rect 8021 29492 8033 29495
rect 7708 29464 8033 29492
rect 7708 29452 7714 29464
rect 8021 29461 8033 29464
rect 8067 29461 8079 29495
rect 8021 29455 8079 29461
rect 9122 29452 9128 29504
rect 9180 29492 9186 29504
rect 9493 29495 9551 29501
rect 9493 29492 9505 29495
rect 9180 29464 9505 29492
rect 9180 29452 9186 29464
rect 9493 29461 9505 29464
rect 9539 29461 9551 29495
rect 9493 29455 9551 29461
rect 11698 29452 11704 29504
rect 11756 29492 11762 29504
rect 11974 29492 11980 29504
rect 11756 29464 11980 29492
rect 11756 29452 11762 29464
rect 11974 29452 11980 29464
rect 12032 29452 12038 29504
rect 15470 29492 15476 29504
rect 15431 29464 15476 29492
rect 15470 29452 15476 29464
rect 15528 29452 15534 29504
rect 16942 29452 16948 29504
rect 17000 29492 17006 29504
rect 17144 29501 17172 29532
rect 18322 29520 18328 29532
rect 18380 29520 18386 29572
rect 19797 29563 19855 29569
rect 19797 29529 19809 29563
rect 19843 29560 19855 29563
rect 20254 29560 20260 29572
rect 19843 29532 20260 29560
rect 19843 29529 19855 29532
rect 19797 29523 19855 29529
rect 20254 29520 20260 29532
rect 20312 29520 20318 29572
rect 20530 29520 20536 29572
rect 20588 29560 20594 29572
rect 20809 29563 20867 29569
rect 20809 29560 20821 29563
rect 20588 29532 20821 29560
rect 20588 29520 20594 29532
rect 20809 29529 20821 29532
rect 20855 29529 20867 29563
rect 20809 29523 20867 29529
rect 17037 29495 17095 29501
rect 17037 29492 17049 29495
rect 17000 29464 17049 29492
rect 17000 29452 17006 29464
rect 17037 29461 17049 29464
rect 17083 29461 17095 29495
rect 17037 29455 17095 29461
rect 17129 29495 17187 29501
rect 17129 29461 17141 29495
rect 17175 29492 17187 29495
rect 17402 29492 17408 29504
rect 17175 29464 17408 29492
rect 17175 29461 17187 29464
rect 17129 29455 17187 29461
rect 17402 29452 17408 29464
rect 17460 29452 17466 29504
rect 17954 29452 17960 29504
rect 18012 29492 18018 29504
rect 18141 29495 18199 29501
rect 18141 29492 18153 29495
rect 18012 29464 18153 29492
rect 18012 29452 18018 29464
rect 18141 29461 18153 29464
rect 18187 29492 18199 29495
rect 18230 29492 18236 29504
rect 18187 29464 18236 29492
rect 18187 29461 18199 29464
rect 18141 29455 18199 29461
rect 18230 29452 18236 29464
rect 18288 29452 18294 29504
rect 19886 29452 19892 29504
rect 19944 29492 19950 29504
rect 20073 29495 20131 29501
rect 20073 29492 20085 29495
rect 19944 29464 20085 29492
rect 19944 29452 19950 29464
rect 20073 29461 20085 29464
rect 20119 29461 20131 29495
rect 20073 29455 20131 29461
rect 20162 29452 20168 29504
rect 20220 29492 20226 29504
rect 21100 29501 21128 29668
rect 21192 29637 21220 29736
rect 21361 29733 21373 29767
rect 21407 29733 21419 29767
rect 22066 29764 22094 29804
rect 22066 29736 22140 29764
rect 21361 29727 21419 29733
rect 22112 29705 22140 29736
rect 22097 29699 22155 29705
rect 22097 29665 22109 29699
rect 22143 29665 22155 29699
rect 22097 29659 22155 29665
rect 21177 29631 21235 29637
rect 21177 29597 21189 29631
rect 21223 29597 21235 29631
rect 21818 29628 21824 29640
rect 21779 29600 21824 29628
rect 21177 29591 21235 29597
rect 21818 29588 21824 29600
rect 21876 29588 21882 29640
rect 22189 29631 22247 29637
rect 22189 29597 22201 29631
rect 22235 29628 22247 29631
rect 29730 29628 29736 29640
rect 22235 29600 29736 29628
rect 22235 29597 22247 29600
rect 22189 29591 22247 29597
rect 29730 29588 29736 29600
rect 29788 29588 29794 29640
rect 22094 29520 22100 29572
rect 22152 29560 22158 29572
rect 22306 29563 22364 29569
rect 22306 29560 22318 29563
rect 22152 29532 22318 29560
rect 22152 29520 22158 29532
rect 22306 29529 22318 29532
rect 22352 29529 22364 29563
rect 22306 29523 22364 29529
rect 20993 29495 21051 29501
rect 20993 29492 21005 29495
rect 20220 29464 21005 29492
rect 20220 29452 20226 29464
rect 20993 29461 21005 29464
rect 21039 29461 21051 29495
rect 20993 29455 21051 29461
rect 21085 29495 21143 29501
rect 21085 29461 21097 29495
rect 21131 29461 21143 29495
rect 22462 29492 22468 29504
rect 22423 29464 22468 29492
rect 21085 29455 21143 29461
rect 22462 29452 22468 29464
rect 22520 29452 22526 29504
rect 1104 29402 30820 29424
rect 1104 29350 10880 29402
rect 10932 29350 10944 29402
rect 10996 29350 11008 29402
rect 11060 29350 11072 29402
rect 11124 29350 11136 29402
rect 11188 29350 20811 29402
rect 20863 29350 20875 29402
rect 20927 29350 20939 29402
rect 20991 29350 21003 29402
rect 21055 29350 21067 29402
rect 21119 29350 30820 29402
rect 1104 29328 30820 29350
rect 2317 29291 2375 29297
rect 2317 29257 2329 29291
rect 2363 29288 2375 29291
rect 2774 29288 2780 29300
rect 2363 29260 2780 29288
rect 2363 29257 2375 29260
rect 2317 29251 2375 29257
rect 2774 29248 2780 29260
rect 2832 29248 2838 29300
rect 3234 29248 3240 29300
rect 3292 29288 3298 29300
rect 3421 29291 3479 29297
rect 3421 29288 3433 29291
rect 3292 29260 3433 29288
rect 3292 29248 3298 29260
rect 3421 29257 3433 29260
rect 3467 29257 3479 29291
rect 5258 29288 5264 29300
rect 5219 29260 5264 29288
rect 3421 29251 3479 29257
rect 5258 29248 5264 29260
rect 5316 29248 5322 29300
rect 8570 29248 8576 29300
rect 8628 29288 8634 29300
rect 8757 29291 8815 29297
rect 8757 29288 8769 29291
rect 8628 29260 8769 29288
rect 8628 29248 8634 29260
rect 8757 29257 8769 29260
rect 8803 29257 8815 29291
rect 9122 29288 9128 29300
rect 9083 29260 9128 29288
rect 8757 29251 8815 29257
rect 9122 29248 9128 29260
rect 9180 29248 9186 29300
rect 11885 29291 11943 29297
rect 11885 29257 11897 29291
rect 11931 29288 11943 29291
rect 12066 29288 12072 29300
rect 11931 29260 12072 29288
rect 11931 29257 11943 29260
rect 11885 29251 11943 29257
rect 12066 29248 12072 29260
rect 12124 29248 12130 29300
rect 13170 29288 13176 29300
rect 13131 29260 13176 29288
rect 13170 29248 13176 29260
rect 13228 29248 13234 29300
rect 14642 29288 14648 29300
rect 14603 29260 14648 29288
rect 14642 29248 14648 29260
rect 14700 29248 14706 29300
rect 17126 29288 17132 29300
rect 17039 29260 17132 29288
rect 12621 29223 12679 29229
rect 12621 29189 12633 29223
rect 12667 29220 12679 29223
rect 12710 29220 12716 29232
rect 12667 29192 12716 29220
rect 12667 29189 12679 29192
rect 12621 29183 12679 29189
rect 12710 29180 12716 29192
rect 12768 29180 12774 29232
rect 13541 29223 13599 29229
rect 13541 29189 13553 29223
rect 13587 29220 13599 29223
rect 15470 29220 15476 29232
rect 13587 29192 15476 29220
rect 13587 29189 13599 29192
rect 13541 29183 13599 29189
rect 15470 29180 15476 29192
rect 15528 29220 15534 29232
rect 16025 29223 16083 29229
rect 15528 29192 15976 29220
rect 15528 29180 15534 29192
rect 1673 29155 1731 29161
rect 1673 29121 1685 29155
rect 1719 29121 1731 29155
rect 2130 29152 2136 29164
rect 2091 29124 2136 29152
rect 1673 29115 1731 29121
rect 1688 29084 1716 29115
rect 2130 29112 2136 29124
rect 2188 29112 2194 29164
rect 3602 29152 3608 29164
rect 3563 29124 3608 29152
rect 3602 29112 3608 29124
rect 3660 29112 3666 29164
rect 4062 29112 4068 29164
rect 4120 29152 4126 29164
rect 4249 29155 4307 29161
rect 4249 29152 4261 29155
rect 4120 29124 4261 29152
rect 4120 29112 4126 29124
rect 4249 29121 4261 29124
rect 4295 29152 4307 29155
rect 5077 29155 5135 29161
rect 5077 29152 5089 29155
rect 4295 29124 5089 29152
rect 4295 29121 4307 29124
rect 4249 29115 4307 29121
rect 5077 29121 5089 29124
rect 5123 29121 5135 29155
rect 7006 29152 7012 29164
rect 6967 29124 7012 29152
rect 5077 29115 5135 29121
rect 7006 29112 7012 29124
rect 7064 29112 7070 29164
rect 8021 29155 8079 29161
rect 8021 29121 8033 29155
rect 8067 29152 8079 29155
rect 8202 29152 8208 29164
rect 8067 29124 8208 29152
rect 8067 29121 8079 29124
rect 8021 29115 8079 29121
rect 8202 29112 8208 29124
rect 8260 29112 8266 29164
rect 9048 29124 9352 29152
rect 4706 29084 4712 29096
rect 1688 29056 4712 29084
rect 4706 29044 4712 29056
rect 4764 29044 4770 29096
rect 5534 29044 5540 29096
rect 5592 29084 5598 29096
rect 7101 29087 7159 29093
rect 7101 29084 7113 29087
rect 5592 29056 7113 29084
rect 5592 29044 5598 29056
rect 7101 29053 7113 29056
rect 7147 29053 7159 29087
rect 7101 29047 7159 29053
rect 7190 29044 7196 29096
rect 7248 29084 7254 29096
rect 9048 29084 9076 29124
rect 9214 29084 9220 29096
rect 7248 29056 9076 29084
rect 9175 29056 9220 29084
rect 7248 29044 7254 29056
rect 9214 29044 9220 29056
rect 9272 29044 9278 29096
rect 9324 29093 9352 29124
rect 10042 29112 10048 29164
rect 10100 29152 10106 29164
rect 10137 29155 10195 29161
rect 10137 29152 10149 29155
rect 10100 29124 10149 29152
rect 10100 29112 10106 29124
rect 10137 29121 10149 29124
rect 10183 29121 10195 29155
rect 10137 29115 10195 29121
rect 11977 29155 12035 29161
rect 11977 29121 11989 29155
rect 12023 29152 12035 29155
rect 12023 29124 12434 29152
rect 12023 29121 12035 29124
rect 11977 29115 12035 29121
rect 9309 29087 9367 29093
rect 9309 29053 9321 29087
rect 9355 29053 9367 29087
rect 12406 29084 12434 29124
rect 12526 29112 12532 29164
rect 12584 29112 12590 29164
rect 12728 29152 12756 29180
rect 13311 29155 13369 29161
rect 13311 29152 13323 29155
rect 12728 29124 13323 29152
rect 13311 29121 13323 29124
rect 13357 29121 13369 29155
rect 13311 29115 13369 29121
rect 13446 29112 13452 29164
rect 13504 29152 13510 29164
rect 13669 29155 13727 29161
rect 13669 29152 13681 29155
rect 13504 29124 13549 29152
rect 13504 29112 13510 29124
rect 13648 29121 13681 29152
rect 13715 29121 13727 29155
rect 13648 29115 13727 29121
rect 13817 29155 13875 29161
rect 13817 29121 13829 29155
rect 13863 29121 13875 29155
rect 14734 29152 14740 29164
rect 14695 29124 14740 29152
rect 13817 29115 13875 29121
rect 12544 29084 12572 29112
rect 12406 29056 12756 29084
rect 9309 29047 9367 29053
rect 1486 29016 1492 29028
rect 1447 28988 1492 29016
rect 1486 28976 1492 28988
rect 1544 28976 1550 29028
rect 7834 29016 7840 29028
rect 7795 28988 7840 29016
rect 7834 28976 7840 28988
rect 7892 28976 7898 29028
rect 8386 28976 8392 29028
rect 8444 29016 8450 29028
rect 9953 29019 10011 29025
rect 9953 29016 9965 29019
rect 8444 28988 9965 29016
rect 8444 28976 8450 28988
rect 9953 28985 9965 28988
rect 9999 28985 10011 29019
rect 9953 28979 10011 28985
rect 12437 29019 12495 29025
rect 12437 28985 12449 29019
rect 12483 29016 12495 29019
rect 12526 29016 12532 29028
rect 12483 28988 12532 29016
rect 12483 28985 12495 28988
rect 12437 28979 12495 28985
rect 12526 28976 12532 28988
rect 12584 28976 12590 29028
rect 12728 29016 12756 29056
rect 12802 29044 12808 29096
rect 12860 29084 12866 29096
rect 13648 29084 13676 29115
rect 12860 29056 13676 29084
rect 13832 29084 13860 29115
rect 14734 29112 14740 29124
rect 14792 29112 14798 29164
rect 15948 29161 15976 29192
rect 16025 29189 16037 29223
rect 16071 29220 16083 29223
rect 16942 29220 16948 29232
rect 16071 29192 16948 29220
rect 16071 29189 16083 29192
rect 16025 29183 16083 29189
rect 16942 29180 16948 29192
rect 17000 29180 17006 29232
rect 15933 29155 15991 29161
rect 15933 29121 15945 29155
rect 15979 29121 15991 29155
rect 16666 29152 16672 29164
rect 16627 29124 16672 29152
rect 15933 29115 15991 29121
rect 16666 29112 16672 29124
rect 16724 29112 16730 29164
rect 16850 29152 16856 29164
rect 16811 29124 16856 29152
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 17052 29161 17080 29260
rect 17126 29248 17132 29260
rect 17184 29288 17190 29300
rect 20993 29291 21051 29297
rect 17184 29260 18368 29288
rect 17184 29248 17190 29260
rect 17402 29180 17408 29232
rect 17460 29220 17466 29232
rect 18340 29220 18368 29260
rect 20993 29257 21005 29291
rect 21039 29288 21051 29291
rect 21818 29288 21824 29300
rect 21039 29260 21824 29288
rect 21039 29257 21051 29260
rect 20993 29251 21051 29257
rect 21818 29248 21824 29260
rect 21876 29248 21882 29300
rect 22373 29291 22431 29297
rect 22373 29257 22385 29291
rect 22419 29257 22431 29291
rect 22373 29251 22431 29257
rect 21542 29220 21548 29232
rect 17460 29192 18276 29220
rect 18340 29192 21548 29220
rect 17460 29180 17466 29192
rect 17037 29155 17095 29161
rect 17037 29121 17049 29155
rect 17083 29121 17095 29155
rect 17218 29152 17224 29164
rect 17179 29124 17224 29152
rect 17037 29115 17095 29121
rect 17218 29112 17224 29124
rect 17276 29112 17282 29164
rect 17770 29152 17776 29164
rect 17328 29124 17776 29152
rect 13998 29084 14004 29096
rect 13832 29056 14004 29084
rect 12860 29044 12866 29056
rect 13998 29044 14004 29056
rect 14056 29084 14062 29096
rect 15102 29084 15108 29096
rect 14056 29056 15108 29084
rect 14056 29044 14062 29056
rect 15102 29044 15108 29056
rect 15160 29044 15166 29096
rect 16945 29087 17003 29093
rect 16945 29053 16957 29087
rect 16991 29084 17003 29087
rect 17328 29084 17356 29124
rect 17770 29112 17776 29124
rect 17828 29112 17834 29164
rect 18046 29152 18052 29164
rect 18007 29124 18052 29152
rect 18046 29112 18052 29124
rect 18104 29112 18110 29164
rect 18248 29161 18276 29192
rect 21542 29180 21548 29192
rect 21600 29180 21606 29232
rect 22388 29220 22416 29251
rect 23078 29223 23136 29229
rect 23078 29220 23090 29223
rect 22388 29192 23090 29220
rect 23078 29189 23090 29192
rect 23124 29189 23136 29223
rect 23078 29183 23136 29189
rect 18233 29155 18291 29161
rect 18233 29121 18245 29155
rect 18279 29121 18291 29155
rect 18233 29115 18291 29121
rect 18322 29112 18328 29164
rect 18380 29152 18386 29164
rect 18380 29124 18425 29152
rect 18380 29112 18386 29124
rect 20162 29112 20168 29164
rect 20220 29152 20226 29164
rect 20717 29155 20775 29161
rect 20717 29152 20729 29155
rect 20220 29124 20729 29152
rect 20220 29112 20226 29124
rect 20717 29121 20729 29124
rect 20763 29121 20775 29155
rect 20717 29115 20775 29121
rect 22189 29155 22247 29161
rect 22189 29121 22201 29155
rect 22235 29152 22247 29155
rect 22462 29152 22468 29164
rect 22235 29124 22468 29152
rect 22235 29121 22247 29124
rect 22189 29115 22247 29121
rect 22462 29112 22468 29124
rect 22520 29112 22526 29164
rect 22554 29112 22560 29164
rect 22612 29152 22618 29164
rect 22833 29155 22891 29161
rect 22833 29152 22845 29155
rect 22612 29124 22845 29152
rect 22612 29112 22618 29124
rect 22833 29121 22845 29124
rect 22879 29121 22891 29155
rect 22833 29115 22891 29121
rect 29825 29155 29883 29161
rect 29825 29121 29837 29155
rect 29871 29152 29883 29155
rect 30190 29152 30196 29164
rect 29871 29124 30196 29152
rect 29871 29121 29883 29124
rect 29825 29115 29883 29121
rect 30190 29112 30196 29124
rect 30248 29112 30254 29164
rect 16991 29056 17356 29084
rect 17405 29087 17463 29093
rect 16991 29053 17003 29056
rect 16945 29047 17003 29053
rect 17405 29053 17417 29087
rect 17451 29084 17463 29087
rect 17957 29087 18015 29093
rect 17957 29084 17969 29087
rect 17451 29056 17969 29084
rect 17451 29053 17463 29056
rect 17405 29047 17463 29053
rect 17957 29053 17969 29056
rect 18003 29053 18015 29087
rect 20530 29084 20536 29096
rect 20491 29056 20536 29084
rect 17957 29047 18015 29053
rect 20530 29044 20536 29056
rect 20588 29044 20594 29096
rect 20622 29044 20628 29096
rect 20680 29084 20686 29096
rect 20809 29087 20867 29093
rect 20680 29056 20725 29084
rect 20680 29044 20686 29056
rect 20809 29053 20821 29087
rect 20855 29084 20867 29087
rect 21450 29084 21456 29096
rect 20855 29056 21456 29084
rect 20855 29053 20867 29056
rect 20809 29047 20867 29053
rect 21450 29044 21456 29056
rect 21508 29084 21514 29096
rect 21726 29084 21732 29096
rect 21508 29056 21732 29084
rect 21508 29044 21514 29056
rect 21726 29044 21732 29056
rect 21784 29044 21790 29096
rect 13170 29016 13176 29028
rect 12728 28988 13176 29016
rect 13170 28976 13176 28988
rect 13228 28976 13234 29028
rect 17862 29016 17868 29028
rect 17823 28988 17868 29016
rect 17862 28976 17868 28988
rect 17920 28976 17926 29028
rect 24213 29019 24271 29025
rect 24213 28985 24225 29019
rect 24259 29016 24271 29019
rect 29822 29016 29828 29028
rect 24259 28988 29828 29016
rect 24259 28985 24271 28988
rect 24213 28979 24271 28985
rect 29822 28976 29828 28988
rect 29880 28976 29886 29028
rect 30006 29016 30012 29028
rect 29967 28988 30012 29016
rect 30006 28976 30012 28988
rect 30064 28976 30070 29028
rect 3786 28908 3792 28960
rect 3844 28948 3850 28960
rect 4065 28951 4123 28957
rect 4065 28948 4077 28951
rect 3844 28920 4077 28948
rect 3844 28908 3850 28920
rect 4065 28917 4077 28920
rect 4111 28917 4123 28951
rect 6638 28948 6644 28960
rect 6599 28920 6644 28948
rect 4065 28911 4123 28917
rect 6638 28908 6644 28920
rect 6696 28908 6702 28960
rect 1104 28858 30820 28880
rect 1104 28806 5915 28858
rect 5967 28806 5979 28858
rect 6031 28806 6043 28858
rect 6095 28806 6107 28858
rect 6159 28806 6171 28858
rect 6223 28806 15846 28858
rect 15898 28806 15910 28858
rect 15962 28806 15974 28858
rect 16026 28806 16038 28858
rect 16090 28806 16102 28858
rect 16154 28806 25776 28858
rect 25828 28806 25840 28858
rect 25892 28806 25904 28858
rect 25956 28806 25968 28858
rect 26020 28806 26032 28858
rect 26084 28806 30820 28858
rect 1104 28784 30820 28806
rect 3973 28747 4031 28753
rect 3973 28713 3985 28747
rect 4019 28744 4031 28747
rect 4154 28744 4160 28756
rect 4019 28716 4160 28744
rect 4019 28713 4031 28716
rect 3973 28707 4031 28713
rect 4154 28704 4160 28716
rect 4212 28704 4218 28756
rect 5169 28747 5227 28753
rect 5169 28713 5181 28747
rect 5215 28744 5227 28747
rect 5534 28744 5540 28756
rect 5215 28716 5540 28744
rect 5215 28713 5227 28716
rect 5169 28707 5227 28713
rect 5534 28704 5540 28716
rect 5592 28704 5598 28756
rect 5813 28747 5871 28753
rect 5813 28713 5825 28747
rect 5859 28744 5871 28747
rect 7006 28744 7012 28756
rect 5859 28716 7012 28744
rect 5859 28713 5871 28716
rect 5813 28707 5871 28713
rect 7006 28704 7012 28716
rect 7064 28704 7070 28756
rect 11330 28744 11336 28756
rect 11243 28716 11336 28744
rect 11330 28704 11336 28716
rect 11388 28744 11394 28756
rect 12618 28744 12624 28756
rect 11388 28716 12624 28744
rect 11388 28704 11394 28716
rect 12618 28704 12624 28716
rect 12676 28704 12682 28756
rect 14642 28744 14648 28756
rect 12820 28716 14648 28744
rect 7558 28676 7564 28688
rect 5644 28648 7564 28676
rect 2685 28611 2743 28617
rect 2685 28608 2697 28611
rect 1688 28580 2697 28608
rect 1688 28549 1716 28580
rect 2685 28577 2697 28580
rect 2731 28577 2743 28611
rect 2685 28571 2743 28577
rect 1673 28543 1731 28549
rect 1673 28509 1685 28543
rect 1719 28509 1731 28543
rect 2590 28540 2596 28552
rect 2551 28512 2596 28540
rect 1673 28503 1731 28509
rect 2590 28500 2596 28512
rect 2648 28500 2654 28552
rect 2777 28543 2835 28549
rect 2777 28509 2789 28543
rect 2823 28540 2835 28543
rect 3605 28543 3663 28549
rect 3605 28540 3617 28543
rect 2823 28512 3617 28540
rect 2823 28509 2835 28512
rect 2777 28503 2835 28509
rect 3605 28509 3617 28512
rect 3651 28509 3663 28543
rect 3786 28540 3792 28552
rect 3747 28512 3792 28540
rect 3605 28503 3663 28509
rect 3786 28500 3792 28512
rect 3844 28500 3850 28552
rect 4982 28540 4988 28552
rect 4943 28512 4988 28540
rect 4982 28500 4988 28512
rect 5040 28500 5046 28552
rect 5644 28549 5672 28648
rect 7558 28636 7564 28648
rect 7616 28636 7622 28688
rect 12069 28679 12127 28685
rect 12069 28645 12081 28679
rect 12115 28676 12127 28679
rect 12434 28676 12440 28688
rect 12115 28648 12440 28676
rect 12115 28645 12127 28648
rect 12069 28639 12127 28645
rect 12434 28636 12440 28648
rect 12492 28676 12498 28688
rect 12710 28676 12716 28688
rect 12492 28648 12716 28676
rect 12492 28636 12498 28648
rect 12710 28636 12716 28648
rect 12768 28636 12774 28688
rect 7009 28611 7067 28617
rect 7009 28577 7021 28611
rect 7055 28608 7067 28611
rect 7190 28608 7196 28620
rect 7055 28580 7196 28608
rect 7055 28577 7067 28580
rect 7009 28571 7067 28577
rect 7190 28568 7196 28580
rect 7248 28608 7254 28620
rect 7466 28608 7472 28620
rect 7248 28580 7472 28608
rect 7248 28568 7254 28580
rect 7466 28568 7472 28580
rect 7524 28608 7530 28620
rect 8113 28611 8171 28617
rect 8113 28608 8125 28611
rect 7524 28580 8125 28608
rect 7524 28568 7530 28580
rect 8113 28577 8125 28580
rect 8159 28577 8171 28611
rect 8113 28571 8171 28577
rect 9674 28568 9680 28620
rect 9732 28608 9738 28620
rect 9953 28611 10011 28617
rect 9953 28608 9965 28611
rect 9732 28580 9965 28608
rect 9732 28568 9738 28580
rect 9953 28577 9965 28580
rect 9999 28577 10011 28611
rect 12820 28608 12848 28716
rect 14642 28704 14648 28716
rect 14700 28704 14706 28756
rect 16485 28747 16543 28753
rect 16485 28713 16497 28747
rect 16531 28744 16543 28747
rect 16850 28744 16856 28756
rect 16531 28716 16856 28744
rect 16531 28713 16543 28716
rect 16485 28707 16543 28713
rect 16850 28704 16856 28716
rect 16908 28704 16914 28756
rect 22002 28704 22008 28756
rect 22060 28744 22066 28756
rect 22649 28747 22707 28753
rect 22649 28744 22661 28747
rect 22060 28716 22661 28744
rect 22060 28704 22066 28716
rect 22649 28713 22661 28716
rect 22695 28713 22707 28747
rect 22649 28707 22707 28713
rect 14737 28679 14795 28685
rect 14737 28645 14749 28679
rect 14783 28676 14795 28679
rect 15102 28676 15108 28688
rect 14783 28648 15108 28676
rect 14783 28645 14795 28648
rect 14737 28639 14795 28645
rect 15102 28636 15108 28648
rect 15160 28636 15166 28688
rect 16206 28636 16212 28688
rect 16264 28676 16270 28688
rect 16264 28648 21312 28676
rect 16264 28636 16270 28648
rect 14458 28608 14464 28620
rect 9953 28571 10011 28577
rect 12728 28580 12848 28608
rect 13004 28580 14464 28608
rect 5629 28543 5687 28549
rect 5629 28509 5641 28543
rect 5675 28509 5687 28543
rect 5629 28503 5687 28509
rect 5810 28500 5816 28552
rect 5868 28540 5874 28552
rect 6733 28543 6791 28549
rect 6733 28540 6745 28543
rect 5868 28512 6745 28540
rect 5868 28500 5874 28512
rect 6733 28509 6745 28512
rect 6779 28509 6791 28543
rect 6733 28503 6791 28509
rect 7929 28543 7987 28549
rect 7929 28509 7941 28543
rect 7975 28540 7987 28543
rect 8386 28540 8392 28552
rect 7975 28512 8392 28540
rect 7975 28509 7987 28512
rect 7929 28503 7987 28509
rect 8386 28500 8392 28512
rect 8444 28500 8450 28552
rect 9125 28543 9183 28549
rect 9125 28509 9137 28543
rect 9171 28540 9183 28543
rect 9306 28540 9312 28552
rect 9171 28512 9312 28540
rect 9171 28509 9183 28512
rect 9125 28503 9183 28509
rect 9306 28500 9312 28512
rect 9364 28540 9370 28552
rect 9490 28540 9496 28552
rect 9364 28512 9496 28540
rect 9364 28500 9370 28512
rect 9490 28500 9496 28512
rect 9548 28500 9554 28552
rect 12728 28549 12756 28580
rect 12713 28543 12771 28549
rect 12713 28509 12725 28543
rect 12759 28509 12771 28543
rect 12713 28503 12771 28509
rect 12802 28500 12808 28552
rect 12860 28540 12866 28552
rect 13004 28549 13032 28580
rect 14458 28568 14464 28580
rect 14516 28568 14522 28620
rect 16942 28608 16948 28620
rect 16903 28580 16948 28608
rect 16942 28568 16948 28580
rect 17000 28568 17006 28620
rect 17129 28611 17187 28617
rect 17129 28577 17141 28611
rect 17175 28577 17187 28611
rect 17129 28571 17187 28577
rect 12989 28543 13047 28549
rect 12860 28512 12905 28540
rect 12860 28500 12866 28512
rect 12989 28509 13001 28543
rect 13035 28509 13047 28543
rect 12989 28503 13047 28509
rect 13178 28543 13236 28549
rect 13178 28509 13190 28543
rect 13224 28509 13236 28543
rect 14734 28540 14740 28552
rect 13178 28503 13236 28509
rect 14568 28512 14740 28540
rect 2130 28432 2136 28484
rect 2188 28472 2194 28484
rect 10220 28475 10278 28481
rect 2188 28444 7604 28472
rect 2188 28432 2194 28444
rect 1486 28404 1492 28416
rect 1447 28376 1492 28404
rect 1486 28364 1492 28376
rect 1544 28364 1550 28416
rect 3605 28407 3663 28413
rect 3605 28373 3617 28407
rect 3651 28404 3663 28407
rect 6365 28407 6423 28413
rect 6365 28404 6377 28407
rect 3651 28376 6377 28404
rect 3651 28373 3663 28376
rect 3605 28367 3663 28373
rect 6365 28373 6377 28376
rect 6411 28373 6423 28407
rect 6365 28367 6423 28373
rect 6822 28364 6828 28416
rect 6880 28404 6886 28416
rect 7576 28413 7604 28444
rect 10220 28441 10232 28475
rect 10266 28472 10278 28475
rect 10318 28472 10324 28484
rect 10266 28444 10324 28472
rect 10266 28441 10278 28444
rect 10220 28435 10278 28441
rect 10318 28432 10324 28444
rect 10376 28432 10382 28484
rect 10410 28432 10416 28484
rect 10468 28472 10474 28484
rect 11885 28475 11943 28481
rect 11885 28472 11897 28475
rect 10468 28444 11897 28472
rect 10468 28432 10474 28444
rect 11885 28441 11897 28444
rect 11931 28441 11943 28475
rect 13078 28472 13084 28484
rect 13039 28444 13084 28472
rect 11885 28435 11943 28441
rect 13078 28432 13084 28444
rect 13136 28432 13142 28484
rect 7561 28407 7619 28413
rect 6880 28376 6925 28404
rect 6880 28364 6886 28376
rect 7561 28373 7573 28407
rect 7607 28373 7619 28407
rect 7561 28367 7619 28373
rect 8018 28364 8024 28416
rect 8076 28404 8082 28416
rect 9030 28404 9036 28416
rect 8076 28376 8121 28404
rect 8991 28376 9036 28404
rect 8076 28364 8082 28376
rect 9030 28364 9036 28376
rect 9088 28364 9094 28416
rect 11238 28364 11244 28416
rect 11296 28404 11302 28416
rect 13188 28404 13216 28503
rect 13998 28432 14004 28484
rect 14056 28472 14062 28484
rect 14568 28481 14596 28512
rect 14734 28500 14740 28512
rect 14792 28540 14798 28552
rect 15381 28543 15439 28549
rect 15381 28540 15393 28543
rect 14792 28512 15393 28540
rect 14792 28500 14798 28512
rect 15381 28509 15393 28512
rect 15427 28509 15439 28543
rect 17144 28540 17172 28571
rect 17678 28568 17684 28620
rect 17736 28608 17742 28620
rect 18046 28608 18052 28620
rect 17736 28580 18052 28608
rect 17736 28568 17742 28580
rect 18046 28568 18052 28580
rect 18104 28568 18110 28620
rect 18138 28568 18144 28620
rect 18196 28608 18202 28620
rect 18233 28611 18291 28617
rect 18233 28608 18245 28611
rect 18196 28580 18245 28608
rect 18196 28568 18202 28580
rect 18233 28577 18245 28580
rect 18279 28577 18291 28611
rect 18233 28571 18291 28577
rect 18322 28568 18328 28620
rect 18380 28608 18386 28620
rect 21284 28617 21312 28648
rect 21269 28611 21327 28617
rect 18380 28580 20576 28608
rect 18380 28568 18386 28580
rect 18414 28540 18420 28552
rect 17144 28512 18420 28540
rect 15381 28503 15439 28509
rect 18414 28500 18420 28512
rect 18472 28540 18478 28552
rect 18874 28540 18880 28552
rect 18472 28512 18880 28540
rect 18472 28500 18478 28512
rect 18874 28500 18880 28512
rect 18932 28500 18938 28552
rect 19904 28549 19932 28580
rect 19889 28543 19947 28549
rect 19889 28509 19901 28543
rect 19935 28509 19947 28543
rect 19889 28503 19947 28509
rect 20441 28543 20499 28549
rect 20441 28509 20453 28543
rect 20487 28509 20499 28543
rect 20548 28540 20576 28580
rect 21269 28577 21281 28611
rect 21315 28577 21327 28611
rect 21269 28571 21327 28577
rect 22094 28540 22100 28552
rect 20548 28512 22100 28540
rect 20441 28503 20499 28509
rect 14553 28475 14611 28481
rect 14553 28472 14565 28475
rect 14056 28444 14565 28472
rect 14056 28432 14062 28444
rect 14553 28441 14565 28444
rect 14599 28441 14611 28475
rect 15194 28472 15200 28484
rect 15155 28444 15200 28472
rect 14553 28435 14611 28441
rect 15194 28432 15200 28444
rect 15252 28432 15258 28484
rect 15565 28475 15623 28481
rect 15565 28441 15577 28475
rect 15611 28472 15623 28475
rect 20456 28472 20484 28503
rect 22094 28500 22100 28512
rect 22152 28500 22158 28552
rect 15611 28444 20484 28472
rect 15611 28441 15623 28444
rect 15565 28435 15623 28441
rect 20530 28432 20536 28484
rect 20588 28472 20594 28484
rect 21514 28475 21572 28481
rect 21514 28472 21526 28475
rect 20588 28444 21526 28472
rect 20588 28432 20594 28444
rect 21514 28441 21526 28444
rect 21560 28441 21572 28475
rect 21514 28435 21572 28441
rect 13354 28404 13360 28416
rect 11296 28376 13216 28404
rect 13315 28376 13360 28404
rect 11296 28364 11302 28376
rect 13354 28364 13360 28376
rect 13412 28364 13418 28416
rect 16850 28404 16856 28416
rect 16811 28376 16856 28404
rect 16850 28364 16856 28376
rect 16908 28364 16914 28416
rect 18046 28364 18052 28416
rect 18104 28404 18110 28416
rect 18325 28407 18383 28413
rect 18325 28404 18337 28407
rect 18104 28376 18337 28404
rect 18104 28364 18110 28376
rect 18325 28373 18337 28376
rect 18371 28373 18383 28407
rect 18325 28367 18383 28373
rect 18506 28364 18512 28416
rect 18564 28404 18570 28416
rect 18693 28407 18751 28413
rect 18693 28404 18705 28407
rect 18564 28376 18705 28404
rect 18564 28364 18570 28376
rect 18693 28373 18705 28376
rect 18739 28373 18751 28407
rect 18693 28367 18751 28373
rect 19702 28364 19708 28416
rect 19760 28404 19766 28416
rect 19889 28407 19947 28413
rect 19889 28404 19901 28407
rect 19760 28376 19901 28404
rect 19760 28364 19766 28376
rect 19889 28373 19901 28376
rect 19935 28404 19947 28407
rect 20438 28404 20444 28416
rect 19935 28376 20444 28404
rect 19935 28373 19947 28376
rect 19889 28367 19947 28373
rect 20438 28364 20444 28376
rect 20496 28364 20502 28416
rect 20622 28404 20628 28416
rect 20535 28376 20628 28404
rect 20622 28364 20628 28376
rect 20680 28404 20686 28416
rect 29086 28404 29092 28416
rect 20680 28376 29092 28404
rect 20680 28364 20686 28376
rect 29086 28364 29092 28376
rect 29144 28364 29150 28416
rect 1104 28314 30820 28336
rect 1104 28262 10880 28314
rect 10932 28262 10944 28314
rect 10996 28262 11008 28314
rect 11060 28262 11072 28314
rect 11124 28262 11136 28314
rect 11188 28262 20811 28314
rect 20863 28262 20875 28314
rect 20927 28262 20939 28314
rect 20991 28262 21003 28314
rect 21055 28262 21067 28314
rect 21119 28262 30820 28314
rect 1104 28240 30820 28262
rect 4706 28200 4712 28212
rect 4667 28172 4712 28200
rect 4706 28160 4712 28172
rect 4764 28160 4770 28212
rect 4982 28160 4988 28212
rect 5040 28200 5046 28212
rect 6822 28200 6828 28212
rect 5040 28172 6684 28200
rect 6783 28172 6828 28200
rect 5040 28160 5046 28172
rect 3878 28132 3884 28144
rect 3068 28104 3884 28132
rect 1673 28067 1731 28073
rect 1673 28033 1685 28067
rect 1719 28033 1731 28067
rect 2130 28064 2136 28076
rect 2091 28036 2136 28064
rect 1673 28027 1731 28033
rect 1688 27996 1716 28027
rect 2130 28024 2136 28036
rect 2188 28024 2194 28076
rect 3068 28073 3096 28104
rect 3878 28092 3884 28104
rect 3936 28092 3942 28144
rect 4065 28135 4123 28141
rect 4065 28101 4077 28135
rect 4111 28132 4123 28135
rect 5350 28132 5356 28144
rect 4111 28104 5356 28132
rect 4111 28101 4123 28104
rect 4065 28095 4123 28101
rect 5350 28092 5356 28104
rect 5408 28092 5414 28144
rect 5445 28135 5503 28141
rect 5445 28101 5457 28135
rect 5491 28132 5503 28135
rect 5718 28132 5724 28144
rect 5491 28104 5724 28132
rect 5491 28101 5503 28104
rect 5445 28095 5503 28101
rect 5718 28092 5724 28104
rect 5776 28092 5782 28144
rect 6656 28132 6684 28172
rect 6822 28160 6828 28172
rect 6880 28160 6886 28212
rect 7469 28203 7527 28209
rect 7469 28169 7481 28203
rect 7515 28200 7527 28203
rect 8018 28200 8024 28212
rect 7515 28172 8024 28200
rect 7515 28169 7527 28172
rect 7469 28163 7527 28169
rect 8018 28160 8024 28172
rect 8076 28160 8082 28212
rect 8754 28200 8760 28212
rect 8405 28172 8760 28200
rect 7190 28132 7196 28144
rect 6656 28104 7196 28132
rect 7190 28092 7196 28104
rect 7248 28092 7254 28144
rect 7282 28092 7288 28144
rect 7340 28132 7346 28144
rect 8405 28132 8433 28172
rect 8754 28160 8760 28172
rect 8812 28160 8818 28212
rect 9214 28200 9220 28212
rect 9175 28172 9220 28200
rect 9214 28160 9220 28172
rect 9272 28160 9278 28212
rect 10318 28200 10324 28212
rect 10279 28172 10324 28200
rect 10318 28160 10324 28172
rect 10376 28160 10382 28212
rect 14458 28200 14464 28212
rect 14419 28172 14464 28200
rect 14458 28160 14464 28172
rect 14516 28160 14522 28212
rect 16117 28203 16175 28209
rect 16117 28169 16129 28203
rect 16163 28200 16175 28203
rect 16666 28200 16672 28212
rect 16163 28172 16672 28200
rect 16163 28169 16175 28172
rect 16117 28163 16175 28169
rect 16666 28160 16672 28172
rect 16724 28160 16730 28212
rect 16850 28160 16856 28212
rect 16908 28200 16914 28212
rect 17037 28203 17095 28209
rect 17037 28200 17049 28203
rect 16908 28172 17049 28200
rect 16908 28160 16914 28172
rect 17037 28169 17049 28172
rect 17083 28169 17095 28203
rect 20530 28200 20536 28212
rect 20491 28172 20536 28200
rect 17037 28163 17095 28169
rect 20530 28160 20536 28172
rect 20588 28160 20594 28212
rect 21910 28200 21916 28212
rect 20640 28172 21916 28200
rect 10873 28135 10931 28141
rect 10873 28132 10885 28135
rect 7340 28104 7788 28132
rect 7340 28092 7346 28104
rect 2317 28067 2375 28073
rect 2317 28033 2329 28067
rect 2363 28033 2375 28067
rect 2317 28027 2375 28033
rect 3053 28067 3111 28073
rect 3053 28033 3065 28067
rect 3099 28033 3111 28067
rect 3053 28027 3111 28033
rect 4617 28067 4675 28073
rect 4617 28033 4629 28067
rect 4663 28033 4675 28067
rect 4617 28027 4675 28033
rect 4801 28067 4859 28073
rect 4801 28033 4813 28067
rect 4847 28064 4859 28067
rect 6638 28064 6644 28076
rect 4847 28036 6644 28064
rect 4847 28033 4859 28036
rect 4801 28027 4859 28033
rect 2225 27999 2283 28005
rect 2225 27996 2237 27999
rect 1688 27968 2237 27996
rect 2225 27965 2237 27968
rect 2271 27965 2283 27999
rect 2332 27996 2360 28027
rect 2590 27996 2596 28008
rect 2332 27968 2596 27996
rect 2225 27959 2283 27965
rect 2590 27956 2596 27968
rect 2648 27996 2654 28008
rect 4632 27996 4660 28027
rect 6638 28024 6644 28036
rect 6696 28024 6702 28076
rect 7006 28064 7012 28076
rect 6967 28036 7012 28064
rect 7006 28024 7012 28036
rect 7064 28024 7070 28076
rect 7760 28073 7788 28104
rect 8036 28104 8433 28132
rect 8680 28104 10885 28132
rect 7653 28067 7711 28073
rect 7653 28033 7665 28067
rect 7699 28033 7711 28067
rect 7653 28027 7711 28033
rect 7745 28067 7803 28073
rect 7745 28033 7757 28067
rect 7791 28064 7803 28067
rect 7926 28064 7932 28076
rect 7791 28036 7932 28064
rect 7791 28033 7803 28036
rect 7745 28027 7803 28033
rect 2648 27968 4660 27996
rect 7668 27996 7696 28027
rect 7926 28024 7932 28036
rect 7984 28024 7990 28076
rect 8036 28073 8064 28104
rect 8021 28067 8079 28073
rect 8021 28033 8033 28067
rect 8067 28033 8079 28067
rect 8021 28027 8079 28033
rect 8110 28024 8116 28076
rect 8168 28064 8174 28076
rect 8168 28036 8433 28064
rect 8168 28024 8174 28036
rect 8202 27996 8208 28008
rect 7668 27968 8208 27996
rect 2648 27956 2654 27968
rect 8202 27956 8208 27968
rect 8260 27956 8266 28008
rect 8405 27996 8433 28036
rect 8478 28024 8484 28076
rect 8536 28064 8542 28076
rect 8680 28073 8708 28104
rect 10873 28101 10885 28104
rect 10919 28101 10931 28135
rect 10873 28095 10931 28101
rect 12345 28135 12403 28141
rect 12345 28101 12357 28135
rect 12391 28132 12403 28135
rect 12802 28132 12808 28144
rect 12391 28104 12808 28132
rect 12391 28101 12403 28104
rect 12345 28095 12403 28101
rect 12802 28092 12808 28104
rect 12860 28092 12866 28144
rect 14090 28132 14096 28144
rect 13096 28104 14096 28132
rect 8665 28067 8723 28073
rect 8536 28036 8581 28064
rect 8536 28024 8542 28036
rect 8665 28033 8677 28067
rect 8711 28033 8723 28067
rect 9030 28064 9036 28076
rect 8991 28036 9036 28064
rect 8665 28027 8723 28033
rect 9030 28024 9036 28036
rect 9088 28024 9094 28076
rect 9122 28024 9128 28076
rect 9180 28064 9186 28076
rect 9677 28067 9735 28073
rect 9677 28064 9689 28067
rect 9180 28036 9689 28064
rect 9180 28024 9186 28036
rect 9677 28033 9689 28036
rect 9723 28033 9735 28067
rect 9677 28027 9735 28033
rect 9770 28067 9828 28073
rect 9770 28033 9782 28067
rect 9816 28033 9828 28067
rect 9770 28027 9828 28033
rect 9953 28067 10011 28073
rect 9953 28033 9965 28067
rect 9999 28033 10011 28067
rect 9953 28027 10011 28033
rect 8757 27999 8815 28005
rect 8757 27996 8769 27999
rect 8405 27968 8769 27996
rect 8757 27965 8769 27968
rect 8803 27965 8815 27999
rect 8757 27959 8815 27965
rect 8849 27999 8907 28005
rect 8849 27965 8861 27999
rect 8895 27965 8907 27999
rect 8849 27959 8907 27965
rect 5626 27928 5632 27940
rect 5587 27900 5632 27928
rect 5626 27888 5632 27900
rect 5684 27888 5690 27940
rect 5810 27888 5816 27940
rect 5868 27928 5874 27940
rect 5868 27900 8064 27928
rect 5868 27888 5874 27900
rect 1486 27860 1492 27872
rect 1447 27832 1492 27860
rect 1486 27820 1492 27832
rect 1544 27820 1550 27872
rect 2866 27860 2872 27872
rect 2779 27832 2872 27860
rect 2866 27820 2872 27832
rect 2924 27860 2930 27872
rect 3694 27860 3700 27872
rect 2924 27832 3700 27860
rect 2924 27820 2930 27832
rect 3694 27820 3700 27832
rect 3752 27820 3758 27872
rect 7374 27820 7380 27872
rect 7432 27860 7438 27872
rect 7929 27863 7987 27869
rect 7929 27860 7941 27863
rect 7432 27832 7941 27860
rect 7432 27820 7438 27832
rect 7929 27829 7941 27832
rect 7975 27829 7987 27863
rect 8036 27860 8064 27900
rect 8110 27888 8116 27940
rect 8168 27928 8174 27940
rect 8864 27928 8892 27959
rect 9306 27956 9312 28008
rect 9364 27996 9370 28008
rect 9784 27996 9812 28027
rect 9364 27968 9812 27996
rect 9968 27996 9996 28027
rect 10042 28024 10048 28076
rect 10100 28064 10106 28076
rect 10226 28073 10232 28076
rect 10183 28067 10232 28073
rect 10100 28036 10145 28064
rect 10100 28024 10106 28036
rect 10183 28033 10195 28067
rect 10229 28033 10232 28067
rect 10183 28027 10232 28033
rect 10226 28024 10232 28027
rect 10284 28024 10290 28076
rect 10965 28067 11023 28073
rect 10965 28033 10977 28067
rect 11011 28064 11023 28067
rect 11330 28064 11336 28076
rect 11011 28036 11336 28064
rect 11011 28033 11023 28036
rect 10965 28027 11023 28033
rect 10980 27996 11008 28027
rect 11330 28024 11336 28036
rect 11388 28024 11394 28076
rect 11517 28067 11575 28073
rect 11517 28033 11529 28067
rect 11563 28064 11575 28067
rect 11606 28064 11612 28076
rect 11563 28036 11612 28064
rect 11563 28033 11575 28036
rect 11517 28027 11575 28033
rect 11606 28024 11612 28036
rect 11664 28024 11670 28076
rect 13096 28073 13124 28104
rect 14090 28092 14096 28104
rect 14148 28092 14154 28144
rect 17497 28135 17555 28141
rect 17497 28101 17509 28135
rect 17543 28132 17555 28135
rect 17586 28132 17592 28144
rect 17543 28104 17592 28132
rect 17543 28101 17555 28104
rect 17497 28095 17555 28101
rect 17586 28092 17592 28104
rect 17644 28092 17650 28144
rect 20640 28141 20668 28172
rect 21910 28160 21916 28172
rect 21968 28160 21974 28212
rect 29730 28160 29736 28212
rect 29788 28200 29794 28212
rect 30009 28203 30067 28209
rect 30009 28200 30021 28203
rect 29788 28172 30021 28200
rect 29788 28160 29794 28172
rect 30009 28169 30021 28172
rect 30055 28169 30067 28203
rect 30009 28163 30067 28169
rect 20625 28135 20683 28141
rect 20625 28101 20637 28135
rect 20671 28101 20683 28135
rect 20625 28095 20683 28101
rect 21266 28092 21272 28144
rect 21324 28132 21330 28144
rect 22002 28132 22008 28144
rect 21324 28104 22008 28132
rect 21324 28092 21330 28104
rect 22002 28092 22008 28104
rect 22060 28092 22066 28144
rect 13354 28073 13360 28076
rect 13081 28067 13139 28073
rect 13081 28033 13093 28067
rect 13127 28033 13139 28067
rect 13348 28064 13360 28073
rect 13315 28036 13360 28064
rect 13081 28027 13139 28033
rect 13348 28027 13360 28036
rect 13354 28024 13360 28027
rect 13412 28024 13418 28076
rect 14642 28024 14648 28076
rect 14700 28064 14706 28076
rect 14921 28067 14979 28073
rect 14921 28064 14933 28067
rect 14700 28036 14933 28064
rect 14700 28024 14706 28036
rect 14921 28033 14933 28036
rect 14967 28033 14979 28067
rect 15746 28064 15752 28076
rect 15707 28036 15752 28064
rect 14921 28027 14979 28033
rect 15746 28024 15752 28036
rect 15804 28024 15810 28076
rect 15933 28067 15991 28073
rect 15933 28033 15945 28067
rect 15979 28064 15991 28067
rect 16206 28064 16212 28076
rect 15979 28036 16212 28064
rect 15979 28033 15991 28036
rect 15933 28027 15991 28033
rect 16206 28024 16212 28036
rect 16264 28024 16270 28076
rect 17402 28064 17408 28076
rect 17363 28036 17408 28064
rect 17402 28024 17408 28036
rect 17460 28024 17466 28076
rect 18322 28024 18328 28076
rect 18380 28064 18386 28076
rect 18601 28067 18659 28073
rect 18601 28064 18613 28067
rect 18380 28036 18613 28064
rect 18380 28024 18386 28036
rect 18601 28033 18613 28036
rect 18647 28033 18659 28067
rect 18601 28027 18659 28033
rect 18690 28024 18696 28076
rect 18748 28064 18754 28076
rect 18966 28064 18972 28076
rect 18748 28036 18793 28064
rect 18927 28036 18972 28064
rect 18748 28024 18754 28036
rect 18966 28024 18972 28036
rect 19024 28024 19030 28076
rect 19334 28024 19340 28076
rect 19392 28064 19398 28076
rect 20349 28067 20407 28073
rect 20349 28064 20361 28067
rect 19392 28036 20361 28064
rect 19392 28024 19398 28036
rect 20349 28033 20361 28036
rect 20395 28033 20407 28067
rect 20349 28027 20407 28033
rect 20441 28067 20499 28073
rect 20441 28033 20453 28067
rect 20487 28033 20499 28067
rect 20714 28064 20720 28076
rect 20675 28036 20720 28064
rect 20441 28027 20499 28033
rect 9968 27968 11008 27996
rect 9364 27956 9370 27968
rect 16390 27956 16396 28008
rect 16448 27996 16454 28008
rect 17589 27999 17647 28005
rect 17589 27996 17601 27999
rect 16448 27968 17601 27996
rect 16448 27956 16454 27968
rect 17589 27965 17601 27968
rect 17635 27996 17647 27999
rect 17678 27996 17684 28008
rect 17635 27968 17684 27996
rect 17635 27965 17647 27968
rect 17589 27959 17647 27965
rect 17678 27956 17684 27968
rect 17736 27956 17742 28008
rect 20456 27996 20484 28027
rect 20714 28024 20720 28036
rect 20772 28024 20778 28076
rect 20806 28024 20812 28076
rect 20864 28064 20870 28076
rect 21821 28067 21879 28073
rect 20864 28036 20909 28064
rect 20864 28024 20870 28036
rect 21821 28033 21833 28067
rect 21867 28064 21879 28067
rect 22094 28064 22100 28076
rect 21867 28036 22100 28064
rect 21867 28033 21879 28036
rect 21821 28027 21879 28033
rect 22094 28024 22100 28036
rect 22152 28024 22158 28076
rect 22189 28067 22247 28073
rect 22189 28033 22201 28067
rect 22235 28064 22247 28067
rect 22370 28064 22376 28076
rect 22235 28036 22376 28064
rect 22235 28033 22247 28036
rect 22189 28027 22247 28033
rect 22370 28024 22376 28036
rect 22428 28024 22434 28076
rect 29822 28064 29828 28076
rect 29783 28036 29828 28064
rect 29822 28024 29828 28036
rect 29880 28024 29886 28076
rect 21542 27996 21548 28008
rect 20456 27968 21548 27996
rect 21542 27956 21548 27968
rect 21600 27956 21606 28008
rect 9490 27928 9496 27940
rect 8168 27900 8892 27928
rect 8956 27900 9496 27928
rect 8168 27888 8174 27900
rect 8956 27860 8984 27900
rect 9490 27888 9496 27900
rect 9548 27928 9554 27940
rect 10962 27928 10968 27940
rect 9548 27900 10968 27928
rect 9548 27888 9554 27900
rect 10962 27888 10968 27900
rect 11020 27888 11026 27940
rect 12158 27928 12164 27940
rect 12119 27900 12164 27928
rect 12158 27888 12164 27900
rect 12216 27888 12222 27940
rect 8036 27832 8984 27860
rect 7929 27823 7987 27829
rect 9122 27820 9128 27872
rect 9180 27860 9186 27872
rect 11609 27863 11667 27869
rect 11609 27860 11621 27863
rect 9180 27832 11621 27860
rect 9180 27820 9186 27832
rect 11609 27829 11621 27832
rect 11655 27829 11667 27863
rect 11609 27823 11667 27829
rect 15013 27863 15071 27869
rect 15013 27829 15025 27863
rect 15059 27860 15071 27863
rect 15286 27860 15292 27872
rect 15059 27832 15292 27860
rect 15059 27829 15071 27832
rect 15013 27823 15071 27829
rect 15286 27820 15292 27832
rect 15344 27820 15350 27872
rect 18414 27860 18420 27872
rect 18375 27832 18420 27860
rect 18414 27820 18420 27832
rect 18472 27820 18478 27872
rect 18877 27863 18935 27869
rect 18877 27829 18889 27863
rect 18923 27860 18935 27863
rect 19426 27860 19432 27872
rect 18923 27832 19432 27860
rect 18923 27829 18935 27832
rect 18877 27823 18935 27829
rect 19426 27820 19432 27832
rect 19484 27820 19490 27872
rect 1104 27770 30820 27792
rect 1104 27718 5915 27770
rect 5967 27718 5979 27770
rect 6031 27718 6043 27770
rect 6095 27718 6107 27770
rect 6159 27718 6171 27770
rect 6223 27718 15846 27770
rect 15898 27718 15910 27770
rect 15962 27718 15974 27770
rect 16026 27718 16038 27770
rect 16090 27718 16102 27770
rect 16154 27718 25776 27770
rect 25828 27718 25840 27770
rect 25892 27718 25904 27770
rect 25956 27718 25968 27770
rect 26020 27718 26032 27770
rect 26084 27718 30820 27770
rect 1104 27696 30820 27718
rect 5810 27656 5816 27668
rect 5771 27628 5816 27656
rect 5810 27616 5816 27628
rect 5868 27616 5874 27668
rect 7006 27616 7012 27668
rect 7064 27656 7070 27668
rect 7285 27659 7343 27665
rect 7285 27656 7297 27659
rect 7064 27628 7297 27656
rect 7064 27616 7070 27628
rect 7285 27625 7297 27628
rect 7331 27625 7343 27659
rect 7285 27619 7343 27625
rect 7374 27616 7380 27668
rect 7432 27656 7438 27668
rect 7469 27659 7527 27665
rect 7469 27656 7481 27659
rect 7432 27628 7481 27656
rect 7432 27616 7438 27628
rect 7469 27625 7481 27628
rect 7515 27625 7527 27659
rect 13630 27656 13636 27668
rect 7469 27619 7527 27625
rect 7760 27628 13636 27656
rect 6546 27588 6552 27600
rect 6507 27560 6552 27588
rect 6546 27548 6552 27560
rect 6604 27548 6610 27600
rect 2792 27492 4568 27520
rect 2590 27452 2596 27464
rect 2551 27424 2596 27452
rect 2590 27412 2596 27424
rect 2648 27412 2654 27464
rect 2792 27461 2820 27492
rect 2777 27455 2835 27461
rect 2777 27421 2789 27455
rect 2823 27421 2835 27455
rect 2777 27415 2835 27421
rect 4338 27412 4344 27464
rect 4396 27452 4402 27464
rect 4433 27455 4491 27461
rect 4433 27452 4445 27455
rect 4396 27424 4445 27452
rect 4396 27412 4402 27424
rect 4433 27421 4445 27424
rect 4479 27421 4491 27455
rect 4540 27452 4568 27492
rect 4540 27424 6868 27452
rect 4433 27415 4491 27421
rect 4700 27387 4758 27393
rect 4700 27353 4712 27387
rect 4746 27384 4758 27387
rect 4890 27384 4896 27396
rect 4746 27356 4896 27384
rect 4746 27353 4758 27356
rect 4700 27347 4758 27353
rect 4890 27344 4896 27356
rect 4948 27344 4954 27396
rect 6730 27384 6736 27396
rect 6691 27356 6736 27384
rect 6730 27344 6736 27356
rect 6788 27344 6794 27396
rect 6840 27384 6868 27424
rect 7098 27412 7104 27464
rect 7156 27452 7162 27464
rect 7760 27461 7788 27628
rect 13630 27616 13636 27628
rect 13688 27616 13694 27668
rect 16117 27659 16175 27665
rect 16117 27625 16129 27659
rect 16163 27656 16175 27659
rect 16206 27656 16212 27668
rect 16163 27628 16212 27656
rect 16163 27625 16175 27628
rect 16117 27619 16175 27625
rect 16206 27616 16212 27628
rect 16264 27616 16270 27668
rect 18966 27616 18972 27668
rect 19024 27656 19030 27668
rect 19245 27659 19303 27665
rect 19245 27656 19257 27659
rect 19024 27628 19257 27656
rect 19024 27616 19030 27628
rect 19245 27625 19257 27628
rect 19291 27625 19303 27659
rect 19245 27619 19303 27625
rect 20806 27616 20812 27668
rect 20864 27656 20870 27668
rect 21085 27659 21143 27665
rect 21085 27656 21097 27659
rect 20864 27628 21097 27656
rect 20864 27616 20870 27628
rect 21085 27625 21097 27628
rect 21131 27625 21143 27659
rect 21085 27619 21143 27625
rect 8297 27591 8355 27597
rect 8297 27557 8309 27591
rect 8343 27588 8355 27591
rect 8386 27588 8392 27600
rect 8343 27560 8392 27588
rect 8343 27557 8355 27560
rect 8297 27551 8355 27557
rect 8386 27548 8392 27560
rect 8444 27548 8450 27600
rect 9490 27548 9496 27600
rect 9548 27548 9554 27600
rect 9769 27591 9827 27597
rect 9769 27557 9781 27591
rect 9815 27588 9827 27591
rect 9858 27588 9864 27600
rect 9815 27560 9864 27588
rect 9815 27557 9827 27560
rect 9769 27551 9827 27557
rect 9858 27548 9864 27560
rect 9916 27548 9922 27600
rect 10781 27591 10839 27597
rect 10781 27557 10793 27591
rect 10827 27588 10839 27591
rect 11238 27588 11244 27600
rect 10827 27560 11244 27588
rect 10827 27557 10839 27560
rect 10781 27551 10839 27557
rect 11238 27548 11244 27560
rect 11296 27548 11302 27600
rect 14274 27548 14280 27600
rect 14332 27588 14338 27600
rect 14461 27591 14519 27597
rect 14461 27588 14473 27591
rect 14332 27560 14473 27588
rect 14332 27548 14338 27560
rect 14461 27557 14473 27560
rect 14507 27557 14519 27591
rect 14461 27551 14519 27557
rect 18690 27548 18696 27600
rect 18748 27588 18754 27600
rect 18748 27560 20576 27588
rect 18748 27548 18754 27560
rect 9508 27520 9536 27548
rect 10689 27523 10747 27529
rect 10689 27520 10701 27523
rect 9508 27492 10701 27520
rect 10689 27489 10701 27492
rect 10735 27489 10747 27523
rect 10689 27483 10747 27489
rect 14829 27523 14887 27529
rect 14829 27489 14841 27523
rect 14875 27520 14887 27523
rect 15381 27523 15439 27529
rect 15381 27520 15393 27523
rect 14875 27492 15393 27520
rect 14875 27489 14887 27492
rect 14829 27483 14887 27489
rect 15381 27489 15393 27492
rect 15427 27489 15439 27523
rect 15381 27483 15439 27489
rect 15565 27523 15623 27529
rect 15565 27489 15577 27523
rect 15611 27520 15623 27523
rect 15654 27520 15660 27532
rect 15611 27492 15660 27520
rect 15611 27489 15623 27492
rect 15565 27483 15623 27489
rect 15654 27480 15660 27492
rect 15712 27480 15718 27532
rect 16390 27480 16396 27532
rect 16448 27520 16454 27532
rect 16669 27523 16727 27529
rect 16669 27520 16681 27523
rect 16448 27492 16681 27520
rect 16448 27480 16454 27492
rect 16669 27489 16681 27492
rect 16715 27489 16727 27523
rect 17402 27520 17408 27532
rect 16669 27483 16727 27489
rect 16776 27492 17408 27520
rect 7745 27455 7803 27461
rect 7745 27452 7757 27455
rect 7156 27424 7757 27452
rect 7156 27412 7162 27424
rect 7745 27421 7757 27424
rect 7791 27421 7803 27455
rect 7745 27415 7803 27421
rect 8389 27455 8447 27461
rect 8389 27421 8401 27455
rect 8435 27452 8447 27455
rect 8662 27452 8668 27464
rect 8435 27424 8668 27452
rect 8435 27421 8447 27424
rect 8389 27415 8447 27421
rect 8662 27412 8668 27424
rect 8720 27412 8726 27464
rect 9030 27412 9036 27464
rect 9088 27452 9094 27464
rect 9306 27461 9312 27464
rect 9125 27455 9183 27461
rect 9125 27452 9137 27455
rect 9088 27424 9137 27452
rect 9088 27412 9094 27424
rect 9125 27421 9137 27424
rect 9171 27421 9183 27455
rect 9125 27415 9183 27421
rect 9273 27455 9312 27461
rect 9273 27421 9285 27455
rect 9273 27415 9312 27421
rect 9306 27412 9312 27415
rect 9364 27412 9370 27464
rect 9674 27461 9680 27464
rect 9631 27455 9680 27461
rect 9631 27421 9643 27455
rect 9677 27421 9680 27455
rect 9631 27415 9680 27421
rect 9674 27412 9680 27415
rect 9732 27452 9738 27464
rect 10226 27452 10232 27464
rect 9732 27424 10232 27452
rect 9732 27412 9738 27424
rect 10226 27412 10232 27424
rect 10284 27412 10290 27464
rect 10318 27412 10324 27464
rect 10376 27452 10382 27464
rect 10873 27455 10931 27461
rect 10873 27452 10885 27455
rect 10376 27424 10885 27452
rect 10376 27412 10382 27424
rect 10873 27421 10885 27424
rect 10919 27421 10931 27455
rect 10873 27415 10931 27421
rect 10962 27412 10968 27464
rect 11020 27452 11026 27464
rect 11422 27452 11428 27464
rect 11020 27424 11065 27452
rect 11383 27424 11428 27452
rect 11020 27412 11026 27424
rect 11422 27412 11428 27424
rect 11480 27412 11486 27464
rect 14366 27452 14372 27464
rect 14327 27424 14372 27452
rect 14366 27412 14372 27424
rect 14424 27412 14430 27464
rect 14550 27412 14556 27464
rect 14608 27452 14614 27464
rect 14645 27455 14703 27461
rect 14645 27452 14657 27455
rect 14608 27424 14657 27452
rect 14608 27412 14614 27424
rect 14645 27421 14657 27424
rect 14691 27421 14703 27455
rect 15286 27452 15292 27464
rect 15247 27424 15292 27452
rect 14645 27415 14703 27421
rect 15286 27412 15292 27424
rect 15344 27412 15350 27464
rect 16485 27455 16543 27461
rect 16485 27421 16497 27455
rect 16531 27452 16543 27455
rect 16776 27452 16804 27492
rect 17402 27480 17408 27492
rect 17460 27480 17466 27532
rect 17678 27480 17684 27532
rect 17736 27520 17742 27532
rect 18233 27523 18291 27529
rect 18233 27520 18245 27523
rect 17736 27492 18245 27520
rect 17736 27480 17742 27492
rect 18233 27489 18245 27492
rect 18279 27489 18291 27523
rect 18233 27483 18291 27489
rect 18966 27480 18972 27532
rect 19024 27520 19030 27532
rect 19797 27523 19855 27529
rect 19797 27520 19809 27523
rect 19024 27492 19809 27520
rect 19024 27480 19030 27492
rect 19797 27489 19809 27492
rect 19843 27489 19855 27523
rect 19797 27483 19855 27489
rect 16531 27424 16804 27452
rect 16531 27421 16543 27424
rect 16485 27415 16543 27421
rect 16850 27412 16856 27464
rect 16908 27452 16914 27464
rect 17313 27455 17371 27461
rect 17313 27452 17325 27455
rect 16908 27424 17325 27452
rect 16908 27412 16914 27424
rect 17313 27421 17325 27424
rect 17359 27421 17371 27455
rect 17313 27415 17371 27421
rect 17494 27412 17500 27464
rect 17552 27452 17558 27464
rect 17957 27455 18015 27461
rect 17957 27452 17969 27455
rect 17552 27424 17969 27452
rect 17552 27412 17558 27424
rect 17957 27421 17969 27424
rect 18003 27421 18015 27455
rect 18138 27452 18144 27464
rect 18099 27424 18144 27452
rect 17957 27415 18015 27421
rect 18138 27412 18144 27424
rect 18196 27412 18202 27464
rect 18325 27455 18383 27461
rect 18325 27421 18337 27455
rect 18371 27421 18383 27455
rect 18506 27452 18512 27464
rect 18467 27424 18512 27452
rect 18325 27415 18383 27421
rect 8570 27384 8576 27396
rect 6840 27356 8576 27384
rect 8570 27344 8576 27356
rect 8628 27344 8634 27396
rect 8680 27384 8708 27412
rect 9401 27387 9459 27393
rect 9401 27384 9413 27387
rect 8680 27356 9413 27384
rect 9401 27353 9413 27356
rect 9447 27353 9459 27387
rect 9401 27347 9459 27353
rect 9493 27387 9551 27393
rect 9493 27353 9505 27387
rect 9539 27353 9551 27387
rect 9493 27347 9551 27353
rect 1670 27276 1676 27328
rect 1728 27316 1734 27328
rect 2685 27319 2743 27325
rect 2685 27316 2697 27319
rect 1728 27288 2697 27316
rect 1728 27276 1734 27288
rect 2685 27285 2697 27288
rect 2731 27285 2743 27319
rect 2685 27279 2743 27285
rect 6270 27276 6276 27328
rect 6328 27316 6334 27328
rect 8386 27316 8392 27328
rect 6328 27288 8392 27316
rect 6328 27276 6334 27288
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 8846 27276 8852 27328
rect 8904 27316 8910 27328
rect 9508 27316 9536 27347
rect 11514 27344 11520 27396
rect 11572 27384 11578 27396
rect 11670 27387 11728 27393
rect 11670 27384 11682 27387
rect 11572 27356 11682 27384
rect 11572 27344 11578 27356
rect 11670 27353 11682 27356
rect 11716 27353 11728 27387
rect 18340 27384 18368 27415
rect 18506 27412 18512 27424
rect 18564 27412 18570 27464
rect 19058 27412 19064 27464
rect 19116 27452 19122 27464
rect 20441 27455 20499 27461
rect 20441 27452 20453 27455
rect 19116 27424 20453 27452
rect 19116 27412 19122 27424
rect 20441 27421 20453 27424
rect 20487 27421 20499 27455
rect 20548 27452 20576 27560
rect 20714 27548 20720 27600
rect 20772 27588 20778 27600
rect 21174 27588 21180 27600
rect 20772 27560 21180 27588
rect 20772 27548 20778 27560
rect 21174 27548 21180 27560
rect 21232 27588 21238 27600
rect 21637 27591 21695 27597
rect 21637 27588 21649 27591
rect 21232 27560 21649 27588
rect 21232 27548 21238 27560
rect 21637 27557 21649 27560
rect 21683 27557 21695 27591
rect 21637 27551 21695 27557
rect 20806 27520 20812 27532
rect 20767 27492 20812 27520
rect 20806 27480 20812 27492
rect 20864 27480 20870 27532
rect 20625 27455 20683 27461
rect 20625 27452 20637 27455
rect 20548 27424 20637 27452
rect 20441 27415 20499 27421
rect 20625 27421 20637 27424
rect 20671 27421 20683 27455
rect 20625 27415 20683 27421
rect 20717 27455 20775 27461
rect 20717 27421 20729 27455
rect 20763 27421 20775 27455
rect 20717 27415 20775 27421
rect 20901 27455 20959 27461
rect 20901 27421 20913 27455
rect 20947 27452 20959 27455
rect 21266 27452 21272 27464
rect 20947 27424 21272 27452
rect 20947 27421 20959 27424
rect 20901 27415 20959 27421
rect 18782 27384 18788 27396
rect 18340 27356 18788 27384
rect 11670 27347 11728 27353
rect 18524 27328 18552 27356
rect 18782 27344 18788 27356
rect 18840 27344 18846 27396
rect 19150 27344 19156 27396
rect 19208 27384 19214 27396
rect 19705 27387 19763 27393
rect 19705 27384 19717 27387
rect 19208 27356 19717 27384
rect 19208 27344 19214 27356
rect 19705 27353 19717 27356
rect 19751 27353 19763 27387
rect 19705 27347 19763 27353
rect 20530 27344 20536 27396
rect 20588 27384 20594 27396
rect 20732 27384 20760 27415
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 21542 27452 21548 27464
rect 21503 27424 21548 27452
rect 21542 27412 21548 27424
rect 21600 27412 21606 27464
rect 29362 27412 29368 27464
rect 29420 27452 29426 27464
rect 29825 27455 29883 27461
rect 29825 27452 29837 27455
rect 29420 27424 29837 27452
rect 29420 27412 29426 27424
rect 29825 27421 29837 27424
rect 29871 27421 29883 27455
rect 29825 27415 29883 27421
rect 20588 27356 20760 27384
rect 20588 27344 20594 27356
rect 8904 27288 9536 27316
rect 8904 27276 8910 27288
rect 12710 27276 12716 27328
rect 12768 27316 12774 27328
rect 12805 27319 12863 27325
rect 12805 27316 12817 27319
rect 12768 27288 12817 27316
rect 12768 27276 12774 27288
rect 12805 27285 12817 27288
rect 12851 27285 12863 27319
rect 15562 27316 15568 27328
rect 15523 27288 15568 27316
rect 12805 27279 12863 27285
rect 15562 27276 15568 27288
rect 15620 27276 15626 27328
rect 16577 27319 16635 27325
rect 16577 27285 16589 27319
rect 16623 27316 16635 27319
rect 16666 27316 16672 27328
rect 16623 27288 16672 27316
rect 16623 27285 16635 27288
rect 16577 27279 16635 27285
rect 16666 27276 16672 27288
rect 16724 27276 16730 27328
rect 17402 27316 17408 27328
rect 17363 27288 17408 27316
rect 17402 27276 17408 27288
rect 17460 27276 17466 27328
rect 18506 27276 18512 27328
rect 18564 27276 18570 27328
rect 18598 27276 18604 27328
rect 18656 27316 18662 27328
rect 18693 27319 18751 27325
rect 18693 27316 18705 27319
rect 18656 27288 18705 27316
rect 18656 27276 18662 27288
rect 18693 27285 18705 27288
rect 18739 27285 18751 27319
rect 18693 27279 18751 27285
rect 19058 27276 19064 27328
rect 19116 27316 19122 27328
rect 19613 27319 19671 27325
rect 19613 27316 19625 27319
rect 19116 27288 19625 27316
rect 19116 27276 19122 27288
rect 19613 27285 19625 27288
rect 19659 27285 19671 27319
rect 30006 27316 30012 27328
rect 29967 27288 30012 27316
rect 19613 27279 19671 27285
rect 30006 27276 30012 27288
rect 30064 27276 30070 27328
rect 1104 27226 30820 27248
rect 1104 27174 10880 27226
rect 10932 27174 10944 27226
rect 10996 27174 11008 27226
rect 11060 27174 11072 27226
rect 11124 27174 11136 27226
rect 11188 27174 20811 27226
rect 20863 27174 20875 27226
rect 20927 27174 20939 27226
rect 20991 27174 21003 27226
rect 21055 27174 21067 27226
rect 21119 27174 30820 27226
rect 1104 27152 30820 27174
rect 5813 27115 5871 27121
rect 5813 27081 5825 27115
rect 5859 27112 5871 27115
rect 8202 27112 8208 27124
rect 5859 27084 8208 27112
rect 5859 27081 5871 27084
rect 5813 27075 5871 27081
rect 8202 27072 8208 27084
rect 8260 27072 8266 27124
rect 8386 27072 8392 27124
rect 8444 27112 8450 27124
rect 10318 27112 10324 27124
rect 8444 27084 10324 27112
rect 8444 27072 8450 27084
rect 10318 27072 10324 27084
rect 10376 27112 10382 27124
rect 10686 27112 10692 27124
rect 10376 27084 10692 27112
rect 10376 27072 10382 27084
rect 10686 27072 10692 27084
rect 10744 27072 10750 27124
rect 10778 27072 10784 27124
rect 10836 27112 10842 27124
rect 10873 27115 10931 27121
rect 10873 27112 10885 27115
rect 10836 27084 10885 27112
rect 10836 27072 10842 27084
rect 10873 27081 10885 27084
rect 10919 27081 10931 27115
rect 16666 27112 16672 27124
rect 16627 27084 16672 27112
rect 10873 27075 10931 27081
rect 16666 27072 16672 27084
rect 16724 27072 16730 27124
rect 20530 27112 20536 27124
rect 20491 27084 20536 27112
rect 20530 27072 20536 27084
rect 20588 27072 20594 27124
rect 4338 27044 4344 27056
rect 3344 27016 4344 27044
rect 1670 26976 1676 26988
rect 1631 26948 1676 26976
rect 1670 26936 1676 26948
rect 1728 26936 1734 26988
rect 3344 26985 3372 27016
rect 4338 27004 4344 27016
rect 4396 27004 4402 27056
rect 6730 27004 6736 27056
rect 6788 27044 6794 27056
rect 8481 27047 8539 27053
rect 8481 27044 8493 27047
rect 6788 27016 8493 27044
rect 6788 27004 6794 27016
rect 8481 27013 8493 27016
rect 8527 27013 8539 27047
rect 8481 27007 8539 27013
rect 8665 27047 8723 27053
rect 8665 27013 8677 27047
rect 8711 27044 8723 27047
rect 10410 27044 10416 27056
rect 8711 27016 10416 27044
rect 8711 27013 8723 27016
rect 8665 27007 8723 27013
rect 10410 27004 10416 27016
rect 10468 27004 10474 27056
rect 15562 27004 15568 27056
rect 15620 27044 15626 27056
rect 15933 27047 15991 27053
rect 15933 27044 15945 27047
rect 15620 27016 15945 27044
rect 15620 27004 15626 27016
rect 15933 27013 15945 27016
rect 15979 27013 15991 27047
rect 18966 27044 18972 27056
rect 15933 27007 15991 27013
rect 18156 27016 18972 27044
rect 3602 26985 3608 26988
rect 3329 26979 3387 26985
rect 3329 26945 3341 26979
rect 3375 26945 3387 26979
rect 3329 26939 3387 26945
rect 3596 26939 3608 26985
rect 3660 26976 3666 26988
rect 3660 26948 3696 26976
rect 3602 26936 3608 26939
rect 3660 26936 3666 26948
rect 4982 26936 4988 26988
rect 5040 26976 5046 26988
rect 5353 26979 5411 26985
rect 5353 26976 5365 26979
rect 5040 26948 5365 26976
rect 5040 26936 5046 26948
rect 5353 26945 5365 26948
rect 5399 26945 5411 26979
rect 5353 26939 5411 26945
rect 5629 26979 5687 26985
rect 5629 26945 5641 26979
rect 5675 26976 5687 26979
rect 5810 26976 5816 26988
rect 5675 26948 5816 26976
rect 5675 26945 5687 26948
rect 5629 26939 5687 26945
rect 5810 26936 5816 26948
rect 5868 26936 5874 26988
rect 6641 26979 6699 26985
rect 6641 26945 6653 26979
rect 6687 26945 6699 26979
rect 6641 26939 6699 26945
rect 7469 26979 7527 26985
rect 7469 26945 7481 26979
rect 7515 26976 7527 26979
rect 7558 26976 7564 26988
rect 7515 26948 7564 26976
rect 7515 26945 7527 26948
rect 7469 26939 7527 26945
rect 5442 26908 5448 26920
rect 4724 26880 5448 26908
rect 1486 26840 1492 26852
rect 1447 26812 1492 26840
rect 1486 26800 1492 26812
rect 1544 26800 1550 26852
rect 4724 26784 4752 26880
rect 5442 26868 5448 26880
rect 5500 26908 5506 26920
rect 6656 26908 6684 26939
rect 7558 26936 7564 26948
rect 7616 26936 7622 26988
rect 7837 26979 7895 26985
rect 7837 26945 7849 26979
rect 7883 26976 7895 26979
rect 7926 26976 7932 26988
rect 7883 26948 7932 26976
rect 7883 26945 7895 26948
rect 7837 26939 7895 26945
rect 7926 26936 7932 26948
rect 7984 26936 7990 26988
rect 8021 26979 8079 26985
rect 8021 26945 8033 26979
rect 8067 26976 8079 26979
rect 8067 26948 8248 26976
rect 8067 26945 8079 26948
rect 8021 26939 8079 26945
rect 5500 26880 6684 26908
rect 5500 26868 5506 26880
rect 7374 26868 7380 26920
rect 7432 26908 7438 26920
rect 7653 26911 7711 26917
rect 7653 26908 7665 26911
rect 7432 26880 7665 26908
rect 7432 26868 7438 26880
rect 7653 26877 7665 26880
rect 7699 26877 7711 26911
rect 7653 26871 7711 26877
rect 7745 26911 7803 26917
rect 7745 26877 7757 26911
rect 7791 26908 7803 26911
rect 8110 26908 8116 26920
rect 7791 26880 8116 26908
rect 7791 26877 7803 26880
rect 7745 26871 7803 26877
rect 8110 26868 8116 26880
rect 8168 26868 8174 26920
rect 5537 26843 5595 26849
rect 5537 26809 5549 26843
rect 5583 26840 5595 26843
rect 5718 26840 5724 26852
rect 5583 26812 5724 26840
rect 5583 26809 5595 26812
rect 5537 26803 5595 26809
rect 5718 26800 5724 26812
rect 5776 26840 5782 26852
rect 6270 26840 6276 26852
rect 5776 26812 6276 26840
rect 5776 26800 5782 26812
rect 6270 26800 6276 26812
rect 6328 26800 6334 26852
rect 6733 26843 6791 26849
rect 6733 26809 6745 26843
rect 6779 26840 6791 26843
rect 7926 26840 7932 26852
rect 6779 26812 7932 26840
rect 6779 26809 6791 26812
rect 6733 26803 6791 26809
rect 7926 26800 7932 26812
rect 7984 26800 7990 26852
rect 8018 26800 8024 26852
rect 8076 26840 8082 26852
rect 8220 26840 8248 26948
rect 8938 26936 8944 26988
rect 8996 26976 9002 26988
rect 9766 26985 9772 26988
rect 9493 26979 9551 26985
rect 9493 26976 9505 26979
rect 8996 26948 9505 26976
rect 8996 26936 9002 26948
rect 9493 26945 9505 26948
rect 9539 26945 9551 26979
rect 9493 26939 9551 26945
rect 9760 26939 9772 26985
rect 9824 26976 9830 26988
rect 9824 26948 9860 26976
rect 9766 26936 9772 26939
rect 9824 26936 9830 26948
rect 10318 26936 10324 26988
rect 10376 26976 10382 26988
rect 11517 26979 11575 26985
rect 11517 26976 11529 26979
rect 10376 26948 11529 26976
rect 10376 26936 10382 26948
rect 11517 26945 11529 26948
rect 11563 26945 11575 26979
rect 11517 26939 11575 26945
rect 12618 26936 12624 26988
rect 12676 26976 12682 26988
rect 12785 26979 12843 26985
rect 12785 26976 12797 26979
rect 12676 26948 12797 26976
rect 12676 26936 12682 26948
rect 12785 26945 12797 26948
rect 12831 26945 12843 26979
rect 14737 26979 14795 26985
rect 14737 26976 14749 26979
rect 12785 26939 12843 26945
rect 14660 26948 14749 26976
rect 11422 26868 11428 26920
rect 11480 26908 11486 26920
rect 12529 26911 12587 26917
rect 12529 26908 12541 26911
rect 11480 26880 12541 26908
rect 11480 26868 11486 26880
rect 12529 26877 12541 26880
rect 12575 26877 12587 26911
rect 14366 26908 14372 26920
rect 12529 26871 12587 26877
rect 13924 26880 14372 26908
rect 11609 26843 11667 26849
rect 11609 26840 11621 26843
rect 8076 26812 8248 26840
rect 10428 26812 11621 26840
rect 8076 26800 8082 26812
rect 4706 26772 4712 26784
rect 4667 26744 4712 26772
rect 4706 26732 4712 26744
rect 4764 26732 4770 26784
rect 6822 26732 6828 26784
rect 6880 26772 6886 26784
rect 7285 26775 7343 26781
rect 7285 26772 7297 26775
rect 6880 26744 7297 26772
rect 6880 26732 6886 26744
rect 7285 26741 7297 26744
rect 7331 26741 7343 26775
rect 7285 26735 7343 26741
rect 9674 26732 9680 26784
rect 9732 26772 9738 26784
rect 10428 26772 10456 26812
rect 11609 26809 11621 26812
rect 11655 26809 11667 26843
rect 11609 26803 11667 26809
rect 9732 26744 10456 26772
rect 9732 26732 9738 26744
rect 12434 26732 12440 26784
rect 12492 26772 12498 26784
rect 13924 26781 13952 26880
rect 14366 26868 14372 26880
rect 14424 26908 14430 26920
rect 14660 26908 14688 26948
rect 14737 26945 14749 26948
rect 14783 26945 14795 26979
rect 15010 26976 15016 26988
rect 14971 26948 15016 26976
rect 14737 26939 14795 26945
rect 15010 26936 15016 26948
rect 15068 26936 15074 26988
rect 15102 26936 15108 26988
rect 15160 26976 15166 26988
rect 15289 26979 15347 26985
rect 15160 26948 15205 26976
rect 15160 26936 15166 26948
rect 15289 26945 15301 26979
rect 15335 26976 15347 26979
rect 15749 26979 15807 26985
rect 15749 26976 15761 26979
rect 15335 26948 15761 26976
rect 15335 26945 15347 26948
rect 15289 26939 15347 26945
rect 15749 26945 15761 26948
rect 15795 26945 15807 26979
rect 15749 26939 15807 26945
rect 16117 26979 16175 26985
rect 16117 26945 16129 26979
rect 16163 26976 16175 26979
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 16163 26948 16865 26976
rect 16163 26945 16175 26948
rect 16117 26939 16175 26945
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 17126 26936 17132 26988
rect 17184 26976 17190 26988
rect 17310 26976 17316 26988
rect 17184 26948 17316 26976
rect 17184 26936 17190 26948
rect 17310 26936 17316 26948
rect 17368 26936 17374 26988
rect 18156 26985 18184 27016
rect 18800 26988 18828 27016
rect 18966 27004 18972 27016
rect 19024 27004 19030 27056
rect 20070 27004 20076 27056
rect 20128 27044 20134 27056
rect 22005 27047 22063 27053
rect 20128 27016 20208 27044
rect 20128 27004 20134 27016
rect 17497 26979 17555 26985
rect 17497 26945 17509 26979
rect 17543 26976 17555 26979
rect 17957 26979 18015 26985
rect 17957 26976 17969 26979
rect 17543 26948 17969 26976
rect 17543 26945 17555 26948
rect 17497 26939 17555 26945
rect 17957 26945 17969 26948
rect 18003 26945 18015 26979
rect 17957 26939 18015 26945
rect 18141 26979 18199 26985
rect 18141 26945 18153 26979
rect 18187 26945 18199 26979
rect 18141 26939 18199 26945
rect 18230 26936 18236 26988
rect 18288 26976 18294 26988
rect 18414 26976 18420 26988
rect 18288 26948 18333 26976
rect 18375 26948 18420 26976
rect 18288 26936 18294 26948
rect 18414 26936 18420 26948
rect 18472 26936 18478 26988
rect 18598 26976 18604 26988
rect 18559 26948 18604 26976
rect 18598 26936 18604 26948
rect 18656 26936 18662 26988
rect 18782 26936 18788 26988
rect 18840 26936 18846 26988
rect 19334 26936 19340 26988
rect 19392 26976 19398 26988
rect 20180 26985 20208 27016
rect 22005 27013 22017 27047
rect 22051 27044 22063 27047
rect 22278 27044 22284 27056
rect 22051 27016 22284 27044
rect 22051 27013 22063 27016
rect 22005 27007 22063 27013
rect 22278 27004 22284 27016
rect 22336 27004 22342 27056
rect 19429 26979 19487 26985
rect 19429 26976 19441 26979
rect 19392 26948 19441 26976
rect 19392 26936 19398 26948
rect 19429 26945 19441 26948
rect 19475 26945 19487 26979
rect 19429 26939 19487 26945
rect 20165 26979 20223 26985
rect 20165 26945 20177 26979
rect 20211 26945 20223 26979
rect 20165 26939 20223 26945
rect 20349 26979 20407 26985
rect 20349 26945 20361 26979
rect 20395 26945 20407 26979
rect 22189 26979 22247 26985
rect 22189 26976 22201 26979
rect 20349 26939 20407 26945
rect 22112 26948 22201 26976
rect 14424 26880 14688 26908
rect 14424 26868 14430 26880
rect 15654 26868 15660 26920
rect 15712 26908 15718 26920
rect 19150 26908 19156 26920
rect 15712 26880 19156 26908
rect 15712 26868 15718 26880
rect 19150 26868 19156 26880
rect 19208 26908 19214 26920
rect 20073 26911 20131 26917
rect 20073 26908 20085 26911
rect 19208 26880 20085 26908
rect 19208 26868 19214 26880
rect 20073 26877 20085 26880
rect 20119 26877 20131 26911
rect 20364 26908 20392 26939
rect 22112 26920 22140 26948
rect 22189 26945 22201 26948
rect 22235 26945 22247 26979
rect 22189 26939 22247 26945
rect 22094 26908 22100 26920
rect 20364 26880 22100 26908
rect 20073 26871 20131 26877
rect 22094 26868 22100 26880
rect 22152 26868 22158 26920
rect 14274 26800 14280 26852
rect 14332 26840 14338 26852
rect 14829 26843 14887 26849
rect 14829 26840 14841 26843
rect 14332 26812 14841 26840
rect 14332 26800 14338 26812
rect 14829 26809 14841 26812
rect 14875 26809 14887 26843
rect 14829 26803 14887 26809
rect 18046 26800 18052 26852
rect 18104 26840 18110 26852
rect 18230 26840 18236 26852
rect 18104 26812 18236 26840
rect 18104 26800 18110 26812
rect 18230 26800 18236 26812
rect 18288 26840 18294 26852
rect 18325 26843 18383 26849
rect 18325 26840 18337 26843
rect 18288 26812 18337 26840
rect 18288 26800 18294 26812
rect 18325 26809 18337 26812
rect 18371 26840 18383 26843
rect 19058 26840 19064 26852
rect 18371 26812 19064 26840
rect 18371 26809 18383 26812
rect 18325 26803 18383 26809
rect 19058 26800 19064 26812
rect 19116 26800 19122 26852
rect 13909 26775 13967 26781
rect 13909 26772 13921 26775
rect 12492 26744 13921 26772
rect 12492 26732 12498 26744
rect 13909 26741 13921 26744
rect 13955 26741 13967 26775
rect 13909 26735 13967 26741
rect 17405 26775 17463 26781
rect 17405 26741 17417 26775
rect 17451 26772 17463 26775
rect 17678 26772 17684 26784
rect 17451 26744 17684 26772
rect 17451 26741 17463 26744
rect 17405 26735 17463 26741
rect 17678 26732 17684 26744
rect 17736 26732 17742 26784
rect 19426 26732 19432 26784
rect 19484 26772 19490 26784
rect 19521 26775 19579 26781
rect 19521 26772 19533 26775
rect 19484 26744 19533 26772
rect 19484 26732 19490 26744
rect 19521 26741 19533 26744
rect 19567 26741 19579 26775
rect 19521 26735 19579 26741
rect 21634 26732 21640 26784
rect 21692 26772 21698 26784
rect 21821 26775 21879 26781
rect 21821 26772 21833 26775
rect 21692 26744 21833 26772
rect 21692 26732 21698 26744
rect 21821 26741 21833 26744
rect 21867 26741 21879 26775
rect 21821 26735 21879 26741
rect 1104 26682 30820 26704
rect 1104 26630 5915 26682
rect 5967 26630 5979 26682
rect 6031 26630 6043 26682
rect 6095 26630 6107 26682
rect 6159 26630 6171 26682
rect 6223 26630 15846 26682
rect 15898 26630 15910 26682
rect 15962 26630 15974 26682
rect 16026 26630 16038 26682
rect 16090 26630 16102 26682
rect 16154 26630 25776 26682
rect 25828 26630 25840 26682
rect 25892 26630 25904 26682
rect 25956 26630 25968 26682
rect 26020 26630 26032 26682
rect 26084 26630 30820 26682
rect 1104 26608 30820 26630
rect 4890 26568 4896 26580
rect 4851 26540 4896 26568
rect 4890 26528 4896 26540
rect 4948 26528 4954 26580
rect 6914 26568 6920 26580
rect 5000 26540 6920 26568
rect 4614 26460 4620 26512
rect 4672 26500 4678 26512
rect 5000 26500 5028 26540
rect 6914 26528 6920 26540
rect 6972 26568 6978 26580
rect 6972 26540 7144 26568
rect 6972 26528 6978 26540
rect 4672 26472 5028 26500
rect 4672 26460 4678 26472
rect 5442 26460 5448 26512
rect 5500 26500 5506 26512
rect 5997 26503 6055 26509
rect 5997 26500 6009 26503
rect 5500 26472 6009 26500
rect 5500 26460 5506 26472
rect 5997 26469 6009 26472
rect 6043 26469 6055 26503
rect 5997 26463 6055 26469
rect 6089 26503 6147 26509
rect 6089 26469 6101 26503
rect 6135 26500 6147 26503
rect 6270 26500 6276 26512
rect 6135 26472 6276 26500
rect 6135 26469 6147 26472
rect 6089 26463 6147 26469
rect 6270 26460 6276 26472
rect 6328 26460 6334 26512
rect 7009 26503 7067 26509
rect 7009 26469 7021 26503
rect 7055 26469 7067 26503
rect 7116 26500 7144 26540
rect 7558 26528 7564 26580
rect 7616 26568 7622 26580
rect 7926 26568 7932 26580
rect 7616 26540 7932 26568
rect 7616 26528 7622 26540
rect 7926 26528 7932 26540
rect 7984 26528 7990 26580
rect 8036 26540 9720 26568
rect 8036 26500 8064 26540
rect 7116 26472 8064 26500
rect 7009 26463 7067 26469
rect 7024 26432 7052 26463
rect 8386 26460 8392 26512
rect 8444 26500 8450 26512
rect 9582 26500 9588 26512
rect 8444 26472 9588 26500
rect 8444 26460 8450 26472
rect 9582 26460 9588 26472
rect 9640 26460 9646 26512
rect 9692 26500 9720 26540
rect 9766 26528 9772 26580
rect 9824 26568 9830 26580
rect 9861 26571 9919 26577
rect 9861 26568 9873 26571
rect 9824 26540 9873 26568
rect 9824 26528 9830 26540
rect 9861 26537 9873 26540
rect 9907 26537 9919 26571
rect 10410 26568 10416 26580
rect 10371 26540 10416 26568
rect 9861 26531 9919 26537
rect 10410 26528 10416 26540
rect 10468 26528 10474 26580
rect 12894 26568 12900 26580
rect 11072 26540 12900 26568
rect 10042 26500 10048 26512
rect 9692 26472 10048 26500
rect 10042 26460 10048 26472
rect 10100 26460 10106 26512
rect 7469 26435 7527 26441
rect 7469 26432 7481 26435
rect 2884 26404 7052 26432
rect 7300 26404 7481 26432
rect 1673 26367 1731 26373
rect 1673 26333 1685 26367
rect 1719 26333 1731 26367
rect 1673 26327 1731 26333
rect 1688 26296 1716 26327
rect 2590 26324 2596 26376
rect 2648 26364 2654 26376
rect 2884 26373 2912 26404
rect 2685 26367 2743 26373
rect 2685 26364 2697 26367
rect 2648 26336 2697 26364
rect 2648 26324 2654 26336
rect 2685 26333 2697 26336
rect 2731 26333 2743 26367
rect 2685 26327 2743 26333
rect 2869 26367 2927 26373
rect 2869 26333 2881 26367
rect 2915 26333 2927 26367
rect 4246 26364 4252 26376
rect 4207 26336 4252 26364
rect 2869 26327 2927 26333
rect 4246 26324 4252 26336
rect 4304 26324 4310 26376
rect 4342 26367 4400 26373
rect 4342 26333 4354 26367
rect 4388 26333 4400 26367
rect 4614 26364 4620 26376
rect 4575 26336 4620 26364
rect 4342 26327 4400 26333
rect 2958 26296 2964 26308
rect 1688 26268 2964 26296
rect 2958 26256 2964 26268
rect 3016 26256 3022 26308
rect 4356 26296 4384 26327
rect 4614 26324 4620 26336
rect 4672 26324 4678 26376
rect 4798 26373 4804 26376
rect 4755 26367 4804 26373
rect 4755 26333 4767 26367
rect 4801 26333 4804 26367
rect 4755 26327 4804 26333
rect 4798 26324 4804 26327
rect 4856 26324 4862 26376
rect 5258 26324 5264 26376
rect 5316 26364 5322 26376
rect 5905 26367 5963 26373
rect 5905 26364 5917 26367
rect 5316 26336 5917 26364
rect 5316 26324 5322 26336
rect 5905 26333 5917 26336
rect 5951 26333 5963 26367
rect 5905 26327 5963 26333
rect 6181 26367 6239 26373
rect 6181 26333 6193 26367
rect 6227 26333 6239 26367
rect 6181 26327 6239 26333
rect 4264 26268 4384 26296
rect 4525 26299 4583 26305
rect 4264 26240 4292 26268
rect 4525 26265 4537 26299
rect 4571 26296 4583 26299
rect 5810 26296 5816 26308
rect 4571 26268 5816 26296
rect 4571 26265 4583 26268
rect 4525 26259 4583 26265
rect 5810 26256 5816 26268
rect 5868 26296 5874 26308
rect 6196 26296 6224 26327
rect 6822 26324 6828 26376
rect 6880 26364 6886 26376
rect 7300 26364 7328 26404
rect 7469 26401 7481 26404
rect 7515 26401 7527 26435
rect 7469 26395 7527 26401
rect 7558 26392 7564 26444
rect 7616 26432 7622 26444
rect 7616 26404 7661 26432
rect 7616 26392 7622 26404
rect 8662 26392 8668 26444
rect 8720 26432 8726 26444
rect 9030 26432 9036 26444
rect 8720 26404 9036 26432
rect 8720 26392 8726 26404
rect 9030 26392 9036 26404
rect 9088 26432 9094 26444
rect 10778 26432 10784 26444
rect 9088 26404 9260 26432
rect 9088 26392 9094 26404
rect 6880 26336 7328 26364
rect 7377 26367 7435 26373
rect 6880 26324 6886 26336
rect 7377 26333 7389 26367
rect 7423 26362 7435 26367
rect 7834 26364 7840 26376
rect 7484 26362 7840 26364
rect 7423 26336 7840 26362
rect 7423 26334 7512 26336
rect 7423 26333 7435 26334
rect 7377 26327 7435 26333
rect 7834 26324 7840 26336
rect 7892 26324 7898 26376
rect 7926 26324 7932 26376
rect 7984 26364 7990 26376
rect 8297 26367 8355 26373
rect 8297 26364 8309 26367
rect 7984 26336 8309 26364
rect 7984 26324 7990 26336
rect 8297 26333 8309 26336
rect 8343 26333 8355 26367
rect 8297 26327 8355 26333
rect 8389 26367 8447 26373
rect 8389 26333 8401 26367
rect 8435 26364 8447 26367
rect 8938 26364 8944 26376
rect 8435 26336 8944 26364
rect 8435 26333 8447 26336
rect 8389 26327 8447 26333
rect 8938 26324 8944 26336
rect 8996 26324 9002 26376
rect 9232 26373 9260 26404
rect 9508 26404 10784 26432
rect 9217 26367 9275 26373
rect 9217 26333 9229 26367
rect 9263 26333 9275 26367
rect 9217 26327 9275 26333
rect 9306 26324 9312 26376
rect 9364 26364 9370 26376
rect 9508 26373 9536 26404
rect 10778 26392 10784 26404
rect 10836 26392 10842 26444
rect 9493 26367 9551 26373
rect 9364 26336 9409 26364
rect 9364 26324 9370 26336
rect 9493 26333 9505 26367
rect 9539 26333 9551 26367
rect 9493 26327 9551 26333
rect 9723 26367 9781 26373
rect 9723 26333 9735 26367
rect 9769 26364 9781 26367
rect 10226 26364 10232 26376
rect 9769 26336 10232 26364
rect 9769 26333 9781 26336
rect 9723 26327 9781 26333
rect 10226 26324 10232 26336
rect 10284 26324 10290 26376
rect 10505 26367 10563 26373
rect 10505 26333 10517 26367
rect 10551 26364 10563 26367
rect 11072 26364 11100 26540
rect 12894 26528 12900 26540
rect 12952 26528 12958 26580
rect 14274 26568 14280 26580
rect 14187 26540 14280 26568
rect 14274 26528 14280 26540
rect 14332 26528 14338 26580
rect 14642 26568 14648 26580
rect 14603 26540 14648 26568
rect 14642 26528 14648 26540
rect 14700 26528 14706 26580
rect 15010 26528 15016 26580
rect 15068 26568 15074 26580
rect 15197 26571 15255 26577
rect 15197 26568 15209 26571
rect 15068 26540 15209 26568
rect 15068 26528 15074 26540
rect 15197 26537 15209 26540
rect 15243 26537 15255 26571
rect 17494 26568 17500 26580
rect 17455 26540 17500 26568
rect 15197 26531 15255 26537
rect 11149 26503 11207 26509
rect 11149 26469 11161 26503
rect 11195 26500 11207 26503
rect 11238 26500 11244 26512
rect 11195 26472 11244 26500
rect 11195 26469 11207 26472
rect 11149 26463 11207 26469
rect 11238 26460 11244 26472
rect 11296 26460 11302 26512
rect 12066 26500 12072 26512
rect 11900 26472 12072 26500
rect 10551 26336 11100 26364
rect 11241 26367 11299 26373
rect 10551 26333 10563 26336
rect 10505 26327 10563 26333
rect 11241 26333 11253 26367
rect 11287 26364 11299 26367
rect 11330 26364 11336 26376
rect 11287 26336 11336 26364
rect 11287 26333 11299 26336
rect 11241 26327 11299 26333
rect 11330 26324 11336 26336
rect 11388 26324 11394 26376
rect 11900 26373 11928 26472
rect 12066 26460 12072 26472
rect 12124 26460 12130 26512
rect 12158 26460 12164 26512
rect 12216 26460 12222 26512
rect 12618 26500 12624 26512
rect 12579 26472 12624 26500
rect 12618 26460 12624 26472
rect 12676 26460 12682 26512
rect 12710 26460 12716 26512
rect 12768 26500 12774 26512
rect 14292 26500 14320 26528
rect 12768 26472 14688 26500
rect 12768 26460 12774 26472
rect 12176 26432 12204 26460
rect 14550 26432 14556 26444
rect 12084 26404 12204 26432
rect 14292 26404 14556 26432
rect 12084 26373 12112 26404
rect 11885 26367 11943 26373
rect 11885 26333 11897 26367
rect 11931 26333 11943 26367
rect 11885 26327 11943 26333
rect 12069 26367 12127 26373
rect 12069 26333 12081 26367
rect 12115 26333 12127 26367
rect 12069 26327 12127 26333
rect 12161 26367 12219 26373
rect 12161 26333 12173 26367
rect 12207 26333 12219 26367
rect 12161 26327 12219 26333
rect 12253 26367 12311 26373
rect 12253 26333 12265 26367
rect 12299 26333 12311 26367
rect 12434 26364 12440 26376
rect 12395 26336 12440 26364
rect 12253 26327 12311 26333
rect 5868 26268 6224 26296
rect 6365 26299 6423 26305
rect 5868 26256 5874 26268
rect 6365 26265 6377 26299
rect 6411 26296 6423 26299
rect 9582 26296 9588 26308
rect 6411 26268 9444 26296
rect 9543 26268 9588 26296
rect 6411 26265 6423 26268
rect 6365 26259 6423 26265
rect 1486 26228 1492 26240
rect 1447 26200 1492 26228
rect 1486 26188 1492 26200
rect 1544 26188 1550 26240
rect 2774 26188 2780 26240
rect 2832 26228 2838 26240
rect 2832 26200 2877 26228
rect 2832 26188 2838 26200
rect 4246 26188 4252 26240
rect 4304 26188 4310 26240
rect 7282 26188 7288 26240
rect 7340 26228 7346 26240
rect 7926 26228 7932 26240
rect 7340 26200 7932 26228
rect 7340 26188 7346 26200
rect 7926 26188 7932 26200
rect 7984 26188 7990 26240
rect 9416 26228 9444 26268
rect 9582 26256 9588 26268
rect 9640 26256 9646 26308
rect 12176 26296 12204 26327
rect 9692 26268 12204 26296
rect 12268 26296 12296 26327
rect 12434 26324 12440 26336
rect 12492 26324 12498 26376
rect 12802 26324 12808 26376
rect 12860 26364 12866 26376
rect 14292 26373 14320 26404
rect 14550 26392 14556 26404
rect 14608 26392 14614 26444
rect 13265 26367 13323 26373
rect 13265 26364 13277 26367
rect 12860 26336 13277 26364
rect 12860 26324 12866 26336
rect 13265 26333 13277 26336
rect 13311 26333 13323 26367
rect 13265 26327 13323 26333
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26333 14335 26367
rect 14277 26327 14335 26333
rect 14461 26367 14519 26373
rect 14461 26333 14473 26367
rect 14507 26333 14519 26367
rect 14660 26364 14688 26472
rect 15105 26367 15163 26373
rect 15105 26364 15117 26367
rect 14660 26336 15117 26364
rect 14461 26327 14519 26333
rect 15105 26333 15117 26336
rect 15151 26333 15163 26367
rect 15212 26364 15240 26531
rect 17494 26528 17500 26540
rect 17552 26528 17558 26580
rect 17957 26571 18015 26577
rect 17957 26537 17969 26571
rect 18003 26568 18015 26571
rect 18138 26568 18144 26580
rect 18003 26540 18144 26568
rect 18003 26537 18015 26540
rect 17957 26531 18015 26537
rect 18138 26528 18144 26540
rect 18196 26528 18202 26580
rect 20714 26528 20720 26580
rect 20772 26568 20778 26580
rect 20809 26571 20867 26577
rect 20809 26568 20821 26571
rect 20772 26540 20821 26568
rect 20772 26528 20778 26540
rect 20809 26537 20821 26540
rect 20855 26537 20867 26571
rect 20809 26531 20867 26537
rect 19334 26460 19340 26512
rect 19392 26500 19398 26512
rect 20625 26503 20683 26509
rect 20625 26500 20637 26503
rect 19392 26472 20637 26500
rect 19392 26460 19398 26472
rect 20625 26469 20637 26472
rect 20671 26469 20683 26503
rect 22094 26500 22100 26512
rect 20625 26463 20683 26469
rect 21008 26472 22100 26500
rect 15562 26392 15568 26444
rect 15620 26432 15626 26444
rect 17310 26432 17316 26444
rect 15620 26404 15976 26432
rect 15620 26392 15626 26404
rect 15948 26373 15976 26404
rect 17144 26404 17316 26432
rect 15749 26367 15807 26373
rect 15749 26364 15761 26367
rect 15212 26336 15761 26364
rect 15105 26327 15163 26333
rect 15749 26333 15761 26336
rect 15795 26333 15807 26367
rect 15749 26327 15807 26333
rect 15933 26367 15991 26373
rect 15933 26333 15945 26367
rect 15979 26333 15991 26367
rect 15933 26327 15991 26333
rect 12526 26296 12532 26308
rect 12268 26268 12532 26296
rect 9692 26228 9720 26268
rect 12526 26256 12532 26268
rect 12584 26256 12590 26308
rect 12986 26256 12992 26308
rect 13044 26296 13050 26308
rect 13081 26299 13139 26305
rect 13081 26296 13093 26299
rect 13044 26268 13093 26296
rect 13044 26256 13050 26268
rect 13081 26265 13093 26268
rect 13127 26265 13139 26299
rect 13081 26259 13139 26265
rect 14366 26256 14372 26308
rect 14424 26296 14430 26308
rect 14476 26296 14504 26327
rect 14424 26268 14504 26296
rect 15841 26299 15899 26305
rect 14424 26256 14430 26268
rect 15841 26265 15853 26299
rect 15887 26296 15899 26299
rect 17034 26296 17040 26308
rect 15887 26268 17040 26296
rect 15887 26265 15899 26268
rect 15841 26259 15899 26265
rect 17034 26256 17040 26268
rect 17092 26256 17098 26308
rect 17144 26305 17172 26404
rect 17310 26392 17316 26404
rect 17368 26392 17374 26444
rect 18046 26392 18052 26444
rect 18104 26432 18110 26444
rect 18509 26435 18567 26441
rect 18509 26432 18521 26435
rect 18104 26404 18521 26432
rect 18104 26392 18110 26404
rect 18509 26401 18521 26404
rect 18555 26432 18567 26435
rect 18782 26432 18788 26444
rect 18555 26404 18788 26432
rect 18555 26401 18567 26404
rect 18509 26395 18567 26401
rect 18782 26392 18788 26404
rect 18840 26392 18846 26444
rect 17494 26324 17500 26376
rect 17552 26364 17558 26376
rect 21008 26373 21036 26472
rect 22094 26460 22100 26472
rect 22152 26500 22158 26512
rect 23017 26503 23075 26509
rect 23017 26500 23029 26503
rect 22152 26472 23029 26500
rect 22152 26460 22158 26472
rect 23017 26469 23029 26472
rect 23063 26469 23075 26503
rect 23017 26463 23075 26469
rect 21634 26432 21640 26444
rect 21595 26404 21640 26432
rect 21634 26392 21640 26404
rect 21692 26392 21698 26444
rect 21913 26435 21971 26441
rect 21913 26401 21925 26435
rect 21959 26432 21971 26435
rect 22370 26432 22376 26444
rect 21959 26404 22376 26432
rect 21959 26401 21971 26404
rect 21913 26395 21971 26401
rect 22066 26376 22094 26404
rect 22370 26392 22376 26404
rect 22428 26392 22434 26444
rect 19245 26367 19303 26373
rect 19245 26364 19257 26367
rect 17552 26336 19257 26364
rect 17552 26324 17558 26336
rect 19245 26333 19257 26336
rect 19291 26333 19303 26367
rect 19245 26327 19303 26333
rect 20901 26367 20959 26373
rect 20901 26333 20913 26367
rect 20947 26333 20959 26367
rect 20901 26327 20959 26333
rect 20993 26367 21051 26373
rect 20993 26333 21005 26367
rect 21039 26333 21051 26367
rect 22066 26336 22100 26376
rect 20993 26327 21051 26333
rect 17129 26299 17187 26305
rect 17129 26265 17141 26299
rect 17175 26265 17187 26299
rect 17310 26296 17316 26308
rect 17271 26268 17316 26296
rect 17129 26259 17187 26265
rect 9416 26200 9720 26228
rect 16942 26188 16948 26240
rect 17000 26228 17006 26240
rect 17144 26228 17172 26259
rect 17310 26256 17316 26268
rect 17368 26256 17374 26308
rect 18417 26299 18475 26305
rect 18417 26265 18429 26299
rect 18463 26296 18475 26299
rect 18690 26296 18696 26308
rect 18463 26268 18696 26296
rect 18463 26265 18475 26268
rect 18417 26259 18475 26265
rect 18690 26256 18696 26268
rect 18748 26296 18754 26308
rect 19337 26299 19395 26305
rect 19337 26296 19349 26299
rect 18748 26268 19349 26296
rect 18748 26256 18754 26268
rect 19337 26265 19349 26268
rect 19383 26265 19395 26299
rect 20916 26296 20944 26327
rect 22094 26324 22100 26336
rect 22152 26324 22158 26376
rect 23106 26364 23112 26376
rect 23067 26336 23112 26364
rect 23106 26324 23112 26336
rect 23164 26324 23170 26376
rect 21266 26296 21272 26308
rect 20916 26268 21272 26296
rect 19337 26259 19395 26265
rect 21266 26256 21272 26268
rect 21324 26296 21330 26308
rect 22002 26296 22008 26308
rect 21324 26268 22008 26296
rect 21324 26256 21330 26268
rect 22002 26256 22008 26268
rect 22060 26256 22066 26308
rect 17000 26200 17172 26228
rect 17000 26188 17006 26200
rect 18230 26188 18236 26240
rect 18288 26228 18294 26240
rect 18325 26231 18383 26237
rect 18325 26228 18337 26231
rect 18288 26200 18337 26228
rect 18288 26188 18294 26200
rect 18325 26197 18337 26200
rect 18371 26197 18383 26231
rect 18325 26191 18383 26197
rect 1104 26138 30820 26160
rect 1104 26086 10880 26138
rect 10932 26086 10944 26138
rect 10996 26086 11008 26138
rect 11060 26086 11072 26138
rect 11124 26086 11136 26138
rect 11188 26086 20811 26138
rect 20863 26086 20875 26138
rect 20927 26086 20939 26138
rect 20991 26086 21003 26138
rect 21055 26086 21067 26138
rect 21119 26086 30820 26138
rect 1104 26064 30820 26086
rect 2777 26027 2835 26033
rect 2777 25993 2789 26027
rect 2823 26024 2835 26027
rect 2958 26024 2964 26036
rect 2823 25996 2964 26024
rect 2823 25993 2835 25996
rect 2777 25987 2835 25993
rect 2958 25984 2964 25996
rect 3016 25984 3022 26036
rect 3602 25984 3608 26036
rect 3660 26024 3666 26036
rect 3789 26027 3847 26033
rect 3789 26024 3801 26027
rect 3660 25996 3801 26024
rect 3660 25984 3666 25996
rect 3789 25993 3801 25996
rect 3835 25993 3847 26027
rect 4430 26024 4436 26036
rect 3789 25987 3847 25993
rect 3988 25996 4436 26024
rect 1673 25891 1731 25897
rect 1673 25857 1685 25891
rect 1719 25857 1731 25891
rect 2682 25888 2688 25900
rect 2643 25860 2688 25888
rect 1673 25851 1731 25857
rect 1688 25820 1716 25851
rect 2682 25848 2688 25860
rect 2740 25848 2746 25900
rect 3988 25897 4016 25996
rect 4430 25984 4436 25996
rect 4488 26024 4494 26036
rect 4798 26024 4804 26036
rect 4488 25996 4804 26024
rect 4488 25984 4494 25996
rect 4798 25984 4804 25996
rect 4856 25984 4862 26036
rect 5810 26024 5816 26036
rect 5000 25996 5816 26024
rect 4157 25959 4215 25965
rect 4157 25925 4169 25959
rect 4203 25956 4215 25959
rect 4706 25956 4712 25968
rect 4203 25928 4712 25956
rect 4203 25925 4215 25928
rect 4157 25919 4215 25925
rect 4706 25916 4712 25928
rect 4764 25916 4770 25968
rect 2869 25891 2927 25897
rect 2869 25857 2881 25891
rect 2915 25857 2927 25891
rect 2869 25851 2927 25857
rect 3968 25891 4026 25897
rect 3968 25857 3980 25891
rect 4014 25857 4026 25891
rect 3968 25851 4026 25857
rect 2774 25820 2780 25832
rect 1688 25792 2780 25820
rect 2774 25780 2780 25792
rect 2832 25780 2838 25832
rect 2884 25820 2912 25851
rect 4062 25848 4068 25900
rect 4120 25888 4126 25900
rect 4120 25860 4165 25888
rect 4120 25848 4126 25860
rect 4246 25848 4252 25900
rect 4304 25897 4310 25900
rect 4304 25891 4343 25897
rect 4331 25857 4343 25891
rect 4304 25851 4343 25857
rect 4433 25891 4491 25897
rect 4433 25857 4445 25891
rect 4479 25888 4491 25891
rect 4522 25888 4528 25900
rect 4479 25860 4528 25888
rect 4479 25857 4491 25860
rect 4433 25851 4491 25857
rect 4304 25848 4310 25851
rect 4522 25848 4528 25860
rect 4580 25848 4586 25900
rect 4890 25888 4896 25900
rect 4803 25860 4896 25888
rect 4890 25848 4896 25860
rect 4948 25888 4954 25900
rect 5000 25888 5028 25996
rect 5810 25984 5816 25996
rect 5868 25984 5874 26036
rect 7098 25984 7104 26036
rect 7156 26024 7162 26036
rect 7466 26024 7472 26036
rect 7156 25996 7472 26024
rect 7156 25984 7162 25996
rect 7466 25984 7472 25996
rect 7524 25984 7530 26036
rect 7745 26027 7803 26033
rect 7745 25993 7757 26027
rect 7791 26024 7803 26027
rect 8018 26024 8024 26036
rect 7791 25996 8024 26024
rect 7791 25993 7803 25996
rect 7745 25987 7803 25993
rect 8018 25984 8024 25996
rect 8076 25984 8082 26036
rect 8941 26027 8999 26033
rect 8941 26024 8953 26027
rect 8128 25996 8953 26024
rect 5721 25959 5779 25965
rect 5721 25925 5733 25959
rect 5767 25956 5779 25959
rect 6546 25956 6552 25968
rect 5767 25928 6552 25956
rect 5767 25925 5779 25928
rect 5721 25919 5779 25925
rect 6546 25916 6552 25928
rect 6604 25916 6610 25968
rect 8128 25956 8156 25996
rect 8941 25993 8953 25996
rect 8987 25993 8999 26027
rect 8941 25987 8999 25993
rect 9214 25984 9220 26036
rect 9272 26024 9278 26036
rect 9309 26027 9367 26033
rect 9309 26024 9321 26027
rect 9272 25996 9321 26024
rect 9272 25984 9278 25996
rect 9309 25993 9321 25996
rect 9355 25993 9367 26027
rect 9309 25987 9367 25993
rect 9401 26027 9459 26033
rect 9401 25993 9413 26027
rect 9447 26024 9459 26027
rect 9582 26024 9588 26036
rect 9447 25996 9588 26024
rect 9447 25993 9459 25996
rect 9401 25987 9459 25993
rect 9582 25984 9588 25996
rect 9640 25984 9646 26036
rect 11514 26024 11520 26036
rect 11475 25996 11520 26024
rect 11514 25984 11520 25996
rect 11572 25984 11578 26036
rect 14921 26027 14979 26033
rect 14921 25993 14933 26027
rect 14967 26024 14979 26027
rect 15102 26024 15108 26036
rect 14967 25996 15108 26024
rect 14967 25993 14979 25996
rect 14921 25987 14979 25993
rect 15102 25984 15108 25996
rect 15160 25984 15166 26036
rect 16669 26027 16727 26033
rect 16669 25993 16681 26027
rect 16715 25993 16727 26027
rect 16669 25987 16727 25993
rect 10229 25959 10287 25965
rect 10229 25956 10241 25959
rect 6656 25928 8156 25956
rect 8312 25928 10241 25956
rect 4948 25860 5028 25888
rect 4948 25848 4954 25860
rect 5074 25848 5080 25900
rect 5132 25888 5138 25900
rect 6365 25891 6423 25897
rect 6365 25888 6377 25891
rect 5132 25860 6377 25888
rect 5132 25848 5138 25860
rect 6365 25857 6377 25860
rect 6411 25857 6423 25891
rect 6365 25851 6423 25857
rect 6656 25820 6684 25928
rect 6917 25891 6975 25897
rect 6917 25857 6929 25891
rect 6963 25888 6975 25891
rect 7742 25888 7748 25900
rect 6963 25860 7748 25888
rect 6963 25857 6975 25860
rect 6917 25851 6975 25857
rect 7742 25848 7748 25860
rect 7800 25848 7806 25900
rect 7929 25891 7987 25897
rect 7929 25857 7941 25891
rect 7975 25857 7987 25891
rect 7929 25851 7987 25857
rect 7006 25820 7012 25832
rect 2884 25792 6684 25820
rect 6967 25792 7012 25820
rect 7006 25780 7012 25792
rect 7064 25780 7070 25832
rect 7193 25823 7251 25829
rect 7193 25789 7205 25823
rect 7239 25820 7251 25823
rect 7558 25820 7564 25832
rect 7239 25792 7564 25820
rect 7239 25789 7251 25792
rect 7193 25783 7251 25789
rect 7558 25780 7564 25792
rect 7616 25820 7622 25832
rect 7834 25820 7840 25832
rect 7616 25792 7840 25820
rect 7616 25780 7622 25792
rect 7834 25780 7840 25792
rect 7892 25780 7898 25832
rect 4985 25755 5043 25761
rect 4985 25721 4997 25755
rect 5031 25752 5043 25755
rect 6822 25752 6828 25764
rect 5031 25724 6828 25752
rect 5031 25721 5043 25724
rect 4985 25715 5043 25721
rect 6822 25712 6828 25724
rect 6880 25712 6886 25764
rect 7944 25752 7972 25851
rect 8018 25848 8024 25900
rect 8076 25888 8082 25900
rect 8312 25897 8340 25928
rect 10229 25925 10241 25928
rect 10275 25925 10287 25959
rect 12710 25956 12716 25968
rect 10229 25919 10287 25925
rect 11716 25928 12716 25956
rect 8297 25891 8355 25897
rect 8076 25860 8121 25888
rect 8076 25848 8082 25860
rect 8297 25857 8309 25891
rect 8343 25857 8355 25891
rect 8297 25851 8355 25857
rect 8956 25860 9628 25888
rect 8202 25780 8208 25832
rect 8260 25820 8266 25832
rect 8956 25820 8984 25860
rect 8260 25792 8984 25820
rect 8260 25780 8266 25792
rect 9398 25780 9404 25832
rect 9456 25820 9462 25832
rect 9493 25823 9551 25829
rect 9493 25820 9505 25823
rect 9456 25792 9505 25820
rect 9456 25780 9462 25792
rect 9493 25789 9505 25792
rect 9539 25789 9551 25823
rect 9600 25820 9628 25860
rect 9950 25848 9956 25900
rect 10008 25888 10014 25900
rect 10321 25891 10379 25897
rect 10321 25888 10333 25891
rect 10008 25860 10333 25888
rect 10008 25848 10014 25860
rect 10321 25857 10333 25860
rect 10367 25857 10379 25891
rect 10321 25851 10379 25857
rect 10778 25848 10784 25900
rect 10836 25888 10842 25900
rect 11716 25897 11744 25928
rect 12710 25916 12716 25928
rect 12768 25916 12774 25968
rect 13814 25956 13820 25968
rect 12820 25928 13820 25956
rect 10965 25891 11023 25897
rect 10965 25888 10977 25891
rect 10836 25860 10977 25888
rect 10836 25848 10842 25860
rect 10965 25857 10977 25860
rect 11011 25857 11023 25891
rect 10965 25851 11023 25857
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25857 11759 25891
rect 11977 25891 12035 25897
rect 11977 25888 11989 25891
rect 11701 25851 11759 25857
rect 11808 25860 11989 25888
rect 11808 25820 11836 25860
rect 11977 25857 11989 25860
rect 12023 25857 12035 25891
rect 11977 25851 12035 25857
rect 12069 25891 12127 25897
rect 12069 25857 12081 25891
rect 12115 25888 12127 25891
rect 12158 25888 12164 25900
rect 12115 25860 12164 25888
rect 12115 25857 12127 25860
rect 12069 25851 12127 25857
rect 12158 25848 12164 25860
rect 12216 25848 12222 25900
rect 12253 25891 12311 25897
rect 12253 25857 12265 25891
rect 12299 25888 12311 25891
rect 12342 25888 12348 25900
rect 12299 25860 12348 25888
rect 12299 25857 12311 25860
rect 12253 25851 12311 25857
rect 12342 25848 12348 25860
rect 12400 25848 12406 25900
rect 9600 25792 11836 25820
rect 11885 25823 11943 25829
rect 9493 25783 9551 25789
rect 11885 25789 11897 25823
rect 11931 25789 11943 25823
rect 12526 25820 12532 25832
rect 11885 25783 11943 25789
rect 12176 25792 12532 25820
rect 10873 25755 10931 25761
rect 10873 25752 10885 25755
rect 7944 25724 9444 25752
rect 1486 25684 1492 25696
rect 1447 25656 1492 25684
rect 1486 25644 1492 25656
rect 1544 25644 1550 25696
rect 5629 25687 5687 25693
rect 5629 25653 5641 25687
rect 5675 25684 5687 25687
rect 5810 25684 5816 25696
rect 5675 25656 5816 25684
rect 5675 25653 5687 25656
rect 5629 25647 5687 25653
rect 5810 25644 5816 25656
rect 5868 25644 5874 25696
rect 6365 25687 6423 25693
rect 6365 25653 6377 25687
rect 6411 25684 6423 25687
rect 6549 25687 6607 25693
rect 6549 25684 6561 25687
rect 6411 25656 6561 25684
rect 6411 25653 6423 25656
rect 6365 25647 6423 25653
rect 6549 25653 6561 25656
rect 6595 25653 6607 25687
rect 6549 25647 6607 25653
rect 7926 25644 7932 25696
rect 7984 25684 7990 25696
rect 8205 25687 8263 25693
rect 8205 25684 8217 25687
rect 7984 25656 8217 25684
rect 7984 25644 7990 25656
rect 8205 25653 8217 25656
rect 8251 25653 8263 25687
rect 9416 25684 9444 25724
rect 9646 25724 10885 25752
rect 9646 25684 9674 25724
rect 10873 25721 10885 25724
rect 10919 25721 10931 25755
rect 11900 25752 11928 25783
rect 12176 25752 12204 25792
rect 12526 25780 12532 25792
rect 12584 25780 12590 25832
rect 12820 25752 12848 25928
rect 13814 25916 13820 25928
rect 13872 25916 13878 25968
rect 15746 25956 15752 25968
rect 15707 25928 15752 25956
rect 15746 25916 15752 25928
rect 15804 25916 15810 25968
rect 15933 25959 15991 25965
rect 15933 25925 15945 25959
rect 15979 25956 15991 25959
rect 16684 25956 16712 25987
rect 17034 25984 17040 26036
rect 17092 26024 17098 26036
rect 17129 26027 17187 26033
rect 17129 26024 17141 26027
rect 17092 25996 17141 26024
rect 17092 25984 17098 25996
rect 17129 25993 17141 25996
rect 17175 25993 17187 26027
rect 18322 26024 18328 26036
rect 18283 25996 18328 26024
rect 17129 25987 17187 25993
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 19334 26024 19340 26036
rect 19260 25996 19340 26024
rect 15979 25928 16712 25956
rect 18693 25959 18751 25965
rect 15979 25925 15991 25928
rect 15933 25919 15991 25925
rect 18693 25925 18705 25959
rect 18739 25956 18751 25959
rect 18782 25956 18788 25968
rect 18739 25928 18788 25956
rect 18739 25925 18751 25928
rect 18693 25919 18751 25925
rect 18782 25916 18788 25928
rect 18840 25916 18846 25968
rect 13354 25848 13360 25900
rect 13412 25888 13418 25900
rect 13918 25891 13976 25897
rect 13918 25888 13930 25891
rect 13412 25860 13930 25888
rect 13412 25848 13418 25860
rect 13918 25857 13930 25860
rect 13964 25857 13976 25891
rect 13918 25851 13976 25857
rect 14366 25848 14372 25900
rect 14424 25888 14430 25900
rect 14829 25891 14887 25897
rect 14829 25888 14841 25891
rect 14424 25860 14841 25888
rect 14424 25848 14430 25860
rect 14829 25857 14841 25860
rect 14875 25857 14887 25891
rect 14829 25851 14887 25857
rect 14185 25823 14243 25829
rect 14185 25789 14197 25823
rect 14231 25820 14243 25823
rect 15194 25820 15200 25832
rect 14231 25792 15200 25820
rect 14231 25789 14243 25792
rect 14185 25783 14243 25789
rect 15194 25780 15200 25792
rect 15252 25780 15258 25832
rect 15764 25820 15792 25916
rect 16482 25848 16488 25900
rect 16540 25888 16546 25900
rect 17037 25891 17095 25897
rect 17037 25888 17049 25891
rect 16540 25860 17049 25888
rect 16540 25848 16546 25860
rect 17037 25857 17049 25860
rect 17083 25857 17095 25891
rect 19260 25888 19288 25996
rect 19334 25984 19340 25996
rect 19392 26024 19398 26036
rect 19518 26024 19524 26036
rect 19392 25996 19524 26024
rect 19392 25984 19398 25996
rect 19518 25984 19524 25996
rect 19576 25984 19582 26036
rect 22278 26024 22284 26036
rect 20732 25996 22284 26024
rect 17037 25851 17095 25857
rect 17144 25860 19288 25888
rect 17144 25820 17172 25860
rect 19334 25848 19340 25900
rect 19392 25888 19398 25900
rect 19613 25891 19671 25897
rect 19613 25888 19625 25891
rect 19392 25860 19625 25888
rect 19392 25848 19398 25860
rect 19613 25857 19625 25860
rect 19659 25857 19671 25891
rect 19613 25851 19671 25857
rect 20533 25891 20591 25897
rect 20533 25857 20545 25891
rect 20579 25888 20591 25891
rect 20622 25888 20628 25900
rect 20579 25860 20628 25888
rect 20579 25857 20591 25860
rect 20533 25851 20591 25857
rect 20622 25848 20628 25860
rect 20680 25848 20686 25900
rect 20732 25897 20760 25996
rect 22278 25984 22284 25996
rect 22336 26024 22342 26036
rect 23198 26024 23204 26036
rect 22336 25996 23204 26024
rect 22336 25984 22342 25996
rect 23198 25984 23204 25996
rect 23256 25984 23262 26036
rect 20898 25956 20904 25968
rect 20811 25928 20904 25956
rect 20824 25897 20852 25928
rect 20898 25916 20904 25928
rect 20956 25956 20962 25968
rect 21174 25956 21180 25968
rect 20956 25928 21180 25956
rect 20956 25916 20962 25928
rect 21174 25916 21180 25928
rect 21232 25916 21238 25968
rect 20717 25891 20775 25897
rect 20717 25857 20729 25891
rect 20763 25857 20775 25891
rect 20717 25851 20775 25857
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25857 20867 25891
rect 21082 25888 21088 25900
rect 21043 25860 21088 25888
rect 20809 25851 20867 25857
rect 21082 25848 21088 25860
rect 21140 25848 21146 25900
rect 21450 25848 21456 25900
rect 21508 25888 21514 25900
rect 22077 25891 22135 25897
rect 22077 25888 22089 25891
rect 21508 25860 22089 25888
rect 21508 25848 21514 25860
rect 22077 25857 22089 25860
rect 22123 25857 22135 25891
rect 22077 25851 22135 25857
rect 15764 25792 17172 25820
rect 17313 25823 17371 25829
rect 17313 25789 17325 25823
rect 17359 25820 17371 25823
rect 18046 25820 18052 25832
rect 17359 25792 18052 25820
rect 17359 25789 17371 25792
rect 17313 25783 17371 25789
rect 18046 25780 18052 25792
rect 18104 25780 18110 25832
rect 18690 25780 18696 25832
rect 18748 25820 18754 25832
rect 18785 25823 18843 25829
rect 18785 25820 18797 25823
rect 18748 25792 18797 25820
rect 18748 25780 18754 25792
rect 18785 25789 18797 25792
rect 18831 25789 18843 25823
rect 18785 25783 18843 25789
rect 18874 25780 18880 25832
rect 18932 25820 18938 25832
rect 19886 25820 19892 25832
rect 18932 25792 18977 25820
rect 19847 25792 19892 25820
rect 18932 25780 18938 25792
rect 19886 25780 19892 25792
rect 19944 25780 19950 25832
rect 19981 25823 20039 25829
rect 19981 25789 19993 25823
rect 20027 25820 20039 25823
rect 20346 25820 20352 25832
rect 20027 25792 20352 25820
rect 20027 25789 20039 25792
rect 19981 25783 20039 25789
rect 20346 25780 20352 25792
rect 20404 25780 20410 25832
rect 20901 25823 20959 25829
rect 20901 25789 20913 25823
rect 20947 25820 20959 25823
rect 21174 25820 21180 25832
rect 20947 25792 21180 25820
rect 20947 25789 20959 25792
rect 20901 25783 20959 25789
rect 21174 25780 21180 25792
rect 21232 25780 21238 25832
rect 21818 25820 21824 25832
rect 21779 25792 21824 25820
rect 21818 25780 21824 25792
rect 21876 25780 21882 25832
rect 17494 25752 17500 25764
rect 11900 25724 12204 25752
rect 12406 25724 12848 25752
rect 14936 25724 17500 25752
rect 10873 25715 10931 25721
rect 9416 25656 9674 25684
rect 8205 25647 8263 25653
rect 9950 25644 9956 25696
rect 10008 25684 10014 25696
rect 12406 25684 12434 25724
rect 10008 25656 12434 25684
rect 10008 25644 10014 25656
rect 12618 25644 12624 25696
rect 12676 25684 12682 25696
rect 12805 25687 12863 25693
rect 12805 25684 12817 25687
rect 12676 25656 12817 25684
rect 12676 25644 12682 25656
rect 12805 25653 12817 25656
rect 12851 25684 12863 25687
rect 14936 25684 14964 25724
rect 17494 25712 17500 25724
rect 17552 25712 17558 25764
rect 12851 25656 14964 25684
rect 12851 25653 12863 25656
rect 12805 25647 12863 25653
rect 15746 25644 15752 25696
rect 15804 25684 15810 25696
rect 16117 25687 16175 25693
rect 16117 25684 16129 25687
rect 15804 25656 16129 25684
rect 15804 25644 15810 25656
rect 16117 25653 16129 25656
rect 16163 25653 16175 25687
rect 16117 25647 16175 25653
rect 19426 25644 19432 25696
rect 19484 25684 19490 25696
rect 19705 25687 19763 25693
rect 19705 25684 19717 25687
rect 19484 25656 19717 25684
rect 19484 25644 19490 25656
rect 19705 25653 19717 25656
rect 19751 25653 19763 25687
rect 19705 25647 19763 25653
rect 20073 25687 20131 25693
rect 20073 25653 20085 25687
rect 20119 25684 20131 25687
rect 20990 25684 20996 25696
rect 20119 25656 20996 25684
rect 20119 25653 20131 25656
rect 20073 25647 20131 25653
rect 20990 25644 20996 25656
rect 21048 25644 21054 25696
rect 21266 25684 21272 25696
rect 21227 25656 21272 25684
rect 21266 25644 21272 25656
rect 21324 25644 21330 25696
rect 22462 25644 22468 25696
rect 22520 25684 22526 25696
rect 23106 25684 23112 25696
rect 22520 25656 23112 25684
rect 22520 25644 22526 25656
rect 23106 25644 23112 25656
rect 23164 25684 23170 25696
rect 23201 25687 23259 25693
rect 23201 25684 23213 25687
rect 23164 25656 23213 25684
rect 23164 25644 23170 25656
rect 23201 25653 23213 25656
rect 23247 25653 23259 25687
rect 23201 25647 23259 25653
rect 1104 25594 30820 25616
rect 1104 25542 5915 25594
rect 5967 25542 5979 25594
rect 6031 25542 6043 25594
rect 6095 25542 6107 25594
rect 6159 25542 6171 25594
rect 6223 25542 15846 25594
rect 15898 25542 15910 25594
rect 15962 25542 15974 25594
rect 16026 25542 16038 25594
rect 16090 25542 16102 25594
rect 16154 25542 25776 25594
rect 25828 25542 25840 25594
rect 25892 25542 25904 25594
rect 25956 25542 25968 25594
rect 26020 25542 26032 25594
rect 26084 25542 30820 25594
rect 1104 25520 30820 25542
rect 4062 25440 4068 25492
rect 4120 25480 4126 25492
rect 6362 25480 6368 25492
rect 4120 25452 6368 25480
rect 4120 25440 4126 25452
rect 6362 25440 6368 25452
rect 6420 25440 6426 25492
rect 6914 25440 6920 25492
rect 6972 25480 6978 25492
rect 7282 25480 7288 25492
rect 6972 25452 7288 25480
rect 6972 25440 6978 25452
rect 7282 25440 7288 25452
rect 7340 25440 7346 25492
rect 7834 25440 7840 25492
rect 7892 25480 7898 25492
rect 9398 25480 9404 25492
rect 7892 25452 9404 25480
rect 7892 25440 7898 25452
rect 9398 25440 9404 25452
rect 9456 25440 9462 25492
rect 11057 25483 11115 25489
rect 11057 25449 11069 25483
rect 11103 25480 11115 25483
rect 11790 25480 11796 25492
rect 11103 25452 11796 25480
rect 11103 25449 11115 25452
rect 11057 25443 11115 25449
rect 11790 25440 11796 25452
rect 11848 25440 11854 25492
rect 12066 25440 12072 25492
rect 12124 25480 12130 25492
rect 12342 25480 12348 25492
rect 12124 25452 12348 25480
rect 12124 25440 12130 25452
rect 12342 25440 12348 25452
rect 12400 25440 12406 25492
rect 12805 25483 12863 25489
rect 12805 25449 12817 25483
rect 12851 25480 12863 25483
rect 13354 25480 13360 25492
rect 12851 25452 13360 25480
rect 12851 25449 12863 25452
rect 12805 25443 12863 25449
rect 13354 25440 13360 25452
rect 13412 25440 13418 25492
rect 16390 25440 16396 25492
rect 16448 25480 16454 25492
rect 16666 25480 16672 25492
rect 16448 25452 16672 25480
rect 16448 25440 16454 25452
rect 16666 25440 16672 25452
rect 16724 25440 16730 25492
rect 16758 25440 16764 25492
rect 16816 25480 16822 25492
rect 17034 25480 17040 25492
rect 16816 25452 17040 25480
rect 16816 25440 16822 25452
rect 17034 25440 17040 25452
rect 17092 25440 17098 25492
rect 17310 25440 17316 25492
rect 17368 25480 17374 25492
rect 17773 25483 17831 25489
rect 17773 25480 17785 25483
rect 17368 25452 17785 25480
rect 17368 25440 17374 25452
rect 17773 25449 17785 25452
rect 17819 25449 17831 25483
rect 19610 25480 19616 25492
rect 19571 25452 19616 25480
rect 17773 25443 17831 25449
rect 19610 25440 19616 25452
rect 19668 25440 19674 25492
rect 21361 25483 21419 25489
rect 21361 25449 21373 25483
rect 21407 25480 21419 25483
rect 21450 25480 21456 25492
rect 21407 25452 21456 25480
rect 21407 25449 21419 25452
rect 21361 25443 21419 25449
rect 21450 25440 21456 25452
rect 21508 25440 21514 25492
rect 23198 25480 23204 25492
rect 23159 25452 23204 25480
rect 23198 25440 23204 25452
rect 23256 25440 23262 25492
rect 5629 25415 5687 25421
rect 5629 25381 5641 25415
rect 5675 25412 5687 25415
rect 5718 25412 5724 25424
rect 5675 25384 5724 25412
rect 5675 25381 5687 25384
rect 5629 25375 5687 25381
rect 5718 25372 5724 25384
rect 5776 25372 5782 25424
rect 7558 25412 7564 25424
rect 7471 25384 7564 25412
rect 7558 25372 7564 25384
rect 7616 25412 7622 25424
rect 10318 25412 10324 25424
rect 7616 25384 10324 25412
rect 7616 25372 7622 25384
rect 10318 25372 10324 25384
rect 10376 25372 10382 25424
rect 10778 25412 10784 25424
rect 10739 25384 10784 25412
rect 10778 25372 10784 25384
rect 10836 25372 10842 25424
rect 14829 25415 14887 25421
rect 14829 25381 14841 25415
rect 14875 25412 14887 25415
rect 15194 25412 15200 25424
rect 14875 25384 15200 25412
rect 14875 25381 14887 25384
rect 14829 25375 14887 25381
rect 15194 25372 15200 25384
rect 15252 25412 15258 25424
rect 15654 25412 15660 25424
rect 15252 25384 15660 25412
rect 15252 25372 15258 25384
rect 15654 25372 15660 25384
rect 15712 25412 15718 25424
rect 15712 25384 21864 25412
rect 15712 25372 15718 25384
rect 21836 25356 21864 25384
rect 7926 25304 7932 25356
rect 7984 25344 7990 25356
rect 9401 25347 9459 25353
rect 9401 25344 9413 25347
rect 7984 25316 9413 25344
rect 7984 25304 7990 25316
rect 9401 25313 9413 25316
rect 9447 25313 9459 25347
rect 9401 25307 9459 25313
rect 10502 25304 10508 25356
rect 10560 25344 10566 25356
rect 10689 25347 10747 25353
rect 10689 25344 10701 25347
rect 10560 25316 10701 25344
rect 10560 25304 10566 25316
rect 10689 25313 10701 25316
rect 10735 25313 10747 25347
rect 10689 25307 10747 25313
rect 11882 25304 11888 25356
rect 11940 25344 11946 25356
rect 12342 25344 12348 25356
rect 11940 25316 12348 25344
rect 11940 25304 11946 25316
rect 12342 25304 12348 25316
rect 12400 25304 12406 25356
rect 12437 25347 12495 25353
rect 12437 25313 12449 25347
rect 12483 25344 12495 25347
rect 12526 25344 12532 25356
rect 12483 25316 12532 25344
rect 12483 25313 12495 25316
rect 12437 25307 12495 25313
rect 12526 25304 12532 25316
rect 12584 25304 12590 25356
rect 13538 25304 13544 25356
rect 13596 25344 13602 25356
rect 13596 25316 16620 25344
rect 13596 25304 13602 25316
rect 4249 25279 4307 25285
rect 4249 25245 4261 25279
rect 4295 25276 4307 25279
rect 4338 25276 4344 25288
rect 4295 25248 4344 25276
rect 4295 25245 4307 25248
rect 4249 25239 4307 25245
rect 4338 25236 4344 25248
rect 4396 25276 4402 25288
rect 5810 25276 5816 25288
rect 4396 25248 5816 25276
rect 4396 25236 4402 25248
rect 5810 25236 5816 25248
rect 5868 25276 5874 25288
rect 6181 25279 6239 25285
rect 6181 25276 6193 25279
rect 5868 25248 6193 25276
rect 5868 25236 5874 25248
rect 6181 25245 6193 25248
rect 6227 25276 6239 25279
rect 6227 25248 6684 25276
rect 6227 25245 6239 25248
rect 6181 25239 6239 25245
rect 6656 25220 6684 25248
rect 6914 25236 6920 25288
rect 6972 25276 6978 25288
rect 8297 25279 8355 25285
rect 8297 25276 8309 25279
rect 6972 25248 8309 25276
rect 6972 25236 6978 25248
rect 8297 25245 8309 25248
rect 8343 25245 8355 25279
rect 9122 25276 9128 25288
rect 9083 25248 9128 25276
rect 8297 25239 8355 25245
rect 9122 25236 9128 25248
rect 9180 25236 9186 25288
rect 9217 25279 9275 25285
rect 9217 25245 9229 25279
rect 9263 25245 9275 25279
rect 9217 25239 9275 25245
rect 9493 25279 9551 25285
rect 9493 25245 9505 25279
rect 9539 25276 9551 25279
rect 9674 25276 9680 25288
rect 9539 25248 9680 25276
rect 9539 25245 9551 25248
rect 9493 25239 9551 25245
rect 4516 25211 4574 25217
rect 4516 25177 4528 25211
rect 4562 25208 4574 25211
rect 4798 25208 4804 25220
rect 4562 25180 4804 25208
rect 4562 25177 4574 25180
rect 4516 25171 4574 25177
rect 4798 25168 4804 25180
rect 4856 25168 4862 25220
rect 6454 25217 6460 25220
rect 6448 25171 6460 25217
rect 6512 25208 6518 25220
rect 6512 25180 6548 25208
rect 6454 25168 6460 25171
rect 6512 25168 6518 25180
rect 6638 25168 6644 25220
rect 6696 25168 6702 25220
rect 8018 25168 8024 25220
rect 8076 25208 8082 25220
rect 9232 25208 9260 25239
rect 9674 25236 9680 25248
rect 9732 25236 9738 25288
rect 10597 25279 10655 25285
rect 10597 25245 10609 25279
rect 10643 25245 10655 25279
rect 10597 25239 10655 25245
rect 10873 25279 10931 25285
rect 10873 25245 10885 25279
rect 10919 25276 10931 25279
rect 11606 25276 11612 25288
rect 10919 25248 11612 25276
rect 10919 25245 10931 25248
rect 10873 25239 10931 25245
rect 8076 25180 9260 25208
rect 8076 25168 8082 25180
rect 8202 25140 8208 25152
rect 8163 25112 8208 25140
rect 8202 25100 8208 25112
rect 8260 25100 8266 25152
rect 8570 25100 8576 25152
rect 8628 25140 8634 25152
rect 8941 25143 8999 25149
rect 8941 25140 8953 25143
rect 8628 25112 8953 25140
rect 8628 25100 8634 25112
rect 8941 25109 8953 25112
rect 8987 25109 8999 25143
rect 10612 25140 10640 25239
rect 11606 25236 11612 25248
rect 11664 25236 11670 25288
rect 12066 25276 12072 25288
rect 12027 25248 12072 25276
rect 12066 25236 12072 25248
rect 12124 25236 12130 25288
rect 12253 25279 12311 25285
rect 12253 25245 12265 25279
rect 12299 25245 12311 25279
rect 12618 25276 12624 25288
rect 12579 25248 12624 25276
rect 12253 25239 12311 25245
rect 11330 25168 11336 25220
rect 11388 25208 11394 25220
rect 12268 25208 12296 25239
rect 12618 25236 12624 25248
rect 12676 25236 12682 25288
rect 13262 25276 13268 25288
rect 13223 25248 13268 25276
rect 13262 25236 13268 25248
rect 13320 25236 13326 25288
rect 13354 25236 13360 25288
rect 13412 25276 13418 25288
rect 13412 25248 13457 25276
rect 13412 25236 13418 25248
rect 15286 25236 15292 25288
rect 15344 25276 15350 25288
rect 16592 25276 16620 25316
rect 16666 25304 16672 25356
rect 16724 25344 16730 25356
rect 18046 25344 18052 25356
rect 16724 25316 18052 25344
rect 16724 25304 16730 25316
rect 18046 25304 18052 25316
rect 18104 25344 18110 25356
rect 18325 25347 18383 25353
rect 18325 25344 18337 25347
rect 18104 25316 18337 25344
rect 18104 25304 18110 25316
rect 18325 25313 18337 25316
rect 18371 25313 18383 25347
rect 18325 25307 18383 25313
rect 19889 25347 19947 25353
rect 19889 25313 19901 25347
rect 19935 25344 19947 25347
rect 20070 25344 20076 25356
rect 19935 25316 20076 25344
rect 19935 25313 19947 25316
rect 19889 25307 19947 25313
rect 20070 25304 20076 25316
rect 20128 25304 20134 25356
rect 20990 25344 20996 25356
rect 20951 25316 20996 25344
rect 20990 25304 20996 25316
rect 21048 25304 21054 25356
rect 21818 25344 21824 25356
rect 21779 25316 21824 25344
rect 21818 25304 21824 25316
rect 21876 25304 21882 25356
rect 19518 25276 19524 25288
rect 15344 25248 15389 25276
rect 16592 25248 19380 25276
rect 19479 25248 19524 25276
rect 15344 25236 15350 25248
rect 11388 25180 12296 25208
rect 11388 25168 11394 25180
rect 12986 25168 12992 25220
rect 13044 25208 13050 25220
rect 14645 25211 14703 25217
rect 14645 25208 14657 25211
rect 13044 25180 14657 25208
rect 13044 25168 13050 25180
rect 14645 25177 14657 25180
rect 14691 25177 14703 25211
rect 16945 25211 17003 25217
rect 16945 25208 16957 25211
rect 14645 25171 14703 25177
rect 16776 25180 16957 25208
rect 11514 25140 11520 25152
rect 10612 25112 11520 25140
rect 8941 25103 8999 25109
rect 11514 25100 11520 25112
rect 11572 25100 11578 25152
rect 15378 25140 15384 25152
rect 15339 25112 15384 25140
rect 15378 25100 15384 25112
rect 15436 25100 15442 25152
rect 16482 25100 16488 25152
rect 16540 25140 16546 25152
rect 16776 25140 16804 25180
rect 16945 25177 16957 25180
rect 16991 25177 17003 25211
rect 16945 25171 17003 25177
rect 18046 25168 18052 25220
rect 18104 25208 18110 25220
rect 18233 25211 18291 25217
rect 18233 25208 18245 25211
rect 18104 25180 18245 25208
rect 18104 25168 18110 25180
rect 18233 25177 18245 25180
rect 18279 25177 18291 25211
rect 19352 25208 19380 25248
rect 19518 25236 19524 25248
rect 19576 25236 19582 25288
rect 19981 25279 20039 25285
rect 19981 25245 19993 25279
rect 20027 25276 20039 25279
rect 20530 25276 20536 25288
rect 20027 25248 20536 25276
rect 20027 25245 20039 25248
rect 19981 25239 20039 25245
rect 20530 25236 20536 25248
rect 20588 25236 20594 25288
rect 20622 25236 20628 25288
rect 20680 25276 20686 25288
rect 20809 25279 20867 25285
rect 20680 25248 20773 25276
rect 20680 25236 20686 25248
rect 20809 25245 20821 25279
rect 20855 25245 20867 25279
rect 20809 25239 20867 25245
rect 20640 25208 20668 25236
rect 19352 25180 20668 25208
rect 18233 25171 18291 25177
rect 16540 25112 16804 25140
rect 16853 25143 16911 25149
rect 16540 25100 16546 25112
rect 16853 25109 16865 25143
rect 16899 25140 16911 25143
rect 17034 25140 17040 25152
rect 16899 25112 17040 25140
rect 16899 25109 16911 25112
rect 16853 25103 16911 25109
rect 17034 25100 17040 25112
rect 17092 25100 17098 25152
rect 17218 25100 17224 25152
rect 17276 25140 17282 25152
rect 17313 25143 17371 25149
rect 17313 25140 17325 25143
rect 17276 25112 17325 25140
rect 17276 25100 17282 25112
rect 17313 25109 17325 25112
rect 17359 25109 17371 25143
rect 18138 25140 18144 25152
rect 18099 25112 18144 25140
rect 17313 25103 17371 25109
rect 18138 25100 18144 25112
rect 18196 25100 18202 25152
rect 20165 25143 20223 25149
rect 20165 25109 20177 25143
rect 20211 25140 20223 25143
rect 20346 25140 20352 25152
rect 20211 25112 20352 25140
rect 20211 25109 20223 25112
rect 20165 25103 20223 25109
rect 20346 25100 20352 25112
rect 20404 25100 20410 25152
rect 20824 25140 20852 25239
rect 20898 25236 20904 25288
rect 20956 25276 20962 25288
rect 20956 25248 21001 25276
rect 20956 25236 20962 25248
rect 21082 25236 21088 25288
rect 21140 25276 21146 25288
rect 21177 25279 21235 25285
rect 21177 25276 21189 25279
rect 21140 25248 21189 25276
rect 21140 25236 21146 25248
rect 21177 25245 21189 25248
rect 21223 25245 21235 25279
rect 21177 25239 21235 25245
rect 21192 25208 21220 25239
rect 21266 25236 21272 25288
rect 21324 25276 21330 25288
rect 22077 25279 22135 25285
rect 22077 25276 22089 25279
rect 21324 25248 22089 25276
rect 21324 25236 21330 25248
rect 22077 25245 22089 25248
rect 22123 25245 22135 25279
rect 22077 25239 22135 25245
rect 29178 25236 29184 25288
rect 29236 25276 29242 25288
rect 29825 25279 29883 25285
rect 29825 25276 29837 25279
rect 29236 25248 29837 25276
rect 29236 25236 29242 25248
rect 29825 25245 29837 25248
rect 29871 25245 29883 25279
rect 29825 25239 29883 25245
rect 21542 25208 21548 25220
rect 21192 25180 21548 25208
rect 21542 25168 21548 25180
rect 21600 25168 21606 25220
rect 22462 25140 22468 25152
rect 20824 25112 22468 25140
rect 22462 25100 22468 25112
rect 22520 25100 22526 25152
rect 30006 25140 30012 25152
rect 29967 25112 30012 25140
rect 30006 25100 30012 25112
rect 30064 25100 30070 25152
rect 1104 25050 30820 25072
rect 1104 24998 10880 25050
rect 10932 24998 10944 25050
rect 10996 24998 11008 25050
rect 11060 24998 11072 25050
rect 11124 24998 11136 25050
rect 11188 24998 20811 25050
rect 20863 24998 20875 25050
rect 20927 24998 20939 25050
rect 20991 24998 21003 25050
rect 21055 24998 21067 25050
rect 21119 24998 30820 25050
rect 1104 24976 30820 24998
rect 4798 24936 4804 24948
rect 4759 24908 4804 24936
rect 4798 24896 4804 24908
rect 4856 24896 4862 24948
rect 7650 24936 7656 24948
rect 7611 24908 7656 24936
rect 7650 24896 7656 24908
rect 7708 24896 7714 24948
rect 9309 24939 9367 24945
rect 9309 24905 9321 24939
rect 9355 24936 9367 24939
rect 9582 24936 9588 24948
rect 9355 24908 9588 24936
rect 9355 24905 9367 24908
rect 9309 24899 9367 24905
rect 9582 24896 9588 24908
rect 9640 24896 9646 24948
rect 10686 24896 10692 24948
rect 10744 24936 10750 24948
rect 11698 24936 11704 24948
rect 10744 24908 11704 24936
rect 10744 24896 10750 24908
rect 11698 24896 11704 24908
rect 11756 24936 11762 24948
rect 12158 24936 12164 24948
rect 11756 24908 12164 24936
rect 11756 24896 11762 24908
rect 12158 24896 12164 24908
rect 12216 24896 12222 24948
rect 12897 24939 12955 24945
rect 12897 24905 12909 24939
rect 12943 24936 12955 24939
rect 13262 24936 13268 24948
rect 12943 24908 13268 24936
rect 12943 24905 12955 24908
rect 12897 24899 12955 24905
rect 8404 24840 8892 24868
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24769 1731 24803
rect 2682 24800 2688 24812
rect 2643 24772 2688 24800
rect 1673 24763 1731 24769
rect 1688 24732 1716 24763
rect 2682 24760 2688 24772
rect 2740 24760 2746 24812
rect 2869 24803 2927 24809
rect 2869 24769 2881 24803
rect 2915 24769 2927 24803
rect 2869 24763 2927 24769
rect 4065 24803 4123 24809
rect 4065 24769 4077 24803
rect 4111 24800 4123 24803
rect 4154 24800 4160 24812
rect 4111 24772 4160 24800
rect 4111 24769 4123 24772
rect 4065 24763 4123 24769
rect 2777 24735 2835 24741
rect 2777 24732 2789 24735
rect 1688 24704 2789 24732
rect 2777 24701 2789 24704
rect 2823 24701 2835 24735
rect 2777 24695 2835 24701
rect 1486 24664 1492 24676
rect 1447 24636 1492 24664
rect 1486 24624 1492 24636
rect 1544 24624 1550 24676
rect 2884 24596 2912 24763
rect 4154 24760 4160 24772
rect 4212 24760 4218 24812
rect 4249 24803 4307 24809
rect 4249 24769 4261 24803
rect 4295 24800 4307 24803
rect 4522 24800 4528 24812
rect 4295 24772 4528 24800
rect 4295 24769 4307 24772
rect 4249 24763 4307 24769
rect 4522 24760 4528 24772
rect 4580 24760 4586 24812
rect 4617 24803 4675 24809
rect 4617 24769 4629 24803
rect 4663 24800 4675 24803
rect 4890 24800 4896 24812
rect 4663 24772 4896 24800
rect 4663 24769 4675 24772
rect 4617 24763 4675 24769
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 5721 24803 5779 24809
rect 5721 24769 5733 24803
rect 5767 24800 5779 24803
rect 6365 24803 6423 24809
rect 6365 24800 6377 24803
rect 5767 24772 6377 24800
rect 5767 24769 5779 24772
rect 5721 24763 5779 24769
rect 6365 24769 6377 24772
rect 6411 24769 6423 24803
rect 6365 24763 6423 24769
rect 6730 24760 6736 24812
rect 6788 24800 6794 24812
rect 6788 24772 6833 24800
rect 6788 24760 6794 24772
rect 7374 24760 7380 24812
rect 7432 24800 7438 24812
rect 7650 24800 7656 24812
rect 7432 24772 7656 24800
rect 7432 24760 7438 24772
rect 7650 24760 7656 24772
rect 7708 24800 7714 24812
rect 8404 24800 8432 24840
rect 8570 24800 8576 24812
rect 7708 24772 8432 24800
rect 8531 24772 8576 24800
rect 7708 24760 7714 24772
rect 8570 24760 8576 24772
rect 8628 24760 8634 24812
rect 8757 24803 8815 24809
rect 8757 24769 8769 24803
rect 8803 24769 8815 24803
rect 8864 24800 8892 24840
rect 10152 24840 10916 24868
rect 8941 24803 8999 24809
rect 8941 24800 8953 24803
rect 8864 24772 8953 24800
rect 8757 24763 8815 24769
rect 8941 24769 8953 24772
rect 8987 24769 8999 24803
rect 8941 24763 8999 24769
rect 9125 24803 9183 24809
rect 9125 24769 9137 24803
rect 9171 24800 9183 24803
rect 10152 24800 10180 24840
rect 9171 24772 10180 24800
rect 9171 24769 9183 24772
rect 9125 24763 9183 24769
rect 4338 24732 4344 24744
rect 4299 24704 4344 24732
rect 4338 24692 4344 24704
rect 4396 24692 4402 24744
rect 4430 24692 4436 24744
rect 4488 24732 4494 24744
rect 4488 24704 4533 24732
rect 4488 24692 4494 24704
rect 6822 24692 6828 24744
rect 6880 24732 6886 24744
rect 7742 24732 7748 24744
rect 6880 24704 7604 24732
rect 7703 24704 7748 24732
rect 6880 24692 6886 24704
rect 4062 24624 4068 24676
rect 4120 24664 4126 24676
rect 5537 24667 5595 24673
rect 5537 24664 5549 24667
rect 4120 24636 5549 24664
rect 4120 24624 4126 24636
rect 5537 24633 5549 24636
rect 5583 24633 5595 24667
rect 7285 24667 7343 24673
rect 7285 24664 7297 24667
rect 5537 24627 5595 24633
rect 5644 24636 7297 24664
rect 5644 24596 5672 24636
rect 7285 24633 7297 24636
rect 7331 24633 7343 24667
rect 7576 24664 7604 24704
rect 7742 24692 7748 24704
rect 7800 24692 7806 24744
rect 7834 24692 7840 24744
rect 7892 24732 7898 24744
rect 7892 24704 7937 24732
rect 7892 24692 7898 24704
rect 8772 24664 8800 24763
rect 10226 24760 10232 24812
rect 10284 24800 10290 24812
rect 10413 24803 10471 24809
rect 10284 24772 10329 24800
rect 10284 24760 10290 24772
rect 10413 24769 10425 24803
rect 10459 24769 10471 24803
rect 10413 24763 10471 24769
rect 10505 24803 10563 24809
rect 10505 24769 10517 24803
rect 10551 24800 10563 24803
rect 10686 24800 10692 24812
rect 10551 24772 10692 24800
rect 10551 24769 10563 24772
rect 10505 24763 10563 24769
rect 8849 24735 8907 24741
rect 8849 24701 8861 24735
rect 8895 24701 8907 24735
rect 8849 24695 8907 24701
rect 7576 24636 8800 24664
rect 7285 24627 7343 24633
rect 2884 24568 5672 24596
rect 6365 24599 6423 24605
rect 6365 24565 6377 24599
rect 6411 24596 6423 24599
rect 6641 24599 6699 24605
rect 6641 24596 6653 24599
rect 6411 24568 6653 24596
rect 6411 24565 6423 24568
rect 6365 24559 6423 24565
rect 6641 24565 6653 24568
rect 6687 24596 6699 24599
rect 7098 24596 7104 24608
rect 6687 24568 7104 24596
rect 6687 24565 6699 24568
rect 6641 24559 6699 24565
rect 7098 24556 7104 24568
rect 7156 24556 7162 24608
rect 8110 24556 8116 24608
rect 8168 24596 8174 24608
rect 8864 24596 8892 24695
rect 10318 24692 10324 24744
rect 10376 24732 10382 24744
rect 10428 24732 10456 24763
rect 10686 24760 10692 24772
rect 10744 24760 10750 24812
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24769 10839 24803
rect 10888 24800 10916 24840
rect 11238 24800 11244 24812
rect 10888 24772 11244 24800
rect 10781 24763 10839 24769
rect 10376 24704 10456 24732
rect 10597 24735 10655 24741
rect 10376 24692 10382 24704
rect 10597 24701 10609 24735
rect 10643 24732 10655 24735
rect 10643 24704 10732 24732
rect 10643 24701 10655 24704
rect 10597 24695 10655 24701
rect 10704 24676 10732 24704
rect 10686 24624 10692 24676
rect 10744 24624 10750 24676
rect 8168 24568 8892 24596
rect 10796 24596 10824 24763
rect 11238 24760 11244 24772
rect 11296 24760 11302 24812
rect 11422 24760 11428 24812
rect 11480 24800 11486 24812
rect 11517 24803 11575 24809
rect 11517 24800 11529 24803
rect 11480 24772 11529 24800
rect 11480 24760 11486 24772
rect 11517 24769 11529 24772
rect 11563 24769 11575 24803
rect 11773 24803 11831 24809
rect 11773 24800 11785 24803
rect 11517 24763 11575 24769
rect 11624 24772 11785 24800
rect 10965 24735 11023 24741
rect 10965 24701 10977 24735
rect 11011 24732 11023 24735
rect 11624 24732 11652 24772
rect 11773 24769 11785 24772
rect 11819 24769 11831 24803
rect 11773 24763 11831 24769
rect 11011 24704 11652 24732
rect 11011 24701 11023 24704
rect 10965 24695 11023 24701
rect 12912 24596 12940 24899
rect 13262 24896 13268 24908
rect 13320 24896 13326 24948
rect 13630 24896 13636 24948
rect 13688 24936 13694 24948
rect 17126 24936 17132 24948
rect 13688 24908 17132 24936
rect 13688 24896 13694 24908
rect 17126 24896 17132 24908
rect 17184 24896 17190 24948
rect 17862 24936 17868 24948
rect 17823 24908 17868 24936
rect 17862 24896 17868 24908
rect 17920 24896 17926 24948
rect 19886 24936 19892 24948
rect 19847 24908 19892 24936
rect 19886 24896 19892 24908
rect 19944 24936 19950 24948
rect 20993 24939 21051 24945
rect 19944 24908 20392 24936
rect 19944 24896 19950 24908
rect 15197 24871 15255 24877
rect 15197 24837 15209 24871
rect 15243 24868 15255 24871
rect 15243 24840 15792 24868
rect 15243 24837 15255 24840
rect 15197 24831 15255 24837
rect 14734 24800 14740 24812
rect 14695 24772 14740 24800
rect 14734 24760 14740 24772
rect 14792 24760 14798 24812
rect 14829 24803 14887 24809
rect 14829 24769 14841 24803
rect 14875 24769 14887 24803
rect 14829 24763 14887 24769
rect 15013 24803 15071 24809
rect 15013 24769 15025 24803
rect 15059 24800 15071 24803
rect 15562 24800 15568 24812
rect 15059 24772 15568 24800
rect 15059 24769 15071 24772
rect 15013 24763 15071 24769
rect 14844 24732 14872 24763
rect 15562 24760 15568 24772
rect 15620 24760 15626 24812
rect 15657 24803 15715 24809
rect 15657 24769 15669 24803
rect 15703 24769 15715 24803
rect 15764 24800 15792 24840
rect 17494 24828 17500 24880
rect 17552 24868 17558 24880
rect 18874 24868 18880 24880
rect 17552 24840 18880 24868
rect 17552 24828 17558 24840
rect 18874 24828 18880 24840
rect 18932 24828 18938 24880
rect 20364 24877 20392 24908
rect 20993 24905 21005 24939
rect 21039 24936 21051 24939
rect 21174 24936 21180 24948
rect 21039 24908 21180 24936
rect 21039 24905 21051 24908
rect 20993 24899 21051 24905
rect 21174 24896 21180 24908
rect 21232 24896 21238 24948
rect 20349 24871 20407 24877
rect 20349 24837 20361 24871
rect 20395 24837 20407 24871
rect 20349 24831 20407 24837
rect 20530 24828 20536 24880
rect 20588 24868 20594 24880
rect 21726 24868 21732 24880
rect 20588 24840 21732 24868
rect 20588 24828 20594 24840
rect 18046 24800 18052 24812
rect 15764 24772 18052 24800
rect 15657 24763 15715 24769
rect 15286 24732 15292 24744
rect 14844 24704 15292 24732
rect 15028 24676 15056 24704
rect 15286 24692 15292 24704
rect 15344 24692 15350 24744
rect 15470 24732 15476 24744
rect 15396 24704 15476 24732
rect 15010 24624 15016 24676
rect 15068 24624 15074 24676
rect 10796 24568 12940 24596
rect 8168 24556 8174 24568
rect 15102 24556 15108 24608
rect 15160 24596 15166 24608
rect 15396 24596 15424 24704
rect 15470 24692 15476 24704
rect 15528 24732 15534 24744
rect 15672 24732 15700 24763
rect 18046 24760 18052 24772
rect 18104 24760 18110 24812
rect 19061 24803 19119 24809
rect 19061 24769 19073 24803
rect 19107 24800 19119 24803
rect 19334 24800 19340 24812
rect 19107 24772 19340 24800
rect 19107 24769 19119 24772
rect 19061 24763 19119 24769
rect 19334 24760 19340 24772
rect 19392 24760 19398 24812
rect 19613 24803 19671 24809
rect 19613 24769 19625 24803
rect 19659 24769 19671 24803
rect 19613 24763 19671 24769
rect 19705 24803 19763 24809
rect 19705 24769 19717 24803
rect 19751 24800 19763 24803
rect 19978 24800 19984 24812
rect 19751 24772 19984 24800
rect 19751 24769 19763 24772
rect 19705 24763 19763 24769
rect 15528 24704 15700 24732
rect 15528 24692 15534 24704
rect 16942 24692 16948 24744
rect 17000 24732 17006 24744
rect 17589 24735 17647 24741
rect 17589 24732 17601 24735
rect 17000 24704 17601 24732
rect 17000 24692 17006 24704
rect 17589 24701 17601 24704
rect 17635 24701 17647 24735
rect 17589 24695 17647 24701
rect 17773 24735 17831 24741
rect 17773 24701 17785 24735
rect 17819 24732 17831 24735
rect 17862 24732 17868 24744
rect 17819 24704 17868 24732
rect 17819 24701 17831 24704
rect 17773 24695 17831 24701
rect 17862 24692 17868 24704
rect 17920 24692 17926 24744
rect 19150 24692 19156 24744
rect 19208 24732 19214 24744
rect 19628 24732 19656 24763
rect 19978 24760 19984 24772
rect 20036 24800 20042 24812
rect 20162 24800 20168 24812
rect 20036 24772 20168 24800
rect 20036 24760 20042 24772
rect 20162 24760 20168 24772
rect 20220 24760 20226 24812
rect 20824 24809 20852 24840
rect 21726 24828 21732 24840
rect 21784 24828 21790 24880
rect 20809 24803 20867 24809
rect 20809 24769 20821 24803
rect 20855 24769 20867 24803
rect 20809 24763 20867 24769
rect 19208 24704 19656 24732
rect 19889 24735 19947 24741
rect 19208 24692 19214 24704
rect 19889 24701 19901 24735
rect 19935 24701 19947 24735
rect 19889 24695 19947 24701
rect 19610 24624 19616 24676
rect 19668 24664 19674 24676
rect 19904 24664 19932 24695
rect 20530 24692 20536 24744
rect 20588 24732 20594 24744
rect 20625 24735 20683 24741
rect 20625 24732 20637 24735
rect 20588 24704 20637 24732
rect 20588 24692 20594 24704
rect 20625 24701 20637 24704
rect 20671 24701 20683 24735
rect 20625 24695 20683 24701
rect 19668 24636 19932 24664
rect 19668 24624 19674 24636
rect 15160 24568 15424 24596
rect 15160 24556 15166 24568
rect 15470 24556 15476 24608
rect 15528 24596 15534 24608
rect 15749 24599 15807 24605
rect 15749 24596 15761 24599
rect 15528 24568 15761 24596
rect 15528 24556 15534 24568
rect 15749 24565 15761 24568
rect 15795 24565 15807 24599
rect 15749 24559 15807 24565
rect 18233 24599 18291 24605
rect 18233 24565 18245 24599
rect 18279 24596 18291 24599
rect 18874 24596 18880 24608
rect 18279 24568 18880 24596
rect 18279 24565 18291 24568
rect 18233 24559 18291 24565
rect 18874 24556 18880 24568
rect 18932 24556 18938 24608
rect 18966 24556 18972 24608
rect 19024 24596 19030 24608
rect 20438 24596 20444 24608
rect 19024 24568 19069 24596
rect 20399 24568 20444 24596
rect 19024 24556 19030 24568
rect 20438 24556 20444 24568
rect 20496 24556 20502 24608
rect 1104 24506 30820 24528
rect 1104 24454 5915 24506
rect 5967 24454 5979 24506
rect 6031 24454 6043 24506
rect 6095 24454 6107 24506
rect 6159 24454 6171 24506
rect 6223 24454 15846 24506
rect 15898 24454 15910 24506
rect 15962 24454 15974 24506
rect 16026 24454 16038 24506
rect 16090 24454 16102 24506
rect 16154 24454 25776 24506
rect 25828 24454 25840 24506
rect 25892 24454 25904 24506
rect 25956 24454 25968 24506
rect 26020 24454 26032 24506
rect 26084 24454 30820 24506
rect 1104 24432 30820 24454
rect 5074 24392 5080 24404
rect 3712 24364 5080 24392
rect 2777 24259 2835 24265
rect 2777 24256 2789 24259
rect 1688 24228 2789 24256
rect 1688 24197 1716 24228
rect 2777 24225 2789 24228
rect 2823 24225 2835 24259
rect 2777 24219 2835 24225
rect 1673 24191 1731 24197
rect 1673 24157 1685 24191
rect 1719 24157 1731 24191
rect 2682 24188 2688 24200
rect 2595 24160 2688 24188
rect 1673 24151 1731 24157
rect 2682 24148 2688 24160
rect 2740 24148 2746 24200
rect 2869 24191 2927 24197
rect 2869 24157 2881 24191
rect 2915 24188 2927 24191
rect 3712 24188 3740 24364
rect 5074 24352 5080 24364
rect 5132 24352 5138 24404
rect 6365 24395 6423 24401
rect 6365 24361 6377 24395
rect 6411 24392 6423 24395
rect 6454 24392 6460 24404
rect 6411 24364 6460 24392
rect 6411 24361 6423 24364
rect 6365 24355 6423 24361
rect 6454 24352 6460 24364
rect 6512 24352 6518 24404
rect 6638 24352 6644 24404
rect 6696 24392 6702 24404
rect 6696 24364 7696 24392
rect 6696 24352 6702 24364
rect 4338 24284 4344 24336
rect 4396 24284 4402 24336
rect 4522 24284 4528 24336
rect 4580 24324 4586 24336
rect 5902 24324 5908 24336
rect 4580 24296 5908 24324
rect 4580 24284 4586 24296
rect 5902 24284 5908 24296
rect 5960 24284 5966 24336
rect 7558 24324 7564 24336
rect 7208 24296 7564 24324
rect 4249 24259 4307 24265
rect 4249 24225 4261 24259
rect 4295 24256 4307 24259
rect 4356 24256 4384 24284
rect 5166 24256 5172 24268
rect 4295 24228 5172 24256
rect 4295 24225 4307 24228
rect 4249 24219 4307 24225
rect 5166 24216 5172 24228
rect 5224 24216 5230 24268
rect 5920 24256 5948 24284
rect 5828 24228 5948 24256
rect 5997 24259 6055 24265
rect 2915 24160 3740 24188
rect 3973 24191 4031 24197
rect 2915 24157 2927 24160
rect 2869 24151 2927 24157
rect 3973 24157 3985 24191
rect 4019 24157 4031 24191
rect 3973 24151 4031 24157
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24157 4215 24191
rect 4338 24188 4344 24200
rect 4299 24160 4344 24188
rect 4157 24151 4215 24157
rect 2700 24120 2728 24148
rect 3510 24120 3516 24132
rect 2700 24092 3516 24120
rect 3510 24080 3516 24092
rect 3568 24080 3574 24132
rect 1486 24052 1492 24064
rect 1447 24024 1492 24052
rect 1486 24012 1492 24024
rect 1544 24012 1550 24064
rect 3786 24052 3792 24064
rect 3747 24024 3792 24052
rect 3786 24012 3792 24024
rect 3844 24012 3850 24064
rect 3988 24052 4016 24151
rect 4172 24120 4200 24151
rect 4338 24148 4344 24160
rect 4396 24148 4402 24200
rect 4522 24188 4528 24200
rect 4483 24160 4528 24188
rect 4522 24148 4528 24160
rect 4580 24148 4586 24200
rect 4985 24191 5043 24197
rect 4985 24157 4997 24191
rect 5031 24190 5043 24191
rect 5031 24188 5120 24190
rect 5258 24188 5264 24200
rect 5031 24162 5264 24188
rect 5031 24157 5043 24162
rect 5092 24160 5264 24162
rect 4985 24151 5043 24157
rect 5258 24148 5264 24160
rect 5316 24148 5322 24200
rect 5534 24148 5540 24200
rect 5592 24188 5598 24200
rect 5828 24197 5856 24228
rect 5997 24225 6009 24259
rect 6043 24256 6055 24259
rect 6546 24256 6552 24268
rect 6043 24228 6552 24256
rect 6043 24225 6055 24228
rect 5997 24219 6055 24225
rect 6546 24216 6552 24228
rect 6604 24216 6610 24268
rect 5629 24191 5687 24197
rect 5629 24188 5641 24191
rect 5592 24160 5641 24188
rect 5592 24148 5598 24160
rect 5629 24157 5641 24160
rect 5675 24157 5687 24191
rect 5629 24151 5687 24157
rect 5813 24191 5871 24197
rect 5813 24157 5825 24191
rect 5859 24157 5871 24191
rect 5813 24151 5871 24157
rect 5902 24148 5908 24200
rect 5960 24188 5966 24200
rect 6181 24191 6239 24197
rect 5960 24160 6005 24188
rect 5960 24148 5966 24160
rect 6181 24157 6193 24191
rect 6227 24188 6239 24191
rect 7208 24188 7236 24296
rect 7558 24284 7564 24296
rect 7616 24284 7622 24336
rect 7668 24324 7696 24364
rect 7742 24352 7748 24404
rect 7800 24392 7806 24404
rect 8113 24395 8171 24401
rect 8113 24392 8125 24395
rect 7800 24364 8125 24392
rect 7800 24352 7806 24364
rect 8113 24361 8125 24364
rect 8159 24361 8171 24395
rect 8113 24355 8171 24361
rect 10686 24352 10692 24404
rect 10744 24392 10750 24404
rect 11974 24392 11980 24404
rect 10744 24364 11980 24392
rect 10744 24352 10750 24364
rect 11974 24352 11980 24364
rect 12032 24352 12038 24404
rect 14277 24395 14335 24401
rect 14277 24361 14289 24395
rect 14323 24392 14335 24395
rect 14734 24392 14740 24404
rect 14323 24364 14740 24392
rect 14323 24361 14335 24364
rect 14277 24355 14335 24361
rect 14734 24352 14740 24364
rect 14792 24352 14798 24404
rect 17862 24392 17868 24404
rect 15028 24364 15608 24392
rect 17823 24364 17868 24392
rect 7668 24296 9812 24324
rect 7653 24259 7711 24265
rect 7653 24225 7665 24259
rect 7699 24256 7711 24259
rect 8110 24256 8116 24268
rect 7699 24228 8116 24256
rect 7699 24225 7711 24228
rect 7653 24219 7711 24225
rect 8110 24216 8116 24228
rect 8168 24216 8174 24268
rect 9784 24265 9812 24296
rect 9769 24259 9827 24265
rect 9769 24225 9781 24259
rect 9815 24225 9827 24259
rect 9769 24219 9827 24225
rect 10778 24216 10784 24268
rect 10836 24256 10842 24268
rect 12342 24256 12348 24268
rect 10836 24228 12204 24256
rect 12303 24228 12348 24256
rect 10836 24216 10842 24228
rect 7374 24188 7380 24200
rect 6227 24160 7236 24188
rect 7335 24160 7380 24188
rect 6227 24157 6239 24160
rect 6181 24151 6239 24157
rect 7374 24148 7380 24160
rect 7432 24148 7438 24200
rect 7561 24191 7619 24197
rect 7561 24157 7573 24191
rect 7607 24157 7619 24191
rect 7561 24151 7619 24157
rect 4246 24120 4252 24132
rect 4172 24092 4252 24120
rect 4246 24080 4252 24092
rect 4304 24120 4310 24132
rect 4430 24120 4436 24132
rect 4304 24092 4436 24120
rect 4304 24080 4310 24092
rect 4430 24080 4436 24092
rect 4488 24080 4494 24132
rect 5077 24123 5135 24129
rect 5077 24089 5089 24123
rect 5123 24120 5135 24123
rect 7576 24120 7604 24151
rect 7742 24148 7748 24200
rect 7800 24188 7806 24200
rect 7929 24191 7987 24197
rect 7800 24160 7845 24188
rect 7800 24148 7806 24160
rect 7929 24157 7941 24191
rect 7975 24188 7987 24191
rect 9033 24191 9091 24197
rect 9033 24188 9045 24191
rect 7975 24160 9045 24188
rect 7975 24157 7987 24160
rect 7929 24151 7987 24157
rect 9033 24157 9045 24160
rect 9079 24157 9091 24191
rect 9033 24151 9091 24157
rect 9122 24148 9128 24200
rect 9180 24188 9186 24200
rect 12066 24188 12072 24200
rect 9180 24160 9225 24188
rect 12027 24160 12072 24188
rect 9180 24148 9186 24160
rect 12066 24148 12072 24160
rect 12124 24148 12130 24200
rect 12176 24188 12204 24228
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 12437 24259 12495 24265
rect 12437 24225 12449 24259
rect 12483 24256 12495 24259
rect 12526 24256 12532 24268
rect 12483 24228 12532 24256
rect 12483 24225 12495 24228
rect 12437 24219 12495 24225
rect 12526 24216 12532 24228
rect 12584 24216 12590 24268
rect 15028 24256 15056 24364
rect 15580 24336 15608 24364
rect 17862 24352 17868 24364
rect 17920 24352 17926 24404
rect 18966 24392 18972 24404
rect 18432 24364 18972 24392
rect 15378 24324 15384 24336
rect 14844 24228 15056 24256
rect 15120 24296 15384 24324
rect 12253 24191 12311 24197
rect 12253 24188 12265 24191
rect 12176 24160 12265 24188
rect 12253 24157 12265 24160
rect 12299 24157 12311 24191
rect 12253 24151 12311 24157
rect 5123 24092 7604 24120
rect 5123 24089 5135 24092
rect 5077 24083 5135 24089
rect 9858 24080 9864 24132
rect 9916 24120 9922 24132
rect 10014 24123 10072 24129
rect 10014 24120 10026 24123
rect 9916 24092 10026 24120
rect 9916 24080 9922 24092
rect 10014 24089 10026 24092
rect 10060 24089 10072 24123
rect 10014 24083 10072 24089
rect 12158 24080 12164 24132
rect 12216 24120 12222 24132
rect 12360 24120 12388 24216
rect 12621 24191 12679 24197
rect 12621 24157 12633 24191
rect 12667 24188 12679 24191
rect 14185 24191 14243 24197
rect 14185 24188 14197 24191
rect 12667 24160 14197 24188
rect 12667 24157 12679 24160
rect 12621 24151 12679 24157
rect 14185 24157 14197 24160
rect 14231 24188 14243 24191
rect 14274 24188 14280 24200
rect 14231 24160 14280 24188
rect 14231 24157 14243 24160
rect 14185 24151 14243 24157
rect 14274 24148 14280 24160
rect 14332 24148 14338 24200
rect 14369 24191 14427 24197
rect 14369 24157 14381 24191
rect 14415 24188 14427 24191
rect 14642 24188 14648 24200
rect 14415 24160 14648 24188
rect 14415 24157 14427 24160
rect 14369 24151 14427 24157
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 14844 24197 14872 24228
rect 14829 24191 14887 24197
rect 14829 24157 14841 24191
rect 14875 24157 14887 24191
rect 14829 24151 14887 24157
rect 14977 24191 15035 24197
rect 14977 24157 14989 24191
rect 15023 24188 15035 24191
rect 15120 24188 15148 24296
rect 15378 24284 15384 24296
rect 15436 24284 15442 24336
rect 15562 24284 15568 24336
rect 15620 24324 15626 24336
rect 18432 24324 18460 24364
rect 18966 24352 18972 24364
rect 19024 24352 19030 24404
rect 19610 24352 19616 24404
rect 19668 24392 19674 24404
rect 19797 24395 19855 24401
rect 19797 24392 19809 24395
rect 19668 24364 19809 24392
rect 19668 24352 19674 24364
rect 19797 24361 19809 24364
rect 19843 24361 19855 24395
rect 19797 24355 19855 24361
rect 15620 24296 18460 24324
rect 15620 24284 15626 24296
rect 15470 24256 15476 24268
rect 15212 24228 15476 24256
rect 15212 24197 15240 24228
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 16025 24259 16083 24265
rect 16025 24225 16037 24259
rect 16071 24256 16083 24259
rect 16390 24256 16396 24268
rect 16071 24228 16396 24256
rect 16071 24225 16083 24228
rect 16025 24219 16083 24225
rect 15023 24160 15148 24188
rect 15197 24191 15255 24197
rect 15023 24157 15035 24160
rect 14977 24151 15035 24157
rect 15197 24157 15209 24191
rect 15243 24157 15255 24191
rect 15197 24151 15255 24157
rect 15294 24191 15352 24197
rect 15294 24157 15306 24191
rect 15340 24157 15352 24191
rect 15294 24151 15352 24157
rect 15102 24120 15108 24132
rect 12216 24092 12388 24120
rect 15063 24092 15108 24120
rect 12216 24080 12222 24092
rect 15102 24080 15108 24092
rect 15160 24080 15166 24132
rect 4154 24052 4160 24064
rect 3988 24024 4160 24052
rect 4154 24012 4160 24024
rect 4212 24052 4218 24064
rect 5258 24052 5264 24064
rect 4212 24024 5264 24052
rect 4212 24012 4218 24024
rect 5258 24012 5264 24024
rect 5316 24012 5322 24064
rect 5994 24012 6000 24064
rect 6052 24052 6058 24064
rect 8570 24052 8576 24064
rect 6052 24024 8576 24052
rect 6052 24012 6058 24024
rect 8570 24012 8576 24024
rect 8628 24012 8634 24064
rect 11149 24055 11207 24061
rect 11149 24021 11161 24055
rect 11195 24052 11207 24055
rect 11330 24052 11336 24064
rect 11195 24024 11336 24052
rect 11195 24021 11207 24024
rect 11149 24015 11207 24021
rect 11330 24012 11336 24024
rect 11388 24052 11394 24064
rect 11606 24052 11612 24064
rect 11388 24024 11612 24052
rect 11388 24012 11394 24024
rect 11606 24012 11612 24024
rect 11664 24012 11670 24064
rect 12805 24055 12863 24061
rect 12805 24021 12817 24055
rect 12851 24052 12863 24055
rect 13170 24052 13176 24064
rect 12851 24024 13176 24052
rect 12851 24021 12863 24024
rect 12805 24015 12863 24021
rect 13170 24012 13176 24024
rect 13228 24012 13234 24064
rect 15010 24012 15016 24064
rect 15068 24052 15074 24064
rect 15304 24052 15332 24151
rect 15562 24148 15568 24200
rect 15620 24188 15626 24200
rect 16040 24188 16068 24219
rect 16390 24216 16396 24228
rect 16448 24216 16454 24268
rect 17313 24259 17371 24265
rect 17313 24225 17325 24259
rect 17359 24256 17371 24259
rect 18322 24256 18328 24268
rect 17359 24228 18328 24256
rect 17359 24225 17371 24228
rect 17313 24219 17371 24225
rect 18322 24216 18328 24228
rect 18380 24216 18386 24268
rect 15620 24160 16068 24188
rect 15620 24148 15626 24160
rect 17402 24148 17408 24200
rect 17460 24188 17466 24200
rect 18432 24197 18460 24296
rect 18598 24284 18604 24336
rect 18656 24284 18662 24336
rect 18616 24197 18644 24284
rect 21910 24216 21916 24268
rect 21968 24256 21974 24268
rect 22281 24259 22339 24265
rect 22281 24256 22293 24259
rect 21968 24228 22293 24256
rect 21968 24216 21974 24228
rect 22281 24225 22293 24228
rect 22327 24225 22339 24259
rect 22462 24256 22468 24268
rect 22423 24228 22468 24256
rect 22281 24219 22339 24225
rect 22462 24216 22468 24228
rect 22520 24216 22526 24268
rect 17497 24191 17555 24197
rect 17497 24188 17509 24191
rect 17460 24160 17509 24188
rect 17460 24148 17466 24160
rect 17497 24157 17509 24160
rect 17543 24157 17555 24191
rect 17497 24151 17555 24157
rect 18417 24191 18475 24197
rect 18417 24157 18429 24191
rect 18463 24157 18475 24191
rect 18417 24151 18475 24157
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24157 18659 24191
rect 18601 24151 18659 24157
rect 19889 24191 19947 24197
rect 19889 24157 19901 24191
rect 19935 24157 19947 24191
rect 20346 24188 20352 24200
rect 20307 24160 20352 24188
rect 19889 24151 19947 24157
rect 16209 24123 16267 24129
rect 16209 24089 16221 24123
rect 16255 24120 16267 24123
rect 16390 24120 16396 24132
rect 16255 24092 16396 24120
rect 16255 24089 16267 24092
rect 16209 24083 16267 24089
rect 16390 24080 16396 24092
rect 16448 24080 16454 24132
rect 16942 24080 16948 24132
rect 17000 24120 17006 24132
rect 19904 24120 19932 24151
rect 20346 24148 20352 24160
rect 20404 24148 20410 24200
rect 21634 24120 21640 24132
rect 17000 24092 18644 24120
rect 19904 24092 21640 24120
rect 17000 24080 17006 24092
rect 15068 24024 15332 24052
rect 15473 24055 15531 24061
rect 15068 24012 15074 24024
rect 15473 24021 15485 24055
rect 15519 24052 15531 24055
rect 16114 24052 16120 24064
rect 15519 24024 16120 24052
rect 15519 24021 15531 24024
rect 15473 24015 15531 24021
rect 16114 24012 16120 24024
rect 16172 24012 16178 24064
rect 16301 24055 16359 24061
rect 16301 24021 16313 24055
rect 16347 24052 16359 24055
rect 16482 24052 16488 24064
rect 16347 24024 16488 24052
rect 16347 24021 16359 24024
rect 16301 24015 16359 24021
rect 16482 24012 16488 24024
rect 16540 24012 16546 24064
rect 16574 24012 16580 24064
rect 16632 24052 16638 24064
rect 16669 24055 16727 24061
rect 16669 24052 16681 24055
rect 16632 24024 16681 24052
rect 16632 24012 16638 24024
rect 16669 24021 16681 24024
rect 16715 24021 16727 24055
rect 16669 24015 16727 24021
rect 17126 24012 17132 24064
rect 17184 24052 17190 24064
rect 17405 24055 17463 24061
rect 17405 24052 17417 24055
rect 17184 24024 17417 24052
rect 17184 24012 17190 24024
rect 17405 24021 17417 24024
rect 17451 24021 17463 24055
rect 17405 24015 17463 24021
rect 18322 24012 18328 24064
rect 18380 24052 18386 24064
rect 18509 24055 18567 24061
rect 18509 24052 18521 24055
rect 18380 24024 18521 24052
rect 18380 24012 18386 24024
rect 18509 24021 18521 24024
rect 18555 24021 18567 24055
rect 18616 24052 18644 24092
rect 21634 24080 21640 24092
rect 21692 24080 21698 24132
rect 22189 24123 22247 24129
rect 22189 24089 22201 24123
rect 22235 24120 22247 24123
rect 22278 24120 22284 24132
rect 22235 24092 22284 24120
rect 22235 24089 22247 24092
rect 22189 24083 22247 24089
rect 22278 24080 22284 24092
rect 22336 24080 22342 24132
rect 20441 24055 20499 24061
rect 20441 24052 20453 24055
rect 18616 24024 20453 24052
rect 18509 24015 18567 24021
rect 20441 24021 20453 24024
rect 20487 24021 20499 24055
rect 20441 24015 20499 24021
rect 21450 24012 21456 24064
rect 21508 24052 21514 24064
rect 21821 24055 21879 24061
rect 21821 24052 21833 24055
rect 21508 24024 21833 24052
rect 21508 24012 21514 24024
rect 21821 24021 21833 24024
rect 21867 24021 21879 24055
rect 21821 24015 21879 24021
rect 1104 23962 30820 23984
rect 1104 23910 10880 23962
rect 10932 23910 10944 23962
rect 10996 23910 11008 23962
rect 11060 23910 11072 23962
rect 11124 23910 11136 23962
rect 11188 23910 20811 23962
rect 20863 23910 20875 23962
rect 20927 23910 20939 23962
rect 20991 23910 21003 23962
rect 21055 23910 21067 23962
rect 21119 23910 30820 23962
rect 1104 23888 30820 23910
rect 4154 23848 4160 23860
rect 4115 23820 4160 23848
rect 4154 23808 4160 23820
rect 4212 23808 4218 23860
rect 7282 23808 7288 23860
rect 7340 23808 7346 23860
rect 7374 23808 7380 23860
rect 7432 23848 7438 23860
rect 7653 23851 7711 23857
rect 7653 23848 7665 23851
rect 7432 23820 7665 23848
rect 7432 23808 7438 23820
rect 7653 23817 7665 23820
rect 7699 23817 7711 23851
rect 9674 23848 9680 23860
rect 7653 23811 7711 23817
rect 7852 23820 9680 23848
rect 2866 23780 2872 23792
rect 2779 23752 2872 23780
rect 2792 23721 2820 23752
rect 2866 23740 2872 23752
rect 2924 23780 2930 23792
rect 4062 23780 4068 23792
rect 2924 23752 4068 23780
rect 2924 23740 2930 23752
rect 4062 23740 4068 23752
rect 4120 23740 4126 23792
rect 4982 23780 4988 23792
rect 4816 23752 4988 23780
rect 2777 23715 2835 23721
rect 2777 23681 2789 23715
rect 2823 23681 2835 23715
rect 2777 23675 2835 23681
rect 3044 23715 3102 23721
rect 3044 23681 3056 23715
rect 3090 23712 3102 23715
rect 3786 23712 3792 23724
rect 3090 23684 3792 23712
rect 3090 23681 3102 23684
rect 3044 23675 3102 23681
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 4816 23721 4844 23752
rect 4982 23740 4988 23752
rect 5040 23740 5046 23792
rect 5902 23740 5908 23792
rect 5960 23780 5966 23792
rect 7300 23780 7328 23808
rect 7558 23780 7564 23792
rect 5960 23752 6684 23780
rect 7300 23752 7564 23780
rect 5960 23740 5966 23752
rect 6656 23724 6684 23752
rect 7558 23740 7564 23752
rect 7616 23740 7622 23792
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23681 4859 23715
rect 4801 23675 4859 23681
rect 5169 23715 5227 23721
rect 5169 23681 5181 23715
rect 5215 23712 5227 23715
rect 5353 23715 5411 23721
rect 5215 23684 5304 23712
rect 5215 23681 5227 23684
rect 5169 23675 5227 23681
rect 1394 23644 1400 23656
rect 1355 23616 1400 23644
rect 1394 23604 1400 23616
rect 1452 23604 1458 23656
rect 1673 23647 1731 23653
rect 1673 23613 1685 23647
rect 1719 23644 1731 23647
rect 2314 23644 2320 23656
rect 1719 23616 2320 23644
rect 1719 23613 1731 23616
rect 1673 23607 1731 23613
rect 2314 23604 2320 23616
rect 2372 23604 2378 23656
rect 4246 23604 4252 23656
rect 4304 23644 4310 23656
rect 4890 23644 4896 23656
rect 4304 23616 4896 23644
rect 4304 23604 4310 23616
rect 4890 23604 4896 23616
rect 4948 23644 4954 23656
rect 4985 23647 5043 23653
rect 4985 23644 4997 23647
rect 4948 23616 4997 23644
rect 4948 23604 4954 23616
rect 4985 23613 4997 23616
rect 5031 23613 5043 23647
rect 4985 23607 5043 23613
rect 5074 23604 5080 23656
rect 5132 23644 5138 23656
rect 5276 23644 5304 23684
rect 5353 23681 5365 23715
rect 5399 23712 5411 23715
rect 5534 23712 5540 23724
rect 5399 23684 5540 23712
rect 5399 23681 5411 23684
rect 5353 23675 5411 23681
rect 5534 23672 5540 23684
rect 5592 23712 5598 23724
rect 6365 23715 6423 23721
rect 6365 23712 6377 23715
rect 5592 23684 6377 23712
rect 5592 23672 5598 23684
rect 6365 23681 6377 23684
rect 6411 23712 6423 23715
rect 6454 23712 6460 23724
rect 6411 23684 6460 23712
rect 6411 23681 6423 23684
rect 6365 23675 6423 23681
rect 6454 23672 6460 23684
rect 6512 23672 6518 23724
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23681 6607 23715
rect 6549 23675 6607 23681
rect 5718 23644 5724 23656
rect 5132 23616 5177 23644
rect 5276 23616 5724 23644
rect 5132 23604 5138 23616
rect 5718 23604 5724 23616
rect 5776 23604 5782 23656
rect 4338 23536 4344 23588
rect 4396 23576 4402 23588
rect 6564 23576 6592 23675
rect 6638 23672 6644 23724
rect 6696 23712 6702 23724
rect 6696 23684 6789 23712
rect 6696 23672 6702 23684
rect 6914 23672 6920 23724
rect 6972 23712 6978 23724
rect 7282 23712 7288 23724
rect 6972 23684 7288 23712
rect 6972 23672 6978 23684
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 7852 23721 7880 23820
rect 9674 23808 9680 23820
rect 9732 23808 9738 23860
rect 9858 23848 9864 23860
rect 9819 23820 9864 23848
rect 9858 23808 9864 23820
rect 9916 23808 9922 23860
rect 10226 23808 10232 23860
rect 10284 23848 10290 23860
rect 11606 23848 11612 23860
rect 10284 23820 11612 23848
rect 10284 23808 10290 23820
rect 11606 23808 11612 23820
rect 11664 23848 11670 23860
rect 12250 23848 12256 23860
rect 11664 23820 12256 23848
rect 11664 23808 11670 23820
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 14274 23848 14280 23860
rect 14235 23820 14280 23848
rect 14274 23808 14280 23820
rect 14332 23848 14338 23860
rect 14734 23848 14740 23860
rect 14332 23820 14740 23848
rect 14332 23808 14338 23820
rect 14734 23808 14740 23820
rect 14792 23808 14798 23860
rect 18322 23808 18328 23860
rect 18380 23848 18386 23860
rect 18509 23851 18567 23857
rect 18509 23848 18521 23851
rect 18380 23820 18521 23848
rect 18380 23808 18386 23820
rect 18509 23817 18521 23820
rect 18555 23817 18567 23851
rect 20070 23848 20076 23860
rect 20031 23820 20076 23848
rect 18509 23811 18567 23817
rect 20070 23808 20076 23820
rect 20128 23808 20134 23860
rect 22278 23848 22284 23860
rect 21100 23820 22284 23848
rect 8570 23740 8576 23792
rect 8628 23780 8634 23792
rect 11330 23780 11336 23792
rect 8628 23752 9352 23780
rect 8628 23740 8634 23752
rect 7837 23715 7895 23721
rect 7837 23681 7849 23715
rect 7883 23681 7895 23715
rect 7837 23675 7895 23681
rect 7929 23715 7987 23721
rect 7929 23681 7941 23715
rect 7975 23712 7987 23715
rect 8018 23712 8024 23724
rect 7975 23684 8024 23712
rect 7975 23681 7987 23684
rect 7929 23675 7987 23681
rect 8018 23672 8024 23684
rect 8076 23672 8082 23724
rect 8202 23712 8208 23724
rect 8163 23684 8208 23712
rect 8202 23672 8208 23684
rect 8260 23672 8266 23724
rect 9125 23715 9183 23721
rect 9125 23681 9137 23715
rect 9171 23712 9183 23715
rect 9214 23712 9220 23724
rect 9171 23684 9220 23712
rect 9171 23681 9183 23684
rect 9125 23675 9183 23681
rect 9214 23672 9220 23684
rect 9272 23672 9278 23724
rect 9324 23721 9352 23752
rect 9692 23752 11336 23780
rect 9309 23715 9367 23721
rect 9309 23681 9321 23715
rect 9355 23681 9367 23715
rect 9490 23712 9496 23724
rect 9451 23684 9496 23712
rect 9309 23675 9367 23681
rect 9490 23672 9496 23684
rect 9548 23672 9554 23724
rect 9692 23721 9720 23752
rect 11330 23740 11336 23752
rect 11388 23740 11394 23792
rect 11422 23740 11428 23792
rect 11480 23780 11486 23792
rect 11701 23783 11759 23789
rect 11701 23780 11713 23783
rect 11480 23752 11713 23780
rect 11480 23740 11486 23752
rect 11701 23749 11713 23752
rect 11747 23749 11759 23783
rect 11701 23743 11759 23749
rect 11885 23783 11943 23789
rect 11885 23749 11897 23783
rect 11931 23780 11943 23783
rect 12986 23780 12992 23792
rect 11931 23752 12992 23780
rect 11931 23749 11943 23752
rect 11885 23743 11943 23749
rect 9677 23715 9735 23721
rect 9677 23681 9689 23715
rect 9723 23681 9735 23715
rect 10502 23712 10508 23724
rect 10463 23684 10508 23712
rect 9677 23675 9735 23681
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 11716 23712 11744 23743
rect 12986 23740 12992 23752
rect 13044 23740 13050 23792
rect 13170 23789 13176 23792
rect 13164 23780 13176 23789
rect 13131 23752 13176 23780
rect 13164 23743 13176 23752
rect 13170 23740 13176 23743
rect 13228 23740 13234 23792
rect 15102 23740 15108 23792
rect 15160 23780 15166 23792
rect 16298 23780 16304 23792
rect 15160 23752 16304 23780
rect 15160 23740 15166 23752
rect 16298 23740 16304 23752
rect 16356 23740 16362 23792
rect 19334 23740 19340 23792
rect 19392 23780 19398 23792
rect 20346 23780 20352 23792
rect 19392 23752 20352 23780
rect 19392 23740 19398 23752
rect 20346 23740 20352 23752
rect 20404 23740 20410 23792
rect 12342 23712 12348 23724
rect 11716 23684 12348 23712
rect 12342 23672 12348 23684
rect 12400 23712 12406 23724
rect 12897 23715 12955 23721
rect 12897 23712 12909 23715
rect 12400 23684 12909 23712
rect 12400 23672 12406 23684
rect 12897 23681 12909 23684
rect 12943 23681 12955 23715
rect 12897 23675 12955 23681
rect 14274 23672 14280 23724
rect 14332 23712 14338 23724
rect 14737 23715 14795 23721
rect 14737 23712 14749 23715
rect 14332 23684 14749 23712
rect 14332 23672 14338 23684
rect 14737 23681 14749 23684
rect 14783 23681 14795 23715
rect 14737 23675 14795 23681
rect 15749 23715 15807 23721
rect 15749 23681 15761 23715
rect 15795 23712 15807 23715
rect 16482 23712 16488 23724
rect 15795 23684 16488 23712
rect 15795 23681 15807 23684
rect 15749 23675 15807 23681
rect 16482 23672 16488 23684
rect 16540 23672 16546 23724
rect 16666 23712 16672 23724
rect 16627 23684 16672 23712
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 17126 23712 17132 23724
rect 17087 23684 17132 23712
rect 17126 23672 17132 23684
rect 17184 23672 17190 23724
rect 17497 23715 17555 23721
rect 17497 23681 17509 23715
rect 17543 23712 17555 23715
rect 17770 23712 17776 23724
rect 17543 23684 17776 23712
rect 17543 23681 17555 23684
rect 17497 23675 17555 23681
rect 17770 23672 17776 23684
rect 17828 23672 17834 23724
rect 17862 23672 17868 23724
rect 17920 23712 17926 23724
rect 20257 23715 20315 23721
rect 20257 23712 20269 23715
rect 17920 23684 20269 23712
rect 17920 23672 17926 23684
rect 20257 23681 20269 23684
rect 20303 23681 20315 23715
rect 20438 23712 20444 23724
rect 20399 23684 20444 23712
rect 20257 23675 20315 23681
rect 6733 23647 6791 23653
rect 6733 23613 6745 23647
rect 6779 23613 6791 23647
rect 9398 23644 9404 23656
rect 9311 23616 9404 23644
rect 6733 23607 6791 23613
rect 4396 23548 6592 23576
rect 4396 23536 4402 23548
rect 4614 23508 4620 23520
rect 4575 23480 4620 23508
rect 4614 23468 4620 23480
rect 4672 23468 4678 23520
rect 6564 23508 6592 23548
rect 6638 23536 6644 23588
rect 6696 23576 6702 23588
rect 6748 23576 6776 23607
rect 9398 23604 9404 23616
rect 9456 23644 9462 23656
rect 9582 23644 9588 23656
rect 9456 23616 9588 23644
rect 9456 23604 9462 23616
rect 9582 23604 9588 23616
rect 9640 23604 9646 23656
rect 9766 23604 9772 23656
rect 9824 23644 9830 23656
rect 10042 23644 10048 23656
rect 9824 23616 10048 23644
rect 9824 23604 9830 23616
rect 10042 23604 10048 23616
rect 10100 23644 10106 23656
rect 10413 23647 10471 23653
rect 10413 23644 10425 23647
rect 10100 23616 10425 23644
rect 10100 23604 10106 23616
rect 10413 23613 10425 23616
rect 10459 23613 10471 23647
rect 15470 23644 15476 23656
rect 15431 23616 15476 23644
rect 10413 23607 10471 23613
rect 15470 23604 15476 23616
rect 15528 23604 15534 23656
rect 15562 23604 15568 23656
rect 15620 23644 15626 23656
rect 15657 23647 15715 23653
rect 15657 23644 15669 23647
rect 15620 23616 15669 23644
rect 15620 23604 15626 23616
rect 15657 23613 15669 23616
rect 15703 23613 15715 23647
rect 15657 23607 15715 23613
rect 16114 23604 16120 23656
rect 16172 23644 16178 23656
rect 17218 23644 17224 23656
rect 16172 23616 17080 23644
rect 17179 23616 17224 23644
rect 16172 23604 16178 23616
rect 8662 23576 8668 23588
rect 6696 23548 6776 23576
rect 6840 23548 8668 23576
rect 6696 23536 6702 23548
rect 6840 23508 6868 23548
rect 8662 23536 8668 23548
rect 8720 23536 8726 23588
rect 14829 23579 14887 23585
rect 14829 23545 14841 23579
rect 14875 23576 14887 23579
rect 16390 23576 16396 23588
rect 14875 23548 16396 23576
rect 14875 23545 14887 23548
rect 14829 23539 14887 23545
rect 16390 23536 16396 23548
rect 16448 23536 16454 23588
rect 17052 23576 17080 23616
rect 17218 23604 17224 23616
rect 17276 23604 17282 23656
rect 17402 23644 17408 23656
rect 17363 23616 17408 23644
rect 17402 23604 17408 23616
rect 17460 23604 17466 23656
rect 18598 23644 18604 23656
rect 18559 23616 18604 23644
rect 18598 23604 18604 23616
rect 18656 23604 18662 23656
rect 18785 23647 18843 23653
rect 18785 23613 18797 23647
rect 18831 23644 18843 23647
rect 19150 23644 19156 23656
rect 18831 23616 19156 23644
rect 18831 23613 18843 23616
rect 18785 23607 18843 23613
rect 19150 23604 19156 23616
rect 19208 23604 19214 23656
rect 20272 23644 20300 23675
rect 20438 23672 20444 23684
rect 20496 23672 20502 23724
rect 21100 23721 21128 23820
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 21910 23780 21916 23792
rect 21871 23752 21916 23780
rect 21910 23740 21916 23752
rect 21968 23740 21974 23792
rect 21085 23715 21143 23721
rect 21085 23681 21097 23715
rect 21131 23681 21143 23715
rect 21085 23675 21143 23681
rect 22097 23715 22155 23721
rect 22097 23681 22109 23715
rect 22143 23712 22155 23715
rect 22830 23712 22836 23724
rect 22143 23684 22836 23712
rect 22143 23681 22155 23684
rect 22097 23675 22155 23681
rect 22830 23672 22836 23684
rect 22888 23672 22894 23724
rect 20530 23644 20536 23656
rect 20272 23616 20536 23644
rect 20530 23604 20536 23616
rect 20588 23604 20594 23656
rect 20714 23604 20720 23656
rect 20772 23644 20778 23656
rect 21177 23647 21235 23653
rect 21177 23644 21189 23647
rect 20772 23616 21189 23644
rect 20772 23604 20778 23616
rect 21177 23613 21189 23616
rect 21223 23613 21235 23647
rect 22646 23644 22652 23656
rect 22607 23616 22652 23644
rect 21177 23607 21235 23613
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 22922 23644 22928 23656
rect 22883 23616 22928 23644
rect 22922 23604 22928 23616
rect 22980 23604 22986 23656
rect 20622 23576 20628 23588
rect 17052 23548 20628 23576
rect 20622 23536 20628 23548
rect 20680 23536 20686 23588
rect 6564 23480 6868 23508
rect 6914 23468 6920 23520
rect 6972 23508 6978 23520
rect 7101 23511 7159 23517
rect 7101 23508 7113 23511
rect 6972 23480 7113 23508
rect 6972 23468 6978 23480
rect 7101 23477 7113 23480
rect 7147 23477 7159 23511
rect 7101 23471 7159 23477
rect 7926 23468 7932 23520
rect 7984 23508 7990 23520
rect 8113 23511 8171 23517
rect 8113 23508 8125 23511
rect 7984 23480 8125 23508
rect 7984 23468 7990 23480
rect 8113 23477 8125 23480
rect 8159 23477 8171 23511
rect 8113 23471 8171 23477
rect 8938 23468 8944 23520
rect 8996 23508 9002 23520
rect 9766 23508 9772 23520
rect 8996 23480 9772 23508
rect 8996 23468 9002 23480
rect 9766 23468 9772 23480
rect 9824 23468 9830 23520
rect 16117 23511 16175 23517
rect 16117 23477 16129 23511
rect 16163 23508 16175 23511
rect 16206 23508 16212 23520
rect 16163 23480 16212 23508
rect 16163 23477 16175 23480
rect 16117 23471 16175 23477
rect 16206 23468 16212 23480
rect 16264 23468 16270 23520
rect 16298 23468 16304 23520
rect 16356 23508 16362 23520
rect 16761 23511 16819 23517
rect 16761 23508 16773 23511
rect 16356 23480 16773 23508
rect 16356 23468 16362 23480
rect 16761 23477 16773 23480
rect 16807 23477 16819 23511
rect 18138 23508 18144 23520
rect 18099 23480 18144 23508
rect 16761 23471 16819 23477
rect 18138 23468 18144 23480
rect 18196 23468 18202 23520
rect 19518 23468 19524 23520
rect 19576 23508 19582 23520
rect 20257 23511 20315 23517
rect 20257 23508 20269 23511
rect 19576 23480 20269 23508
rect 19576 23468 19582 23480
rect 20257 23477 20269 23480
rect 20303 23477 20315 23511
rect 20257 23471 20315 23477
rect 1104 23418 30820 23440
rect 1104 23366 5915 23418
rect 5967 23366 5979 23418
rect 6031 23366 6043 23418
rect 6095 23366 6107 23418
rect 6159 23366 6171 23418
rect 6223 23366 15846 23418
rect 15898 23366 15910 23418
rect 15962 23366 15974 23418
rect 16026 23366 16038 23418
rect 16090 23366 16102 23418
rect 16154 23366 25776 23418
rect 25828 23366 25840 23418
rect 25892 23366 25904 23418
rect 25956 23366 25968 23418
rect 26020 23366 26032 23418
rect 26084 23366 30820 23418
rect 1104 23344 30820 23366
rect 4982 23264 4988 23316
rect 5040 23304 5046 23316
rect 5442 23304 5448 23316
rect 5040 23276 5448 23304
rect 5040 23264 5046 23276
rect 5442 23264 5448 23276
rect 5500 23264 5506 23316
rect 5718 23264 5724 23316
rect 5776 23304 5782 23316
rect 7282 23304 7288 23316
rect 5776 23276 7144 23304
rect 7243 23276 7288 23304
rect 5776 23264 5782 23276
rect 7116 23236 7144 23276
rect 7282 23264 7288 23276
rect 7340 23304 7346 23316
rect 7650 23304 7656 23316
rect 7340 23276 7656 23304
rect 7340 23264 7346 23276
rect 7650 23264 7656 23276
rect 7708 23264 7714 23316
rect 11514 23304 11520 23316
rect 10336 23276 11520 23304
rect 7116 23208 9444 23236
rect 4062 23168 4068 23180
rect 4023 23140 4068 23168
rect 4062 23128 4068 23140
rect 4120 23128 4126 23180
rect 5810 23128 5816 23180
rect 5868 23168 5874 23180
rect 5905 23171 5963 23177
rect 5905 23168 5917 23171
rect 5868 23140 5917 23168
rect 5868 23128 5874 23140
rect 5905 23137 5917 23140
rect 5951 23137 5963 23171
rect 5905 23131 5963 23137
rect 7282 23128 7288 23180
rect 7340 23168 7346 23180
rect 7834 23168 7840 23180
rect 7340 23140 7840 23168
rect 7340 23128 7346 23140
rect 7834 23128 7840 23140
rect 7892 23128 7898 23180
rect 1397 23103 1455 23109
rect 1397 23069 1409 23103
rect 1443 23069 1455 23103
rect 2038 23100 2044 23112
rect 1999 23072 2044 23100
rect 1397 23063 1455 23069
rect 1412 23032 1440 23063
rect 2038 23060 2044 23072
rect 2096 23060 2102 23112
rect 4332 23103 4390 23109
rect 4332 23069 4344 23103
rect 4378 23100 4390 23103
rect 4614 23100 4620 23112
rect 4378 23072 4620 23100
rect 4378 23069 4390 23072
rect 4332 23063 4390 23069
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 6172 23103 6230 23109
rect 6172 23069 6184 23103
rect 6218 23100 6230 23103
rect 6914 23100 6920 23112
rect 6218 23072 6920 23100
rect 6218 23069 6230 23072
rect 6172 23063 6230 23069
rect 6914 23060 6920 23072
rect 6972 23060 6978 23112
rect 7745 23103 7803 23109
rect 7745 23069 7757 23103
rect 7791 23100 7803 23103
rect 9214 23100 9220 23112
rect 7791 23072 7972 23100
rect 9175 23072 9220 23100
rect 7791 23069 7803 23072
rect 7745 23063 7803 23069
rect 2774 23032 2780 23044
rect 1412 23004 2780 23032
rect 2774 22992 2780 23004
rect 2832 22992 2838 23044
rect 1581 22967 1639 22973
rect 1581 22933 1593 22967
rect 1627 22964 1639 22967
rect 1670 22964 1676 22976
rect 1627 22936 1676 22964
rect 1627 22933 1639 22936
rect 1581 22927 1639 22933
rect 1670 22924 1676 22936
rect 1728 22924 1734 22976
rect 2225 22967 2283 22973
rect 2225 22933 2237 22967
rect 2271 22964 2283 22967
rect 4246 22964 4252 22976
rect 2271 22936 4252 22964
rect 2271 22933 2283 22936
rect 2225 22927 2283 22933
rect 4246 22924 4252 22936
rect 4304 22924 4310 22976
rect 7834 22964 7840 22976
rect 7795 22936 7840 22964
rect 7834 22924 7840 22936
rect 7892 22924 7898 22976
rect 7944 22964 7972 23072
rect 9214 23060 9220 23072
rect 9272 23060 9278 23112
rect 9416 23109 9444 23208
rect 9490 23196 9496 23248
rect 9548 23236 9554 23248
rect 9548 23208 9628 23236
rect 9548 23196 9554 23208
rect 9600 23177 9628 23208
rect 9585 23171 9643 23177
rect 9585 23137 9597 23171
rect 9631 23137 9643 23171
rect 9585 23131 9643 23137
rect 9401 23103 9459 23109
rect 9401 23069 9413 23103
rect 9447 23069 9459 23103
rect 9401 23063 9459 23069
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23069 9551 23103
rect 9493 23063 9551 23069
rect 9769 23103 9827 23109
rect 9769 23069 9781 23103
rect 9815 23100 9827 23103
rect 10336 23100 10364 23276
rect 11514 23264 11520 23276
rect 11572 23264 11578 23316
rect 13078 23304 13084 23316
rect 12406 23276 13084 23304
rect 12406 23236 12434 23276
rect 13078 23264 13084 23276
rect 13136 23264 13142 23316
rect 14921 23307 14979 23313
rect 14921 23273 14933 23307
rect 14967 23304 14979 23307
rect 15010 23304 15016 23316
rect 14967 23276 15016 23304
rect 14967 23273 14979 23276
rect 14921 23267 14979 23273
rect 15010 23264 15016 23276
rect 15068 23264 15074 23316
rect 15473 23307 15531 23313
rect 15473 23273 15485 23307
rect 15519 23304 15531 23307
rect 15562 23304 15568 23316
rect 15519 23276 15568 23304
rect 15519 23273 15531 23276
rect 15473 23267 15531 23273
rect 15562 23264 15568 23276
rect 15620 23264 15626 23316
rect 16666 23264 16672 23316
rect 16724 23304 16730 23316
rect 16761 23307 16819 23313
rect 16761 23304 16773 23307
rect 16724 23276 16773 23304
rect 16724 23264 16730 23276
rect 16761 23273 16773 23276
rect 16807 23273 16819 23307
rect 19518 23304 19524 23316
rect 19479 23276 19524 23304
rect 16761 23267 16819 23273
rect 19518 23264 19524 23276
rect 19576 23264 19582 23316
rect 22557 23307 22615 23313
rect 22557 23273 22569 23307
rect 22603 23304 22615 23307
rect 22646 23304 22652 23316
rect 22603 23276 22652 23304
rect 22603 23273 22615 23276
rect 22557 23267 22615 23273
rect 22646 23264 22652 23276
rect 22704 23264 22710 23316
rect 22186 23236 22192 23248
rect 11256 23208 12434 23236
rect 21744 23208 22192 23236
rect 11256 23177 11284 23208
rect 11241 23171 11299 23177
rect 11241 23137 11253 23171
rect 11287 23137 11299 23171
rect 11698 23168 11704 23180
rect 11241 23131 11299 23137
rect 11348 23140 11704 23168
rect 9815 23072 10364 23100
rect 9815 23069 9827 23072
rect 9769 23063 9827 23069
rect 9508 23032 9536 23063
rect 10410 23060 10416 23112
rect 10468 23100 10474 23112
rect 10873 23103 10931 23109
rect 10873 23100 10885 23103
rect 10468 23072 10885 23100
rect 10468 23060 10474 23072
rect 10873 23069 10885 23072
rect 10919 23069 10931 23103
rect 10873 23063 10931 23069
rect 11057 23103 11115 23109
rect 11057 23069 11069 23103
rect 11103 23069 11115 23103
rect 11057 23063 11115 23069
rect 11149 23103 11207 23109
rect 11149 23069 11161 23103
rect 11195 23100 11207 23103
rect 11348 23100 11376 23140
rect 11698 23128 11704 23140
rect 11756 23128 11762 23180
rect 12158 23128 12164 23180
rect 12216 23168 12222 23180
rect 12345 23171 12403 23177
rect 12345 23168 12357 23171
rect 12216 23140 12357 23168
rect 12216 23128 12222 23140
rect 12345 23137 12357 23140
rect 12391 23137 12403 23171
rect 12345 23131 12403 23137
rect 12437 23171 12495 23177
rect 12437 23137 12449 23171
rect 12483 23168 12495 23171
rect 12526 23168 12532 23180
rect 12483 23140 12532 23168
rect 12483 23137 12495 23140
rect 12437 23131 12495 23137
rect 12526 23128 12532 23140
rect 12584 23128 12590 23180
rect 14274 23168 14280 23180
rect 12636 23140 14280 23168
rect 11195 23072 11376 23100
rect 11425 23103 11483 23109
rect 11195 23069 11207 23072
rect 11149 23063 11207 23069
rect 11425 23069 11437 23103
rect 11471 23069 11483 23103
rect 12066 23100 12072 23112
rect 12027 23072 12072 23100
rect 11425 23063 11483 23069
rect 9582 23032 9588 23044
rect 9508 23004 9588 23032
rect 9582 22992 9588 23004
rect 9640 22992 9646 23044
rect 11072 23032 11100 23063
rect 9692 23004 11100 23032
rect 11440 23032 11468 23063
rect 12066 23060 12072 23072
rect 12124 23060 12130 23112
rect 12250 23100 12256 23112
rect 12211 23072 12256 23100
rect 12250 23060 12256 23072
rect 12308 23060 12314 23112
rect 12636 23109 12664 23140
rect 14274 23128 14280 23140
rect 14332 23128 14338 23180
rect 16393 23171 16451 23177
rect 16393 23137 16405 23171
rect 16439 23168 16451 23171
rect 16666 23168 16672 23180
rect 16439 23140 16672 23168
rect 16439 23137 16451 23140
rect 16393 23131 16451 23137
rect 16666 23128 16672 23140
rect 16724 23128 16730 23180
rect 17034 23128 17040 23180
rect 17092 23168 17098 23180
rect 20714 23168 20720 23180
rect 17092 23140 19472 23168
rect 17092 23128 17098 23140
rect 12621 23103 12679 23109
rect 12621 23069 12633 23103
rect 12667 23069 12679 23103
rect 12621 23063 12679 23069
rect 13722 23060 13728 23112
rect 13780 23100 13786 23112
rect 15381 23103 15439 23109
rect 15381 23100 15393 23103
rect 13780 23072 15393 23100
rect 13780 23060 13786 23072
rect 15381 23069 15393 23072
rect 15427 23069 15439 23103
rect 15381 23063 15439 23069
rect 15746 23060 15752 23112
rect 15804 23100 15810 23112
rect 16025 23103 16083 23109
rect 16025 23100 16037 23103
rect 15804 23072 16037 23100
rect 15804 23060 15810 23072
rect 16025 23069 16037 23072
rect 16071 23069 16083 23103
rect 16206 23100 16212 23112
rect 16167 23072 16212 23100
rect 16025 23063 16083 23069
rect 16206 23060 16212 23072
rect 16264 23060 16270 23112
rect 16301 23103 16359 23109
rect 16301 23069 16313 23103
rect 16347 23069 16359 23103
rect 16574 23100 16580 23112
rect 16535 23072 16580 23100
rect 16301 23063 16359 23069
rect 12986 23032 12992 23044
rect 11440 23004 12992 23032
rect 8018 22964 8024 22976
rect 7944 22936 8024 22964
rect 8018 22924 8024 22936
rect 8076 22964 8082 22976
rect 9692 22964 9720 23004
rect 12986 22992 12992 23004
rect 13044 22992 13050 23044
rect 14550 23032 14556 23044
rect 14511 23004 14556 23032
rect 14550 22992 14556 23004
rect 14608 22992 14614 23044
rect 14734 23032 14740 23044
rect 14695 23004 14740 23032
rect 14734 22992 14740 23004
rect 14792 22992 14798 23044
rect 16316 23032 16344 23063
rect 16574 23060 16580 23072
rect 16632 23060 16638 23112
rect 17052 23032 17080 23128
rect 18141 23103 18199 23109
rect 18141 23069 18153 23103
rect 18187 23100 18199 23103
rect 18966 23100 18972 23112
rect 18187 23072 18972 23100
rect 18187 23069 18199 23072
rect 18141 23063 18199 23069
rect 18966 23060 18972 23072
rect 19024 23100 19030 23112
rect 19150 23100 19156 23112
rect 19024 23072 19156 23100
rect 19024 23060 19030 23072
rect 19150 23060 19156 23072
rect 19208 23060 19214 23112
rect 19444 23109 19472 23140
rect 20364 23140 20720 23168
rect 19429 23103 19487 23109
rect 19429 23069 19441 23103
rect 19475 23100 19487 23103
rect 19702 23100 19708 23112
rect 19475 23072 19708 23100
rect 19475 23069 19487 23072
rect 19429 23063 19487 23069
rect 19702 23060 19708 23072
rect 19760 23060 19766 23112
rect 20070 23100 20076 23112
rect 20031 23072 20076 23100
rect 20070 23060 20076 23072
rect 20128 23060 20134 23112
rect 20254 23100 20260 23112
rect 20215 23072 20260 23100
rect 20254 23060 20260 23072
rect 20312 23060 20318 23112
rect 20364 23109 20392 23140
rect 20714 23128 20720 23140
rect 20772 23168 20778 23180
rect 21266 23168 21272 23180
rect 20772 23140 21272 23168
rect 20772 23128 20778 23140
rect 21266 23128 21272 23140
rect 21324 23128 21330 23180
rect 21450 23168 21456 23180
rect 21411 23140 21456 23168
rect 21450 23128 21456 23140
rect 21508 23128 21514 23180
rect 20349 23103 20407 23109
rect 20349 23069 20361 23103
rect 20395 23069 20407 23103
rect 20349 23063 20407 23069
rect 20441 23103 20499 23109
rect 20441 23069 20453 23103
rect 20487 23100 20499 23103
rect 21174 23100 21180 23112
rect 20487 23072 21180 23100
rect 20487 23069 20499 23072
rect 20441 23063 20499 23069
rect 21174 23060 21180 23072
rect 21232 23060 21238 23112
rect 21361 23103 21419 23109
rect 21361 23069 21373 23103
rect 21407 23100 21419 23103
rect 21744 23100 21772 23208
rect 22186 23196 22192 23208
rect 22244 23196 22250 23248
rect 21913 23171 21971 23177
rect 21913 23137 21925 23171
rect 21959 23168 21971 23171
rect 22370 23168 22376 23180
rect 21959 23140 22376 23168
rect 21959 23137 21971 23140
rect 21913 23131 21971 23137
rect 22370 23128 22376 23140
rect 22428 23168 22434 23180
rect 22922 23168 22928 23180
rect 22428 23140 22928 23168
rect 22428 23128 22434 23140
rect 22922 23128 22928 23140
rect 22980 23128 22986 23180
rect 21407 23072 21772 23100
rect 21407 23069 21419 23072
rect 21361 23063 21419 23069
rect 22186 23060 22192 23112
rect 22244 23100 22250 23112
rect 23569 23103 23627 23109
rect 23569 23100 23581 23103
rect 22244 23072 23581 23100
rect 22244 23060 22250 23072
rect 23569 23069 23581 23072
rect 23615 23069 23627 23103
rect 23569 23063 23627 23069
rect 29454 23060 29460 23112
rect 29512 23100 29518 23112
rect 29825 23103 29883 23109
rect 29825 23100 29837 23103
rect 29512 23072 29837 23100
rect 29512 23060 29518 23072
rect 29825 23069 29837 23072
rect 29871 23069 29883 23103
rect 29825 23063 29883 23069
rect 16316 23004 17080 23032
rect 20530 22992 20536 23044
rect 20588 23032 20594 23044
rect 20588 23004 21772 23032
rect 20588 22992 20594 23004
rect 8076 22936 9720 22964
rect 9953 22967 10011 22973
rect 8076 22924 8082 22936
rect 9953 22933 9965 22967
rect 9999 22964 10011 22967
rect 10042 22964 10048 22976
rect 9999 22936 10048 22964
rect 9999 22933 10011 22936
rect 9953 22927 10011 22933
rect 10042 22924 10048 22936
rect 10100 22924 10106 22976
rect 11609 22967 11667 22973
rect 11609 22933 11621 22967
rect 11655 22964 11667 22967
rect 11790 22964 11796 22976
rect 11655 22936 11796 22964
rect 11655 22933 11667 22936
rect 11609 22927 11667 22933
rect 11790 22924 11796 22936
rect 11848 22924 11854 22976
rect 12802 22964 12808 22976
rect 12763 22936 12808 22964
rect 12802 22924 12808 22936
rect 12860 22924 12866 22976
rect 18325 22967 18383 22973
rect 18325 22933 18337 22967
rect 18371 22964 18383 22967
rect 19150 22964 19156 22976
rect 18371 22936 19156 22964
rect 18371 22933 18383 22936
rect 18325 22927 18383 22933
rect 19150 22924 19156 22936
rect 19208 22924 19214 22976
rect 20714 22964 20720 22976
rect 20675 22936 20720 22964
rect 20714 22924 20720 22936
rect 20772 22924 20778 22976
rect 21744 22973 21772 23004
rect 22278 22992 22284 23044
rect 22336 23032 22342 23044
rect 22741 23035 22799 23041
rect 22741 23032 22753 23035
rect 22336 23004 22753 23032
rect 22336 22992 22342 23004
rect 22741 23001 22753 23004
rect 22787 23001 22799 23035
rect 22922 23032 22928 23044
rect 22883 23004 22928 23032
rect 22741 22995 22799 23001
rect 22922 22992 22928 23004
rect 22980 22992 22986 23044
rect 21729 22967 21787 22973
rect 21729 22933 21741 22967
rect 21775 22933 21787 22967
rect 23382 22964 23388 22976
rect 23343 22936 23388 22964
rect 21729 22927 21787 22933
rect 23382 22924 23388 22936
rect 23440 22924 23446 22976
rect 30006 22964 30012 22976
rect 29967 22936 30012 22964
rect 30006 22924 30012 22936
rect 30064 22924 30070 22976
rect 1104 22874 30820 22896
rect 1104 22822 10880 22874
rect 10932 22822 10944 22874
rect 10996 22822 11008 22874
rect 11060 22822 11072 22874
rect 11124 22822 11136 22874
rect 11188 22822 20811 22874
rect 20863 22822 20875 22874
rect 20927 22822 20939 22874
rect 20991 22822 21003 22874
rect 21055 22822 21067 22874
rect 21119 22822 30820 22874
rect 1104 22800 30820 22822
rect 7006 22720 7012 22772
rect 7064 22760 7070 22772
rect 7653 22763 7711 22769
rect 7653 22760 7665 22763
rect 7064 22732 7665 22760
rect 7064 22720 7070 22732
rect 7653 22729 7665 22732
rect 7699 22729 7711 22763
rect 7653 22723 7711 22729
rect 9122 22720 9128 22772
rect 9180 22760 9186 22772
rect 9398 22760 9404 22772
rect 9180 22732 9404 22760
rect 9180 22720 9186 22732
rect 9398 22720 9404 22732
rect 9456 22760 9462 22772
rect 12250 22760 12256 22772
rect 9456 22732 12256 22760
rect 9456 22720 9462 22732
rect 12250 22720 12256 22732
rect 12308 22720 12314 22772
rect 13722 22720 13728 22772
rect 13780 22760 13786 22772
rect 13817 22763 13875 22769
rect 13817 22760 13829 22763
rect 13780 22732 13829 22760
rect 13780 22720 13786 22732
rect 13817 22729 13829 22732
rect 13863 22729 13875 22763
rect 14274 22760 14280 22772
rect 14235 22732 14280 22760
rect 13817 22723 13875 22729
rect 14274 22720 14280 22732
rect 14332 22720 14338 22772
rect 15746 22720 15752 22772
rect 15804 22760 15810 22772
rect 16298 22760 16304 22772
rect 15804 22732 16304 22760
rect 15804 22720 15810 22732
rect 16298 22720 16304 22732
rect 16356 22720 16362 22772
rect 16390 22720 16396 22772
rect 16448 22760 16454 22772
rect 16945 22763 17003 22769
rect 16945 22760 16957 22763
rect 16448 22732 16957 22760
rect 16448 22720 16454 22732
rect 16945 22729 16957 22732
rect 16991 22729 17003 22763
rect 17402 22760 17408 22772
rect 17363 22732 17408 22760
rect 16945 22723 17003 22729
rect 17402 22720 17408 22732
rect 17460 22720 17466 22772
rect 18598 22720 18604 22772
rect 18656 22760 18662 22772
rect 18969 22763 19027 22769
rect 18969 22760 18981 22763
rect 18656 22732 18981 22760
rect 18656 22720 18662 22732
rect 18969 22729 18981 22732
rect 19015 22729 19027 22763
rect 19794 22760 19800 22772
rect 19707 22732 19800 22760
rect 18969 22723 19027 22729
rect 19794 22720 19800 22732
rect 19852 22760 19858 22772
rect 20070 22760 20076 22772
rect 19852 22732 20076 22760
rect 19852 22720 19858 22732
rect 20070 22720 20076 22732
rect 20128 22720 20134 22772
rect 21174 22720 21180 22772
rect 21232 22760 21238 22772
rect 22002 22760 22008 22772
rect 21232 22732 22008 22760
rect 21232 22720 21238 22732
rect 22002 22720 22008 22732
rect 22060 22720 22066 22772
rect 22186 22760 22192 22772
rect 22147 22732 22192 22760
rect 22186 22720 22192 22732
rect 22244 22720 22250 22772
rect 22922 22760 22928 22772
rect 22664 22732 22928 22760
rect 9214 22692 9220 22704
rect 6380 22664 9220 22692
rect 1397 22627 1455 22633
rect 1397 22593 1409 22627
rect 1443 22593 1455 22627
rect 1397 22587 1455 22593
rect 1412 22556 1440 22587
rect 1854 22584 1860 22636
rect 1912 22624 1918 22636
rect 2225 22627 2283 22633
rect 2225 22624 2237 22627
rect 1912 22596 2237 22624
rect 1912 22584 1918 22596
rect 2225 22593 2237 22596
rect 2271 22593 2283 22627
rect 2225 22587 2283 22593
rect 2685 22627 2743 22633
rect 2685 22593 2697 22627
rect 2731 22624 2743 22627
rect 2958 22624 2964 22636
rect 2731 22596 2964 22624
rect 2731 22593 2743 22596
rect 2685 22587 2743 22593
rect 2958 22584 2964 22596
rect 3016 22584 3022 22636
rect 4985 22627 5043 22633
rect 4985 22593 4997 22627
rect 5031 22624 5043 22627
rect 5074 22624 5080 22636
rect 5031 22596 5080 22624
rect 5031 22593 5043 22596
rect 4985 22587 5043 22593
rect 5074 22584 5080 22596
rect 5132 22584 5138 22636
rect 3142 22556 3148 22568
rect 1412 22528 3148 22556
rect 3142 22516 3148 22528
rect 3200 22516 3206 22568
rect 5258 22556 5264 22568
rect 5219 22528 5264 22556
rect 5258 22516 5264 22528
rect 5316 22516 5322 22568
rect 5718 22516 5724 22568
rect 5776 22556 5782 22568
rect 6380 22565 6408 22664
rect 9214 22652 9220 22664
rect 9272 22652 9278 22704
rect 12802 22652 12808 22704
rect 12860 22692 12866 22704
rect 15390 22695 15448 22701
rect 15390 22692 15402 22695
rect 12860 22664 15402 22692
rect 12860 22652 12866 22664
rect 15390 22661 15402 22664
rect 15436 22661 15448 22695
rect 15390 22655 15448 22661
rect 18141 22695 18199 22701
rect 18141 22661 18153 22695
rect 18187 22692 18199 22695
rect 19334 22692 19340 22704
rect 18187 22664 19340 22692
rect 18187 22661 18199 22664
rect 18141 22655 18199 22661
rect 19334 22652 19340 22664
rect 19392 22652 19398 22704
rect 19610 22652 19616 22704
rect 19668 22692 19674 22704
rect 20349 22695 20407 22701
rect 20349 22692 20361 22695
rect 19668 22664 20361 22692
rect 19668 22652 19674 22664
rect 20349 22661 20361 22664
rect 20395 22692 20407 22695
rect 20530 22692 20536 22704
rect 20395 22664 20536 22692
rect 20395 22661 20407 22664
rect 20349 22655 20407 22661
rect 20530 22652 20536 22664
rect 20588 22652 20594 22704
rect 21821 22695 21879 22701
rect 21821 22661 21833 22695
rect 21867 22692 21879 22695
rect 22462 22692 22468 22704
rect 21867 22664 22468 22692
rect 21867 22661 21879 22664
rect 21821 22655 21879 22661
rect 22462 22652 22468 22664
rect 22520 22692 22526 22704
rect 22664 22692 22692 22732
rect 22922 22720 22928 22732
rect 22980 22720 22986 22772
rect 22830 22692 22836 22704
rect 22520 22664 22692 22692
rect 22791 22664 22836 22692
rect 22520 22652 22526 22664
rect 22830 22652 22836 22664
rect 22888 22652 22894 22704
rect 23014 22692 23020 22704
rect 22927 22664 23020 22692
rect 23014 22652 23020 22664
rect 23072 22692 23078 22704
rect 23382 22692 23388 22704
rect 23072 22664 23388 22692
rect 23072 22652 23078 22664
rect 23382 22652 23388 22664
rect 23440 22652 23446 22704
rect 6454 22584 6460 22636
rect 6512 22624 6518 22636
rect 6641 22627 6699 22633
rect 6641 22624 6653 22627
rect 6512 22596 6653 22624
rect 6512 22584 6518 22596
rect 6641 22593 6653 22596
rect 6687 22593 6699 22627
rect 7834 22624 7840 22636
rect 7795 22596 7840 22624
rect 6641 22587 6699 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 8202 22624 8208 22636
rect 8163 22596 8208 22624
rect 8202 22584 8208 22596
rect 8260 22584 8266 22636
rect 8389 22627 8447 22633
rect 8389 22593 8401 22627
rect 8435 22624 8447 22627
rect 9122 22624 9128 22636
rect 8435 22596 9128 22624
rect 8435 22593 8447 22596
rect 8389 22587 8447 22593
rect 9122 22584 9128 22596
rect 9180 22584 9186 22636
rect 9490 22584 9496 22636
rect 9548 22624 9554 22636
rect 9953 22627 10011 22633
rect 9953 22624 9965 22627
rect 9548 22596 9965 22624
rect 9548 22584 9554 22596
rect 9953 22593 9965 22596
rect 9999 22593 10011 22627
rect 9953 22587 10011 22593
rect 12342 22584 12348 22636
rect 12400 22624 12406 22636
rect 12437 22627 12495 22633
rect 12437 22624 12449 22627
rect 12400 22596 12449 22624
rect 12400 22584 12406 22596
rect 12437 22593 12449 22596
rect 12483 22593 12495 22627
rect 12437 22587 12495 22593
rect 12526 22584 12532 22636
rect 12584 22624 12590 22636
rect 12693 22627 12751 22633
rect 12693 22624 12705 22627
rect 12584 22596 12705 22624
rect 12584 22584 12590 22596
rect 12693 22593 12705 22596
rect 12739 22593 12751 22627
rect 15654 22624 15660 22636
rect 15615 22596 15660 22624
rect 12693 22587 12751 22593
rect 15654 22584 15660 22596
rect 15712 22584 15718 22636
rect 17034 22624 17040 22636
rect 16995 22596 17040 22624
rect 17034 22584 17040 22596
rect 17092 22584 17098 22636
rect 18322 22624 18328 22636
rect 18283 22596 18328 22624
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 19150 22624 19156 22636
rect 19111 22596 19156 22624
rect 19150 22584 19156 22596
rect 19208 22584 19214 22636
rect 19889 22627 19947 22633
rect 19889 22593 19901 22627
rect 19935 22624 19947 22627
rect 19978 22624 19984 22636
rect 19935 22596 19984 22624
rect 19935 22593 19947 22596
rect 19889 22587 19947 22593
rect 19978 22584 19984 22596
rect 20036 22584 20042 22636
rect 20714 22624 20720 22636
rect 20675 22596 20720 22624
rect 20714 22584 20720 22596
rect 20772 22584 20778 22636
rect 21266 22584 21272 22636
rect 21324 22624 21330 22636
rect 21994 22627 22052 22633
rect 21994 22624 22006 22627
rect 21324 22596 22006 22624
rect 21324 22584 21330 22596
rect 21994 22593 22006 22596
rect 22040 22593 22052 22627
rect 21994 22587 22052 22593
rect 6365 22559 6423 22565
rect 6365 22556 6377 22559
rect 5776 22528 6377 22556
rect 5776 22516 5782 22528
rect 6365 22525 6377 22528
rect 6411 22525 6423 22559
rect 6365 22519 6423 22525
rect 7926 22516 7932 22568
rect 7984 22556 7990 22568
rect 8021 22559 8079 22565
rect 8021 22556 8033 22559
rect 7984 22528 8033 22556
rect 7984 22516 7990 22528
rect 8021 22525 8033 22528
rect 8067 22525 8079 22559
rect 8021 22519 8079 22525
rect 8113 22559 8171 22565
rect 8113 22525 8125 22559
rect 8159 22556 8171 22559
rect 8294 22556 8300 22568
rect 8159 22528 8300 22556
rect 8159 22525 8171 22528
rect 8113 22519 8171 22525
rect 8036 22488 8064 22519
rect 8294 22516 8300 22528
rect 8352 22516 8358 22568
rect 10229 22559 10287 22565
rect 10229 22525 10241 22559
rect 10275 22556 10287 22559
rect 10318 22556 10324 22568
rect 10275 22528 10324 22556
rect 10275 22525 10287 22528
rect 10229 22519 10287 22525
rect 10318 22516 10324 22528
rect 10376 22516 10382 22568
rect 16853 22559 16911 22565
rect 16853 22525 16865 22559
rect 16899 22556 16911 22559
rect 17402 22556 17408 22568
rect 16899 22528 17408 22556
rect 16899 22525 16911 22528
rect 16853 22519 16911 22525
rect 17402 22516 17408 22528
rect 17460 22516 17466 22568
rect 18414 22516 18420 22568
rect 18472 22556 18478 22568
rect 20533 22559 20591 22565
rect 20533 22556 20545 22559
rect 18472 22528 20545 22556
rect 18472 22516 18478 22528
rect 20533 22525 20545 22528
rect 20579 22525 20591 22559
rect 22649 22559 22707 22565
rect 22649 22556 22661 22559
rect 20533 22519 20591 22525
rect 20640 22528 22661 22556
rect 8938 22488 8944 22500
rect 8036 22460 8944 22488
rect 8938 22448 8944 22460
rect 8996 22448 9002 22500
rect 19702 22448 19708 22500
rect 19760 22488 19766 22500
rect 20640 22488 20668 22528
rect 22649 22525 22661 22528
rect 22695 22525 22707 22559
rect 22649 22519 22707 22525
rect 19760 22460 20668 22488
rect 20717 22491 20775 22497
rect 19760 22448 19766 22460
rect 20717 22457 20729 22491
rect 20763 22488 20775 22491
rect 21542 22488 21548 22500
rect 20763 22460 21548 22488
rect 20763 22457 20775 22460
rect 20717 22451 20775 22457
rect 21542 22448 21548 22460
rect 21600 22448 21606 22500
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 1762 22380 1768 22432
rect 1820 22420 1826 22432
rect 2041 22423 2099 22429
rect 2041 22420 2053 22423
rect 1820 22392 2053 22420
rect 1820 22380 1826 22392
rect 2041 22389 2053 22392
rect 2087 22389 2099 22423
rect 2041 22383 2099 22389
rect 2869 22423 2927 22429
rect 2869 22389 2881 22423
rect 2915 22420 2927 22423
rect 3970 22420 3976 22432
rect 2915 22392 3976 22420
rect 2915 22389 2927 22392
rect 2869 22383 2927 22389
rect 3970 22380 3976 22392
rect 4028 22380 4034 22432
rect 18509 22423 18567 22429
rect 18509 22389 18521 22423
rect 18555 22420 18567 22423
rect 19058 22420 19064 22432
rect 18555 22392 19064 22420
rect 18555 22389 18567 22392
rect 18509 22383 18567 22389
rect 19058 22380 19064 22392
rect 19116 22380 19122 22432
rect 1104 22330 30820 22352
rect 1104 22278 5915 22330
rect 5967 22278 5979 22330
rect 6031 22278 6043 22330
rect 6095 22278 6107 22330
rect 6159 22278 6171 22330
rect 6223 22278 15846 22330
rect 15898 22278 15910 22330
rect 15962 22278 15974 22330
rect 16026 22278 16038 22330
rect 16090 22278 16102 22330
rect 16154 22278 25776 22330
rect 25828 22278 25840 22330
rect 25892 22278 25904 22330
rect 25956 22278 25968 22330
rect 26020 22278 26032 22330
rect 26084 22278 30820 22330
rect 1104 22256 30820 22278
rect 7374 22176 7380 22228
rect 7432 22216 7438 22228
rect 8386 22216 8392 22228
rect 7432 22188 8392 22216
rect 7432 22176 7438 22188
rect 8386 22176 8392 22188
rect 8444 22176 8450 22228
rect 11149 22219 11207 22225
rect 11149 22185 11161 22219
rect 11195 22216 11207 22219
rect 11514 22216 11520 22228
rect 11195 22188 11520 22216
rect 11195 22185 11207 22188
rect 11149 22179 11207 22185
rect 11514 22176 11520 22188
rect 11572 22176 11578 22228
rect 12986 22216 12992 22228
rect 12947 22188 12992 22216
rect 12986 22176 12992 22188
rect 13044 22176 13050 22228
rect 17957 22219 18015 22225
rect 17957 22185 17969 22219
rect 18003 22216 18015 22219
rect 18322 22216 18328 22228
rect 18003 22188 18328 22216
rect 18003 22185 18015 22188
rect 17957 22179 18015 22185
rect 18322 22176 18328 22188
rect 18380 22176 18386 22228
rect 20714 22176 20720 22228
rect 20772 22216 20778 22228
rect 20901 22219 20959 22225
rect 20901 22216 20913 22219
rect 20772 22188 20913 22216
rect 20772 22176 20778 22188
rect 20901 22185 20913 22188
rect 20947 22185 20959 22219
rect 20901 22179 20959 22185
rect 22094 22176 22100 22228
rect 22152 22216 22158 22228
rect 22557 22219 22615 22225
rect 22557 22216 22569 22219
rect 22152 22188 22569 22216
rect 22152 22176 22158 22188
rect 22557 22185 22569 22188
rect 22603 22216 22615 22219
rect 22830 22216 22836 22228
rect 22603 22188 22836 22216
rect 22603 22185 22615 22188
rect 22557 22179 22615 22185
rect 22830 22176 22836 22188
rect 22888 22176 22894 22228
rect 7558 22108 7564 22160
rect 7616 22148 7622 22160
rect 8110 22148 8116 22160
rect 7616 22120 8116 22148
rect 7616 22108 7622 22120
rect 8110 22108 8116 22120
rect 8168 22108 8174 22160
rect 8662 22108 8668 22160
rect 8720 22148 8726 22160
rect 8720 22120 9674 22148
rect 8720 22108 8726 22120
rect 9646 22092 9674 22120
rect 15470 22108 15476 22160
rect 15528 22148 15534 22160
rect 15838 22148 15844 22160
rect 15528 22120 15844 22148
rect 15528 22108 15534 22120
rect 15838 22108 15844 22120
rect 15896 22108 15902 22160
rect 17862 22148 17868 22160
rect 16316 22120 17868 22148
rect 4617 22083 4675 22089
rect 4617 22049 4629 22083
rect 4663 22080 4675 22083
rect 4982 22080 4988 22092
rect 4663 22052 4988 22080
rect 4663 22049 4675 22052
rect 4617 22043 4675 22049
rect 4982 22040 4988 22052
rect 5040 22040 5046 22092
rect 6641 22083 6699 22089
rect 6641 22049 6653 22083
rect 6687 22080 6699 22083
rect 8202 22080 8208 22092
rect 6687 22052 8208 22080
rect 6687 22049 6699 22052
rect 6641 22043 6699 22049
rect 8202 22040 8208 22052
rect 8260 22040 8266 22092
rect 8294 22040 8300 22092
rect 8352 22080 8358 22092
rect 9033 22083 9091 22089
rect 9033 22080 9045 22083
rect 8352 22052 9045 22080
rect 8352 22040 8358 22052
rect 9033 22049 9045 22052
rect 9079 22049 9091 22083
rect 9646 22052 9680 22092
rect 9033 22043 9091 22049
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 15381 22083 15439 22089
rect 15381 22049 15393 22083
rect 15427 22080 15439 22083
rect 15562 22080 15568 22092
rect 15427 22052 15568 22080
rect 15427 22049 15439 22052
rect 15381 22043 15439 22049
rect 15562 22040 15568 22052
rect 15620 22040 15626 22092
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 2866 22012 2872 22024
rect 1903 21984 2872 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 2866 21972 2872 21984
rect 2924 21972 2930 22024
rect 4709 22015 4767 22021
rect 4709 21981 4721 22015
rect 4755 21981 4767 22015
rect 4709 21975 4767 21981
rect 2130 21953 2136 21956
rect 2124 21907 2136 21953
rect 2188 21944 2194 21956
rect 4724 21944 4752 21975
rect 5442 21972 5448 22024
rect 5500 22012 5506 22024
rect 6549 22015 6607 22021
rect 6549 22012 6561 22015
rect 5500 21984 6561 22012
rect 5500 21972 5506 21984
rect 6549 21981 6561 21984
rect 6595 21981 6607 22015
rect 6549 21975 6607 21981
rect 7098 21972 7104 22024
rect 7156 22012 7162 22024
rect 7377 22015 7435 22021
rect 7377 22012 7389 22015
rect 7156 21984 7389 22012
rect 7156 21972 7162 21984
rect 7377 21981 7389 21984
rect 7423 21981 7435 22015
rect 7377 21975 7435 21981
rect 7558 21972 7564 22024
rect 7616 22012 7622 22024
rect 7616 21984 9352 22012
rect 7616 21972 7622 21984
rect 5258 21944 5264 21956
rect 2188 21916 2224 21944
rect 4724 21916 5264 21944
rect 2130 21904 2136 21907
rect 2188 21904 2194 21916
rect 5258 21904 5264 21916
rect 5316 21944 5322 21956
rect 8021 21947 8079 21953
rect 8021 21944 8033 21947
rect 5316 21916 8033 21944
rect 5316 21904 5322 21916
rect 8021 21913 8033 21916
rect 8067 21913 8079 21947
rect 8021 21907 8079 21913
rect 8205 21947 8263 21953
rect 8205 21913 8217 21947
rect 8251 21913 8263 21947
rect 8205 21907 8263 21913
rect 3050 21836 3056 21888
rect 3108 21876 3114 21888
rect 3237 21879 3295 21885
rect 3237 21876 3249 21879
rect 3108 21848 3249 21876
rect 3108 21836 3114 21848
rect 3237 21845 3249 21848
rect 3283 21845 3295 21879
rect 3237 21839 3295 21845
rect 6730 21836 6736 21888
rect 6788 21876 6794 21888
rect 7469 21879 7527 21885
rect 7469 21876 7481 21879
rect 6788 21848 7481 21876
rect 6788 21836 6794 21848
rect 7469 21845 7481 21848
rect 7515 21876 7527 21879
rect 7834 21876 7840 21888
rect 7515 21848 7840 21876
rect 7515 21845 7527 21848
rect 7469 21839 7527 21845
rect 7834 21836 7840 21848
rect 7892 21836 7898 21888
rect 8220 21876 8248 21907
rect 8294 21904 8300 21956
rect 8352 21944 8358 21956
rect 8389 21947 8447 21953
rect 8389 21944 8401 21947
rect 8352 21916 8401 21944
rect 8352 21904 8358 21916
rect 8389 21913 8401 21916
rect 8435 21913 8447 21947
rect 8389 21907 8447 21913
rect 9217 21947 9275 21953
rect 9217 21913 9229 21947
rect 9263 21913 9275 21947
rect 9324 21944 9352 21984
rect 9398 21972 9404 22024
rect 9456 22012 9462 22024
rect 10042 22021 10048 22024
rect 9769 22015 9827 22021
rect 9769 22012 9781 22015
rect 9456 21984 9781 22012
rect 9456 21972 9462 21984
rect 9769 21981 9781 21984
rect 9815 21981 9827 22015
rect 9769 21975 9827 21981
rect 10036 21975 10048 22021
rect 10100 22012 10106 22024
rect 10100 21984 10136 22012
rect 10042 21972 10048 21975
rect 10100 21972 10106 21984
rect 11514 21972 11520 22024
rect 11572 22012 11578 22024
rect 11609 22015 11667 22021
rect 11609 22012 11621 22015
rect 11572 21984 11621 22012
rect 11572 21972 11578 21984
rect 11609 21981 11621 21984
rect 11655 22012 11667 22015
rect 12342 22012 12348 22024
rect 11655 21984 12348 22012
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 12342 21972 12348 21984
rect 12400 21972 12406 22024
rect 15470 22012 15476 22024
rect 15528 22021 15534 22024
rect 15388 21984 15476 22012
rect 15470 21972 15476 21984
rect 15528 22012 15536 22021
rect 16316 22012 16344 22120
rect 17862 22108 17868 22120
rect 17920 22108 17926 22160
rect 19150 22148 19156 22160
rect 17972 22120 19156 22148
rect 16574 22080 16580 22092
rect 16535 22052 16580 22080
rect 16574 22040 16580 22052
rect 16632 22040 16638 22092
rect 16945 22083 17003 22089
rect 16945 22049 16957 22083
rect 16991 22080 17003 22083
rect 17218 22080 17224 22092
rect 16991 22052 17224 22080
rect 16991 22049 17003 22052
rect 16945 22043 17003 22049
rect 17218 22040 17224 22052
rect 17276 22080 17282 22092
rect 17972 22080 18000 22120
rect 19150 22108 19156 22120
rect 19208 22108 19214 22160
rect 17276 22052 18000 22080
rect 17276 22040 17282 22052
rect 18046 22040 18052 22092
rect 18104 22080 18110 22092
rect 18417 22083 18475 22089
rect 18417 22080 18429 22083
rect 18104 22052 18429 22080
rect 18104 22040 18110 22052
rect 18417 22049 18429 22052
rect 18463 22049 18475 22083
rect 18598 22080 18604 22092
rect 18559 22052 18604 22080
rect 18417 22043 18475 22049
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 19242 22040 19248 22092
rect 19300 22080 19306 22092
rect 19705 22083 19763 22089
rect 19705 22080 19717 22083
rect 19300 22052 19717 22080
rect 19300 22040 19306 22052
rect 19705 22049 19717 22052
rect 19751 22049 19763 22083
rect 19886 22080 19892 22092
rect 19847 22052 19892 22080
rect 19705 22043 19763 22049
rect 19886 22040 19892 22052
rect 19944 22040 19950 22092
rect 20533 22083 20591 22089
rect 20533 22049 20545 22083
rect 20579 22080 20591 22083
rect 20806 22080 20812 22092
rect 20579 22052 20812 22080
rect 20579 22049 20591 22052
rect 20533 22043 20591 22049
rect 20806 22040 20812 22052
rect 20864 22040 20870 22092
rect 22002 22040 22008 22092
rect 22060 22080 22066 22092
rect 22060 22052 22508 22080
rect 22060 22040 22066 22052
rect 16482 22012 16488 22024
rect 15528 21984 16344 22012
rect 16443 21984 16488 22012
rect 15528 21975 15536 21984
rect 15528 21972 15534 21975
rect 16482 21972 16488 21984
rect 16540 21972 16546 22024
rect 16669 22015 16727 22021
rect 16669 21981 16681 22015
rect 16715 21981 16727 22015
rect 16669 21975 16727 21981
rect 16761 22015 16819 22021
rect 16761 21981 16773 22015
rect 16807 22012 16819 22015
rect 16850 22012 16856 22024
rect 16807 21984 16856 22012
rect 16807 21981 16819 21984
rect 16761 21975 16819 21981
rect 9950 21944 9956 21956
rect 9324 21916 9956 21944
rect 9217 21907 9275 21913
rect 8570 21876 8576 21888
rect 8220 21848 8576 21876
rect 8570 21836 8576 21848
rect 8628 21876 8634 21888
rect 9232 21876 9260 21907
rect 9950 21904 9956 21916
rect 10008 21904 10014 21956
rect 11882 21953 11888 21956
rect 11876 21907 11888 21953
rect 11940 21944 11946 21956
rect 15105 21947 15163 21953
rect 11940 21916 11976 21944
rect 11882 21904 11888 21907
rect 11940 21904 11946 21916
rect 15105 21913 15117 21947
rect 15151 21913 15163 21947
rect 15286 21944 15292 21956
rect 15247 21916 15292 21944
rect 15105 21907 15163 21913
rect 8628 21848 9260 21876
rect 8628 21836 8634 21848
rect 14366 21836 14372 21888
rect 14424 21876 14430 21888
rect 15120 21876 15148 21907
rect 15286 21904 15292 21916
rect 15344 21904 15350 21956
rect 15378 21904 15384 21956
rect 15436 21944 15442 21956
rect 16684 21944 16712 21975
rect 16850 21972 16856 21984
rect 16908 21972 16914 22024
rect 17037 22015 17095 22021
rect 17037 21981 17049 22015
rect 17083 22012 17095 22015
rect 17862 22012 17868 22024
rect 17083 21984 17868 22012
rect 17083 21981 17095 21984
rect 17037 21975 17095 21981
rect 17862 21972 17868 21984
rect 17920 21972 17926 22024
rect 19426 22012 19432 22024
rect 18156 21984 19432 22012
rect 17126 21944 17132 21956
rect 15436 21916 15481 21944
rect 16684 21916 17132 21944
rect 15436 21904 15442 21916
rect 17126 21904 17132 21916
rect 17184 21904 17190 21956
rect 18156 21876 18184 21984
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 19978 21972 19984 22024
rect 20036 22012 20042 22024
rect 20441 22015 20499 22021
rect 20441 22012 20453 22015
rect 20036 21984 20453 22012
rect 20036 21972 20042 21984
rect 20441 21981 20453 21984
rect 20487 21981 20499 22015
rect 20714 22012 20720 22024
rect 20675 21984 20720 22012
rect 20441 21975 20499 21981
rect 20714 21972 20720 21984
rect 20772 21972 20778 22024
rect 21821 22015 21879 22021
rect 21821 21981 21833 22015
rect 21867 22012 21879 22015
rect 22094 22012 22100 22024
rect 21867 21984 22100 22012
rect 21867 21981 21879 21984
rect 21821 21975 21879 21981
rect 22094 21972 22100 21984
rect 22152 21972 22158 22024
rect 22480 22021 22508 22052
rect 22465 22015 22523 22021
rect 22465 21981 22477 22015
rect 22511 21981 22523 22015
rect 22465 21975 22523 21981
rect 18325 21947 18383 21953
rect 18325 21913 18337 21947
rect 18371 21944 18383 21947
rect 19613 21947 19671 21953
rect 19613 21944 19625 21947
rect 18371 21916 19625 21944
rect 18371 21913 18383 21916
rect 18325 21907 18383 21913
rect 19613 21913 19625 21916
rect 19659 21944 19671 21947
rect 19702 21944 19708 21956
rect 19659 21916 19708 21944
rect 19659 21913 19671 21916
rect 19613 21907 19671 21913
rect 19702 21904 19708 21916
rect 19760 21904 19766 21956
rect 21450 21904 21456 21956
rect 21508 21944 21514 21956
rect 21637 21947 21695 21953
rect 21637 21944 21649 21947
rect 21508 21916 21649 21944
rect 21508 21904 21514 21916
rect 21637 21913 21649 21916
rect 21683 21913 21695 21947
rect 21637 21907 21695 21913
rect 22005 21947 22063 21953
rect 22005 21913 22017 21947
rect 22051 21944 22063 21947
rect 22370 21944 22376 21956
rect 22051 21916 22376 21944
rect 22051 21913 22063 21916
rect 22005 21907 22063 21913
rect 22370 21904 22376 21916
rect 22428 21904 22434 21956
rect 14424 21848 18184 21876
rect 19245 21879 19303 21885
rect 14424 21836 14430 21848
rect 19245 21845 19257 21879
rect 19291 21876 19303 21879
rect 19518 21876 19524 21888
rect 19291 21848 19524 21876
rect 19291 21845 19303 21848
rect 19245 21839 19303 21845
rect 19518 21836 19524 21848
rect 19576 21836 19582 21888
rect 1104 21786 30820 21808
rect 1104 21734 10880 21786
rect 10932 21734 10944 21786
rect 10996 21734 11008 21786
rect 11060 21734 11072 21786
rect 11124 21734 11136 21786
rect 11188 21734 20811 21786
rect 20863 21734 20875 21786
rect 20927 21734 20939 21786
rect 20991 21734 21003 21786
rect 21055 21734 21067 21786
rect 21119 21734 30820 21786
rect 1104 21712 30820 21734
rect 7653 21675 7711 21681
rect 7653 21641 7665 21675
rect 7699 21672 7711 21675
rect 7742 21672 7748 21684
rect 7699 21644 7748 21672
rect 7699 21641 7711 21644
rect 7653 21635 7711 21641
rect 7742 21632 7748 21644
rect 7800 21632 7806 21684
rect 8202 21632 8208 21684
rect 8260 21632 8266 21684
rect 8941 21675 8999 21681
rect 8941 21641 8953 21675
rect 8987 21672 8999 21675
rect 10781 21675 10839 21681
rect 8987 21644 9700 21672
rect 8987 21641 8999 21644
rect 8941 21635 8999 21641
rect 2866 21604 2872 21616
rect 1964 21576 2872 21604
rect 1964 21545 1992 21576
rect 2866 21564 2872 21576
rect 2924 21564 2930 21616
rect 5442 21564 5448 21616
rect 5500 21604 5506 21616
rect 6733 21607 6791 21613
rect 6733 21604 6745 21607
rect 5500 21576 6745 21604
rect 5500 21564 5506 21576
rect 6733 21573 6745 21576
rect 6779 21604 6791 21607
rect 7558 21604 7564 21616
rect 6779 21576 7564 21604
rect 6779 21573 6791 21576
rect 6733 21567 6791 21573
rect 7558 21564 7564 21576
rect 7616 21564 7622 21616
rect 8220 21604 8248 21632
rect 9672 21613 9700 21644
rect 10781 21641 10793 21675
rect 10827 21641 10839 21675
rect 10781 21635 10839 21641
rect 12253 21675 12311 21681
rect 12253 21641 12265 21675
rect 12299 21672 12311 21675
rect 12526 21672 12532 21684
rect 12299 21644 12532 21672
rect 12299 21641 12311 21644
rect 12253 21635 12311 21641
rect 8573 21607 8631 21613
rect 8573 21604 8585 21607
rect 8220 21576 8585 21604
rect 8573 21573 8585 21576
rect 8619 21573 8631 21607
rect 8573 21567 8631 21573
rect 9657 21607 9715 21613
rect 9657 21573 9669 21607
rect 9703 21573 9715 21607
rect 9657 21567 9715 21573
rect 2222 21545 2228 21548
rect 1949 21539 2007 21545
rect 1949 21505 1961 21539
rect 1995 21505 2007 21539
rect 1949 21499 2007 21505
rect 2216 21499 2228 21545
rect 2280 21536 2286 21548
rect 6546 21545 6552 21548
rect 3789 21539 3847 21545
rect 3789 21536 3801 21539
rect 2280 21508 2316 21536
rect 3344 21508 3801 21536
rect 2222 21496 2228 21499
rect 2280 21496 2286 21508
rect 2958 21292 2964 21344
rect 3016 21332 3022 21344
rect 3344 21341 3372 21508
rect 3789 21505 3801 21508
rect 3835 21505 3847 21539
rect 6544 21536 6552 21545
rect 6507 21508 6552 21536
rect 3789 21499 3847 21505
rect 6544 21499 6552 21508
rect 6546 21496 6552 21499
rect 6604 21496 6610 21548
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21505 6699 21539
rect 6641 21499 6699 21505
rect 6454 21428 6460 21480
rect 6512 21468 6518 21480
rect 6656 21468 6684 21499
rect 6822 21496 6828 21548
rect 6880 21545 6886 21548
rect 6880 21539 6919 21545
rect 6907 21505 6919 21539
rect 6880 21499 6919 21505
rect 7009 21539 7067 21545
rect 7009 21505 7021 21539
rect 7055 21505 7067 21539
rect 7009 21499 7067 21505
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21536 7803 21539
rect 8202 21536 8208 21548
rect 7791 21508 8208 21536
rect 7791 21505 7803 21508
rect 7745 21499 7803 21505
rect 6880 21496 6886 21499
rect 6512 21440 6684 21468
rect 7024 21468 7052 21499
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 8304 21539 8362 21545
rect 8304 21505 8316 21539
rect 8350 21505 8362 21539
rect 8304 21499 8362 21505
rect 8390 21539 8448 21545
rect 8390 21505 8402 21539
rect 8436 21505 8448 21539
rect 8673 21539 8731 21545
rect 8673 21534 8685 21539
rect 8390 21499 8448 21505
rect 8516 21506 8685 21534
rect 7834 21468 7840 21480
rect 7024 21440 7840 21468
rect 6512 21428 6518 21440
rect 3329 21335 3387 21341
rect 3329 21332 3341 21335
rect 3016 21304 3341 21332
rect 3016 21292 3022 21304
rect 3329 21301 3341 21304
rect 3375 21301 3387 21335
rect 3329 21295 3387 21301
rect 3881 21335 3939 21341
rect 3881 21301 3893 21335
rect 3927 21332 3939 21335
rect 6270 21332 6276 21344
rect 3927 21304 6276 21332
rect 3927 21301 3939 21304
rect 3881 21295 3939 21301
rect 6270 21292 6276 21304
rect 6328 21292 6334 21344
rect 6365 21335 6423 21341
rect 6365 21301 6377 21335
rect 6411 21332 6423 21335
rect 6546 21332 6552 21344
rect 6411 21304 6552 21332
rect 6411 21301 6423 21304
rect 6365 21295 6423 21301
rect 6546 21292 6552 21304
rect 6604 21292 6610 21344
rect 6656 21332 6684 21440
rect 7834 21428 7840 21440
rect 7892 21468 7898 21480
rect 8312 21468 8340 21499
rect 7892 21440 8340 21468
rect 7892 21428 7898 21440
rect 8404 21412 8432 21499
rect 8386 21360 8392 21412
rect 8444 21360 8450 21412
rect 8516 21400 8544 21506
rect 8673 21505 8685 21506
rect 8719 21505 8731 21539
rect 8673 21499 8731 21505
rect 8803 21539 8861 21545
rect 8803 21505 8815 21539
rect 8849 21536 8861 21539
rect 9214 21536 9220 21548
rect 8849 21508 9220 21536
rect 8849 21505 8861 21508
rect 8803 21499 8861 21505
rect 9214 21496 9220 21508
rect 9272 21496 9278 21548
rect 9490 21496 9496 21548
rect 9548 21534 9554 21548
rect 10502 21536 10508 21548
rect 9646 21534 10508 21536
rect 9548 21508 10508 21534
rect 9548 21506 9674 21508
rect 9548 21496 9554 21506
rect 10502 21496 10508 21508
rect 10560 21536 10566 21548
rect 10796 21536 10824 21635
rect 12526 21632 12532 21644
rect 12584 21632 12590 21684
rect 14921 21675 14979 21681
rect 14921 21641 14933 21675
rect 14967 21672 14979 21675
rect 15286 21672 15292 21684
rect 14967 21644 15292 21672
rect 14967 21641 14979 21644
rect 14921 21635 14979 21641
rect 15286 21632 15292 21644
rect 15344 21632 15350 21684
rect 16482 21632 16488 21684
rect 16540 21672 16546 21684
rect 17405 21675 17463 21681
rect 17405 21672 17417 21675
rect 16540 21644 17417 21672
rect 16540 21632 16546 21644
rect 17405 21641 17417 21644
rect 17451 21641 17463 21675
rect 17862 21672 17868 21684
rect 17823 21644 17868 21672
rect 17405 21635 17463 21641
rect 17862 21632 17868 21644
rect 17920 21632 17926 21684
rect 18138 21632 18144 21684
rect 18196 21672 18202 21684
rect 18325 21675 18383 21681
rect 18325 21672 18337 21675
rect 18196 21644 18337 21672
rect 18196 21632 18202 21644
rect 18325 21641 18337 21644
rect 18371 21641 18383 21675
rect 18325 21635 18383 21641
rect 19334 21632 19340 21684
rect 19392 21632 19398 21684
rect 20438 21632 20444 21684
rect 20496 21672 20502 21684
rect 20993 21675 21051 21681
rect 20993 21672 21005 21675
rect 20496 21644 21005 21672
rect 20496 21632 20502 21644
rect 20993 21641 21005 21644
rect 21039 21641 21051 21675
rect 20993 21635 21051 21641
rect 10560 21508 10824 21536
rect 10888 21576 11744 21604
rect 10560 21496 10566 21508
rect 9398 21428 9404 21480
rect 9456 21468 9462 21480
rect 9456 21440 9501 21468
rect 9456 21428 9462 21440
rect 8662 21400 8668 21412
rect 8516 21372 8668 21400
rect 8662 21360 8668 21372
rect 8720 21360 8726 21412
rect 7374 21332 7380 21344
rect 6656 21304 7380 21332
rect 7374 21292 7380 21304
rect 7432 21292 7438 21344
rect 7650 21292 7656 21344
rect 7708 21332 7714 21344
rect 10888 21332 10916 21576
rect 11517 21539 11575 21545
rect 11517 21505 11529 21539
rect 11563 21536 11575 21539
rect 11606 21536 11612 21548
rect 11563 21508 11612 21536
rect 11563 21505 11575 21508
rect 11517 21499 11575 21505
rect 11606 21496 11612 21508
rect 11664 21496 11670 21548
rect 11716 21545 11744 21576
rect 12986 21564 12992 21616
rect 13044 21604 13050 21616
rect 15381 21607 15439 21613
rect 15381 21604 15393 21607
rect 13044 21576 15393 21604
rect 13044 21564 13050 21576
rect 15381 21573 15393 21576
rect 15427 21573 15439 21607
rect 17770 21604 17776 21616
rect 15381 21567 15439 21573
rect 16960 21576 17776 21604
rect 11701 21539 11759 21545
rect 11701 21505 11713 21539
rect 11747 21505 11759 21539
rect 11701 21499 11759 21505
rect 11790 21496 11796 21548
rect 11848 21536 11854 21548
rect 12069 21539 12127 21545
rect 11848 21508 11893 21536
rect 11848 21496 11854 21508
rect 12069 21505 12081 21539
rect 12115 21536 12127 21539
rect 13722 21536 13728 21548
rect 12115 21508 13728 21536
rect 12115 21505 12127 21508
rect 12069 21499 12127 21505
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 15286 21536 15292 21548
rect 15247 21508 15292 21536
rect 15286 21496 15292 21508
rect 15344 21496 15350 21548
rect 15562 21496 15568 21548
rect 15620 21536 15626 21548
rect 16669 21539 16727 21545
rect 16669 21536 16681 21539
rect 15620 21508 16681 21536
rect 15620 21496 15626 21508
rect 16669 21505 16681 21508
rect 16715 21505 16727 21539
rect 16669 21499 16727 21505
rect 16758 21496 16764 21548
rect 16816 21536 16822 21548
rect 16960 21545 16988 21576
rect 17770 21564 17776 21576
rect 17828 21564 17834 21616
rect 19352 21604 19380 21632
rect 20073 21607 20131 21613
rect 20073 21604 20085 21607
rect 18340 21576 20085 21604
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16816 21508 16865 21536
rect 16816 21496 16822 21508
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 16945 21539 17003 21545
rect 16945 21505 16957 21539
rect 16991 21505 17003 21539
rect 17218 21536 17224 21548
rect 17179 21508 17224 21536
rect 16945 21499 17003 21505
rect 17218 21496 17224 21508
rect 17276 21496 17282 21548
rect 17862 21496 17868 21548
rect 17920 21536 17926 21548
rect 18233 21539 18291 21545
rect 18233 21536 18245 21539
rect 17920 21508 18245 21536
rect 17920 21496 17926 21508
rect 18233 21505 18245 21508
rect 18279 21505 18291 21539
rect 18233 21499 18291 21505
rect 11882 21428 11888 21480
rect 11940 21468 11946 21480
rect 15473 21471 15531 21477
rect 11940 21440 11985 21468
rect 11940 21428 11946 21440
rect 15473 21437 15485 21471
rect 15519 21468 15531 21471
rect 15838 21468 15844 21480
rect 15519 21440 15844 21468
rect 15519 21437 15531 21440
rect 15473 21431 15531 21437
rect 15838 21428 15844 21440
rect 15896 21468 15902 21480
rect 16482 21468 16488 21480
rect 15896 21440 16488 21468
rect 15896 21428 15902 21440
rect 16482 21428 16488 21440
rect 16540 21428 16546 21480
rect 17037 21471 17095 21477
rect 17037 21437 17049 21471
rect 17083 21468 17095 21471
rect 18340 21468 18368 21576
rect 20073 21573 20085 21576
rect 20119 21573 20131 21607
rect 20073 21567 20131 21573
rect 19058 21536 19064 21548
rect 19019 21508 19064 21536
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 19234 21539 19292 21545
rect 19234 21536 19246 21539
rect 19168 21508 19246 21536
rect 17083 21440 18368 21468
rect 17083 21437 17095 21440
rect 17037 21431 17095 21437
rect 18414 21428 18420 21480
rect 18472 21468 18478 21480
rect 18598 21468 18604 21480
rect 18472 21440 18604 21468
rect 18472 21428 18478 21440
rect 18598 21428 18604 21440
rect 18656 21468 18662 21480
rect 19168 21468 19196 21508
rect 19234 21505 19246 21508
rect 19280 21505 19292 21539
rect 19234 21499 19292 21505
rect 19334 21496 19340 21548
rect 19392 21536 19398 21548
rect 19392 21508 19437 21536
rect 19392 21496 19398 21508
rect 19518 21496 19524 21548
rect 19576 21536 19582 21548
rect 19613 21539 19671 21545
rect 19613 21536 19625 21539
rect 19576 21508 19625 21536
rect 19576 21496 19582 21508
rect 19613 21505 19625 21508
rect 19659 21505 19671 21539
rect 20254 21536 20260 21548
rect 20215 21508 20260 21536
rect 19613 21499 19671 21505
rect 20254 21496 20260 21508
rect 20312 21496 20318 21548
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21536 21143 21539
rect 21450 21536 21456 21548
rect 21131 21508 21456 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 21450 21496 21456 21508
rect 21508 21496 21514 21548
rect 29825 21539 29883 21545
rect 29825 21505 29837 21539
rect 29871 21536 29883 21539
rect 29914 21536 29920 21548
rect 29871 21508 29920 21536
rect 29871 21505 29883 21508
rect 29825 21499 29883 21505
rect 29914 21496 29920 21508
rect 29972 21496 29978 21548
rect 19886 21468 19892 21480
rect 18656 21440 19892 21468
rect 18656 21428 18662 21440
rect 19886 21428 19892 21440
rect 19944 21428 19950 21480
rect 15102 21360 15108 21412
rect 15160 21400 15166 21412
rect 15562 21400 15568 21412
rect 15160 21372 15568 21400
rect 15160 21360 15166 21372
rect 15562 21360 15568 21372
rect 15620 21360 15626 21412
rect 19150 21360 19156 21412
rect 19208 21400 19214 21412
rect 19208 21372 19564 21400
rect 19208 21360 19214 21372
rect 19536 21344 19564 21372
rect 7708 21304 10916 21332
rect 7708 21292 7714 21304
rect 16942 21292 16948 21344
rect 17000 21332 17006 21344
rect 17862 21332 17868 21344
rect 17000 21304 17868 21332
rect 17000 21292 17006 21304
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 19061 21335 19119 21341
rect 19061 21301 19073 21335
rect 19107 21332 19119 21335
rect 19242 21332 19248 21344
rect 19107 21304 19248 21332
rect 19107 21301 19119 21304
rect 19061 21295 19119 21301
rect 19242 21292 19248 21304
rect 19300 21292 19306 21344
rect 19518 21332 19524 21344
rect 19479 21304 19524 21332
rect 19518 21292 19524 21304
rect 19576 21292 19582 21344
rect 20441 21335 20499 21341
rect 20441 21301 20453 21335
rect 20487 21332 20499 21335
rect 20530 21332 20536 21344
rect 20487 21304 20536 21332
rect 20487 21301 20499 21304
rect 20441 21295 20499 21301
rect 20530 21292 20536 21304
rect 20588 21292 20594 21344
rect 30006 21332 30012 21344
rect 29967 21304 30012 21332
rect 30006 21292 30012 21304
rect 30064 21292 30070 21344
rect 1104 21242 30820 21264
rect 1104 21190 5915 21242
rect 5967 21190 5979 21242
rect 6031 21190 6043 21242
rect 6095 21190 6107 21242
rect 6159 21190 6171 21242
rect 6223 21190 15846 21242
rect 15898 21190 15910 21242
rect 15962 21190 15974 21242
rect 16026 21190 16038 21242
rect 16090 21190 16102 21242
rect 16154 21190 25776 21242
rect 25828 21190 25840 21242
rect 25892 21190 25904 21242
rect 25956 21190 25968 21242
rect 26020 21190 26032 21242
rect 26084 21190 30820 21242
rect 1104 21168 30820 21190
rect 2222 21088 2228 21140
rect 2280 21128 2286 21140
rect 2317 21131 2375 21137
rect 2317 21128 2329 21131
rect 2280 21100 2329 21128
rect 2280 21088 2286 21100
rect 2317 21097 2329 21100
rect 2363 21097 2375 21131
rect 5442 21128 5448 21140
rect 5403 21100 5448 21128
rect 2317 21091 2375 21097
rect 5442 21088 5448 21100
rect 5500 21088 5506 21140
rect 6638 21088 6644 21140
rect 6696 21128 6702 21140
rect 6822 21128 6828 21140
rect 6696 21100 6828 21128
rect 6696 21088 6702 21100
rect 6822 21088 6828 21100
rect 6880 21128 6886 21140
rect 7377 21131 7435 21137
rect 7377 21128 7389 21131
rect 6880 21100 7389 21128
rect 6880 21088 6886 21100
rect 7377 21097 7389 21100
rect 7423 21097 7435 21131
rect 8202 21128 8208 21140
rect 8163 21100 8208 21128
rect 7377 21091 7435 21097
rect 8202 21088 8208 21100
rect 8260 21088 8266 21140
rect 8389 21131 8447 21137
rect 8389 21097 8401 21131
rect 8435 21128 8447 21131
rect 8478 21128 8484 21140
rect 8435 21100 8484 21128
rect 8435 21097 8447 21100
rect 8389 21091 8447 21097
rect 8478 21088 8484 21100
rect 8536 21088 8542 21140
rect 9214 21088 9220 21140
rect 9272 21128 9278 21140
rect 10318 21128 10324 21140
rect 9272 21100 10324 21128
rect 9272 21088 9278 21100
rect 10318 21088 10324 21100
rect 10376 21088 10382 21140
rect 16758 21128 16764 21140
rect 16719 21100 16764 21128
rect 16758 21088 16764 21100
rect 16816 21088 16822 21140
rect 17126 21088 17132 21140
rect 17184 21128 17190 21140
rect 17221 21131 17279 21137
rect 17221 21128 17233 21131
rect 17184 21100 17233 21128
rect 17184 21088 17190 21100
rect 17221 21097 17233 21100
rect 17267 21097 17279 21131
rect 17221 21091 17279 21097
rect 17862 21088 17868 21140
rect 17920 21128 17926 21140
rect 19245 21131 19303 21137
rect 17920 21100 18552 21128
rect 17920 21088 17926 21100
rect 7926 21020 7932 21072
rect 7984 21060 7990 21072
rect 10413 21063 10471 21069
rect 10413 21060 10425 21063
rect 7984 21032 10425 21060
rect 7984 21020 7990 21032
rect 10413 21029 10425 21032
rect 10459 21029 10471 21063
rect 17586 21060 17592 21072
rect 10413 21023 10471 21029
rect 15488 21032 17592 21060
rect 1946 20992 1952 21004
rect 1859 20964 1952 20992
rect 1946 20952 1952 20964
rect 2004 20992 2010 21004
rect 4157 20995 4215 21001
rect 4157 20992 4169 20995
rect 2004 20964 4169 20992
rect 2004 20952 2010 20964
rect 4157 20961 4169 20964
rect 4203 20992 4215 20995
rect 4430 20992 4436 21004
rect 4203 20964 4436 20992
rect 4203 20961 4215 20964
rect 4157 20955 4215 20961
rect 4430 20952 4436 20964
rect 4488 20952 4494 21004
rect 7374 20952 7380 21004
rect 7432 20992 7438 21004
rect 8478 20992 8484 21004
rect 7432 20964 8484 20992
rect 7432 20952 7438 20964
rect 8478 20952 8484 20964
rect 8536 20952 8542 21004
rect 9582 20952 9588 21004
rect 9640 20992 9646 21004
rect 15488 21001 15516 21032
rect 17586 21020 17592 21032
rect 17644 21020 17650 21072
rect 18414 21060 18420 21072
rect 17788 21032 18420 21060
rect 9677 20995 9735 21001
rect 9677 20992 9689 20995
rect 9640 20964 9689 20992
rect 9640 20952 9646 20964
rect 9677 20961 9689 20964
rect 9723 20961 9735 20995
rect 9677 20955 9735 20961
rect 15473 20995 15531 21001
rect 15473 20961 15485 20995
rect 15519 20961 15531 20995
rect 15473 20955 15531 20961
rect 16209 20995 16267 21001
rect 16209 20961 16221 20995
rect 16255 20992 16267 20995
rect 17402 20992 17408 21004
rect 16255 20964 17408 20992
rect 16255 20961 16267 20964
rect 16209 20955 16267 20961
rect 17402 20952 17408 20964
rect 17460 20952 17466 21004
rect 17788 21001 17816 21032
rect 18414 21020 18420 21032
rect 18472 21020 18478 21072
rect 18524 21060 18552 21100
rect 19245 21097 19257 21131
rect 19291 21128 19303 21131
rect 19334 21128 19340 21140
rect 19291 21100 19340 21128
rect 19291 21097 19303 21100
rect 19245 21091 19303 21097
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 19702 21128 19708 21140
rect 19663 21100 19708 21128
rect 19702 21088 19708 21100
rect 19760 21088 19766 21140
rect 20714 21060 20720 21072
rect 18524 21032 20720 21060
rect 20714 21020 20720 21032
rect 20772 21060 20778 21072
rect 21729 21063 21787 21069
rect 21729 21060 21741 21063
rect 20772 21032 21741 21060
rect 20772 21020 20778 21032
rect 21729 21029 21741 21032
rect 21775 21029 21787 21063
rect 21729 21023 21787 21029
rect 17773 20995 17831 21001
rect 17773 20961 17785 20995
rect 17819 20961 17831 20995
rect 17773 20955 17831 20961
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20893 1639 20927
rect 1762 20924 1768 20936
rect 1723 20896 1768 20924
rect 1581 20887 1639 20893
rect 1394 20748 1400 20800
rect 1452 20788 1458 20800
rect 1596 20788 1624 20887
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 1854 20884 1860 20936
rect 1912 20924 1918 20936
rect 2133 20927 2191 20933
rect 1912 20896 1957 20924
rect 1912 20884 1918 20896
rect 2133 20893 2145 20927
rect 2179 20924 2191 20927
rect 2958 20924 2964 20936
rect 2179 20896 2964 20924
rect 2179 20893 2191 20896
rect 2133 20887 2191 20893
rect 2958 20884 2964 20896
rect 3016 20884 3022 20936
rect 3050 20884 3056 20936
rect 3108 20924 3114 20936
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 3108 20896 3153 20924
rect 3344 20896 3801 20924
rect 3108 20884 3114 20896
rect 3344 20868 3372 20896
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3970 20924 3976 20936
rect 3931 20896 3976 20924
rect 3789 20887 3847 20893
rect 3970 20884 3976 20896
rect 4028 20884 4034 20936
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20924 4123 20927
rect 4341 20927 4399 20933
rect 4111 20896 4200 20924
rect 4111 20893 4123 20896
rect 4065 20887 4123 20893
rect 4172 20868 4200 20896
rect 4341 20893 4353 20927
rect 4387 20924 4399 20927
rect 5166 20924 5172 20936
rect 4387 20896 5172 20924
rect 4387 20893 4399 20896
rect 4341 20887 4399 20893
rect 5166 20884 5172 20896
rect 5224 20884 5230 20936
rect 6546 20884 6552 20936
rect 6604 20933 6610 20936
rect 6604 20924 6616 20933
rect 6604 20896 6649 20924
rect 6604 20887 6616 20896
rect 6604 20884 6610 20887
rect 6730 20884 6736 20936
rect 6788 20924 6794 20936
rect 6825 20927 6883 20933
rect 6825 20924 6837 20927
rect 6788 20896 6837 20924
rect 6788 20884 6794 20896
rect 6825 20893 6837 20896
rect 6871 20893 6883 20927
rect 6825 20887 6883 20893
rect 6914 20884 6920 20936
rect 6972 20924 6978 20936
rect 7469 20927 7527 20933
rect 7469 20924 7481 20927
rect 6972 20896 7481 20924
rect 6972 20884 6978 20896
rect 7469 20893 7481 20896
rect 7515 20893 7527 20927
rect 7926 20924 7932 20936
rect 7887 20896 7932 20924
rect 7469 20887 7527 20893
rect 7926 20884 7932 20896
rect 7984 20884 7990 20936
rect 9306 20884 9312 20936
rect 9364 20924 9370 20936
rect 9953 20927 10011 20933
rect 9953 20924 9965 20927
rect 9364 20896 9965 20924
rect 9364 20884 9370 20896
rect 9953 20893 9965 20896
rect 9999 20893 10011 20927
rect 13354 20924 13360 20936
rect 13315 20896 13360 20924
rect 9953 20887 10011 20893
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 13449 20927 13507 20933
rect 13449 20893 13461 20927
rect 13495 20924 13507 20927
rect 16301 20927 16359 20933
rect 16301 20924 16313 20927
rect 13495 20896 16313 20924
rect 13495 20893 13507 20896
rect 13449 20887 13507 20893
rect 16301 20893 16313 20896
rect 16347 20924 16359 20927
rect 17681 20927 17739 20933
rect 17681 20924 17693 20927
rect 16347 20896 17693 20924
rect 16347 20893 16359 20896
rect 16301 20887 16359 20893
rect 17681 20893 17693 20896
rect 17727 20893 17739 20927
rect 17681 20887 17739 20893
rect 3326 20856 3332 20868
rect 2746 20828 3332 20856
rect 2746 20788 2774 20828
rect 3326 20816 3332 20828
rect 3384 20816 3390 20868
rect 4154 20816 4160 20868
rect 4212 20816 4218 20868
rect 7098 20856 7104 20868
rect 4356 20828 7104 20856
rect 1452 20760 2774 20788
rect 3145 20791 3203 20797
rect 1452 20748 1458 20760
rect 3145 20757 3157 20791
rect 3191 20788 3203 20791
rect 4356 20788 4384 20828
rect 7098 20816 7104 20828
rect 7156 20816 7162 20868
rect 9674 20856 9680 20868
rect 9587 20828 9680 20856
rect 9646 20816 9680 20828
rect 9732 20856 9738 20868
rect 10410 20856 10416 20868
rect 9732 20828 10416 20856
rect 9732 20816 9738 20828
rect 10410 20816 10416 20828
rect 10468 20816 10474 20868
rect 10594 20856 10600 20868
rect 10555 20828 10600 20856
rect 10594 20816 10600 20828
rect 10652 20816 10658 20868
rect 15197 20859 15255 20865
rect 15197 20825 15209 20859
rect 15243 20856 15255 20859
rect 15243 20828 15884 20856
rect 15243 20825 15255 20828
rect 15197 20819 15255 20825
rect 4522 20788 4528 20800
rect 3191 20760 4384 20788
rect 4483 20760 4528 20788
rect 3191 20757 3203 20760
rect 3145 20751 3203 20757
rect 4522 20748 4528 20760
rect 4580 20748 4586 20800
rect 6270 20748 6276 20800
rect 6328 20788 6334 20800
rect 6730 20788 6736 20800
rect 6328 20760 6736 20788
rect 6328 20748 6334 20760
rect 6730 20748 6736 20760
rect 6788 20748 6794 20800
rect 8662 20748 8668 20800
rect 8720 20788 8726 20800
rect 9646 20788 9674 20816
rect 14826 20788 14832 20800
rect 8720 20760 9674 20788
rect 14787 20760 14832 20788
rect 8720 20748 8726 20760
rect 14826 20748 14832 20760
rect 14884 20748 14890 20800
rect 15286 20748 15292 20800
rect 15344 20788 15350 20800
rect 15856 20788 15884 20828
rect 16206 20816 16212 20868
rect 16264 20856 16270 20868
rect 16393 20859 16451 20865
rect 16393 20856 16405 20859
rect 16264 20828 16405 20856
rect 16264 20816 16270 20828
rect 16393 20825 16405 20828
rect 16439 20825 16451 20859
rect 16393 20819 16451 20825
rect 16482 20816 16488 20868
rect 16540 20856 16546 20868
rect 17402 20856 17408 20868
rect 16540 20828 17408 20856
rect 16540 20816 16546 20828
rect 17402 20816 17408 20828
rect 17460 20856 17466 20868
rect 17788 20856 17816 20955
rect 18322 20952 18328 21004
rect 18380 20952 18386 21004
rect 19334 20952 19340 21004
rect 19392 20992 19398 21004
rect 19978 20992 19984 21004
rect 19392 20964 19984 20992
rect 19392 20952 19398 20964
rect 19978 20952 19984 20964
rect 20036 20952 20042 21004
rect 20438 20952 20444 21004
rect 20496 20992 20502 21004
rect 21085 20995 21143 21001
rect 21085 20992 21097 20995
rect 20496 20964 21097 20992
rect 20496 20952 20502 20964
rect 21085 20961 21097 20964
rect 21131 20961 21143 20995
rect 21085 20955 21143 20961
rect 18138 20884 18144 20936
rect 18196 20924 18202 20936
rect 18340 20924 18368 20952
rect 18417 20927 18475 20933
rect 18417 20924 18429 20927
rect 18196 20896 18429 20924
rect 18196 20884 18202 20896
rect 18417 20893 18429 20896
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 18601 20927 18659 20933
rect 18601 20893 18613 20927
rect 18647 20924 18659 20927
rect 18966 20924 18972 20936
rect 18647 20896 18972 20924
rect 18647 20893 18659 20896
rect 18601 20887 18659 20893
rect 18966 20884 18972 20896
rect 19024 20924 19030 20936
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 19024 20896 19441 20924
rect 19024 20884 19030 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19794 20924 19800 20936
rect 19755 20896 19800 20924
rect 19521 20887 19579 20893
rect 17460 20828 17816 20856
rect 19536 20856 19564 20887
rect 19794 20884 19800 20896
rect 19852 20884 19858 20936
rect 20993 20927 21051 20933
rect 20993 20893 21005 20927
rect 21039 20924 21051 20927
rect 21358 20924 21364 20936
rect 21039 20896 21364 20924
rect 21039 20893 21051 20896
rect 20993 20887 21051 20893
rect 21358 20884 21364 20896
rect 21416 20884 21422 20936
rect 21913 20927 21971 20933
rect 21913 20893 21925 20927
rect 21959 20924 21971 20927
rect 22002 20924 22008 20936
rect 21959 20896 22008 20924
rect 21959 20893 21971 20896
rect 21913 20887 21971 20893
rect 22002 20884 22008 20896
rect 22060 20884 22066 20936
rect 22097 20927 22155 20933
rect 22097 20893 22109 20927
rect 22143 20924 22155 20927
rect 22370 20924 22376 20936
rect 22143 20896 22376 20924
rect 22143 20893 22155 20896
rect 22097 20887 22155 20893
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 20162 20856 20168 20868
rect 19536 20828 20168 20856
rect 17460 20816 17466 20828
rect 20162 20816 20168 20828
rect 20220 20816 20226 20868
rect 16574 20788 16580 20800
rect 15344 20760 15389 20788
rect 15856 20760 16580 20788
rect 15344 20748 15350 20760
rect 16574 20748 16580 20760
rect 16632 20748 16638 20800
rect 16758 20748 16764 20800
rect 16816 20788 16822 20800
rect 16942 20788 16948 20800
rect 16816 20760 16948 20788
rect 16816 20748 16822 20760
rect 16942 20748 16948 20760
rect 17000 20788 17006 20800
rect 17589 20791 17647 20797
rect 17589 20788 17601 20791
rect 17000 20760 17601 20788
rect 17000 20748 17006 20760
rect 17589 20757 17601 20760
rect 17635 20757 17647 20791
rect 18506 20788 18512 20800
rect 18467 20760 18512 20788
rect 17589 20751 17647 20757
rect 18506 20748 18512 20760
rect 18564 20748 18570 20800
rect 19978 20748 19984 20800
rect 20036 20788 20042 20800
rect 20533 20791 20591 20797
rect 20533 20788 20545 20791
rect 20036 20760 20545 20788
rect 20036 20748 20042 20760
rect 20533 20757 20545 20760
rect 20579 20757 20591 20791
rect 20533 20751 20591 20757
rect 20714 20748 20720 20800
rect 20772 20788 20778 20800
rect 20901 20791 20959 20797
rect 20901 20788 20913 20791
rect 20772 20760 20913 20788
rect 20772 20748 20778 20760
rect 20901 20757 20913 20760
rect 20947 20757 20959 20791
rect 20901 20751 20959 20757
rect 1104 20698 30820 20720
rect 1104 20646 10880 20698
rect 10932 20646 10944 20698
rect 10996 20646 11008 20698
rect 11060 20646 11072 20698
rect 11124 20646 11136 20698
rect 11188 20646 20811 20698
rect 20863 20646 20875 20698
rect 20927 20646 20939 20698
rect 20991 20646 21003 20698
rect 21055 20646 21067 20698
rect 21119 20646 30820 20698
rect 1104 20624 30820 20646
rect 2130 20544 2136 20596
rect 2188 20584 2194 20596
rect 2225 20587 2283 20593
rect 2225 20584 2237 20587
rect 2188 20556 2237 20584
rect 2188 20544 2194 20556
rect 2225 20553 2237 20556
rect 2271 20553 2283 20587
rect 5166 20584 5172 20596
rect 5127 20556 5172 20584
rect 2225 20547 2283 20553
rect 5166 20544 5172 20556
rect 5224 20544 5230 20596
rect 8018 20584 8024 20596
rect 7979 20556 8024 20584
rect 8018 20544 8024 20556
rect 8076 20544 8082 20596
rect 8386 20544 8392 20596
rect 8444 20584 8450 20596
rect 9306 20584 9312 20596
rect 8444 20556 9312 20584
rect 8444 20544 8450 20556
rect 9306 20544 9312 20556
rect 9364 20544 9370 20596
rect 15286 20544 15292 20596
rect 15344 20584 15350 20596
rect 15381 20587 15439 20593
rect 15381 20584 15393 20587
rect 15344 20556 15393 20584
rect 15344 20544 15350 20556
rect 15381 20553 15393 20556
rect 15427 20553 15439 20587
rect 15381 20547 15439 20553
rect 16853 20587 16911 20593
rect 16853 20553 16865 20587
rect 16899 20584 16911 20587
rect 17218 20584 17224 20596
rect 16899 20556 17224 20584
rect 16899 20553 16911 20556
rect 16853 20547 16911 20553
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 18506 20544 18512 20596
rect 18564 20584 18570 20596
rect 19153 20587 19211 20593
rect 19153 20584 19165 20587
rect 18564 20556 19165 20584
rect 18564 20544 18570 20556
rect 19153 20553 19165 20556
rect 19199 20553 19211 20587
rect 19153 20547 19211 20553
rect 19242 20544 19248 20596
rect 19300 20584 19306 20596
rect 20254 20584 20260 20596
rect 19300 20556 19345 20584
rect 20215 20556 20260 20584
rect 19300 20544 19306 20556
rect 20254 20544 20260 20556
rect 20312 20544 20318 20596
rect 20622 20544 20628 20596
rect 20680 20584 20686 20596
rect 20717 20587 20775 20593
rect 20717 20584 20729 20587
rect 20680 20556 20729 20584
rect 20680 20544 20686 20556
rect 20717 20553 20729 20556
rect 20763 20553 20775 20587
rect 22278 20584 22284 20596
rect 22239 20556 22284 20584
rect 20717 20547 20775 20553
rect 22278 20544 22284 20556
rect 22336 20544 22342 20596
rect 1854 20516 1860 20528
rect 1780 20488 1860 20516
rect 1394 20408 1400 20460
rect 1452 20448 1458 20460
rect 1489 20451 1547 20457
rect 1489 20448 1501 20451
rect 1452 20420 1501 20448
rect 1452 20408 1458 20420
rect 1489 20417 1501 20420
rect 1535 20417 1547 20451
rect 1670 20448 1676 20460
rect 1631 20420 1676 20448
rect 1489 20411 1547 20417
rect 1670 20408 1676 20420
rect 1728 20408 1734 20460
rect 1780 20457 1808 20488
rect 1854 20476 1860 20488
rect 1912 20476 1918 20528
rect 3050 20516 3056 20528
rect 2056 20488 3056 20516
rect 2056 20457 2084 20488
rect 3050 20476 3056 20488
rect 3108 20476 3114 20528
rect 4056 20519 4114 20525
rect 4056 20485 4068 20519
rect 4102 20516 4114 20519
rect 4522 20516 4528 20528
rect 4102 20488 4528 20516
rect 4102 20485 4114 20488
rect 4056 20479 4114 20485
rect 4522 20476 4528 20488
rect 4580 20476 4586 20528
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20417 1823 20451
rect 1765 20411 1823 20417
rect 2041 20451 2099 20457
rect 2041 20417 2053 20451
rect 2087 20417 2099 20451
rect 2041 20411 2099 20417
rect 2869 20451 2927 20457
rect 2869 20417 2881 20451
rect 2915 20448 2927 20451
rect 2958 20448 2964 20460
rect 2915 20420 2964 20448
rect 2915 20417 2927 20420
rect 2869 20411 2927 20417
rect 2958 20408 2964 20420
rect 3016 20408 3022 20460
rect 5184 20448 5212 20544
rect 7006 20476 7012 20528
rect 7064 20516 7070 20528
rect 8481 20519 8539 20525
rect 8481 20516 8493 20519
rect 7064 20488 8493 20516
rect 7064 20476 7070 20488
rect 8481 20485 8493 20488
rect 8527 20485 8539 20519
rect 9324 20516 9352 20544
rect 9677 20519 9735 20525
rect 9324 20488 9628 20516
rect 8481 20479 8539 20485
rect 6914 20457 6920 20460
rect 5629 20451 5687 20457
rect 5629 20448 5641 20451
rect 5184 20420 5641 20448
rect 5629 20417 5641 20420
rect 5675 20417 5687 20451
rect 5629 20411 5687 20417
rect 6908 20411 6920 20457
rect 6972 20448 6978 20460
rect 6972 20420 7008 20448
rect 6914 20408 6920 20411
rect 6972 20408 6978 20420
rect 8294 20408 8300 20460
rect 8352 20448 8358 20460
rect 8665 20451 8723 20457
rect 8665 20448 8677 20451
rect 8352 20420 8677 20448
rect 8352 20408 8358 20420
rect 8665 20417 8677 20420
rect 8711 20417 8723 20451
rect 8665 20411 8723 20417
rect 8849 20451 8907 20457
rect 8849 20417 8861 20451
rect 8895 20448 8907 20451
rect 8938 20448 8944 20460
rect 8895 20420 8944 20448
rect 8895 20417 8907 20420
rect 8849 20411 8907 20417
rect 1857 20383 1915 20389
rect 1857 20349 1869 20383
rect 1903 20380 1915 20383
rect 1946 20380 1952 20392
rect 1903 20352 1952 20380
rect 1903 20349 1915 20352
rect 1857 20343 1915 20349
rect 1946 20340 1952 20352
rect 2004 20340 2010 20392
rect 3786 20380 3792 20392
rect 3747 20352 3792 20380
rect 3786 20340 3792 20352
rect 3844 20340 3850 20392
rect 6638 20380 6644 20392
rect 6599 20352 6644 20380
rect 6638 20340 6644 20352
rect 6696 20340 6702 20392
rect 8680 20380 8708 20411
rect 8938 20408 8944 20420
rect 8996 20408 9002 20460
rect 9493 20451 9551 20457
rect 9493 20417 9505 20451
rect 9539 20417 9551 20451
rect 9600 20448 9628 20488
rect 9677 20485 9689 20519
rect 9723 20516 9735 20519
rect 10226 20516 10232 20528
rect 9723 20488 10232 20516
rect 9723 20485 9735 20488
rect 9677 20479 9735 20485
rect 10226 20476 10232 20488
rect 10284 20516 10290 20528
rect 10594 20516 10600 20528
rect 10284 20488 10600 20516
rect 10284 20476 10290 20488
rect 10594 20476 10600 20488
rect 10652 20476 10658 20528
rect 10686 20476 10692 20528
rect 10744 20516 10750 20528
rect 11701 20519 11759 20525
rect 11701 20516 11713 20519
rect 10744 20488 11713 20516
rect 10744 20476 10750 20488
rect 11701 20485 11713 20488
rect 11747 20485 11759 20519
rect 11701 20479 11759 20485
rect 12158 20476 12164 20528
rect 12216 20516 12222 20528
rect 12253 20519 12311 20525
rect 12253 20516 12265 20519
rect 12216 20488 12265 20516
rect 12216 20476 12222 20488
rect 12253 20485 12265 20488
rect 12299 20485 12311 20519
rect 14921 20519 14979 20525
rect 14921 20516 14933 20519
rect 12253 20479 12311 20485
rect 12360 20488 14933 20516
rect 10137 20451 10195 20457
rect 10137 20448 10149 20451
rect 9600 20420 10149 20448
rect 9493 20411 9551 20417
rect 10137 20417 10149 20420
rect 10183 20417 10195 20451
rect 10137 20411 10195 20417
rect 9508 20380 9536 20411
rect 8680 20352 9536 20380
rect 10229 20383 10287 20389
rect 10229 20349 10241 20383
rect 10275 20380 10287 20383
rect 10318 20380 10324 20392
rect 10275 20352 10324 20380
rect 10275 20349 10287 20352
rect 10229 20343 10287 20349
rect 10318 20340 10324 20352
rect 10376 20340 10382 20392
rect 7650 20272 7656 20324
rect 7708 20312 7714 20324
rect 7926 20312 7932 20324
rect 7708 20284 7932 20312
rect 7708 20272 7714 20284
rect 7926 20272 7932 20284
rect 7984 20312 7990 20324
rect 12360 20312 12388 20488
rect 14921 20485 14933 20488
rect 14967 20485 14979 20519
rect 14921 20479 14979 20485
rect 17313 20519 17371 20525
rect 17313 20485 17325 20519
rect 17359 20516 17371 20519
rect 19058 20516 19064 20528
rect 17359 20488 19064 20516
rect 17359 20485 17371 20488
rect 17313 20479 17371 20485
rect 19058 20476 19064 20488
rect 19116 20516 19122 20528
rect 19886 20516 19892 20528
rect 19116 20488 19892 20516
rect 19116 20476 19122 20488
rect 19886 20476 19892 20488
rect 19944 20476 19950 20528
rect 22002 20476 22008 20528
rect 22060 20516 22066 20528
rect 22189 20519 22247 20525
rect 22189 20516 22201 20519
rect 22060 20488 22201 20516
rect 22060 20476 22066 20488
rect 22189 20485 22201 20488
rect 22235 20516 22247 20519
rect 22370 20516 22376 20528
rect 22235 20488 22376 20516
rect 22235 20485 22247 20488
rect 22189 20479 22247 20485
rect 22370 20476 22376 20488
rect 22428 20476 22434 20528
rect 12434 20408 12440 20460
rect 12492 20448 12498 20460
rect 13078 20448 13084 20460
rect 12492 20420 13084 20448
rect 12492 20408 12498 20420
rect 13078 20408 13084 20420
rect 13136 20408 13142 20460
rect 13446 20448 13452 20460
rect 13407 20420 13452 20448
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 13909 20451 13967 20457
rect 13909 20417 13921 20451
rect 13955 20448 13967 20451
rect 15013 20451 15071 20457
rect 13955 20420 14596 20448
rect 13955 20417 13967 20420
rect 13909 20411 13967 20417
rect 14568 20324 14596 20420
rect 15013 20417 15025 20451
rect 15059 20448 15071 20451
rect 15841 20451 15899 20457
rect 15841 20448 15853 20451
rect 15059 20420 15853 20448
rect 15059 20417 15071 20420
rect 15013 20411 15071 20417
rect 15841 20417 15853 20420
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 16117 20451 16175 20457
rect 16117 20417 16129 20451
rect 16163 20448 16175 20451
rect 16206 20448 16212 20460
rect 16163 20420 16212 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 16206 20408 16212 20420
rect 16264 20408 16270 20460
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 17221 20451 17279 20457
rect 17221 20448 17233 20451
rect 16816 20420 17233 20448
rect 16816 20408 16822 20420
rect 17221 20417 17233 20420
rect 17267 20448 17279 20451
rect 17267 20420 17724 20448
rect 17267 20417 17279 20420
rect 17221 20411 17279 20417
rect 14829 20383 14887 20389
rect 14829 20349 14841 20383
rect 14875 20380 14887 20383
rect 14918 20380 14924 20392
rect 14875 20352 14924 20380
rect 14875 20349 14887 20352
rect 14829 20343 14887 20349
rect 14918 20340 14924 20352
rect 14976 20340 14982 20392
rect 17402 20380 17408 20392
rect 17363 20352 17408 20380
rect 17402 20340 17408 20352
rect 17460 20340 17466 20392
rect 17696 20380 17724 20420
rect 17770 20408 17776 20460
rect 17828 20448 17834 20460
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 17828 20420 18061 20448
rect 17828 20408 17834 20420
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 18233 20451 18291 20457
rect 18233 20417 18245 20451
rect 18279 20417 18291 20451
rect 18233 20411 18291 20417
rect 20625 20451 20683 20457
rect 20625 20417 20637 20451
rect 20671 20448 20683 20451
rect 20714 20448 20720 20460
rect 20671 20420 20720 20448
rect 20671 20417 20683 20420
rect 20625 20411 20683 20417
rect 18248 20380 18276 20411
rect 20714 20408 20720 20420
rect 20772 20408 20778 20460
rect 19058 20380 19064 20392
rect 17696 20352 18276 20380
rect 19019 20352 19064 20380
rect 19058 20340 19064 20352
rect 19116 20340 19122 20392
rect 20438 20340 20444 20392
rect 20496 20380 20502 20392
rect 20809 20383 20867 20389
rect 20809 20380 20821 20383
rect 20496 20352 20821 20380
rect 20496 20340 20502 20352
rect 20809 20349 20821 20352
rect 20855 20349 20867 20383
rect 20809 20343 20867 20349
rect 21910 20340 21916 20392
rect 21968 20380 21974 20392
rect 22373 20383 22431 20389
rect 22373 20380 22385 20383
rect 21968 20352 22385 20380
rect 21968 20340 21974 20352
rect 22373 20349 22385 20352
rect 22419 20349 22431 20383
rect 22373 20343 22431 20349
rect 7984 20284 12388 20312
rect 13541 20315 13599 20321
rect 7984 20272 7990 20284
rect 13541 20281 13553 20315
rect 13587 20312 13599 20315
rect 14090 20312 14096 20324
rect 13587 20284 14096 20312
rect 13587 20281 13599 20284
rect 13541 20275 13599 20281
rect 14090 20272 14096 20284
rect 14148 20272 14154 20324
rect 14550 20272 14556 20324
rect 14608 20312 14614 20324
rect 21821 20315 21879 20321
rect 21821 20312 21833 20315
rect 14608 20284 21833 20312
rect 14608 20272 14614 20284
rect 21821 20281 21833 20284
rect 21867 20281 21879 20315
rect 21821 20275 21879 20281
rect 1854 20204 1860 20256
rect 1912 20244 1918 20256
rect 2685 20247 2743 20253
rect 2685 20244 2697 20247
rect 1912 20216 2697 20244
rect 1912 20204 1918 20216
rect 2685 20213 2697 20216
rect 2731 20213 2743 20247
rect 2685 20207 2743 20213
rect 5721 20247 5779 20253
rect 5721 20213 5733 20247
rect 5767 20244 5779 20247
rect 6546 20244 6552 20256
rect 5767 20216 6552 20244
rect 5767 20213 5779 20216
rect 5721 20207 5779 20213
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 8938 20204 8944 20256
rect 8996 20244 9002 20256
rect 9950 20244 9956 20256
rect 8996 20216 9956 20244
rect 8996 20204 9002 20216
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 11606 20244 11612 20256
rect 11567 20216 11612 20244
rect 11606 20204 11612 20216
rect 11664 20204 11670 20256
rect 13262 20204 13268 20256
rect 13320 20244 13326 20256
rect 13633 20247 13691 20253
rect 13633 20244 13645 20247
rect 13320 20216 13645 20244
rect 13320 20204 13326 20216
rect 13633 20213 13645 20216
rect 13679 20213 13691 20247
rect 13633 20207 13691 20213
rect 13771 20247 13829 20253
rect 13771 20213 13783 20247
rect 13817 20244 13829 20247
rect 14458 20244 14464 20256
rect 13817 20216 14464 20244
rect 13817 20213 13829 20216
rect 13771 20207 13829 20213
rect 14458 20204 14464 20216
rect 14516 20204 14522 20256
rect 16942 20204 16948 20256
rect 17000 20244 17006 20256
rect 18417 20247 18475 20253
rect 18417 20244 18429 20247
rect 17000 20216 18429 20244
rect 17000 20204 17006 20216
rect 18417 20213 18429 20216
rect 18463 20213 18475 20247
rect 18417 20207 18475 20213
rect 19426 20204 19432 20256
rect 19484 20244 19490 20256
rect 19613 20247 19671 20253
rect 19613 20244 19625 20247
rect 19484 20216 19625 20244
rect 19484 20204 19490 20216
rect 19613 20213 19625 20216
rect 19659 20213 19671 20247
rect 19613 20207 19671 20213
rect 1104 20154 30820 20176
rect 1104 20102 5915 20154
rect 5967 20102 5979 20154
rect 6031 20102 6043 20154
rect 6095 20102 6107 20154
rect 6159 20102 6171 20154
rect 6223 20102 15846 20154
rect 15898 20102 15910 20154
rect 15962 20102 15974 20154
rect 16026 20102 16038 20154
rect 16090 20102 16102 20154
rect 16154 20102 25776 20154
rect 25828 20102 25840 20154
rect 25892 20102 25904 20154
rect 25956 20102 25968 20154
rect 26020 20102 26032 20154
rect 26084 20102 30820 20154
rect 1104 20080 30820 20102
rect 6914 20000 6920 20052
rect 6972 20040 6978 20052
rect 7101 20043 7159 20049
rect 7101 20040 7113 20043
rect 6972 20012 7113 20040
rect 6972 20000 6978 20012
rect 7101 20009 7113 20012
rect 7147 20009 7159 20043
rect 7101 20003 7159 20009
rect 7190 20000 7196 20052
rect 7248 20040 7254 20052
rect 7561 20043 7619 20049
rect 7561 20040 7573 20043
rect 7248 20012 7573 20040
rect 7248 20000 7254 20012
rect 7561 20009 7573 20012
rect 7607 20009 7619 20043
rect 7561 20003 7619 20009
rect 7929 20043 7987 20049
rect 7929 20009 7941 20043
rect 7975 20009 7987 20043
rect 7929 20003 7987 20009
rect 3234 19972 3240 19984
rect 3147 19944 3240 19972
rect 3234 19932 3240 19944
rect 3292 19972 3298 19984
rect 7006 19972 7012 19984
rect 3292 19944 5396 19972
rect 3292 19932 3298 19944
rect 4430 19904 4436 19916
rect 4391 19876 4436 19904
rect 4430 19864 4436 19876
rect 4488 19864 4494 19916
rect 4540 19876 5304 19904
rect 1857 19839 1915 19845
rect 1857 19805 1869 19839
rect 1903 19836 1915 19839
rect 2866 19836 2872 19848
rect 1903 19808 2872 19836
rect 1903 19805 1915 19808
rect 1857 19799 1915 19805
rect 2866 19796 2872 19808
rect 2924 19796 2930 19848
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19805 4123 19839
rect 4246 19836 4252 19848
rect 4207 19808 4252 19836
rect 4065 19799 4123 19805
rect 2124 19771 2182 19777
rect 2124 19737 2136 19771
rect 2170 19768 2182 19771
rect 2222 19768 2228 19780
rect 2170 19740 2228 19768
rect 2170 19737 2182 19740
rect 2124 19731 2182 19737
rect 2222 19728 2228 19740
rect 2280 19728 2286 19780
rect 4080 19768 4108 19799
rect 4246 19796 4252 19808
rect 4304 19796 4310 19848
rect 4338 19796 4344 19848
rect 4396 19836 4402 19848
rect 4540 19836 4568 19876
rect 4396 19808 4568 19836
rect 4617 19839 4675 19845
rect 4396 19796 4402 19808
rect 4617 19805 4629 19839
rect 4663 19836 4675 19839
rect 5166 19836 5172 19848
rect 4663 19808 5172 19836
rect 4663 19805 4675 19808
rect 4617 19799 4675 19805
rect 5166 19796 5172 19808
rect 5224 19796 5230 19848
rect 4706 19768 4712 19780
rect 4080 19740 4712 19768
rect 4706 19728 4712 19740
rect 4764 19728 4770 19780
rect 5276 19768 5304 19876
rect 5368 19845 5396 19944
rect 6656 19944 7012 19972
rect 5810 19864 5816 19916
rect 5868 19904 5874 19916
rect 6656 19913 6684 19944
rect 7006 19932 7012 19944
rect 7064 19932 7070 19984
rect 7944 19972 7972 20003
rect 9122 20000 9128 20052
rect 9180 20040 9186 20052
rect 9401 20043 9459 20049
rect 9401 20040 9413 20043
rect 9180 20012 9413 20040
rect 9180 20000 9186 20012
rect 9401 20009 9413 20012
rect 9447 20009 9459 20043
rect 9401 20003 9459 20009
rect 9766 20000 9772 20052
rect 9824 20040 9830 20052
rect 9824 20012 10548 20040
rect 9824 20000 9830 20012
rect 8202 19972 8208 19984
rect 7944 19944 8208 19972
rect 8202 19932 8208 19944
rect 8260 19972 8266 19984
rect 9674 19972 9680 19984
rect 8260 19944 9680 19972
rect 8260 19932 8266 19944
rect 9674 19932 9680 19944
rect 9732 19932 9738 19984
rect 9861 19975 9919 19981
rect 9861 19941 9873 19975
rect 9907 19972 9919 19975
rect 10413 19975 10471 19981
rect 10413 19972 10425 19975
rect 9907 19944 10425 19972
rect 9907 19941 9919 19944
rect 9861 19935 9919 19941
rect 10413 19941 10425 19944
rect 10459 19941 10471 19975
rect 10413 19935 10471 19941
rect 6641 19907 6699 19913
rect 5868 19876 6592 19904
rect 5868 19864 5874 19876
rect 5353 19839 5411 19845
rect 5353 19805 5365 19839
rect 5399 19805 5411 19839
rect 6362 19836 6368 19848
rect 6323 19808 6368 19836
rect 5353 19799 5411 19805
rect 6362 19796 6368 19808
rect 6420 19796 6426 19848
rect 6564 19845 6592 19876
rect 6641 19873 6653 19907
rect 6687 19873 6699 19907
rect 6641 19867 6699 19873
rect 6733 19907 6791 19913
rect 6733 19873 6745 19907
rect 6779 19904 6791 19907
rect 6822 19904 6828 19916
rect 6779 19876 6828 19904
rect 6779 19873 6791 19876
rect 6733 19867 6791 19873
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 7190 19864 7196 19916
rect 7248 19904 7254 19916
rect 10318 19904 10324 19916
rect 7248 19876 10324 19904
rect 7248 19864 7254 19876
rect 10318 19864 10324 19876
rect 10376 19864 10382 19916
rect 6549 19839 6607 19845
rect 6549 19805 6561 19839
rect 6595 19805 6607 19839
rect 6549 19799 6607 19805
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19836 6975 19839
rect 7926 19836 7932 19848
rect 6963 19808 7932 19836
rect 6963 19805 6975 19808
rect 6917 19799 6975 19805
rect 6564 19768 6592 19799
rect 7926 19796 7932 19808
rect 7984 19796 7990 19848
rect 8018 19796 8024 19848
rect 8076 19836 8082 19848
rect 8076 19808 8121 19836
rect 8076 19796 8082 19808
rect 8386 19796 8392 19848
rect 8444 19836 8450 19848
rect 8754 19836 8760 19848
rect 8444 19808 8760 19836
rect 8444 19796 8450 19808
rect 8754 19796 8760 19808
rect 8812 19796 8818 19848
rect 9306 19796 9312 19848
rect 9364 19836 9370 19848
rect 9585 19839 9643 19845
rect 9585 19836 9597 19839
rect 9364 19808 9597 19836
rect 9364 19796 9370 19808
rect 9585 19805 9597 19808
rect 9631 19805 9643 19839
rect 9585 19799 9643 19805
rect 9674 19796 9680 19848
rect 9732 19836 9738 19848
rect 9953 19839 10011 19845
rect 9732 19808 9825 19836
rect 9732 19796 9738 19808
rect 9953 19805 9965 19839
rect 9999 19836 10011 19839
rect 10520 19836 10548 20012
rect 12526 20000 12532 20052
rect 12584 20040 12590 20052
rect 12897 20043 12955 20049
rect 12897 20040 12909 20043
rect 12584 20012 12909 20040
rect 12584 20000 12590 20012
rect 12897 20009 12909 20012
rect 12943 20040 12955 20043
rect 13354 20040 13360 20052
rect 12943 20012 13360 20040
rect 12943 20009 12955 20012
rect 12897 20003 12955 20009
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 14384 20012 15976 20040
rect 11422 19972 11428 19984
rect 10612 19944 11428 19972
rect 10612 19913 10640 19944
rect 11422 19932 11428 19944
rect 11480 19932 11486 19984
rect 14384 19981 14412 20012
rect 14369 19975 14427 19981
rect 14369 19941 14381 19975
rect 14415 19941 14427 19975
rect 14369 19935 14427 19941
rect 14458 19932 14464 19984
rect 14516 19972 14522 19984
rect 15948 19972 15976 20012
rect 16206 20000 16212 20052
rect 16264 20040 16270 20052
rect 16669 20043 16727 20049
rect 16669 20040 16681 20043
rect 16264 20012 16681 20040
rect 16264 20000 16270 20012
rect 16669 20009 16681 20012
rect 16715 20009 16727 20043
rect 16669 20003 16727 20009
rect 17218 20000 17224 20052
rect 17276 20040 17282 20052
rect 17862 20040 17868 20052
rect 17276 20012 17868 20040
rect 17276 20000 17282 20012
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 20162 20000 20168 20052
rect 20220 20040 20226 20052
rect 20441 20043 20499 20049
rect 20441 20040 20453 20043
rect 20220 20012 20453 20040
rect 20220 20000 20226 20012
rect 20441 20009 20453 20012
rect 20487 20009 20499 20043
rect 20441 20003 20499 20009
rect 19337 19975 19395 19981
rect 19337 19972 19349 19975
rect 14516 19944 14561 19972
rect 15948 19944 19349 19972
rect 14516 19932 14522 19944
rect 19337 19941 19349 19944
rect 19383 19941 19395 19975
rect 19337 19935 19395 19941
rect 10597 19907 10655 19913
rect 10597 19873 10609 19907
rect 10643 19873 10655 19907
rect 11514 19904 11520 19916
rect 11475 19876 11520 19904
rect 10597 19867 10655 19873
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 14734 19904 14740 19916
rect 14292 19876 14740 19904
rect 10689 19839 10747 19845
rect 10689 19836 10701 19839
rect 9999 19808 10548 19836
rect 10612 19808 10701 19836
rect 9999 19805 10011 19808
rect 9953 19799 10011 19805
rect 8938 19768 8944 19780
rect 5276 19740 6408 19768
rect 6564 19740 8944 19768
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 3418 19700 3424 19712
rect 1728 19672 3424 19700
rect 1728 19660 1734 19672
rect 3418 19660 3424 19672
rect 3476 19660 3482 19712
rect 4798 19700 4804 19712
rect 4759 19672 4804 19700
rect 4798 19660 4804 19672
rect 4856 19660 4862 19712
rect 5445 19703 5503 19709
rect 5445 19669 5457 19703
rect 5491 19700 5503 19703
rect 6270 19700 6276 19712
rect 5491 19672 6276 19700
rect 5491 19669 5503 19672
rect 5445 19663 5503 19669
rect 6270 19660 6276 19672
rect 6328 19660 6334 19712
rect 6380 19700 6408 19740
rect 8938 19728 8944 19740
rect 8996 19728 9002 19780
rect 9692 19768 9720 19796
rect 10612 19780 10640 19808
rect 10689 19805 10701 19808
rect 10735 19836 10747 19839
rect 10965 19839 11023 19845
rect 10965 19836 10977 19839
rect 10735 19808 10977 19836
rect 10735 19805 10747 19808
rect 10689 19799 10747 19805
rect 10965 19805 10977 19808
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19836 11115 19839
rect 13538 19836 13544 19848
rect 11103 19808 12434 19836
rect 13499 19808 13544 19836
rect 11103 19805 11115 19808
rect 11057 19799 11115 19805
rect 9858 19768 9864 19780
rect 9692 19740 9864 19768
rect 9858 19728 9864 19740
rect 9916 19728 9922 19780
rect 10042 19728 10048 19780
rect 10100 19768 10106 19780
rect 10594 19768 10600 19780
rect 10100 19740 10600 19768
rect 10100 19728 10106 19740
rect 10594 19728 10600 19740
rect 10652 19728 10658 19780
rect 11784 19771 11842 19777
rect 11784 19737 11796 19771
rect 11830 19768 11842 19771
rect 12250 19768 12256 19780
rect 11830 19740 12256 19768
rect 11830 19737 11842 19740
rect 11784 19731 11842 19737
rect 12250 19728 12256 19740
rect 12308 19728 12314 19780
rect 12406 19768 12434 19808
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 14090 19836 14096 19848
rect 14051 19808 14096 19836
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14292 19845 14320 19876
rect 14734 19864 14740 19876
rect 14792 19864 14798 19916
rect 15746 19904 15752 19916
rect 15707 19876 15752 19904
rect 15746 19864 15752 19876
rect 15804 19864 15810 19916
rect 16022 19904 16028 19916
rect 15983 19876 16028 19904
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 16666 19864 16672 19916
rect 16724 19904 16730 19916
rect 17586 19904 17592 19916
rect 16724 19876 17592 19904
rect 16724 19864 16730 19876
rect 17586 19864 17592 19876
rect 17644 19904 17650 19916
rect 17957 19907 18015 19913
rect 17957 19904 17969 19907
rect 17644 19876 17969 19904
rect 17644 19864 17650 19876
rect 17957 19873 17969 19876
rect 18003 19904 18015 19907
rect 19058 19904 19064 19916
rect 18003 19876 19064 19904
rect 18003 19873 18015 19876
rect 17957 19867 18015 19873
rect 19058 19864 19064 19876
rect 19116 19864 19122 19916
rect 20180 19904 20208 20000
rect 21634 19932 21640 19984
rect 21692 19972 21698 19984
rect 21729 19975 21787 19981
rect 21729 19972 21741 19975
rect 21692 19944 21741 19972
rect 21692 19932 21698 19944
rect 21729 19941 21741 19944
rect 21775 19941 21787 19975
rect 21729 19935 21787 19941
rect 19444 19876 20208 19904
rect 14277 19839 14335 19845
rect 14277 19805 14289 19839
rect 14323 19805 14335 19839
rect 14550 19836 14556 19848
rect 14511 19808 14556 19836
rect 14277 19799 14335 19805
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 13446 19768 13452 19780
rect 12406 19740 13452 19768
rect 13446 19728 13452 19740
rect 13504 19728 13510 19780
rect 14752 19768 14780 19864
rect 15838 19836 15844 19848
rect 15799 19808 15844 19836
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 15930 19796 15936 19848
rect 15988 19836 15994 19848
rect 16853 19839 16911 19845
rect 15988 19808 16033 19836
rect 15988 19796 15994 19808
rect 16853 19805 16865 19839
rect 16899 19836 16911 19839
rect 16942 19836 16948 19848
rect 16899 19808 16948 19836
rect 16899 19805 16911 19808
rect 16853 19799 16911 19805
rect 16942 19796 16948 19808
rect 17000 19796 17006 19848
rect 17678 19836 17684 19848
rect 17639 19808 17684 19836
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 19444 19845 19472 19876
rect 19429 19839 19487 19845
rect 19429 19805 19441 19839
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 19794 19796 19800 19848
rect 19852 19836 19858 19848
rect 20165 19839 20223 19845
rect 20165 19836 20177 19839
rect 19852 19808 20177 19836
rect 19852 19796 19858 19808
rect 20165 19805 20177 19808
rect 20211 19805 20223 19839
rect 20165 19799 20223 19805
rect 20254 19796 20260 19848
rect 20312 19836 20318 19848
rect 20533 19839 20591 19845
rect 20312 19808 20357 19836
rect 20312 19796 20318 19808
rect 20533 19805 20545 19839
rect 20579 19836 20591 19839
rect 20622 19836 20628 19848
rect 20579 19808 20628 19836
rect 20579 19805 20591 19808
rect 20533 19799 20591 19805
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 21910 19836 21916 19848
rect 21871 19808 21916 19836
rect 21910 19796 21916 19808
rect 21968 19796 21974 19848
rect 22097 19839 22155 19845
rect 22097 19805 22109 19839
rect 22143 19836 22155 19839
rect 22462 19836 22468 19848
rect 22143 19808 22468 19836
rect 22143 19805 22155 19808
rect 22097 19799 22155 19805
rect 22462 19796 22468 19808
rect 22520 19836 22526 19848
rect 23014 19836 23020 19848
rect 22520 19808 23020 19836
rect 22520 19796 22526 19808
rect 23014 19796 23020 19808
rect 23072 19796 23078 19848
rect 18598 19768 18604 19780
rect 14752 19740 15700 19768
rect 7190 19700 7196 19712
rect 6380 19672 7196 19700
rect 7190 19660 7196 19672
rect 7248 19660 7254 19712
rect 8018 19660 8024 19712
rect 8076 19700 8082 19712
rect 11330 19700 11336 19712
rect 8076 19672 11336 19700
rect 8076 19660 8082 19672
rect 11330 19660 11336 19672
rect 11388 19660 11394 19712
rect 14734 19700 14740 19712
rect 14695 19672 14740 19700
rect 14734 19660 14740 19672
rect 14792 19660 14798 19712
rect 15286 19660 15292 19712
rect 15344 19700 15350 19712
rect 15565 19703 15623 19709
rect 15565 19700 15577 19703
rect 15344 19672 15577 19700
rect 15344 19660 15350 19672
rect 15565 19669 15577 19672
rect 15611 19669 15623 19703
rect 15672 19700 15700 19740
rect 17052 19740 18604 19768
rect 17052 19700 17080 19740
rect 18598 19728 18604 19740
rect 18656 19728 18662 19780
rect 15672 19672 17080 19700
rect 15565 19663 15623 19669
rect 17126 19660 17132 19712
rect 17184 19700 17190 19712
rect 17313 19703 17371 19709
rect 17313 19700 17325 19703
rect 17184 19672 17325 19700
rect 17184 19660 17190 19672
rect 17313 19669 17325 19672
rect 17359 19669 17371 19703
rect 17313 19663 17371 19669
rect 17586 19660 17592 19712
rect 17644 19700 17650 19712
rect 17773 19703 17831 19709
rect 17773 19700 17785 19703
rect 17644 19672 17785 19700
rect 17644 19660 17650 19672
rect 17773 19669 17785 19672
rect 17819 19669 17831 19703
rect 17773 19663 17831 19669
rect 19981 19703 20039 19709
rect 19981 19669 19993 19703
rect 20027 19700 20039 19703
rect 20254 19700 20260 19712
rect 20027 19672 20260 19700
rect 20027 19669 20039 19672
rect 19981 19663 20039 19669
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 1104 19610 30820 19632
rect 1104 19558 10880 19610
rect 10932 19558 10944 19610
rect 10996 19558 11008 19610
rect 11060 19558 11072 19610
rect 11124 19558 11136 19610
rect 11188 19558 20811 19610
rect 20863 19558 20875 19610
rect 20927 19558 20939 19610
rect 20991 19558 21003 19610
rect 21055 19558 21067 19610
rect 21119 19558 30820 19610
rect 1104 19536 30820 19558
rect 1302 19456 1308 19508
rect 1360 19496 1366 19508
rect 1360 19468 11928 19496
rect 1360 19456 1366 19468
rect 4608 19431 4666 19437
rect 2240 19400 2774 19428
rect 2240 19369 2268 19400
rect 2498 19369 2504 19372
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19360 1455 19363
rect 2225 19363 2283 19369
rect 1443 19332 2176 19360
rect 1443 19329 1455 19332
rect 1397 19323 1455 19329
rect 1581 19227 1639 19233
rect 1581 19193 1593 19227
rect 1627 19224 1639 19227
rect 1670 19224 1676 19236
rect 1627 19196 1676 19224
rect 1627 19193 1639 19196
rect 1581 19187 1639 19193
rect 1670 19184 1676 19196
rect 1728 19184 1734 19236
rect 2148 19156 2176 19332
rect 2225 19329 2237 19363
rect 2271 19329 2283 19363
rect 2225 19323 2283 19329
rect 2492 19323 2504 19369
rect 2556 19360 2562 19372
rect 2746 19360 2774 19400
rect 4608 19397 4620 19431
rect 4654 19428 4666 19431
rect 4798 19428 4804 19440
rect 4654 19400 4804 19428
rect 4654 19397 4666 19400
rect 4608 19391 4666 19397
rect 4798 19388 4804 19400
rect 4856 19388 4862 19440
rect 8386 19388 8392 19440
rect 8444 19428 8450 19440
rect 8665 19431 8723 19437
rect 8665 19428 8677 19431
rect 8444 19400 8677 19428
rect 8444 19388 8450 19400
rect 8665 19397 8677 19400
rect 8711 19397 8723 19431
rect 9306 19428 9312 19440
rect 9267 19400 9312 19428
rect 8665 19391 8723 19397
rect 9306 19388 9312 19400
rect 9364 19388 9370 19440
rect 10042 19428 10048 19440
rect 10003 19400 10048 19428
rect 10042 19388 10048 19400
rect 10100 19388 10106 19440
rect 10226 19428 10232 19440
rect 10187 19400 10232 19428
rect 10226 19388 10232 19400
rect 10284 19388 10290 19440
rect 11422 19428 11428 19440
rect 10612 19400 11428 19428
rect 2866 19360 2872 19372
rect 2556 19332 2592 19360
rect 2746 19332 2872 19360
rect 2498 19320 2504 19323
rect 2556 19320 2562 19332
rect 2866 19320 2872 19332
rect 2924 19360 2930 19372
rect 3786 19360 3792 19372
rect 2924 19332 3792 19360
rect 2924 19320 2930 19332
rect 3786 19320 3792 19332
rect 3844 19360 3850 19372
rect 4341 19363 4399 19369
rect 4341 19360 4353 19363
rect 3844 19332 4353 19360
rect 3844 19320 3850 19332
rect 4341 19329 4353 19332
rect 4387 19329 4399 19363
rect 4341 19323 4399 19329
rect 5166 19320 5172 19372
rect 5224 19360 5230 19372
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 5224 19332 6377 19360
rect 5224 19320 5230 19332
rect 5736 19233 5764 19332
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 6454 19320 6460 19372
rect 6512 19360 6518 19372
rect 8754 19360 8760 19372
rect 6512 19332 6557 19360
rect 8715 19332 8760 19360
rect 6512 19320 6518 19332
rect 8754 19320 8760 19332
rect 8812 19320 8818 19372
rect 9401 19363 9459 19369
rect 9401 19329 9413 19363
rect 9447 19360 9459 19363
rect 9447 19332 9720 19360
rect 9447 19329 9459 19332
rect 9401 19323 9459 19329
rect 9692 19292 9720 19332
rect 9766 19320 9772 19372
rect 9824 19360 9830 19372
rect 9861 19363 9919 19369
rect 9861 19360 9873 19363
rect 9824 19332 9873 19360
rect 9824 19320 9830 19332
rect 9861 19329 9873 19332
rect 9907 19329 9919 19363
rect 10612 19360 10640 19400
rect 11422 19388 11428 19400
rect 11480 19388 11486 19440
rect 11900 19437 11928 19468
rect 12894 19456 12900 19508
rect 12952 19496 12958 19508
rect 13170 19496 13176 19508
rect 12952 19468 13176 19496
rect 12952 19456 12958 19468
rect 13170 19456 13176 19468
rect 13228 19456 13234 19508
rect 13538 19456 13544 19508
rect 13596 19496 13602 19508
rect 14093 19499 14151 19505
rect 14093 19496 14105 19499
rect 13596 19468 14105 19496
rect 13596 19456 13602 19468
rect 14093 19465 14105 19468
rect 14139 19465 14151 19499
rect 15930 19496 15936 19508
rect 14093 19459 14151 19465
rect 14660 19468 15936 19496
rect 11885 19431 11943 19437
rect 11885 19397 11897 19431
rect 11931 19397 11943 19431
rect 11885 19391 11943 19397
rect 13262 19388 13268 19440
rect 13320 19428 13326 19440
rect 14660 19428 14688 19468
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 16025 19499 16083 19505
rect 16025 19465 16037 19499
rect 16071 19496 16083 19499
rect 16298 19496 16304 19508
rect 16071 19468 16304 19496
rect 16071 19465 16083 19468
rect 16025 19459 16083 19465
rect 16298 19456 16304 19468
rect 16356 19456 16362 19508
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 17586 19496 17592 19508
rect 16816 19468 17448 19496
rect 17547 19468 17592 19496
rect 16816 19456 16822 19468
rect 13320 19400 14688 19428
rect 13320 19388 13326 19400
rect 14734 19388 14740 19440
rect 14792 19428 14798 19440
rect 15206 19431 15264 19437
rect 15206 19428 15218 19431
rect 14792 19400 15218 19428
rect 14792 19388 14798 19400
rect 15206 19397 15218 19400
rect 15252 19397 15264 19431
rect 15206 19391 15264 19397
rect 15304 19400 17356 19428
rect 9861 19323 9919 19329
rect 9968 19332 10640 19360
rect 9968 19292 9996 19332
rect 10686 19320 10692 19372
rect 10744 19320 10750 19372
rect 10778 19320 10784 19372
rect 10836 19360 10842 19372
rect 10965 19363 11023 19369
rect 10965 19360 10977 19363
rect 10836 19332 10977 19360
rect 10836 19320 10842 19332
rect 10965 19329 10977 19332
rect 11011 19329 11023 19363
rect 10965 19323 11023 19329
rect 11330 19320 11336 19372
rect 11388 19360 11394 19372
rect 15304 19360 15332 19400
rect 11388 19332 15332 19360
rect 15473 19363 15531 19369
rect 11388 19320 11394 19332
rect 15473 19329 15485 19363
rect 15519 19360 15531 19363
rect 15654 19360 15660 19372
rect 15519 19332 15660 19360
rect 15519 19329 15531 19332
rect 15473 19323 15531 19329
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 15746 19320 15752 19372
rect 15804 19360 15810 19372
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15804 19332 15945 19360
rect 15804 19320 15810 19332
rect 15933 19329 15945 19332
rect 15979 19329 15991 19363
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 15933 19323 15991 19329
rect 16040 19332 16865 19360
rect 9692 19264 9996 19292
rect 5721 19227 5779 19233
rect 5721 19193 5733 19227
rect 5767 19193 5779 19227
rect 10704 19224 10732 19320
rect 10781 19227 10839 19233
rect 10781 19224 10793 19227
rect 10704 19196 10793 19224
rect 5721 19187 5779 19193
rect 10781 19193 10793 19196
rect 10827 19193 10839 19227
rect 10781 19187 10839 19193
rect 2590 19156 2596 19168
rect 2148 19128 2596 19156
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 2866 19116 2872 19168
rect 2924 19156 2930 19168
rect 3602 19156 3608 19168
rect 2924 19128 3608 19156
rect 2924 19116 2930 19128
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 14182 19116 14188 19168
rect 14240 19156 14246 19168
rect 16040 19156 16068 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19360 17095 19363
rect 17218 19360 17224 19372
rect 17083 19332 17224 19360
rect 17083 19329 17095 19332
rect 17037 19323 17095 19329
rect 17218 19320 17224 19332
rect 17276 19320 17282 19372
rect 17328 19292 17356 19400
rect 17420 19360 17448 19468
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 18782 19496 18788 19508
rect 18743 19468 18788 19496
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 21910 19456 21916 19508
rect 21968 19496 21974 19508
rect 21968 19468 22784 19496
rect 21968 19456 21974 19468
rect 18230 19388 18236 19440
rect 18288 19428 18294 19440
rect 19153 19431 19211 19437
rect 19153 19428 19165 19431
rect 18288 19400 19165 19428
rect 18288 19388 18294 19400
rect 19153 19397 19165 19400
rect 19199 19397 19211 19431
rect 19153 19391 19211 19397
rect 19245 19431 19303 19437
rect 19245 19397 19257 19431
rect 19291 19428 19303 19431
rect 19334 19428 19340 19440
rect 19291 19400 19340 19428
rect 19291 19397 19303 19400
rect 19245 19391 19303 19397
rect 19334 19388 19340 19400
rect 19392 19388 19398 19440
rect 20438 19428 20444 19440
rect 20364 19400 20444 19428
rect 17586 19360 17592 19372
rect 17420 19332 17592 19360
rect 17586 19320 17592 19332
rect 17644 19320 17650 19372
rect 17954 19360 17960 19372
rect 17915 19332 17960 19360
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 19978 19360 19984 19372
rect 19939 19332 19984 19360
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 20254 19360 20260 19372
rect 20215 19332 20260 19360
rect 20254 19320 20260 19332
rect 20312 19320 20318 19372
rect 20364 19369 20392 19400
rect 20438 19388 20444 19400
rect 20496 19388 20502 19440
rect 20622 19388 20628 19440
rect 20680 19428 20686 19440
rect 20680 19400 21220 19428
rect 20680 19388 20686 19400
rect 20349 19363 20407 19369
rect 20349 19329 20361 19363
rect 20395 19329 20407 19363
rect 20530 19360 20536 19372
rect 20491 19332 20536 19360
rect 20349 19323 20407 19329
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17328 19264 18061 19292
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18138 19252 18144 19304
rect 18196 19292 18202 19304
rect 18233 19295 18291 19301
rect 18233 19292 18245 19295
rect 18196 19264 18245 19292
rect 18196 19252 18202 19264
rect 18233 19261 18245 19264
rect 18279 19261 18291 19295
rect 18233 19255 18291 19261
rect 18248 19224 18276 19255
rect 19242 19252 19248 19304
rect 19300 19292 19306 19304
rect 19337 19295 19395 19301
rect 19337 19292 19349 19295
rect 19300 19264 19349 19292
rect 19300 19252 19306 19264
rect 19337 19261 19349 19264
rect 19383 19292 19395 19295
rect 20364 19292 20392 19323
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 21192 19369 21220 19400
rect 22002 19388 22008 19440
rect 22060 19428 22066 19440
rect 22060 19400 22600 19428
rect 22060 19388 22066 19400
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19329 21051 19363
rect 20993 19323 21051 19329
rect 21177 19363 21235 19369
rect 21177 19329 21189 19363
rect 21223 19329 21235 19363
rect 22462 19360 22468 19372
rect 22423 19332 22468 19360
rect 21177 19323 21235 19329
rect 19383 19264 20392 19292
rect 19383 19261 19395 19264
rect 19337 19255 19395 19261
rect 21008 19224 21036 19323
rect 22462 19320 22468 19332
rect 22520 19320 22526 19372
rect 22572 19369 22600 19400
rect 22756 19369 22784 19468
rect 23201 19431 23259 19437
rect 23201 19397 23213 19431
rect 23247 19428 23259 19431
rect 30098 19428 30104 19440
rect 23247 19400 30104 19428
rect 23247 19397 23259 19400
rect 23201 19391 23259 19397
rect 30098 19388 30104 19400
rect 30156 19388 30162 19440
rect 22557 19363 22615 19369
rect 22557 19329 22569 19363
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 22741 19363 22799 19369
rect 22741 19329 22753 19363
rect 22787 19329 22799 19363
rect 29822 19360 29828 19372
rect 29783 19332 29828 19360
rect 22741 19323 22799 19329
rect 29822 19320 29828 19332
rect 29880 19320 29886 19372
rect 18248 19196 21036 19224
rect 16758 19156 16764 19168
rect 14240 19128 16068 19156
rect 16719 19128 16764 19156
rect 14240 19116 14246 19128
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 19518 19116 19524 19168
rect 19576 19156 19582 19168
rect 19978 19156 19984 19168
rect 19576 19128 19984 19156
rect 19576 19116 19582 19128
rect 19978 19116 19984 19128
rect 20036 19156 20042 19168
rect 20073 19159 20131 19165
rect 20073 19156 20085 19159
rect 20036 19128 20085 19156
rect 20036 19116 20042 19128
rect 20073 19125 20085 19128
rect 20119 19125 20131 19159
rect 20073 19119 20131 19125
rect 20165 19159 20223 19165
rect 20165 19125 20177 19159
rect 20211 19156 20223 19159
rect 20346 19156 20352 19168
rect 20211 19128 20352 19156
rect 20211 19125 20223 19128
rect 20165 19119 20223 19125
rect 20346 19116 20352 19128
rect 20404 19116 20410 19168
rect 20438 19116 20444 19168
rect 20496 19156 20502 19168
rect 20993 19159 21051 19165
rect 20993 19156 21005 19159
rect 20496 19128 21005 19156
rect 20496 19116 20502 19128
rect 20993 19125 21005 19128
rect 21039 19125 21051 19159
rect 30006 19156 30012 19168
rect 29967 19128 30012 19156
rect 20993 19119 21051 19125
rect 30006 19116 30012 19128
rect 30064 19116 30070 19168
rect 1104 19066 30820 19088
rect 1104 19014 5915 19066
rect 5967 19014 5979 19066
rect 6031 19014 6043 19066
rect 6095 19014 6107 19066
rect 6159 19014 6171 19066
rect 6223 19014 15846 19066
rect 15898 19014 15910 19066
rect 15962 19014 15974 19066
rect 16026 19014 16038 19066
rect 16090 19014 16102 19066
rect 16154 19014 25776 19066
rect 25828 19014 25840 19066
rect 25892 19014 25904 19066
rect 25956 19014 25968 19066
rect 26020 19014 26032 19066
rect 26084 19014 30820 19066
rect 1104 18992 30820 19014
rect 2222 18952 2228 18964
rect 2183 18924 2228 18952
rect 2222 18912 2228 18924
rect 2280 18912 2286 18964
rect 3786 18912 3792 18964
rect 3844 18952 3850 18964
rect 12250 18952 12256 18964
rect 3844 18924 9444 18952
rect 12211 18924 12256 18952
rect 3844 18912 3850 18924
rect 1670 18884 1676 18896
rect 1583 18856 1676 18884
rect 1596 18816 1624 18856
rect 1670 18844 1676 18856
rect 1728 18884 1734 18896
rect 3326 18884 3332 18896
rect 1728 18856 3332 18884
rect 1728 18844 1734 18856
rect 3326 18844 3332 18856
rect 3384 18884 3390 18896
rect 4019 18887 4077 18893
rect 4019 18884 4031 18887
rect 3384 18856 4031 18884
rect 3384 18844 3390 18856
rect 4019 18853 4031 18856
rect 4065 18853 4077 18887
rect 4019 18847 4077 18853
rect 7852 18856 9352 18884
rect 1762 18816 1768 18828
rect 1504 18788 1624 18816
rect 1723 18788 1768 18816
rect 1504 18757 1532 18788
rect 1762 18776 1768 18788
rect 1820 18776 1826 18828
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18816 1915 18819
rect 1946 18816 1952 18828
rect 1903 18788 1952 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 1946 18776 1952 18788
rect 2004 18776 2010 18828
rect 3602 18776 3608 18828
rect 3660 18816 3666 18828
rect 3660 18788 5488 18816
rect 3660 18776 3666 18788
rect 1489 18751 1547 18757
rect 1489 18717 1501 18751
rect 1535 18717 1547 18751
rect 1489 18711 1547 18717
rect 1578 18708 1584 18760
rect 1636 18748 1642 18760
rect 1673 18751 1731 18757
rect 1673 18748 1685 18751
rect 1636 18720 1685 18748
rect 1636 18708 1642 18720
rect 1673 18717 1685 18720
rect 1719 18717 1731 18751
rect 1673 18711 1731 18717
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18748 2099 18751
rect 3234 18748 3240 18760
rect 2087 18720 3240 18748
rect 2087 18717 2099 18720
rect 2041 18711 2099 18717
rect 3234 18708 3240 18720
rect 3292 18708 3298 18760
rect 3786 18748 3792 18760
rect 3747 18720 3792 18748
rect 3786 18708 3792 18720
rect 3844 18708 3850 18760
rect 5460 18757 5488 18788
rect 6362 18776 6368 18828
rect 6420 18816 6426 18828
rect 7852 18825 7880 18856
rect 6457 18819 6515 18825
rect 6457 18816 6469 18819
rect 6420 18788 6469 18816
rect 6420 18776 6426 18788
rect 6457 18785 6469 18788
rect 6503 18785 6515 18819
rect 6457 18779 6515 18785
rect 7837 18819 7895 18825
rect 7837 18785 7849 18819
rect 7883 18785 7895 18819
rect 7837 18779 7895 18785
rect 7929 18819 7987 18825
rect 7929 18785 7941 18819
rect 7975 18816 7987 18819
rect 9030 18816 9036 18828
rect 7975 18788 9036 18816
rect 7975 18785 7987 18788
rect 7929 18779 7987 18785
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18717 5503 18751
rect 6178 18748 6184 18760
rect 6139 18720 6184 18748
rect 5445 18711 5503 18717
rect 6178 18708 6184 18720
rect 6236 18708 6242 18760
rect 3145 18683 3203 18689
rect 3145 18649 3157 18683
rect 3191 18680 3203 18683
rect 3326 18680 3332 18692
rect 3191 18652 3332 18680
rect 3191 18649 3203 18652
rect 3145 18643 3203 18649
rect 3326 18640 3332 18652
rect 3384 18680 3390 18692
rect 4062 18680 4068 18692
rect 3384 18652 4068 18680
rect 3384 18640 3390 18652
rect 4062 18640 4068 18652
rect 4120 18640 4126 18692
rect 6472 18680 6500 18779
rect 9030 18776 9036 18788
rect 9088 18816 9094 18828
rect 9217 18819 9275 18825
rect 9217 18816 9229 18819
rect 9088 18788 9229 18816
rect 9088 18776 9094 18788
rect 9217 18785 9229 18788
rect 9263 18785 9275 18819
rect 9217 18779 9275 18785
rect 9324 18760 9352 18856
rect 7650 18748 7656 18760
rect 7611 18720 7656 18748
rect 7650 18708 7656 18720
rect 7708 18708 7714 18760
rect 8018 18708 8024 18760
rect 8076 18748 8082 18760
rect 8205 18751 8263 18757
rect 8076 18720 8121 18748
rect 8076 18708 8082 18720
rect 8205 18717 8217 18751
rect 8251 18748 8263 18751
rect 8386 18748 8392 18760
rect 8251 18720 8392 18748
rect 8251 18717 8263 18720
rect 8205 18711 8263 18717
rect 6730 18680 6736 18692
rect 6472 18652 6736 18680
rect 6730 18640 6736 18652
rect 6788 18680 6794 18692
rect 8220 18680 8248 18711
rect 8386 18708 8392 18720
rect 8444 18748 8450 18760
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8444 18720 8953 18748
rect 8444 18708 8450 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9125 18751 9183 18757
rect 9125 18717 9137 18751
rect 9171 18717 9183 18751
rect 9306 18748 9312 18760
rect 9267 18720 9312 18748
rect 9125 18711 9183 18717
rect 6788 18652 8248 18680
rect 6788 18640 6794 18652
rect 8846 18640 8852 18692
rect 8904 18680 8910 18692
rect 9140 18680 9168 18711
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 8904 18652 9168 18680
rect 9416 18680 9444 18924
rect 12250 18912 12256 18924
rect 12308 18912 12314 18964
rect 12434 18912 12440 18964
rect 12492 18952 12498 18964
rect 16758 18952 16764 18964
rect 12492 18924 16764 18952
rect 12492 18912 12498 18924
rect 16758 18912 16764 18924
rect 16816 18912 16822 18964
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 18233 18955 18291 18961
rect 18233 18952 18245 18955
rect 18012 18924 18245 18952
rect 18012 18912 18018 18924
rect 18233 18921 18245 18924
rect 18279 18921 18291 18955
rect 19334 18952 19340 18964
rect 19295 18924 19340 18952
rect 18233 18915 18291 18921
rect 19334 18912 19340 18924
rect 19392 18912 19398 18964
rect 19978 18912 19984 18964
rect 20036 18952 20042 18964
rect 20530 18952 20536 18964
rect 20036 18924 20536 18952
rect 20036 18912 20042 18924
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 29914 18952 29920 18964
rect 29875 18924 29920 18952
rect 29914 18912 29920 18924
rect 29972 18912 29978 18964
rect 11054 18884 11060 18896
rect 11015 18856 11060 18884
rect 11054 18844 11060 18856
rect 11112 18884 11118 18896
rect 11974 18884 11980 18896
rect 11112 18856 11980 18884
rect 11112 18844 11118 18856
rect 11974 18844 11980 18856
rect 12032 18844 12038 18896
rect 14277 18887 14335 18893
rect 14277 18853 14289 18887
rect 14323 18884 14335 18887
rect 14918 18884 14924 18896
rect 14323 18856 14924 18884
rect 14323 18853 14335 18856
rect 14277 18847 14335 18853
rect 14918 18844 14924 18856
rect 14976 18884 14982 18896
rect 14976 18856 17448 18884
rect 14976 18844 14982 18856
rect 11422 18776 11428 18828
rect 11480 18816 11486 18828
rect 11882 18816 11888 18828
rect 11480 18788 11744 18816
rect 11843 18788 11888 18816
rect 11480 18776 11486 18788
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 11517 18751 11575 18757
rect 9548 18720 11008 18748
rect 9548 18708 9554 18720
rect 9416 18652 10088 18680
rect 8904 18640 8910 18652
rect 3050 18612 3056 18624
rect 3011 18584 3056 18612
rect 3050 18572 3056 18584
rect 3108 18572 3114 18624
rect 5534 18612 5540 18624
rect 5495 18584 5540 18612
rect 5534 18572 5540 18584
rect 5592 18572 5598 18624
rect 7466 18612 7472 18624
rect 7427 18584 7472 18612
rect 7466 18572 7472 18584
rect 7524 18572 7530 18624
rect 9677 18615 9735 18621
rect 9677 18581 9689 18615
rect 9723 18612 9735 18615
rect 9950 18612 9956 18624
rect 9723 18584 9956 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 10060 18612 10088 18652
rect 10778 18640 10784 18692
rect 10836 18680 10842 18692
rect 10873 18683 10931 18689
rect 10873 18680 10885 18683
rect 10836 18652 10885 18680
rect 10836 18640 10842 18652
rect 10873 18649 10885 18652
rect 10919 18649 10931 18683
rect 10980 18680 11008 18720
rect 11517 18717 11529 18751
rect 11563 18748 11575 18751
rect 11606 18748 11612 18760
rect 11563 18720 11612 18748
rect 11563 18717 11575 18720
rect 11517 18711 11575 18717
rect 11606 18708 11612 18720
rect 11664 18708 11670 18760
rect 11716 18757 11744 18788
rect 11882 18776 11888 18788
rect 11940 18776 11946 18828
rect 12158 18816 12164 18828
rect 11992 18788 12164 18816
rect 11701 18751 11759 18757
rect 11701 18717 11713 18751
rect 11747 18717 11759 18751
rect 11701 18711 11759 18717
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18748 11851 18751
rect 11992 18748 12020 18788
rect 12158 18776 12164 18788
rect 12216 18776 12222 18828
rect 15028 18825 15056 18856
rect 15013 18819 15071 18825
rect 15013 18785 15025 18819
rect 15059 18785 15071 18819
rect 17034 18816 17040 18828
rect 15013 18779 15071 18785
rect 16316 18788 17040 18816
rect 11839 18720 12020 18748
rect 12069 18751 12127 18757
rect 11839 18717 11851 18720
rect 11793 18711 11851 18717
rect 12069 18717 12081 18751
rect 12115 18748 12127 18751
rect 12526 18748 12532 18760
rect 12115 18720 12532 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 12710 18748 12716 18760
rect 12671 18720 12716 18748
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 14182 18748 14188 18760
rect 14143 18720 14188 18748
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 16316 18757 16344 18788
rect 17034 18776 17040 18788
rect 17092 18776 17098 18828
rect 17310 18816 17316 18828
rect 17271 18788 17316 18816
rect 17310 18776 17316 18788
rect 17368 18776 17374 18828
rect 17420 18816 17448 18856
rect 18046 18844 18052 18896
rect 18104 18884 18110 18896
rect 21637 18887 21695 18893
rect 21637 18884 21649 18887
rect 18104 18856 21649 18884
rect 18104 18844 18110 18856
rect 21637 18853 21649 18856
rect 21683 18853 21695 18887
rect 21637 18847 21695 18853
rect 18138 18816 18144 18828
rect 17420 18788 18144 18816
rect 18138 18776 18144 18788
rect 18196 18776 18202 18828
rect 19058 18776 19064 18828
rect 19116 18816 19122 18828
rect 20438 18816 20444 18828
rect 19116 18788 19380 18816
rect 20399 18788 20444 18816
rect 19116 18776 19122 18788
rect 16301 18751 16359 18757
rect 16301 18717 16313 18751
rect 16347 18717 16359 18751
rect 16301 18711 16359 18717
rect 16942 18708 16948 18760
rect 17000 18748 17006 18760
rect 17589 18751 17647 18757
rect 17589 18748 17601 18751
rect 17000 18720 17601 18748
rect 17000 18708 17006 18720
rect 17589 18717 17601 18720
rect 17635 18717 17647 18751
rect 17589 18711 17647 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18748 18475 18751
rect 18782 18748 18788 18760
rect 18463 18720 18788 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 19245 18751 19303 18757
rect 19245 18717 19257 18751
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 15105 18683 15163 18689
rect 15105 18680 15117 18683
rect 10980 18652 15117 18680
rect 10873 18643 10931 18649
rect 15105 18649 15117 18652
rect 15151 18649 15163 18683
rect 15105 18643 15163 18649
rect 15197 18683 15255 18689
rect 15197 18649 15209 18683
rect 15243 18680 15255 18683
rect 16025 18683 16083 18689
rect 16025 18680 16037 18683
rect 15243 18652 16037 18680
rect 15243 18649 15255 18652
rect 15197 18643 15255 18649
rect 16025 18649 16037 18652
rect 16071 18649 16083 18683
rect 16025 18643 16083 18649
rect 18138 18640 18144 18692
rect 18196 18680 18202 18692
rect 19260 18680 19288 18711
rect 18196 18652 19288 18680
rect 19352 18680 19380 18788
rect 20438 18776 20444 18788
rect 20496 18776 20502 18828
rect 20533 18819 20591 18825
rect 20533 18785 20545 18819
rect 20579 18785 20591 18819
rect 20533 18779 20591 18785
rect 20346 18748 20352 18760
rect 20307 18720 20352 18748
rect 20346 18708 20352 18720
rect 20404 18708 20410 18760
rect 20548 18680 20576 18779
rect 21910 18776 21916 18828
rect 21968 18816 21974 18828
rect 22189 18819 22247 18825
rect 22189 18816 22201 18819
rect 21968 18788 22201 18816
rect 21968 18776 21974 18788
rect 22189 18785 22201 18788
rect 22235 18785 22247 18819
rect 22189 18779 22247 18785
rect 22002 18748 22008 18760
rect 21963 18720 22008 18748
rect 22002 18708 22008 18720
rect 22060 18708 22066 18760
rect 22097 18751 22155 18757
rect 22097 18717 22109 18751
rect 22143 18748 22155 18751
rect 22462 18748 22468 18760
rect 22143 18720 22468 18748
rect 22143 18717 22155 18720
rect 22097 18711 22155 18717
rect 22462 18708 22468 18720
rect 22520 18708 22526 18760
rect 29638 18708 29644 18760
rect 29696 18748 29702 18760
rect 29917 18751 29975 18757
rect 29917 18748 29929 18751
rect 29696 18720 29929 18748
rect 29696 18708 29702 18720
rect 29917 18717 29929 18720
rect 29963 18717 29975 18751
rect 30098 18748 30104 18760
rect 30059 18720 30104 18748
rect 29917 18711 29975 18717
rect 30098 18708 30104 18720
rect 30156 18708 30162 18760
rect 19352 18652 20576 18680
rect 18196 18640 18202 18652
rect 12897 18615 12955 18621
rect 12897 18612 12909 18615
rect 10060 18584 12909 18612
rect 12897 18581 12909 18584
rect 12943 18612 12955 18615
rect 13630 18612 13636 18624
rect 12943 18584 13636 18612
rect 12943 18581 12955 18584
rect 12897 18575 12955 18581
rect 13630 18572 13636 18584
rect 13688 18572 13694 18624
rect 15378 18572 15384 18624
rect 15436 18612 15442 18624
rect 15565 18615 15623 18621
rect 15565 18612 15577 18615
rect 15436 18584 15577 18612
rect 15436 18572 15442 18584
rect 15565 18581 15577 18584
rect 15611 18581 15623 18615
rect 15565 18575 15623 18581
rect 19794 18572 19800 18624
rect 19852 18612 19858 18624
rect 19981 18615 20039 18621
rect 19981 18612 19993 18615
rect 19852 18584 19993 18612
rect 19852 18572 19858 18584
rect 19981 18581 19993 18584
rect 20027 18581 20039 18615
rect 19981 18575 20039 18581
rect 1104 18522 30820 18544
rect 1104 18470 10880 18522
rect 10932 18470 10944 18522
rect 10996 18470 11008 18522
rect 11060 18470 11072 18522
rect 11124 18470 11136 18522
rect 11188 18470 20811 18522
rect 20863 18470 20875 18522
rect 20927 18470 20939 18522
rect 20991 18470 21003 18522
rect 21055 18470 21067 18522
rect 21119 18470 30820 18522
rect 1104 18448 30820 18470
rect 2409 18411 2467 18417
rect 2409 18377 2421 18411
rect 2455 18408 2467 18411
rect 2498 18408 2504 18420
rect 2455 18380 2504 18408
rect 2455 18377 2467 18380
rect 2409 18371 2467 18377
rect 2498 18368 2504 18380
rect 2556 18368 2562 18420
rect 4157 18411 4215 18417
rect 4157 18377 4169 18411
rect 4203 18408 4215 18411
rect 4430 18408 4436 18420
rect 4203 18380 4436 18408
rect 4203 18377 4215 18380
rect 4157 18371 4215 18377
rect 4430 18368 4436 18380
rect 4488 18368 4494 18420
rect 4801 18411 4859 18417
rect 4801 18377 4813 18411
rect 4847 18377 4859 18411
rect 5718 18408 5724 18420
rect 5679 18380 5724 18408
rect 4801 18371 4859 18377
rect 4816 18340 4844 18371
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 7650 18368 7656 18420
rect 7708 18408 7714 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 7708 18380 8309 18408
rect 7708 18368 7714 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 8297 18371 8355 18377
rect 8754 18368 8760 18420
rect 8812 18408 8818 18420
rect 8849 18411 8907 18417
rect 8849 18408 8861 18411
rect 8812 18380 8861 18408
rect 8812 18368 8818 18380
rect 8849 18377 8861 18380
rect 8895 18408 8907 18411
rect 9490 18408 9496 18420
rect 8895 18380 9496 18408
rect 8895 18377 8907 18380
rect 8849 18371 8907 18377
rect 9490 18368 9496 18380
rect 9548 18368 9554 18420
rect 12066 18408 12072 18420
rect 12027 18380 12072 18408
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 15378 18408 15384 18420
rect 15339 18380 15384 18408
rect 15378 18368 15384 18380
rect 15436 18368 15442 18420
rect 18966 18408 18972 18420
rect 18927 18380 18972 18408
rect 18966 18368 18972 18380
rect 19024 18368 19030 18420
rect 19334 18408 19340 18420
rect 19247 18380 19340 18408
rect 19334 18368 19340 18380
rect 19392 18408 19398 18420
rect 19702 18408 19708 18420
rect 19392 18380 19708 18408
rect 19392 18368 19398 18380
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 20533 18411 20591 18417
rect 20533 18377 20545 18411
rect 20579 18408 20591 18411
rect 20622 18408 20628 18420
rect 20579 18380 20628 18408
rect 20579 18377 20591 18380
rect 20533 18371 20591 18377
rect 20622 18368 20628 18380
rect 20680 18368 20686 18420
rect 20714 18368 20720 18420
rect 20772 18408 20778 18420
rect 20901 18411 20959 18417
rect 20901 18408 20913 18411
rect 20772 18380 20913 18408
rect 20772 18368 20778 18380
rect 20901 18377 20913 18380
rect 20947 18408 20959 18411
rect 21821 18411 21879 18417
rect 21821 18408 21833 18411
rect 20947 18380 21833 18408
rect 20947 18377 20959 18380
rect 20901 18371 20959 18377
rect 21821 18377 21833 18380
rect 21867 18377 21879 18411
rect 21821 18371 21879 18377
rect 29822 18368 29828 18420
rect 29880 18408 29886 18420
rect 30009 18411 30067 18417
rect 30009 18408 30021 18411
rect 29880 18380 30021 18408
rect 29880 18368 29886 18380
rect 30009 18377 30021 18380
rect 30055 18377 30067 18411
rect 30009 18371 30067 18377
rect 3436 18312 4844 18340
rect 5629 18343 5687 18349
rect 1670 18272 1676 18284
rect 1631 18244 1676 18272
rect 1670 18232 1676 18244
rect 1728 18232 1734 18284
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 2225 18275 2283 18281
rect 2225 18241 2237 18275
rect 2271 18272 2283 18275
rect 2866 18272 2872 18284
rect 2271 18244 2872 18272
rect 2271 18241 2283 18244
rect 2225 18235 2283 18241
rect 2866 18232 2872 18244
rect 2924 18232 2930 18284
rect 2958 18232 2964 18284
rect 3016 18272 3022 18284
rect 3436 18281 3464 18312
rect 5629 18309 5641 18343
rect 5675 18340 5687 18343
rect 5810 18340 5816 18352
rect 5675 18312 5816 18340
rect 5675 18309 5687 18312
rect 5629 18303 5687 18309
rect 5810 18300 5816 18312
rect 5868 18340 5874 18352
rect 6178 18340 6184 18352
rect 5868 18312 6184 18340
rect 5868 18300 5874 18312
rect 6178 18300 6184 18312
rect 6236 18300 6242 18352
rect 7184 18343 7242 18349
rect 7184 18309 7196 18343
rect 7230 18340 7242 18343
rect 7466 18340 7472 18352
rect 7230 18312 7472 18340
rect 7230 18309 7242 18312
rect 7184 18303 7242 18309
rect 7466 18300 7472 18312
rect 7524 18300 7530 18352
rect 7558 18300 7564 18352
rect 7616 18340 7622 18352
rect 8018 18340 8024 18352
rect 7616 18312 8024 18340
rect 7616 18300 7622 18312
rect 8018 18300 8024 18312
rect 8076 18300 8082 18352
rect 9674 18300 9680 18352
rect 9732 18340 9738 18352
rect 9732 18312 10272 18340
rect 9732 18300 9738 18312
rect 3053 18275 3111 18281
rect 3053 18272 3065 18275
rect 3016 18244 3065 18272
rect 3016 18232 3022 18244
rect 3053 18241 3065 18244
rect 3099 18241 3111 18275
rect 3053 18235 3111 18241
rect 3421 18275 3479 18281
rect 3421 18241 3433 18275
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18272 3663 18275
rect 4062 18272 4068 18284
rect 3651 18244 4068 18272
rect 3651 18241 3663 18244
rect 3605 18235 3663 18241
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 4154 18232 4160 18284
rect 4212 18272 4218 18284
rect 4249 18275 4307 18281
rect 4249 18272 4261 18275
rect 4212 18244 4261 18272
rect 4212 18232 4218 18244
rect 4249 18241 4261 18244
rect 4295 18241 4307 18275
rect 4249 18235 4307 18241
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18241 5043 18275
rect 4985 18235 5043 18241
rect 1762 18164 1768 18216
rect 1820 18204 1826 18216
rect 1949 18207 2007 18213
rect 1949 18204 1961 18207
rect 1820 18176 1961 18204
rect 1820 18164 1826 18176
rect 1949 18173 1961 18176
rect 1995 18173 2007 18207
rect 1949 18167 2007 18173
rect 2041 18207 2099 18213
rect 2041 18173 2053 18207
rect 2087 18204 2099 18207
rect 3142 18204 3148 18216
rect 2087 18176 3148 18204
rect 2087 18173 2099 18176
rect 2041 18167 2099 18173
rect 1964 18136 1992 18167
rect 3142 18164 3148 18176
rect 3200 18204 3206 18216
rect 3237 18207 3295 18213
rect 3237 18204 3249 18207
rect 3200 18176 3249 18204
rect 3200 18164 3206 18176
rect 3237 18173 3249 18176
rect 3283 18173 3295 18207
rect 3237 18167 3295 18173
rect 3329 18207 3387 18213
rect 3329 18173 3341 18207
rect 3375 18173 3387 18207
rect 3329 18167 3387 18173
rect 2590 18136 2596 18148
rect 1964 18108 2596 18136
rect 2590 18096 2596 18108
rect 2648 18136 2654 18148
rect 3344 18136 3372 18167
rect 3878 18164 3884 18216
rect 3936 18204 3942 18216
rect 5000 18204 5028 18235
rect 6638 18232 6644 18284
rect 6696 18272 6702 18284
rect 6917 18275 6975 18281
rect 6917 18272 6929 18275
rect 6696 18244 6929 18272
rect 6696 18232 6702 18244
rect 6917 18241 6929 18244
rect 6963 18241 6975 18275
rect 6917 18235 6975 18241
rect 9950 18232 9956 18284
rect 10008 18281 10014 18284
rect 10244 18281 10272 18312
rect 10778 18300 10784 18352
rect 10836 18340 10842 18352
rect 12710 18340 12716 18352
rect 10836 18312 12716 18340
rect 10836 18300 10842 18312
rect 10980 18281 11008 18312
rect 12710 18300 12716 18312
rect 12768 18340 12774 18352
rect 12805 18343 12863 18349
rect 12805 18340 12817 18343
rect 12768 18312 12817 18340
rect 12768 18300 12774 18312
rect 12805 18309 12817 18312
rect 12851 18309 12863 18343
rect 15286 18340 15292 18352
rect 15247 18312 15292 18340
rect 12805 18303 12863 18309
rect 15286 18300 15292 18312
rect 15344 18300 15350 18352
rect 19429 18343 19487 18349
rect 19429 18309 19441 18343
rect 19475 18340 19487 18343
rect 19518 18340 19524 18352
rect 19475 18312 19524 18340
rect 19475 18309 19487 18312
rect 19429 18303 19487 18309
rect 19518 18300 19524 18312
rect 19576 18300 19582 18352
rect 10008 18272 10020 18281
rect 10229 18275 10287 18281
rect 10008 18244 10053 18272
rect 10008 18235 10020 18244
rect 10229 18241 10241 18275
rect 10275 18241 10287 18275
rect 10229 18235 10287 18241
rect 10965 18275 11023 18281
rect 10965 18241 10977 18275
rect 11011 18241 11023 18275
rect 10965 18235 11023 18241
rect 11977 18275 12035 18281
rect 11977 18241 11989 18275
rect 12023 18241 12035 18275
rect 11977 18235 12035 18241
rect 10008 18232 10014 18235
rect 3936 18176 5028 18204
rect 3936 18164 3942 18176
rect 2648 18108 3372 18136
rect 2648 18096 2654 18108
rect 10594 18096 10600 18148
rect 10652 18136 10658 18148
rect 10781 18139 10839 18145
rect 10781 18136 10793 18139
rect 10652 18108 10793 18136
rect 10652 18096 10658 18108
rect 10781 18105 10793 18108
rect 10827 18136 10839 18139
rect 11992 18136 12020 18235
rect 12618 18232 12624 18284
rect 12676 18272 12682 18284
rect 12897 18275 12955 18281
rect 12897 18272 12909 18275
rect 12676 18244 12909 18272
rect 12676 18232 12682 18244
rect 12897 18241 12909 18244
rect 12943 18272 12955 18275
rect 13998 18272 14004 18284
rect 12943 18244 14004 18272
rect 12943 18241 12955 18244
rect 12897 18235 12955 18241
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 16853 18275 16911 18281
rect 16853 18241 16865 18275
rect 16899 18272 16911 18275
rect 17678 18272 17684 18284
rect 16899 18244 17684 18272
rect 16899 18241 16911 18244
rect 16853 18235 16911 18241
rect 17678 18232 17684 18244
rect 17736 18232 17742 18284
rect 19150 18232 19156 18284
rect 19208 18272 19214 18284
rect 19702 18272 19708 18284
rect 19208 18244 19708 18272
rect 19208 18232 19214 18244
rect 19702 18232 19708 18244
rect 19760 18232 19766 18284
rect 20993 18275 21051 18281
rect 20993 18241 21005 18275
rect 21039 18272 21051 18275
rect 21818 18272 21824 18284
rect 21039 18244 21824 18272
rect 21039 18241 21051 18244
rect 20993 18235 21051 18241
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 22002 18272 22008 18284
rect 21963 18244 22008 18272
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 29270 18232 29276 18284
rect 29328 18272 29334 18284
rect 29917 18275 29975 18281
rect 29917 18272 29929 18275
rect 29328 18244 29929 18272
rect 29328 18232 29334 18244
rect 29917 18241 29929 18244
rect 29963 18241 29975 18275
rect 30098 18272 30104 18284
rect 30059 18244 30104 18272
rect 29917 18235 29975 18241
rect 30098 18232 30104 18244
rect 30156 18232 30162 18284
rect 15565 18207 15623 18213
rect 15565 18173 15577 18207
rect 15611 18204 15623 18207
rect 16666 18204 16672 18216
rect 15611 18176 16672 18204
rect 15611 18173 15623 18176
rect 15565 18167 15623 18173
rect 16666 18164 16672 18176
rect 16724 18164 16730 18216
rect 16758 18164 16764 18216
rect 16816 18204 16822 18216
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 16816 18176 17141 18204
rect 16816 18164 16822 18176
rect 17129 18173 17141 18176
rect 17175 18204 17187 18207
rect 17402 18204 17408 18216
rect 17175 18176 17408 18204
rect 17175 18173 17187 18176
rect 17129 18167 17187 18173
rect 17402 18164 17408 18176
rect 17460 18204 17466 18216
rect 19242 18204 19248 18216
rect 17460 18176 19248 18204
rect 17460 18164 17466 18176
rect 19242 18164 19248 18176
rect 19300 18204 19306 18216
rect 19521 18207 19579 18213
rect 19521 18204 19533 18207
rect 19300 18176 19533 18204
rect 19300 18164 19306 18176
rect 19521 18173 19533 18176
rect 19567 18204 19579 18207
rect 21085 18207 21143 18213
rect 21085 18204 21097 18207
rect 19567 18176 21097 18204
rect 19567 18173 19579 18176
rect 19521 18167 19579 18173
rect 21085 18173 21097 18176
rect 21131 18173 21143 18207
rect 21085 18167 21143 18173
rect 10827 18108 12020 18136
rect 10827 18105 10839 18108
rect 10781 18099 10839 18105
rect 16206 18096 16212 18148
rect 16264 18136 16270 18148
rect 17586 18136 17592 18148
rect 16264 18108 17592 18136
rect 16264 18096 16270 18108
rect 17586 18096 17592 18108
rect 17644 18096 17650 18148
rect 2866 18068 2872 18080
rect 2827 18040 2872 18068
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 5718 18028 5724 18080
rect 5776 18068 5782 18080
rect 6638 18068 6644 18080
rect 5776 18040 6644 18068
rect 5776 18028 5782 18040
rect 6638 18028 6644 18040
rect 6696 18028 6702 18080
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 7834 18068 7840 18080
rect 7340 18040 7840 18068
rect 7340 18028 7346 18040
rect 7834 18028 7840 18040
rect 7892 18028 7898 18080
rect 14642 18028 14648 18080
rect 14700 18068 14706 18080
rect 14921 18071 14979 18077
rect 14921 18068 14933 18071
rect 14700 18040 14933 18068
rect 14700 18028 14706 18040
rect 14921 18037 14933 18040
rect 14967 18037 14979 18071
rect 14921 18031 14979 18037
rect 1104 17978 30820 18000
rect 1104 17926 5915 17978
rect 5967 17926 5979 17978
rect 6031 17926 6043 17978
rect 6095 17926 6107 17978
rect 6159 17926 6171 17978
rect 6223 17926 15846 17978
rect 15898 17926 15910 17978
rect 15962 17926 15974 17978
rect 16026 17926 16038 17978
rect 16090 17926 16102 17978
rect 16154 17926 25776 17978
rect 25828 17926 25840 17978
rect 25892 17926 25904 17978
rect 25956 17926 25968 17978
rect 26020 17926 26032 17978
rect 26084 17926 30820 17978
rect 1104 17904 30820 17926
rect 5810 17824 5816 17876
rect 5868 17864 5874 17876
rect 5997 17867 6055 17873
rect 5997 17864 6009 17867
rect 5868 17836 6009 17864
rect 5868 17824 5874 17836
rect 5997 17833 6009 17836
rect 6043 17833 6055 17867
rect 7926 17864 7932 17876
rect 7887 17836 7932 17864
rect 5997 17827 6055 17833
rect 7926 17824 7932 17836
rect 7984 17824 7990 17876
rect 11238 17824 11244 17876
rect 11296 17864 11302 17876
rect 11333 17867 11391 17873
rect 11333 17864 11345 17867
rect 11296 17836 11345 17864
rect 11296 17824 11302 17836
rect 11333 17833 11345 17836
rect 11379 17833 11391 17867
rect 15473 17867 15531 17873
rect 11333 17827 11391 17833
rect 13188 17836 14504 17864
rect 4614 17796 4620 17808
rect 3804 17768 4620 17796
rect 3804 17740 3832 17768
rect 4614 17756 4620 17768
rect 4672 17756 4678 17808
rect 3786 17728 3792 17740
rect 3747 17700 3792 17728
rect 3786 17688 3792 17700
rect 3844 17688 3850 17740
rect 3970 17688 3976 17740
rect 4028 17728 4034 17740
rect 13188 17728 13216 17836
rect 14476 17808 14504 17836
rect 15473 17833 15485 17867
rect 15519 17864 15531 17867
rect 15746 17864 15752 17876
rect 15519 17836 15752 17864
rect 15519 17833 15531 17836
rect 15473 17827 15531 17833
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 16761 17867 16819 17873
rect 16761 17833 16773 17867
rect 16807 17864 16819 17867
rect 17034 17864 17040 17876
rect 16807 17836 17040 17864
rect 16807 17833 16819 17836
rect 16761 17827 16819 17833
rect 17034 17824 17040 17836
rect 17092 17824 17098 17876
rect 19242 17824 19248 17876
rect 19300 17864 19306 17876
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 19300 17836 19717 17864
rect 19300 17824 19306 17836
rect 19705 17833 19717 17836
rect 19751 17833 19763 17867
rect 19705 17827 19763 17833
rect 20625 17867 20683 17873
rect 20625 17833 20637 17867
rect 20671 17864 20683 17867
rect 22002 17864 22008 17876
rect 20671 17836 22008 17864
rect 20671 17833 20683 17836
rect 20625 17827 20683 17833
rect 22002 17824 22008 17836
rect 22060 17824 22066 17876
rect 13265 17799 13323 17805
rect 13265 17765 13277 17799
rect 13311 17796 13323 17799
rect 14458 17796 14464 17808
rect 13311 17768 14320 17796
rect 14419 17768 14464 17796
rect 13311 17765 13323 17768
rect 13265 17759 13323 17765
rect 14292 17737 14320 17768
rect 14458 17756 14464 17768
rect 14516 17756 14522 17808
rect 18046 17796 18052 17808
rect 14568 17768 18052 17796
rect 13357 17731 13415 17737
rect 13357 17728 13369 17731
rect 4028 17700 5304 17728
rect 4028 17688 4034 17700
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17660 1639 17663
rect 1670 17660 1676 17672
rect 1627 17632 1676 17660
rect 1627 17629 1639 17632
rect 1581 17623 1639 17629
rect 1670 17620 1676 17632
rect 1728 17620 1734 17672
rect 1848 17663 1906 17669
rect 1848 17629 1860 17663
rect 1894 17660 1906 17663
rect 2866 17660 2872 17672
rect 1894 17632 2872 17660
rect 1894 17629 1906 17632
rect 1848 17623 1906 17629
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 4062 17660 4068 17672
rect 4023 17632 4068 17660
rect 4062 17620 4068 17632
rect 4120 17620 4126 17672
rect 5276 17669 5304 17700
rect 6104 17700 6684 17728
rect 13188 17700 13369 17728
rect 6104 17669 6132 17700
rect 5261 17663 5319 17669
rect 5261 17629 5273 17663
rect 5307 17629 5319 17663
rect 5261 17623 5319 17629
rect 6089 17663 6147 17669
rect 6089 17629 6101 17663
rect 6135 17629 6147 17663
rect 6089 17623 6147 17629
rect 6549 17663 6607 17669
rect 6549 17629 6561 17663
rect 6595 17629 6607 17663
rect 6656 17660 6684 17700
rect 13357 17697 13369 17700
rect 13403 17697 13415 17731
rect 13357 17691 13415 17697
rect 13541 17731 13599 17737
rect 13541 17697 13553 17731
rect 13587 17728 13599 17731
rect 14277 17731 14335 17737
rect 13587 17700 14228 17728
rect 13587 17697 13599 17700
rect 13541 17691 13599 17697
rect 7650 17660 7656 17672
rect 6656 17632 7656 17660
rect 6549 17623 6607 17629
rect 3878 17552 3884 17604
rect 3936 17592 3942 17604
rect 6564 17592 6592 17623
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 9953 17663 10011 17669
rect 9953 17660 9965 17663
rect 9732 17632 9965 17660
rect 9732 17620 9738 17632
rect 9953 17629 9965 17632
rect 9999 17629 10011 17663
rect 9953 17623 10011 17629
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17629 12495 17663
rect 12437 17623 12495 17629
rect 12621 17663 12679 17669
rect 12621 17629 12633 17663
rect 12667 17660 12679 17663
rect 12667 17632 13216 17660
rect 12667 17629 12679 17632
rect 12621 17623 12679 17629
rect 3936 17564 6592 17592
rect 6816 17595 6874 17601
rect 3936 17552 3942 17564
rect 6816 17561 6828 17595
rect 6862 17592 6874 17595
rect 7466 17592 7472 17604
rect 6862 17564 7472 17592
rect 6862 17561 6874 17564
rect 6816 17555 6874 17561
rect 7466 17552 7472 17564
rect 7524 17552 7530 17604
rect 9122 17552 9128 17604
rect 9180 17592 9186 17604
rect 10198 17595 10256 17601
rect 10198 17592 10210 17595
rect 9180 17564 10210 17592
rect 9180 17552 9186 17564
rect 10198 17561 10210 17564
rect 10244 17561 10256 17595
rect 12452 17592 12480 17623
rect 13188 17592 13216 17632
rect 13262 17620 13268 17672
rect 13320 17660 13326 17672
rect 14090 17660 14096 17672
rect 13320 17632 13365 17660
rect 14051 17632 14096 17660
rect 13320 17620 13326 17632
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14200 17660 14228 17700
rect 14277 17697 14289 17731
rect 14323 17697 14335 17731
rect 14277 17691 14335 17697
rect 14366 17688 14372 17740
rect 14424 17728 14430 17740
rect 14424 17700 14469 17728
rect 14424 17688 14430 17700
rect 14568 17669 14596 17768
rect 18046 17756 18052 17768
rect 18104 17756 18110 17808
rect 18230 17756 18236 17808
rect 18288 17796 18294 17808
rect 18417 17799 18475 17805
rect 18417 17796 18429 17799
rect 18288 17768 18429 17796
rect 18288 17756 18294 17768
rect 18417 17765 18429 17768
rect 18463 17765 18475 17799
rect 19518 17796 19524 17808
rect 19431 17768 19524 17796
rect 18417 17759 18475 17765
rect 15381 17731 15439 17737
rect 15381 17697 15393 17731
rect 15427 17728 15439 17731
rect 15470 17728 15476 17740
rect 15427 17700 15476 17728
rect 15427 17697 15439 17700
rect 15381 17691 15439 17697
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 15565 17731 15623 17737
rect 15565 17697 15577 17731
rect 15611 17697 15623 17731
rect 15565 17691 15623 17697
rect 16209 17731 16267 17737
rect 16209 17697 16221 17731
rect 16255 17728 16267 17731
rect 16758 17728 16764 17740
rect 16255 17700 16764 17728
rect 16255 17697 16267 17700
rect 16209 17691 16267 17697
rect 14553 17663 14611 17669
rect 14553 17660 14565 17663
rect 14200 17632 14565 17660
rect 14553 17629 14565 17632
rect 14599 17629 14611 17663
rect 14553 17623 14611 17629
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 13538 17592 13544 17604
rect 12452 17564 12664 17592
rect 13188 17564 13544 17592
rect 10198 17555 10256 17561
rect 2958 17524 2964 17536
rect 2919 17496 2964 17524
rect 2958 17484 2964 17496
rect 3016 17484 3022 17536
rect 5074 17524 5080 17536
rect 5035 17496 5080 17524
rect 5074 17484 5080 17496
rect 5132 17484 5138 17536
rect 8754 17484 8760 17536
rect 8812 17524 8818 17536
rect 9214 17524 9220 17536
rect 8812 17496 9220 17524
rect 8812 17484 8818 17496
rect 9214 17484 9220 17496
rect 9272 17484 9278 17536
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 12636 17524 12664 17564
rect 13538 17552 13544 17564
rect 13596 17552 13602 17604
rect 14737 17527 14795 17533
rect 14737 17524 14749 17527
rect 12636 17496 14749 17524
rect 14737 17493 14749 17496
rect 14783 17493 14795 17527
rect 15304 17524 15332 17623
rect 15580 17592 15608 17691
rect 16758 17688 16764 17700
rect 16816 17688 16822 17740
rect 19245 17731 19303 17737
rect 19245 17697 19257 17731
rect 19291 17728 19303 17731
rect 19334 17728 19340 17740
rect 19291 17700 19340 17728
rect 19291 17697 19303 17700
rect 19245 17691 19303 17697
rect 19334 17688 19340 17700
rect 19392 17688 19398 17740
rect 16298 17620 16304 17672
rect 16356 17660 16362 17672
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 16356 17632 16405 17660
rect 16356 17620 16362 17632
rect 16393 17629 16405 17632
rect 16439 17629 16451 17663
rect 17862 17660 17868 17672
rect 17823 17632 17868 17660
rect 16393 17623 16451 17629
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 18138 17660 18144 17672
rect 18099 17632 18144 17660
rect 18138 17620 18144 17632
rect 18196 17620 18202 17672
rect 19444 17669 19472 17768
rect 19518 17756 19524 17768
rect 19576 17796 19582 17808
rect 21821 17799 21879 17805
rect 21821 17796 21833 17799
rect 19576 17768 21833 17796
rect 19576 17756 19582 17768
rect 21821 17765 21833 17768
rect 21867 17765 21879 17799
rect 21821 17759 21879 17765
rect 19536 17700 19932 17728
rect 19536 17669 19564 17700
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17629 18751 17663
rect 18693 17623 18751 17629
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 19521 17663 19579 17669
rect 19521 17629 19533 17663
rect 19567 17629 19579 17663
rect 19521 17623 19579 17629
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 17034 17592 17040 17604
rect 15580 17564 17040 17592
rect 17034 17552 17040 17564
rect 17092 17552 17098 17604
rect 18708 17592 18736 17623
rect 19536 17592 19564 17623
rect 18708 17564 19564 17592
rect 16301 17527 16359 17533
rect 16301 17524 16313 17527
rect 15304 17496 16313 17524
rect 14737 17487 14795 17493
rect 16301 17493 16313 17496
rect 16347 17524 16359 17527
rect 16666 17524 16672 17536
rect 16347 17496 16672 17524
rect 16347 17493 16359 17496
rect 16301 17487 16359 17493
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 19812 17524 19840 17623
rect 19904 17592 19932 17700
rect 20162 17688 20168 17740
rect 20220 17728 20226 17740
rect 20220 17700 20484 17728
rect 20220 17688 20226 17700
rect 19978 17620 19984 17672
rect 20036 17660 20042 17672
rect 20456 17669 20484 17700
rect 20257 17663 20315 17669
rect 20257 17660 20269 17663
rect 20036 17632 20269 17660
rect 20036 17620 20042 17632
rect 20257 17629 20269 17632
rect 20303 17629 20315 17663
rect 20257 17623 20315 17629
rect 20441 17663 20499 17669
rect 20441 17629 20453 17663
rect 20487 17629 20499 17663
rect 20441 17623 20499 17629
rect 20622 17620 20628 17672
rect 20680 17660 20686 17672
rect 21085 17663 21143 17669
rect 21085 17660 21097 17663
rect 20680 17632 21097 17660
rect 20680 17620 20686 17632
rect 21085 17629 21097 17632
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 21266 17620 21272 17672
rect 21324 17660 21330 17672
rect 21729 17663 21787 17669
rect 21729 17660 21741 17663
rect 21324 17632 21741 17660
rect 21324 17620 21330 17632
rect 21729 17629 21741 17632
rect 21775 17629 21787 17663
rect 21729 17623 21787 17629
rect 21177 17595 21235 17601
rect 21177 17592 21189 17595
rect 19904 17564 21189 17592
rect 21177 17561 21189 17564
rect 21223 17561 21235 17595
rect 21177 17555 21235 17561
rect 21266 17524 21272 17536
rect 19812 17496 21272 17524
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 1104 17434 30820 17456
rect 1104 17382 10880 17434
rect 10932 17382 10944 17434
rect 10996 17382 11008 17434
rect 11060 17382 11072 17434
rect 11124 17382 11136 17434
rect 11188 17382 20811 17434
rect 20863 17382 20875 17434
rect 20927 17382 20939 17434
rect 20991 17382 21003 17434
rect 21055 17382 21067 17434
rect 21119 17382 30820 17434
rect 1104 17360 30820 17382
rect 7466 17320 7472 17332
rect 7427 17292 7472 17320
rect 7466 17280 7472 17292
rect 7524 17280 7530 17332
rect 9122 17320 9128 17332
rect 9083 17292 9128 17320
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 9398 17280 9404 17332
rect 9456 17320 9462 17332
rect 9582 17320 9588 17332
rect 9456 17292 9588 17320
rect 9456 17280 9462 17292
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 13262 17280 13268 17332
rect 13320 17320 13326 17332
rect 13722 17320 13728 17332
rect 13320 17292 13728 17320
rect 13320 17280 13326 17292
rect 13722 17280 13728 17292
rect 13780 17280 13786 17332
rect 14550 17280 14556 17332
rect 14608 17320 14614 17332
rect 14829 17323 14887 17329
rect 14829 17320 14841 17323
rect 14608 17292 14841 17320
rect 14608 17280 14614 17292
rect 14829 17289 14841 17292
rect 14875 17320 14887 17323
rect 15194 17320 15200 17332
rect 14875 17292 15200 17320
rect 14875 17289 14887 17292
rect 14829 17283 14887 17289
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 16942 17320 16948 17332
rect 16903 17292 16948 17320
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 19242 17280 19248 17332
rect 19300 17280 19306 17332
rect 20162 17280 20168 17332
rect 20220 17320 20226 17332
rect 20441 17323 20499 17329
rect 20441 17320 20453 17323
rect 20220 17292 20453 17320
rect 20220 17280 20226 17292
rect 20441 17289 20453 17292
rect 20487 17289 20499 17323
rect 20441 17283 20499 17289
rect 21818 17280 21824 17332
rect 21876 17320 21882 17332
rect 21913 17323 21971 17329
rect 21913 17320 21925 17323
rect 21876 17292 21925 17320
rect 21876 17280 21882 17292
rect 21913 17289 21925 17292
rect 21959 17289 21971 17323
rect 21913 17283 21971 17289
rect 8754 17252 8760 17264
rect 8588 17224 8760 17252
rect 1394 17184 1400 17196
rect 1355 17156 1400 17184
rect 1394 17144 1400 17156
rect 1452 17144 1458 17196
rect 2590 17184 2596 17196
rect 2551 17156 2596 17184
rect 2590 17144 2596 17156
rect 2648 17144 2654 17196
rect 4148 17187 4206 17193
rect 4148 17153 4160 17187
rect 4194 17184 4206 17187
rect 4522 17184 4528 17196
rect 4194 17156 4528 17184
rect 4194 17153 4206 17156
rect 4148 17147 4206 17153
rect 4522 17144 4528 17156
rect 4580 17144 4586 17196
rect 6730 17184 6736 17196
rect 6691 17156 6736 17184
rect 6730 17144 6736 17156
rect 6788 17144 6794 17196
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17184 6975 17187
rect 7190 17184 7196 17196
rect 6963 17156 7196 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 7926 17184 7932 17196
rect 7331 17156 7932 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 8386 17184 8392 17196
rect 8347 17156 8392 17184
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 8588 17193 8616 17224
rect 8754 17212 8760 17224
rect 8812 17212 8818 17264
rect 11238 17252 11244 17264
rect 8956 17224 11244 17252
rect 8573 17187 8631 17193
rect 8573 17153 8585 17187
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 8665 17187 8723 17193
rect 8665 17153 8677 17187
rect 8711 17184 8723 17187
rect 8846 17184 8852 17196
rect 8711 17156 8852 17184
rect 8711 17153 8723 17156
rect 8665 17147 8723 17153
rect 8846 17144 8852 17156
rect 8904 17144 8910 17196
rect 8956 17193 8984 17224
rect 11238 17212 11244 17224
rect 11296 17212 11302 17264
rect 11968 17255 12026 17261
rect 11968 17221 11980 17255
rect 12014 17252 12026 17255
rect 12526 17252 12532 17264
rect 12014 17224 12532 17252
rect 12014 17221 12026 17224
rect 11968 17215 12026 17221
rect 12526 17212 12532 17224
rect 12584 17212 12590 17264
rect 13906 17212 13912 17264
rect 13964 17252 13970 17264
rect 14185 17255 14243 17261
rect 13964 17224 14136 17252
rect 13964 17212 13970 17224
rect 8941 17187 8999 17193
rect 8941 17153 8953 17187
rect 8987 17153 8999 17187
rect 8941 17147 8999 17153
rect 10709 17187 10767 17193
rect 10709 17153 10721 17187
rect 10755 17184 10767 17187
rect 10870 17184 10876 17196
rect 10755 17156 10876 17184
rect 10755 17153 10767 17156
rect 10709 17147 10767 17153
rect 10870 17144 10876 17156
rect 10928 17144 10934 17196
rect 13998 17184 14004 17196
rect 13959 17156 14004 17184
rect 13998 17144 14004 17156
rect 14056 17144 14062 17196
rect 14108 17184 14136 17224
rect 14185 17221 14197 17255
rect 14231 17252 14243 17255
rect 15286 17252 15292 17264
rect 14231 17224 15292 17252
rect 14231 17221 14243 17224
rect 14185 17215 14243 17221
rect 15286 17212 15292 17224
rect 15344 17212 15350 17264
rect 17218 17252 17224 17264
rect 16960 17224 17224 17252
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 14108 17156 14749 17184
rect 14737 17153 14749 17156
rect 14783 17184 14795 17187
rect 16960 17184 16988 17224
rect 17218 17212 17224 17224
rect 17276 17212 17282 17264
rect 17589 17255 17647 17261
rect 17589 17221 17601 17255
rect 17635 17252 17647 17255
rect 17862 17252 17868 17264
rect 17635 17224 17868 17252
rect 17635 17221 17647 17224
rect 17589 17215 17647 17221
rect 17862 17212 17868 17224
rect 17920 17252 17926 17264
rect 18417 17255 18475 17261
rect 18417 17252 18429 17255
rect 17920 17224 18429 17252
rect 17920 17212 17926 17224
rect 18417 17221 18429 17224
rect 18463 17221 18475 17255
rect 19260 17252 19288 17280
rect 19334 17252 19340 17264
rect 19260 17224 19340 17252
rect 18417 17215 18475 17221
rect 19334 17212 19340 17224
rect 19392 17212 19398 17264
rect 19560 17224 20024 17252
rect 14783 17156 16988 17184
rect 14783 17153 14795 17156
rect 14737 17147 14795 17153
rect 17034 17144 17040 17196
rect 17092 17184 17098 17196
rect 17129 17187 17187 17193
rect 17129 17184 17141 17187
rect 17092 17156 17141 17184
rect 17092 17144 17098 17156
rect 17129 17153 17141 17156
rect 17175 17184 17187 17187
rect 17770 17184 17776 17196
rect 17175 17156 17776 17184
rect 17175 17153 17187 17156
rect 17129 17147 17187 17153
rect 17770 17144 17776 17156
rect 17828 17184 17834 17196
rect 18049 17187 18107 17193
rect 18049 17184 18061 17187
rect 17828 17156 18061 17184
rect 17828 17144 17834 17156
rect 18049 17153 18061 17156
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 18233 17187 18291 17193
rect 18233 17153 18245 17187
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 3234 17116 3240 17128
rect 2915 17088 3240 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 3234 17076 3240 17088
rect 3292 17076 3298 17128
rect 3694 17076 3700 17128
rect 3752 17116 3758 17128
rect 3878 17116 3884 17128
rect 3752 17088 3884 17116
rect 3752 17076 3758 17088
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17085 7067 17119
rect 7009 17079 7067 17085
rect 7101 17119 7159 17125
rect 7101 17085 7113 17119
rect 7147 17116 7159 17119
rect 8754 17116 8760 17128
rect 7147 17088 8760 17116
rect 7147 17085 7159 17088
rect 7101 17079 7159 17085
rect 7024 17048 7052 17079
rect 8754 17076 8760 17088
rect 8812 17076 8818 17128
rect 8864 17116 8892 17144
rect 9030 17116 9036 17128
rect 8864 17088 9036 17116
rect 8864 17048 8892 17088
rect 9030 17076 9036 17088
rect 9088 17076 9094 17128
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17116 11023 17119
rect 11698 17116 11704 17128
rect 11011 17088 11704 17116
rect 11011 17085 11023 17088
rect 10965 17079 11023 17085
rect 11698 17076 11704 17088
rect 11756 17076 11762 17128
rect 13817 17119 13875 17125
rect 13817 17085 13829 17119
rect 13863 17116 13875 17119
rect 14182 17116 14188 17128
rect 13863 17088 14188 17116
rect 13863 17085 13875 17088
rect 13817 17079 13875 17085
rect 14182 17076 14188 17088
rect 14240 17076 14246 17128
rect 17218 17076 17224 17128
rect 17276 17116 17282 17128
rect 18248 17116 18276 17147
rect 18598 17144 18604 17196
rect 18656 17184 18662 17196
rect 19245 17187 19303 17193
rect 19245 17184 19257 17187
rect 18656 17156 19257 17184
rect 18656 17144 18662 17156
rect 19245 17153 19257 17156
rect 19291 17153 19303 17187
rect 19245 17147 19303 17153
rect 19429 17187 19487 17193
rect 19429 17153 19441 17187
rect 19475 17184 19487 17187
rect 19560 17184 19588 17224
rect 19475 17156 19588 17184
rect 19659 17187 19717 17193
rect 19475 17153 19487 17156
rect 19429 17147 19487 17153
rect 19659 17153 19671 17187
rect 19705 17184 19717 17187
rect 19797 17187 19855 17193
rect 19705 17153 19739 17184
rect 19659 17147 19739 17153
rect 19797 17153 19809 17187
rect 19843 17184 19855 17187
rect 19843 17156 19932 17184
rect 19843 17153 19855 17156
rect 19797 17147 19855 17153
rect 18506 17116 18512 17128
rect 17276 17088 18512 17116
rect 17276 17076 17282 17088
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 19521 17119 19579 17125
rect 19392 17108 19481 17116
rect 19521 17108 19533 17119
rect 19392 17088 19533 17108
rect 19392 17076 19398 17088
rect 19453 17085 19533 17088
rect 19567 17085 19579 17119
rect 19453 17080 19579 17085
rect 19521 17079 19579 17080
rect 7024 17020 8892 17048
rect 19150 17008 19156 17060
rect 19208 17048 19214 17060
rect 19711 17048 19739 17147
rect 19208 17020 19739 17048
rect 19208 17008 19214 17020
rect 19794 17008 19800 17060
rect 19852 17048 19858 17060
rect 19904 17048 19932 17156
rect 19996 17116 20024 17224
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17184 20775 17187
rect 21266 17184 21272 17196
rect 20763 17156 21272 17184
rect 20763 17153 20775 17156
rect 20717 17147 20775 17153
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 21818 17184 21824 17196
rect 21779 17156 21824 17184
rect 21818 17144 21824 17156
rect 21876 17144 21882 17196
rect 29825 17187 29883 17193
rect 29825 17153 29837 17187
rect 29871 17184 29883 17187
rect 29914 17184 29920 17196
rect 29871 17156 29920 17184
rect 29871 17153 29883 17156
rect 29825 17147 29883 17153
rect 29914 17144 29920 17156
rect 29972 17144 29978 17196
rect 20346 17116 20352 17128
rect 19996 17088 20352 17116
rect 20346 17076 20352 17088
rect 20404 17116 20410 17128
rect 20441 17119 20499 17125
rect 20441 17116 20453 17119
rect 20404 17088 20453 17116
rect 20404 17076 20410 17088
rect 20441 17085 20453 17088
rect 20487 17085 20499 17119
rect 20622 17116 20628 17128
rect 20583 17088 20628 17116
rect 20441 17079 20499 17085
rect 20622 17076 20628 17088
rect 20680 17076 20686 17128
rect 19852 17020 19932 17048
rect 19852 17008 19858 17020
rect 1581 16983 1639 16989
rect 1581 16949 1593 16983
rect 1627 16980 1639 16983
rect 2314 16980 2320 16992
rect 1627 16952 2320 16980
rect 1627 16949 1639 16952
rect 1581 16943 1639 16949
rect 2314 16940 2320 16952
rect 2372 16940 2378 16992
rect 4982 16940 4988 16992
rect 5040 16980 5046 16992
rect 5261 16983 5319 16989
rect 5261 16980 5273 16983
rect 5040 16952 5273 16980
rect 5040 16940 5046 16952
rect 5261 16949 5273 16952
rect 5307 16949 5319 16983
rect 5261 16943 5319 16949
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 13081 16983 13139 16989
rect 13081 16980 13093 16983
rect 12860 16952 13093 16980
rect 12860 16940 12866 16952
rect 13081 16949 13093 16952
rect 13127 16949 13139 16983
rect 13081 16943 13139 16949
rect 13722 16940 13728 16992
rect 13780 16980 13786 16992
rect 15102 16980 15108 16992
rect 13780 16952 15108 16980
rect 13780 16940 13786 16952
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 19981 16983 20039 16989
rect 19981 16949 19993 16983
rect 20027 16980 20039 16983
rect 20438 16980 20444 16992
rect 20027 16952 20444 16980
rect 20027 16949 20039 16952
rect 19981 16943 20039 16949
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 30006 16980 30012 16992
rect 29967 16952 30012 16980
rect 30006 16940 30012 16952
rect 30064 16940 30070 16992
rect 1104 16890 30820 16912
rect 1104 16838 5915 16890
rect 5967 16838 5979 16890
rect 6031 16838 6043 16890
rect 6095 16838 6107 16890
rect 6159 16838 6171 16890
rect 6223 16838 15846 16890
rect 15898 16838 15910 16890
rect 15962 16838 15974 16890
rect 16026 16838 16038 16890
rect 16090 16838 16102 16890
rect 16154 16838 25776 16890
rect 25828 16838 25840 16890
rect 25892 16838 25904 16890
rect 25956 16838 25968 16890
rect 26020 16838 26032 16890
rect 26084 16838 30820 16890
rect 1104 16816 30820 16838
rect 2958 16736 2964 16788
rect 3016 16776 3022 16788
rect 3016 16748 6224 16776
rect 3016 16736 3022 16748
rect 3694 16600 3700 16652
rect 3752 16640 3758 16652
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 3752 16612 4353 16640
rect 3752 16600 3758 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 1210 16532 1216 16584
rect 1268 16572 1274 16584
rect 1397 16575 1455 16581
rect 1397 16572 1409 16575
rect 1268 16544 1409 16572
rect 1268 16532 1274 16544
rect 1397 16541 1409 16544
rect 1443 16541 1455 16575
rect 1397 16535 1455 16541
rect 2866 16532 2872 16584
rect 2924 16572 2930 16584
rect 2961 16575 3019 16581
rect 2961 16572 2973 16575
rect 2924 16544 2973 16572
rect 2924 16532 2930 16544
rect 2961 16541 2973 16544
rect 3007 16541 3019 16575
rect 3234 16572 3240 16584
rect 3195 16544 3240 16572
rect 2961 16535 3019 16541
rect 3234 16532 3240 16544
rect 3292 16532 3298 16584
rect 3418 16532 3424 16584
rect 3476 16572 3482 16584
rect 3970 16572 3976 16584
rect 3476 16544 3976 16572
rect 3476 16532 3482 16544
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 6196 16581 6224 16748
rect 10870 16736 10876 16788
rect 10928 16776 10934 16788
rect 10965 16779 11023 16785
rect 10965 16776 10977 16779
rect 10928 16748 10977 16776
rect 10928 16736 10934 16748
rect 10965 16745 10977 16748
rect 11011 16745 11023 16779
rect 10965 16739 11023 16745
rect 13265 16779 13323 16785
rect 13265 16745 13277 16779
rect 13311 16776 13323 16779
rect 14093 16779 14151 16785
rect 13311 16748 13492 16776
rect 13311 16745 13323 16748
rect 13265 16739 13323 16745
rect 13464 16720 13492 16748
rect 14093 16745 14105 16779
rect 14139 16776 14151 16779
rect 14458 16776 14464 16788
rect 14139 16748 14464 16776
rect 14139 16745 14151 16748
rect 14093 16739 14151 16745
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 17218 16776 17224 16788
rect 17179 16748 17224 16776
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 20346 16736 20352 16788
rect 20404 16776 20410 16788
rect 21729 16779 21787 16785
rect 21729 16776 21741 16779
rect 20404 16748 21741 16776
rect 20404 16736 20410 16748
rect 21729 16745 21741 16748
rect 21775 16776 21787 16779
rect 21818 16776 21824 16788
rect 21775 16748 21824 16776
rect 21775 16745 21787 16748
rect 21729 16739 21787 16745
rect 21818 16736 21824 16748
rect 21876 16736 21882 16788
rect 8846 16668 8852 16720
rect 8904 16708 8910 16720
rect 13354 16708 13360 16720
rect 8904 16680 10548 16708
rect 8904 16668 8910 16680
rect 8754 16600 8760 16652
rect 8812 16640 8818 16652
rect 9306 16640 9312 16652
rect 8812 16612 9312 16640
rect 8812 16600 8818 16612
rect 9306 16600 9312 16612
rect 9364 16640 9370 16652
rect 10520 16649 10548 16680
rect 13188 16680 13360 16708
rect 13188 16649 13216 16680
rect 13354 16668 13360 16680
rect 13412 16668 13418 16720
rect 13446 16668 13452 16720
rect 13504 16708 13510 16720
rect 14369 16711 14427 16717
rect 14369 16708 14381 16711
rect 13504 16680 14381 16708
rect 13504 16668 13510 16680
rect 14369 16677 14381 16680
rect 14415 16677 14427 16711
rect 15102 16708 15108 16720
rect 15063 16680 15108 16708
rect 14369 16671 14427 16677
rect 15102 16668 15108 16680
rect 15160 16708 15166 16720
rect 19978 16708 19984 16720
rect 15160 16680 19984 16708
rect 15160 16668 15166 16680
rect 19978 16668 19984 16680
rect 20036 16668 20042 16720
rect 9493 16643 9551 16649
rect 9493 16640 9505 16643
rect 9364 16612 9505 16640
rect 9364 16600 9370 16612
rect 9493 16609 9505 16612
rect 9539 16640 9551 16643
rect 10505 16643 10563 16649
rect 9539 16612 9904 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 6181 16575 6239 16581
rect 6181 16541 6193 16575
rect 6227 16541 6239 16575
rect 6181 16535 6239 16541
rect 6825 16575 6883 16581
rect 6825 16541 6837 16575
rect 6871 16541 6883 16575
rect 6825 16535 6883 16541
rect 9769 16575 9827 16581
rect 9769 16541 9781 16575
rect 9815 16541 9827 16575
rect 9769 16535 9827 16541
rect 4246 16464 4252 16516
rect 4304 16504 4310 16516
rect 4586 16507 4644 16513
rect 4586 16504 4598 16507
rect 4304 16476 4598 16504
rect 4304 16464 4310 16476
rect 4586 16473 4598 16476
rect 4632 16473 4644 16507
rect 6840 16504 6868 16535
rect 4586 16467 4644 16473
rect 5736 16476 6868 16504
rect 5736 16448 5764 16476
rect 9398 16464 9404 16516
rect 9456 16504 9462 16516
rect 9784 16504 9812 16535
rect 9456 16476 9812 16504
rect 9876 16504 9904 16612
rect 10505 16609 10517 16643
rect 10551 16609 10563 16643
rect 10505 16603 10563 16609
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16609 13231 16643
rect 14461 16643 14519 16649
rect 14461 16640 14473 16643
rect 13173 16603 13231 16609
rect 13409 16612 14473 16640
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10229 16575 10287 16581
rect 10229 16572 10241 16575
rect 10192 16544 10241 16572
rect 10192 16532 10198 16544
rect 10229 16541 10241 16544
rect 10275 16541 10287 16575
rect 10410 16572 10416 16584
rect 10371 16544 10416 16572
rect 10229 16535 10287 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16541 10655 16575
rect 10597 16535 10655 16541
rect 10781 16575 10839 16581
rect 10781 16541 10793 16575
rect 10827 16541 10839 16575
rect 11974 16572 11980 16584
rect 11935 16544 11980 16572
rect 10781 16535 10839 16541
rect 10612 16504 10640 16535
rect 9876 16476 10640 16504
rect 9456 16464 9462 16476
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16436 1639 16439
rect 2682 16436 2688 16448
rect 1627 16408 2688 16436
rect 1627 16405 1639 16408
rect 1581 16399 1639 16405
rect 2682 16396 2688 16408
rect 2740 16396 2746 16448
rect 5718 16436 5724 16448
rect 5679 16408 5724 16436
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 6270 16436 6276 16448
rect 6231 16408 6276 16436
rect 6270 16396 6276 16408
rect 6328 16396 6334 16448
rect 6917 16439 6975 16445
rect 6917 16405 6929 16439
rect 6963 16436 6975 16439
rect 7742 16436 7748 16448
rect 6963 16408 7748 16436
rect 6963 16405 6975 16408
rect 6917 16399 6975 16405
rect 7742 16396 7748 16408
rect 7800 16396 7806 16448
rect 9582 16396 9588 16448
rect 9640 16436 9646 16448
rect 10796 16436 10824 16535
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 12802 16532 12808 16584
rect 12860 16572 12866 16584
rect 13409 16581 13437 16612
rect 14461 16609 14473 16612
rect 14507 16609 14519 16643
rect 14461 16603 14519 16609
rect 16942 16600 16948 16652
rect 17000 16640 17006 16652
rect 19610 16640 19616 16652
rect 17000 16612 17264 16640
rect 17000 16600 17006 16612
rect 13394 16575 13452 16581
rect 13394 16574 13406 16575
rect 13280 16572 13406 16574
rect 12860 16546 13406 16572
rect 12860 16544 13308 16546
rect 12860 16532 12866 16544
rect 13394 16541 13406 16546
rect 13440 16541 13452 16575
rect 13394 16535 13452 16541
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16572 13599 16575
rect 13906 16572 13912 16584
rect 13587 16544 13912 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 13906 16532 13912 16544
rect 13964 16532 13970 16584
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16541 14335 16575
rect 14550 16572 14556 16584
rect 14511 16544 14556 16572
rect 14277 16535 14335 16541
rect 12345 16507 12403 16513
rect 12345 16473 12357 16507
rect 12391 16504 12403 16507
rect 13078 16504 13084 16516
rect 12391 16476 13084 16504
rect 12391 16473 12403 16476
rect 12345 16467 12403 16473
rect 13078 16464 13084 16476
rect 13136 16464 13142 16516
rect 14292 16504 14320 16535
rect 14550 16532 14556 16544
rect 14608 16532 14614 16584
rect 15286 16572 15292 16584
rect 15247 16544 15292 16572
rect 15286 16532 15292 16544
rect 15344 16572 15350 16584
rect 16209 16575 16267 16581
rect 16209 16572 16221 16575
rect 15344 16544 16221 16572
rect 15344 16532 15350 16544
rect 16209 16541 16221 16544
rect 16255 16541 16267 16575
rect 16209 16535 16267 16541
rect 16393 16575 16451 16581
rect 16393 16541 16405 16575
rect 16439 16572 16451 16575
rect 16758 16572 16764 16584
rect 16439 16544 16764 16572
rect 16439 16541 16451 16544
rect 16393 16535 16451 16541
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 17034 16572 17040 16584
rect 16995 16544 17040 16572
rect 17034 16532 17040 16544
rect 17092 16532 17098 16584
rect 17236 16581 17264 16612
rect 19444 16612 19616 16640
rect 17221 16575 17279 16581
rect 17221 16541 17233 16575
rect 17267 16572 17279 16575
rect 18138 16572 18144 16584
rect 17267 16544 18144 16572
rect 17267 16541 17279 16544
rect 17221 16535 17279 16541
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 19444 16581 19472 16612
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 19518 16532 19524 16584
rect 19576 16572 19582 16584
rect 20349 16575 20407 16581
rect 20349 16572 20361 16575
rect 19576 16544 20361 16572
rect 19576 16532 19582 16544
rect 20349 16541 20361 16544
rect 20395 16541 20407 16575
rect 20349 16535 20407 16541
rect 20438 16532 20444 16584
rect 20496 16572 20502 16584
rect 20605 16575 20663 16581
rect 20605 16572 20617 16575
rect 20496 16544 20617 16572
rect 20496 16532 20502 16544
rect 20605 16541 20617 16544
rect 20651 16541 20663 16575
rect 20605 16535 20663 16541
rect 13372 16476 14320 16504
rect 16577 16507 16635 16513
rect 13372 16448 13400 16476
rect 16577 16473 16589 16507
rect 16623 16504 16635 16507
rect 19242 16504 19248 16516
rect 16623 16476 19248 16504
rect 16623 16473 16635 16476
rect 16577 16467 16635 16473
rect 9640 16408 10824 16436
rect 9640 16396 9646 16408
rect 11238 16396 11244 16448
rect 11296 16436 11302 16448
rect 12897 16439 12955 16445
rect 12897 16436 12909 16439
rect 11296 16408 12909 16436
rect 11296 16396 11302 16408
rect 12897 16405 12909 16408
rect 12943 16405 12955 16439
rect 12897 16399 12955 16405
rect 13354 16396 13360 16448
rect 13412 16396 13418 16448
rect 16298 16396 16304 16448
rect 16356 16436 16362 16448
rect 16850 16436 16856 16448
rect 16356 16408 16856 16436
rect 16356 16396 16362 16408
rect 16850 16396 16856 16408
rect 16908 16396 16914 16448
rect 17420 16445 17448 16476
rect 19242 16464 19248 16476
rect 19300 16464 19306 16516
rect 17405 16439 17463 16445
rect 17405 16405 17417 16439
rect 17451 16405 17463 16439
rect 17405 16399 17463 16405
rect 18598 16396 18604 16448
rect 18656 16436 18662 16448
rect 19337 16439 19395 16445
rect 19337 16436 19349 16439
rect 18656 16408 19349 16436
rect 18656 16396 18662 16408
rect 19337 16405 19349 16408
rect 19383 16405 19395 16439
rect 19337 16399 19395 16405
rect 1104 16346 30820 16368
rect 1104 16294 10880 16346
rect 10932 16294 10944 16346
rect 10996 16294 11008 16346
rect 11060 16294 11072 16346
rect 11124 16294 11136 16346
rect 11188 16294 20811 16346
rect 20863 16294 20875 16346
rect 20927 16294 20939 16346
rect 20991 16294 21003 16346
rect 21055 16294 21067 16346
rect 21119 16294 30820 16346
rect 1104 16272 30820 16294
rect 3786 16232 3792 16244
rect 3620 16204 3792 16232
rect 1762 16056 1768 16108
rect 1820 16096 1826 16108
rect 1929 16099 1987 16105
rect 1929 16096 1941 16099
rect 1820 16068 1941 16096
rect 1820 16056 1826 16068
rect 1929 16065 1941 16068
rect 1975 16065 1987 16099
rect 1929 16059 1987 16065
rect 3513 16099 3571 16105
rect 3513 16065 3525 16099
rect 3559 16096 3571 16099
rect 3620 16096 3648 16204
rect 3786 16192 3792 16204
rect 3844 16232 3850 16244
rect 4062 16232 4068 16244
rect 3844 16204 4068 16232
rect 3844 16192 3850 16204
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 4246 16232 4252 16244
rect 4207 16204 4252 16232
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 5166 16192 5172 16244
rect 5224 16232 5230 16244
rect 7190 16232 7196 16244
rect 5224 16204 6408 16232
rect 7151 16204 7196 16232
rect 5224 16192 5230 16204
rect 5074 16164 5080 16176
rect 3712 16136 5080 16164
rect 3712 16105 3740 16136
rect 5074 16124 5080 16136
rect 5132 16124 5138 16176
rect 3559 16068 3648 16096
rect 3697 16099 3755 16105
rect 3559 16065 3571 16068
rect 3513 16059 3571 16065
rect 3697 16065 3709 16099
rect 3743 16065 3755 16099
rect 3697 16059 3755 16065
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16065 4123 16099
rect 4982 16096 4988 16108
rect 4943 16068 4988 16096
rect 4065 16059 4123 16065
rect 1670 16028 1676 16040
rect 1631 16000 1676 16028
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 2866 15988 2872 16040
rect 2924 16028 2930 16040
rect 3789 16031 3847 16037
rect 3789 16028 3801 16031
rect 2924 16000 3801 16028
rect 2924 15988 2930 16000
rect 3789 15997 3801 16000
rect 3835 15997 3847 16031
rect 3789 15991 3847 15997
rect 3878 15988 3884 16040
rect 3936 16028 3942 16040
rect 4080 16028 4108 16059
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 6380 16105 6408 16204
rect 7190 16192 7196 16204
rect 7248 16192 7254 16244
rect 9582 16192 9588 16244
rect 9640 16232 9646 16244
rect 10965 16235 11023 16241
rect 10965 16232 10977 16235
rect 9640 16204 10977 16232
rect 9640 16192 9646 16204
rect 10965 16201 10977 16204
rect 11011 16232 11023 16235
rect 11422 16232 11428 16244
rect 11011 16204 11428 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 13725 16235 13783 16241
rect 13725 16201 13737 16235
rect 13771 16232 13783 16235
rect 13998 16232 14004 16244
rect 13771 16204 14004 16232
rect 13771 16201 13783 16204
rect 13725 16195 13783 16201
rect 13998 16192 14004 16204
rect 14056 16192 14062 16244
rect 18138 16192 18144 16244
rect 18196 16232 18202 16244
rect 18325 16235 18383 16241
rect 18325 16232 18337 16235
rect 18196 16204 18337 16232
rect 18196 16192 18202 16204
rect 18325 16201 18337 16204
rect 18371 16201 18383 16235
rect 18325 16195 18383 16201
rect 19058 16192 19064 16244
rect 19116 16232 19122 16244
rect 19116 16204 19656 16232
rect 19116 16192 19122 16204
rect 7101 16167 7159 16173
rect 7101 16133 7113 16167
rect 7147 16164 7159 16167
rect 7466 16164 7472 16176
rect 7147 16136 7472 16164
rect 7147 16133 7159 16136
rect 7101 16127 7159 16133
rect 7466 16124 7472 16136
rect 7524 16164 7530 16176
rect 11238 16164 11244 16176
rect 7524 16136 11244 16164
rect 7524 16124 7530 16136
rect 11238 16124 11244 16136
rect 11296 16124 11302 16176
rect 12713 16167 12771 16173
rect 12713 16133 12725 16167
rect 12759 16164 12771 16167
rect 19518 16164 19524 16176
rect 12759 16136 13584 16164
rect 12759 16133 12771 16136
rect 12713 16127 12771 16133
rect 5629 16099 5687 16105
rect 5629 16065 5641 16099
rect 5675 16096 5687 16099
rect 6365 16099 6423 16105
rect 5675 16068 5856 16096
rect 5675 16065 5687 16068
rect 5629 16059 5687 16065
rect 5718 16028 5724 16040
rect 3936 16000 3981 16028
rect 4080 16000 5724 16028
rect 3936 15988 3942 16000
rect 5718 15988 5724 16000
rect 5776 15988 5782 16040
rect 3053 15963 3111 15969
rect 3053 15960 3065 15963
rect 2746 15932 3065 15960
rect 1946 15852 1952 15904
rect 2004 15892 2010 15904
rect 2746 15892 2774 15932
rect 3053 15929 3065 15932
rect 3099 15960 3111 15963
rect 5828 15960 5856 16068
rect 6365 16065 6377 16099
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 8110 16056 8116 16108
rect 8168 16096 8174 16108
rect 9033 16099 9091 16105
rect 9033 16096 9045 16099
rect 8168 16068 9045 16096
rect 8168 16056 8174 16068
rect 9033 16065 9045 16068
rect 9079 16065 9091 16099
rect 9033 16059 9091 16065
rect 9585 16099 9643 16105
rect 9585 16065 9597 16099
rect 9631 16096 9643 16099
rect 9674 16096 9680 16108
rect 9631 16068 9680 16096
rect 9631 16065 9643 16068
rect 9585 16059 9643 16065
rect 9674 16056 9680 16068
rect 9732 16056 9738 16108
rect 9858 16105 9864 16108
rect 9852 16059 9864 16105
rect 9916 16096 9922 16108
rect 12802 16096 12808 16108
rect 9916 16068 9952 16096
rect 12763 16068 12808 16096
rect 9858 16056 9864 16059
rect 9916 16056 9922 16068
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 13556 16105 13584 16136
rect 16960 16136 19524 16164
rect 13541 16099 13599 16105
rect 13541 16065 13553 16099
rect 13587 16096 13599 16099
rect 14090 16096 14096 16108
rect 13587 16068 14096 16096
rect 13587 16065 13599 16068
rect 13541 16059 13599 16065
rect 14090 16056 14096 16068
rect 14148 16056 14154 16108
rect 14458 16096 14464 16108
rect 14371 16068 14464 16096
rect 14458 16056 14464 16068
rect 14516 16096 14522 16108
rect 16960 16105 16988 16136
rect 19518 16124 19524 16136
rect 19576 16124 19582 16176
rect 17218 16105 17224 16108
rect 16945 16099 17003 16105
rect 16945 16096 16957 16099
rect 14516 16068 16957 16096
rect 14516 16056 14522 16068
rect 16945 16065 16957 16068
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 17212 16059 17224 16105
rect 17276 16096 17282 16108
rect 17276 16068 17312 16096
rect 17218 16056 17224 16059
rect 17276 16056 17282 16068
rect 18230 16056 18236 16108
rect 18288 16096 18294 16108
rect 18877 16099 18935 16105
rect 18877 16096 18889 16099
rect 18288 16068 18889 16096
rect 18288 16056 18294 16068
rect 18877 16065 18889 16068
rect 18923 16065 18935 16099
rect 19058 16096 19064 16108
rect 19019 16068 19064 16096
rect 18877 16059 18935 16065
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 19242 16096 19248 16108
rect 19203 16068 19248 16096
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 19426 16096 19432 16108
rect 19387 16068 19432 16096
rect 19426 16056 19432 16068
rect 19484 16056 19490 16108
rect 19628 16096 19656 16204
rect 29362 16192 29368 16244
rect 29420 16232 29426 16244
rect 30009 16235 30067 16241
rect 30009 16232 30021 16235
rect 29420 16204 30021 16232
rect 29420 16192 29426 16204
rect 30009 16201 30021 16204
rect 30055 16201 30067 16235
rect 30009 16195 30067 16201
rect 20257 16167 20315 16173
rect 20257 16133 20269 16167
rect 20303 16164 20315 16167
rect 20346 16164 20352 16176
rect 20303 16136 20352 16164
rect 20303 16133 20315 16136
rect 20257 16127 20315 16133
rect 20346 16124 20352 16136
rect 20404 16124 20410 16176
rect 21266 16164 21272 16176
rect 20824 16136 21272 16164
rect 20824 16108 20852 16136
rect 21266 16124 21272 16136
rect 21324 16124 21330 16176
rect 20441 16099 20499 16105
rect 20441 16096 20453 16099
rect 19628 16068 20453 16096
rect 20441 16065 20453 16068
rect 20487 16096 20499 16099
rect 20806 16096 20812 16108
rect 20487 16068 20812 16096
rect 20487 16065 20499 16068
rect 20441 16059 20499 16065
rect 20806 16056 20812 16068
rect 20864 16056 20870 16108
rect 21174 16096 21180 16108
rect 21087 16068 21180 16096
rect 21174 16056 21180 16068
rect 21232 16096 21238 16108
rect 21634 16096 21640 16108
rect 21232 16068 21640 16096
rect 21232 16056 21238 16068
rect 21634 16056 21640 16068
rect 21692 16056 21698 16108
rect 28994 16056 29000 16108
rect 29052 16096 29058 16108
rect 29917 16099 29975 16105
rect 29917 16096 29929 16099
rect 29052 16068 29929 16096
rect 29052 16056 29058 16068
rect 29917 16065 29929 16068
rect 29963 16065 29975 16099
rect 30098 16096 30104 16108
rect 30059 16068 30104 16096
rect 29917 16059 29975 16065
rect 30098 16056 30104 16068
rect 30156 16056 30162 16108
rect 8757 16031 8815 16037
rect 8757 15997 8769 16031
rect 8803 16028 8815 16031
rect 8846 16028 8852 16040
rect 8803 16000 8852 16028
rect 8803 15997 8815 16000
rect 8757 15991 8815 15997
rect 8846 15988 8852 16000
rect 8904 15988 8910 16040
rect 13265 16031 13323 16037
rect 13265 15997 13277 16031
rect 13311 16028 13323 16031
rect 13354 16028 13360 16040
rect 13311 16000 13360 16028
rect 13311 15997 13323 16000
rect 13265 15991 13323 15997
rect 13354 15988 13360 16000
rect 13412 15988 13418 16040
rect 14734 16028 14740 16040
rect 14695 16000 14740 16028
rect 14734 15988 14740 16000
rect 14792 15988 14798 16040
rect 19153 16031 19211 16037
rect 19153 15997 19165 16031
rect 19199 16028 19211 16031
rect 19334 16028 19340 16040
rect 19199 16000 19340 16028
rect 19199 15997 19211 16000
rect 19153 15991 19211 15997
rect 19334 15988 19340 16000
rect 19392 15988 19398 16040
rect 6914 15960 6920 15972
rect 3099 15932 5856 15960
rect 6380 15932 6920 15960
rect 3099 15929 3111 15932
rect 3053 15923 3111 15929
rect 5074 15892 5080 15904
rect 2004 15864 2774 15892
rect 5035 15864 5080 15892
rect 2004 15852 2010 15864
rect 5074 15852 5080 15864
rect 5132 15852 5138 15904
rect 5721 15895 5779 15901
rect 5721 15861 5733 15895
rect 5767 15892 5779 15895
rect 6380 15892 6408 15932
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 20073 15963 20131 15969
rect 20073 15960 20085 15963
rect 19352 15932 20085 15960
rect 5767 15864 6408 15892
rect 6457 15895 6515 15901
rect 5767 15861 5779 15864
rect 5721 15855 5779 15861
rect 6457 15861 6469 15895
rect 6503 15892 6515 15895
rect 7006 15892 7012 15904
rect 6503 15864 7012 15892
rect 6503 15861 6515 15864
rect 6457 15855 6515 15861
rect 7006 15852 7012 15864
rect 7064 15852 7070 15904
rect 7190 15852 7196 15904
rect 7248 15892 7254 15904
rect 10502 15892 10508 15904
rect 7248 15864 10508 15892
rect 7248 15852 7254 15864
rect 10502 15852 10508 15864
rect 10560 15852 10566 15904
rect 13262 15852 13268 15904
rect 13320 15892 13326 15904
rect 13357 15895 13415 15901
rect 13357 15892 13369 15895
rect 13320 15864 13369 15892
rect 13320 15852 13326 15864
rect 13357 15861 13369 15864
rect 13403 15892 13415 15895
rect 13446 15892 13452 15904
rect 13403 15864 13452 15892
rect 13403 15861 13415 15864
rect 13357 15855 13415 15861
rect 13446 15852 13452 15864
rect 13504 15852 13510 15904
rect 15102 15852 15108 15904
rect 15160 15892 15166 15904
rect 15841 15895 15899 15901
rect 15841 15892 15853 15895
rect 15160 15864 15853 15892
rect 15160 15852 15166 15864
rect 15841 15861 15853 15864
rect 15887 15892 15899 15895
rect 16206 15892 16212 15904
rect 15887 15864 16212 15892
rect 15887 15861 15899 15864
rect 15841 15855 15899 15861
rect 16206 15852 16212 15864
rect 16264 15852 16270 15904
rect 16758 15852 16764 15904
rect 16816 15892 16822 15904
rect 17310 15892 17316 15904
rect 16816 15864 17316 15892
rect 16816 15852 16822 15864
rect 17310 15852 17316 15864
rect 17368 15892 17374 15904
rect 19352 15892 19380 15932
rect 20073 15929 20085 15932
rect 20119 15929 20131 15963
rect 20073 15923 20131 15929
rect 17368 15864 19380 15892
rect 19613 15895 19671 15901
rect 17368 15852 17374 15864
rect 19613 15861 19625 15895
rect 19659 15892 19671 15895
rect 19702 15892 19708 15904
rect 19659 15864 19708 15892
rect 19659 15861 19671 15864
rect 19613 15855 19671 15861
rect 19702 15852 19708 15864
rect 19760 15852 19766 15904
rect 20714 15852 20720 15904
rect 20772 15892 20778 15904
rect 20993 15895 21051 15901
rect 20993 15892 21005 15895
rect 20772 15864 21005 15892
rect 20772 15852 20778 15864
rect 20993 15861 21005 15864
rect 21039 15861 21051 15895
rect 20993 15855 21051 15861
rect 1104 15802 30820 15824
rect 1104 15750 5915 15802
rect 5967 15750 5979 15802
rect 6031 15750 6043 15802
rect 6095 15750 6107 15802
rect 6159 15750 6171 15802
rect 6223 15750 15846 15802
rect 15898 15750 15910 15802
rect 15962 15750 15974 15802
rect 16026 15750 16038 15802
rect 16090 15750 16102 15802
rect 16154 15750 25776 15802
rect 25828 15750 25840 15802
rect 25892 15750 25904 15802
rect 25956 15750 25968 15802
rect 26020 15750 26032 15802
rect 26084 15750 30820 15802
rect 1104 15728 30820 15750
rect 1762 15688 1768 15700
rect 1723 15660 1768 15688
rect 1762 15648 1768 15660
rect 1820 15648 1826 15700
rect 4522 15688 4528 15700
rect 4483 15660 4528 15688
rect 4522 15648 4528 15660
rect 4580 15648 4586 15700
rect 6454 15688 6460 15700
rect 5828 15660 6460 15688
rect 3142 15620 3148 15632
rect 2148 15592 3148 15620
rect 2148 15561 2176 15592
rect 3142 15580 3148 15592
rect 3200 15620 3206 15632
rect 3200 15592 3924 15620
rect 3200 15580 3206 15592
rect 3896 15564 3924 15592
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15521 2191 15555
rect 2774 15552 2780 15564
rect 2133 15515 2191 15521
rect 2516 15524 2780 15552
rect 1946 15484 1952 15496
rect 1907 15456 1952 15484
rect 1946 15444 1952 15456
rect 2004 15444 2010 15496
rect 2225 15487 2283 15493
rect 2225 15453 2237 15487
rect 2271 15453 2283 15487
rect 2225 15447 2283 15453
rect 2240 15416 2268 15447
rect 2314 15444 2320 15496
rect 2372 15484 2378 15496
rect 2516 15493 2544 15524
rect 2774 15512 2780 15524
rect 2832 15552 2838 15564
rect 2832 15524 3832 15552
rect 2832 15512 2838 15524
rect 3804 15496 3832 15524
rect 3878 15512 3884 15564
rect 3936 15552 3942 15564
rect 4157 15555 4215 15561
rect 4157 15552 4169 15555
rect 3936 15524 4169 15552
rect 3936 15512 3942 15524
rect 4157 15521 4169 15524
rect 4203 15521 4215 15555
rect 4157 15515 4215 15521
rect 2501 15487 2559 15493
rect 2372 15456 2417 15484
rect 2372 15444 2378 15456
rect 2501 15453 2513 15487
rect 2547 15453 2559 15487
rect 3142 15484 3148 15496
rect 3103 15456 3148 15484
rect 2501 15447 2559 15453
rect 3142 15444 3148 15456
rect 3200 15444 3206 15496
rect 3786 15484 3792 15496
rect 3747 15456 3792 15484
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 3970 15484 3976 15496
rect 3931 15456 3976 15484
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 4065 15487 4123 15493
rect 4065 15453 4077 15487
rect 4111 15453 4123 15487
rect 4065 15447 4123 15453
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15484 4399 15487
rect 4982 15484 4988 15496
rect 4387 15456 4988 15484
rect 4387 15453 4399 15456
rect 4341 15447 4399 15453
rect 2866 15416 2872 15428
rect 2240 15388 2872 15416
rect 2866 15376 2872 15388
rect 2924 15416 2930 15428
rect 4080 15416 4108 15447
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 5074 15444 5080 15496
rect 5132 15484 5138 15496
rect 5132 15456 5177 15484
rect 5132 15444 5138 15456
rect 5442 15444 5448 15496
rect 5500 15484 5506 15496
rect 5721 15487 5779 15493
rect 5721 15484 5733 15487
rect 5500 15456 5733 15484
rect 5500 15444 5506 15456
rect 5721 15453 5733 15456
rect 5767 15453 5779 15487
rect 5828 15484 5856 15660
rect 6454 15648 6460 15660
rect 6512 15648 6518 15700
rect 6638 15648 6644 15700
rect 6696 15688 6702 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 6696 15660 8953 15688
rect 6696 15648 6702 15660
rect 8941 15657 8953 15660
rect 8987 15657 8999 15691
rect 8941 15651 8999 15657
rect 9769 15691 9827 15697
rect 9769 15657 9781 15691
rect 9815 15688 9827 15691
rect 9858 15688 9864 15700
rect 9815 15660 9864 15688
rect 9815 15657 9827 15660
rect 9769 15651 9827 15657
rect 7650 15580 7656 15632
rect 7708 15580 7714 15632
rect 8956 15620 8984 15651
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 14553 15691 14611 15697
rect 14553 15657 14565 15691
rect 14599 15688 14611 15691
rect 14734 15688 14740 15700
rect 14599 15660 14740 15688
rect 14599 15657 14611 15660
rect 14553 15651 14611 15657
rect 14734 15648 14740 15660
rect 14792 15648 14798 15700
rect 16117 15691 16175 15697
rect 16117 15657 16129 15691
rect 16163 15688 16175 15691
rect 16298 15688 16304 15700
rect 16163 15660 16304 15688
rect 16163 15657 16175 15660
rect 16117 15651 16175 15657
rect 16298 15648 16304 15660
rect 16356 15648 16362 15700
rect 16408 15660 16988 15688
rect 10134 15620 10140 15632
rect 8956 15592 10140 15620
rect 10134 15580 10140 15592
rect 10192 15580 10198 15632
rect 16408 15620 16436 15660
rect 16850 15620 16856 15632
rect 15028 15592 16436 15620
rect 16776 15592 16856 15620
rect 5997 15555 6055 15561
rect 5997 15521 6009 15555
rect 6043 15552 6055 15555
rect 6638 15552 6644 15564
rect 6043 15524 6644 15552
rect 6043 15521 6055 15524
rect 5997 15515 6055 15521
rect 6638 15512 6644 15524
rect 6696 15512 6702 15564
rect 7668 15552 7696 15580
rect 15028 15564 15056 15592
rect 8754 15552 8760 15564
rect 7576 15524 8760 15552
rect 5905 15487 5963 15493
rect 5905 15484 5917 15487
rect 5828 15456 5917 15484
rect 5721 15447 5779 15453
rect 5905 15453 5917 15456
rect 5951 15453 5963 15487
rect 5905 15447 5963 15453
rect 6089 15487 6147 15493
rect 6089 15453 6101 15487
rect 6135 15453 6147 15487
rect 6089 15447 6147 15453
rect 2924 15388 4108 15416
rect 6104 15416 6132 15447
rect 6178 15444 6184 15496
rect 6236 15484 6242 15496
rect 7576 15493 7604 15524
rect 8754 15512 8760 15524
rect 8812 15512 8818 15564
rect 9398 15552 9404 15564
rect 8864 15524 9404 15552
rect 6273 15487 6331 15493
rect 6273 15484 6285 15487
rect 6236 15456 6285 15484
rect 6236 15444 6242 15456
rect 6273 15453 6285 15456
rect 6319 15453 6331 15487
rect 6273 15447 6331 15453
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15453 7619 15487
rect 7561 15447 7619 15453
rect 7650 15444 7656 15496
rect 7708 15484 7714 15496
rect 8067 15487 8125 15493
rect 7708 15456 7753 15484
rect 7708 15444 7714 15456
rect 8067 15453 8079 15487
rect 8113 15484 8125 15487
rect 8864 15484 8892 15524
rect 9398 15512 9404 15524
rect 9456 15552 9462 15564
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 9456 15524 10333 15552
rect 9456 15512 9462 15524
rect 10321 15521 10333 15524
rect 10367 15521 10379 15555
rect 10321 15515 10379 15521
rect 13449 15555 13507 15561
rect 13449 15521 13461 15555
rect 13495 15552 13507 15555
rect 14090 15552 14096 15564
rect 13495 15524 14096 15552
rect 13495 15521 13507 15524
rect 13449 15515 13507 15521
rect 14090 15512 14096 15524
rect 14148 15512 14154 15564
rect 15010 15552 15016 15564
rect 14923 15524 15016 15552
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 15194 15512 15200 15564
rect 15252 15552 15258 15564
rect 15252 15524 16712 15552
rect 15252 15512 15258 15524
rect 8113 15456 8892 15484
rect 8941 15487 8999 15493
rect 8113 15453 8125 15456
rect 8067 15447 8125 15453
rect 8941 15453 8953 15487
rect 8987 15484 8999 15487
rect 9033 15487 9091 15493
rect 9033 15484 9045 15487
rect 8987 15456 9045 15484
rect 8987 15453 8999 15456
rect 8941 15447 8999 15453
rect 9033 15453 9045 15456
rect 9079 15453 9091 15487
rect 9033 15447 9091 15453
rect 9122 15444 9128 15496
rect 9180 15484 9186 15496
rect 9217 15487 9275 15493
rect 9217 15484 9229 15487
rect 9180 15456 9229 15484
rect 9180 15444 9186 15456
rect 9217 15453 9229 15456
rect 9263 15453 9275 15487
rect 9217 15447 9275 15453
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15453 9367 15487
rect 9582 15484 9588 15496
rect 9543 15456 9588 15484
rect 9309 15447 9367 15453
rect 6730 15416 6736 15428
rect 6104 15388 6736 15416
rect 2924 15376 2930 15388
rect 6730 15376 6736 15388
rect 6788 15376 6794 15428
rect 7374 15376 7380 15428
rect 7432 15416 7438 15428
rect 7837 15419 7895 15425
rect 7837 15416 7849 15419
rect 7432 15388 7849 15416
rect 7432 15376 7438 15388
rect 7837 15385 7849 15388
rect 7883 15385 7895 15419
rect 7837 15379 7895 15385
rect 7926 15376 7932 15428
rect 7984 15416 7990 15428
rect 9324 15416 9352 15447
rect 9582 15444 9588 15456
rect 9640 15444 9646 15496
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 10042 15484 10048 15496
rect 9732 15456 10048 15484
rect 9732 15444 9738 15456
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 12621 15487 12679 15493
rect 12621 15453 12633 15487
rect 12667 15484 12679 15487
rect 13081 15487 13139 15493
rect 13081 15484 13093 15487
rect 12667 15456 13093 15484
rect 12667 15453 12679 15456
rect 12621 15447 12679 15453
rect 13081 15453 13093 15456
rect 13127 15453 13139 15487
rect 13081 15447 13139 15453
rect 13265 15487 13323 15493
rect 13265 15453 13277 15487
rect 13311 15484 13323 15487
rect 13354 15484 13360 15496
rect 13311 15456 13360 15484
rect 13311 15453 13323 15456
rect 13265 15447 13323 15453
rect 10244 15416 10272 15447
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 14734 15484 14740 15496
rect 14695 15456 14740 15484
rect 14734 15444 14740 15456
rect 14792 15444 14798 15496
rect 14921 15487 14979 15493
rect 14921 15453 14933 15487
rect 14967 15453 14979 15487
rect 14921 15447 14979 15453
rect 15101 15485 15159 15491
rect 15101 15451 15113 15485
rect 15147 15462 15159 15485
rect 15289 15487 15347 15493
rect 15147 15451 15240 15462
rect 7984 15388 8029 15416
rect 8128 15388 10272 15416
rect 7984 15376 7990 15388
rect 8128 15360 8156 15388
rect 10318 15376 10324 15428
rect 10376 15416 10382 15428
rect 11238 15416 11244 15428
rect 10376 15388 11244 15416
rect 10376 15376 10382 15388
rect 11238 15376 11244 15388
rect 11296 15376 11302 15428
rect 14936 15416 14964 15447
rect 15101 15445 15240 15451
rect 15289 15453 15301 15487
rect 15335 15484 15347 15487
rect 16574 15484 16580 15496
rect 15335 15456 16580 15484
rect 15335 15453 15347 15456
rect 15289 15447 15347 15453
rect 15120 15434 15240 15445
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 16684 15493 16712 15524
rect 16669 15487 16727 15493
rect 16669 15453 16681 15487
rect 16715 15453 16727 15487
rect 16669 15447 16727 15453
rect 16776 15480 16804 15592
rect 16850 15580 16856 15592
rect 16908 15580 16914 15632
rect 16960 15620 16988 15660
rect 17218 15648 17224 15700
rect 17276 15688 17282 15700
rect 17405 15691 17463 15697
rect 17405 15688 17417 15691
rect 17276 15660 17417 15688
rect 17276 15648 17282 15660
rect 17405 15657 17417 15660
rect 17451 15657 17463 15691
rect 20806 15688 20812 15700
rect 20767 15660 20812 15688
rect 17405 15651 17463 15657
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 29454 15648 29460 15700
rect 29512 15688 29518 15700
rect 29917 15691 29975 15697
rect 29917 15688 29929 15691
rect 29512 15660 29929 15688
rect 29512 15648 29518 15660
rect 29917 15657 29929 15660
rect 29963 15657 29975 15691
rect 29917 15651 29975 15657
rect 16960 15592 17255 15620
rect 16960 15561 16988 15592
rect 16945 15555 17003 15561
rect 16945 15521 16957 15555
rect 16991 15521 17003 15555
rect 17227 15552 17255 15592
rect 19334 15552 19340 15564
rect 17227 15524 19340 15552
rect 16945 15515 17003 15521
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 16841 15487 16899 15493
rect 16841 15480 16853 15487
rect 16776 15453 16853 15480
rect 16887 15453 16899 15487
rect 16776 15452 16899 15453
rect 16841 15447 16899 15452
rect 14844 15388 14964 15416
rect 14844 15360 14872 15388
rect 2958 15348 2964 15360
rect 2919 15320 2964 15348
rect 2958 15308 2964 15320
rect 3016 15308 3022 15360
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 5810 15348 5816 15360
rect 5215 15320 5816 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 5810 15308 5816 15320
rect 5868 15308 5874 15360
rect 6454 15348 6460 15360
rect 6415 15320 6460 15348
rect 6454 15308 6460 15320
rect 6512 15308 6518 15360
rect 7650 15308 7656 15360
rect 7708 15348 7714 15360
rect 8110 15348 8116 15360
rect 7708 15320 8116 15348
rect 7708 15308 7714 15320
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 8205 15351 8263 15357
rect 8205 15317 8217 15351
rect 8251 15348 8263 15351
rect 8754 15348 8760 15360
rect 8251 15320 8760 15348
rect 8251 15317 8263 15320
rect 8205 15311 8263 15317
rect 8754 15308 8760 15320
rect 8812 15308 8818 15360
rect 9306 15308 9312 15360
rect 9364 15348 9370 15360
rect 9674 15348 9680 15360
rect 9364 15320 9680 15348
rect 9364 15308 9370 15320
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 9858 15308 9864 15360
rect 9916 15348 9922 15360
rect 10594 15348 10600 15360
rect 9916 15320 10600 15348
rect 9916 15308 9922 15320
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 12437 15351 12495 15357
rect 12437 15317 12449 15351
rect 12483 15348 12495 15351
rect 12526 15348 12532 15360
rect 12483 15320 12532 15348
rect 12483 15317 12495 15320
rect 12437 15311 12495 15317
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 14826 15308 14832 15360
rect 14884 15308 14890 15360
rect 15102 15308 15108 15360
rect 15160 15348 15166 15360
rect 15212 15348 15240 15434
rect 16025 15419 16083 15425
rect 16025 15385 16037 15419
rect 16071 15416 16083 15419
rect 16390 15416 16396 15428
rect 16071 15388 16396 15416
rect 16071 15385 16083 15388
rect 16025 15379 16083 15385
rect 16390 15376 16396 15388
rect 16448 15376 16454 15428
rect 16684 15416 16712 15447
rect 17034 15444 17040 15496
rect 17092 15484 17098 15496
rect 17092 15456 17137 15484
rect 17092 15444 17098 15456
rect 17218 15444 17224 15496
rect 17276 15484 17282 15496
rect 17276 15456 17321 15484
rect 17276 15444 17282 15456
rect 17402 15444 17408 15496
rect 17460 15484 17466 15496
rect 18598 15484 18604 15496
rect 17460 15456 18460 15484
rect 18559 15456 18604 15484
rect 17460 15444 17466 15456
rect 18230 15416 18236 15428
rect 16684 15388 18236 15416
rect 18230 15376 18236 15388
rect 18288 15376 18294 15428
rect 18432 15416 18460 15456
rect 18598 15444 18604 15456
rect 18656 15444 18662 15496
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15484 19487 15487
rect 19518 15484 19524 15496
rect 19475 15456 19524 15484
rect 19475 15453 19487 15456
rect 19429 15447 19487 15453
rect 19518 15444 19524 15456
rect 19576 15444 19582 15496
rect 19702 15493 19708 15496
rect 19696 15484 19708 15493
rect 19663 15456 19708 15484
rect 19696 15447 19708 15456
rect 19702 15444 19708 15447
rect 19760 15444 19766 15496
rect 21269 15487 21327 15493
rect 21269 15453 21281 15487
rect 21315 15484 21327 15487
rect 21450 15484 21456 15496
rect 21315 15456 21456 15484
rect 21315 15453 21327 15456
rect 21269 15447 21327 15453
rect 21450 15444 21456 15456
rect 21508 15444 21514 15496
rect 29914 15484 29920 15496
rect 29875 15456 29920 15484
rect 29914 15444 29920 15456
rect 29972 15444 29978 15496
rect 30098 15484 30104 15496
rect 30059 15456 30104 15484
rect 30098 15444 30104 15456
rect 30156 15444 30162 15496
rect 18432 15388 21496 15416
rect 15160 15320 15240 15348
rect 15160 15308 15166 15320
rect 16942 15308 16948 15360
rect 17000 15348 17006 15360
rect 18509 15351 18567 15357
rect 18509 15348 18521 15351
rect 17000 15320 18521 15348
rect 17000 15308 17006 15320
rect 18509 15317 18521 15320
rect 18555 15348 18567 15351
rect 19242 15348 19248 15360
rect 18555 15320 19248 15348
rect 18555 15317 18567 15320
rect 18509 15311 18567 15317
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 21468 15357 21496 15388
rect 21453 15351 21511 15357
rect 21453 15317 21465 15351
rect 21499 15348 21511 15351
rect 21818 15348 21824 15360
rect 21499 15320 21824 15348
rect 21499 15317 21511 15320
rect 21453 15311 21511 15317
rect 21818 15308 21824 15320
rect 21876 15308 21882 15360
rect 1104 15258 30820 15280
rect 1104 15206 10880 15258
rect 10932 15206 10944 15258
rect 10996 15206 11008 15258
rect 11060 15206 11072 15258
rect 11124 15206 11136 15258
rect 11188 15206 20811 15258
rect 20863 15206 20875 15258
rect 20927 15206 20939 15258
rect 20991 15206 21003 15258
rect 21055 15206 21067 15258
rect 21119 15206 30820 15258
rect 1104 15184 30820 15206
rect 1486 15104 1492 15156
rect 1544 15144 1550 15156
rect 1544 15116 3280 15144
rect 1544 15104 1550 15116
rect 3050 15076 3056 15088
rect 1964 15048 3056 15076
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 1964 15017 1992 15048
rect 3050 15036 3056 15048
rect 3108 15076 3114 15088
rect 3252 15076 3280 15116
rect 7374 15104 7380 15156
rect 7432 15144 7438 15156
rect 7653 15147 7711 15153
rect 7653 15144 7665 15147
rect 7432 15116 7665 15144
rect 7432 15104 7438 15116
rect 7653 15113 7665 15116
rect 7699 15113 7711 15147
rect 7653 15107 7711 15113
rect 8680 15116 11836 15144
rect 3513 15079 3571 15085
rect 3108 15048 3188 15076
rect 3252 15048 3464 15076
rect 3108 15036 3114 15048
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 14977 2007 15011
rect 2130 15008 2136 15020
rect 2091 14980 2136 15008
rect 1949 14971 2007 14977
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 15008 2375 15011
rect 2498 15008 2504 15020
rect 2363 14980 2504 15008
rect 2363 14977 2375 14980
rect 2317 14971 2375 14977
rect 2498 14968 2504 14980
rect 2556 14968 2562 15020
rect 2774 14968 2780 15020
rect 2832 15008 2838 15020
rect 2958 15008 2964 15020
rect 2832 14980 2877 15008
rect 2919 14980 2964 15008
rect 2832 14968 2838 14980
rect 2958 14968 2964 14980
rect 3016 14968 3022 15020
rect 3160 15017 3188 15048
rect 3145 15011 3203 15017
rect 3145 14977 3157 15011
rect 3191 14977 3203 15011
rect 3145 14971 3203 14977
rect 3329 15011 3387 15017
rect 3329 14977 3341 15011
rect 3375 14977 3387 15011
rect 3436 15008 3464 15048
rect 3513 15045 3525 15079
rect 3559 15076 3571 15079
rect 4218 15079 4276 15085
rect 4218 15076 4230 15079
rect 3559 15048 4230 15076
rect 3559 15045 3571 15048
rect 3513 15039 3571 15045
rect 4218 15045 4230 15048
rect 4264 15045 4276 15079
rect 8680 15076 8708 15116
rect 4218 15039 4276 15045
rect 5644 15048 8708 15076
rect 5644 15008 5672 15048
rect 8754 15036 8760 15088
rect 8812 15085 8818 15088
rect 8812 15076 8824 15085
rect 8812 15048 8857 15076
rect 8812 15039 8824 15048
rect 8812 15036 8818 15039
rect 9582 15036 9588 15088
rect 9640 15076 9646 15088
rect 9738 15079 9796 15085
rect 9738 15076 9750 15079
rect 9640 15048 9750 15076
rect 9640 15036 9646 15048
rect 9738 15045 9750 15048
rect 9784 15045 9796 15079
rect 9738 15039 9796 15045
rect 10042 15036 10048 15088
rect 10100 15076 10106 15088
rect 10318 15076 10324 15088
rect 10100 15048 10324 15076
rect 10100 15036 10106 15048
rect 10318 15036 10324 15048
rect 10376 15036 10382 15088
rect 11808 15085 11836 15116
rect 14826 15104 14832 15156
rect 14884 15144 14890 15156
rect 16942 15144 16948 15156
rect 14884 15116 16948 15144
rect 14884 15104 14890 15116
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17681 15147 17739 15153
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 29914 15144 29920 15156
rect 17727 15116 29920 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 29914 15104 29920 15116
rect 29972 15104 29978 15156
rect 11793 15079 11851 15085
rect 11793 15045 11805 15079
rect 11839 15045 11851 15079
rect 13814 15076 13820 15088
rect 11793 15039 11851 15045
rect 11900 15048 13820 15076
rect 3436 14980 5672 15008
rect 3329 14971 3387 14977
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 1486 14764 1492 14816
rect 1544 14804 1550 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 1544 14776 1593 14804
rect 1544 14764 1550 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 2056 14804 2084 14903
rect 2866 14900 2872 14952
rect 2924 14940 2930 14952
rect 3053 14943 3111 14949
rect 3053 14940 3065 14943
rect 2924 14912 3065 14940
rect 2924 14900 2930 14912
rect 3053 14909 3065 14912
rect 3099 14909 3111 14943
rect 3053 14903 3111 14909
rect 2774 14804 2780 14816
rect 2056 14776 2780 14804
rect 1581 14767 1639 14773
rect 2774 14764 2780 14776
rect 2832 14764 2838 14816
rect 3344 14804 3372 14971
rect 5718 14968 5724 15020
rect 5776 15008 5782 15020
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 5776 14980 6377 15008
rect 5776 14968 5782 14980
rect 6365 14977 6377 14980
rect 6411 14977 6423 15011
rect 6546 15008 6552 15020
rect 6507 14980 6552 15008
rect 6365 14971 6423 14977
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 6638 14968 6644 15020
rect 6696 15008 6702 15020
rect 6914 15008 6920 15020
rect 6696 14980 6741 15008
rect 6875 14980 6920 15008
rect 6696 14968 6702 14980
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 7098 14968 7104 15020
rect 7156 15008 7162 15020
rect 9033 15011 9091 15017
rect 7156 14980 8984 15008
rect 7156 14968 7162 14980
rect 3786 14900 3792 14952
rect 3844 14940 3850 14952
rect 3973 14943 4031 14949
rect 3973 14940 3985 14943
rect 3844 14912 3985 14940
rect 3844 14900 3850 14912
rect 3973 14909 3985 14912
rect 4019 14909 4031 14943
rect 3973 14903 4031 14909
rect 6730 14900 6736 14952
rect 6788 14940 6794 14952
rect 8956 14940 8984 14980
rect 9033 14977 9045 15011
rect 9079 15008 9091 15011
rect 9306 15008 9312 15020
rect 9079 14980 9312 15008
rect 9079 14977 9091 14980
rect 9033 14971 9091 14977
rect 9306 14968 9312 14980
rect 9364 15008 9370 15020
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 9364 14980 9505 15008
rect 9364 14968 9370 14980
rect 9493 14977 9505 14980
rect 9539 14977 9551 15011
rect 11900 15008 11928 15048
rect 13814 15036 13820 15048
rect 13872 15036 13878 15088
rect 17034 15076 17040 15088
rect 14292 15048 14872 15076
rect 9493 14971 9551 14977
rect 9600 14980 11928 15008
rect 12253 15011 12311 15017
rect 9600 14940 9628 14980
rect 12253 14977 12265 15011
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 6788 14912 6833 14940
rect 8956 14912 9628 14940
rect 12268 14940 12296 14971
rect 12342 14968 12348 15020
rect 12400 15017 12406 15020
rect 12400 15011 12449 15017
rect 12400 14977 12403 15011
rect 12437 14977 12449 15011
rect 12400 14971 12449 14977
rect 12400 14968 12406 14971
rect 12526 14968 12532 15020
rect 12584 15008 12590 15020
rect 13262 15008 13268 15020
rect 12584 14980 12629 15008
rect 13223 14980 13268 15008
rect 12584 14968 12590 14980
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 15008 13507 15011
rect 13538 15008 13544 15020
rect 13495 14980 13544 15008
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 13538 14968 13544 14980
rect 13596 15008 13602 15020
rect 14292 15008 14320 15048
rect 14458 15008 14464 15020
rect 13596 14980 14320 15008
rect 14419 14980 14464 15008
rect 13596 14968 13602 14980
rect 14458 14968 14464 14980
rect 14516 14968 14522 15020
rect 14550 14968 14556 15020
rect 14608 15008 14614 15020
rect 14717 15011 14775 15017
rect 14717 15008 14729 15011
rect 14608 14980 14729 15008
rect 14608 14968 14614 14980
rect 14717 14977 14729 14980
rect 14763 14977 14775 15011
rect 14844 15008 14872 15048
rect 16684 15048 17040 15076
rect 16684 15008 16712 15048
rect 17034 15036 17040 15048
rect 17092 15036 17098 15088
rect 18417 15079 18475 15085
rect 18417 15045 18429 15079
rect 18463 15076 18475 15079
rect 18874 15076 18880 15088
rect 18463 15048 18880 15076
rect 18463 15045 18475 15048
rect 18417 15039 18475 15045
rect 18874 15036 18880 15048
rect 18932 15036 18938 15088
rect 19426 15036 19432 15088
rect 19484 15076 19490 15088
rect 19521 15079 19579 15085
rect 19521 15076 19533 15079
rect 19484 15048 19533 15076
rect 19484 15036 19490 15048
rect 19521 15045 19533 15048
rect 19567 15045 19579 15079
rect 19521 15039 19579 15045
rect 20456 15048 22140 15076
rect 17126 15008 17132 15020
rect 14844 14980 16712 15008
rect 17087 14980 17132 15008
rect 14717 14971 14775 14977
rect 17126 14968 17132 14980
rect 17184 14968 17190 15020
rect 17218 14968 17224 15020
rect 17276 15008 17282 15020
rect 17405 15011 17463 15017
rect 17405 15008 17417 15011
rect 17276 14980 17417 15008
rect 17276 14968 17282 14980
rect 17405 14977 17417 14980
rect 17451 14977 17463 15011
rect 17405 14971 17463 14977
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 12802 14940 12808 14952
rect 12268 14912 12808 14940
rect 6788 14900 6794 14912
rect 12802 14900 12808 14912
rect 12860 14940 12866 14952
rect 13280 14940 13308 14968
rect 12860 14912 13308 14940
rect 12860 14900 12866 14912
rect 16298 14900 16304 14952
rect 16356 14940 16362 14952
rect 17512 14940 17540 14971
rect 17862 14968 17868 15020
rect 17920 15008 17926 15020
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 17920 14980 18153 15008
rect 17920 14968 17926 14980
rect 18141 14977 18153 14980
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 18289 15011 18347 15017
rect 18289 14977 18301 15011
rect 18335 15008 18347 15011
rect 18506 15008 18512 15020
rect 18335 14977 18368 15008
rect 18467 14980 18512 15008
rect 18289 14971 18368 14977
rect 17954 14940 17960 14952
rect 16356 14912 17960 14940
rect 16356 14900 16362 14912
rect 17954 14900 17960 14912
rect 18012 14900 18018 14952
rect 18340 14940 18368 14971
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 18598 14968 18604 15020
rect 18656 15017 18662 15020
rect 18656 15008 18664 15017
rect 19337 15011 19395 15017
rect 18656 14980 18701 15008
rect 18656 14971 18664 14980
rect 19337 14977 19349 15011
rect 19383 15008 19395 15011
rect 19610 15008 19616 15020
rect 19383 14980 19616 15008
rect 19383 14977 19395 14980
rect 19337 14971 19395 14977
rect 18656 14968 18662 14971
rect 19352 14940 19380 14971
rect 19610 14968 19616 14980
rect 19668 14968 19674 15020
rect 19794 14968 19800 15020
rect 19852 15008 19858 15020
rect 20456 15017 20484 15048
rect 20441 15011 20499 15017
rect 20441 15008 20453 15011
rect 19852 14980 20453 15008
rect 19852 14968 19858 14980
rect 20441 14977 20453 14980
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 20530 14968 20536 15020
rect 20588 15008 20594 15020
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 20588 14980 20729 15008
rect 20588 14968 20594 14980
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 20809 15011 20867 15017
rect 20809 14977 20821 15011
rect 20855 14977 20867 15011
rect 21818 15008 21824 15020
rect 21779 14980 21824 15008
rect 20809 14971 20867 14977
rect 18340 14912 19380 14940
rect 20622 14900 20628 14952
rect 20680 14940 20686 14952
rect 20824 14940 20852 14971
rect 21818 14968 21824 14980
rect 21876 14968 21882 15020
rect 22112 15017 22140 15048
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 14977 22155 15011
rect 29181 15011 29239 15017
rect 29181 15008 29193 15011
rect 22097 14971 22155 14977
rect 26206 14980 29193 15008
rect 20680 14912 20852 14940
rect 20680 14900 20686 14912
rect 5902 14832 5908 14884
rect 5960 14872 5966 14884
rect 6546 14872 6552 14884
rect 5960 14844 6552 14872
rect 5960 14832 5966 14844
rect 6546 14832 6552 14844
rect 6604 14832 6610 14884
rect 7101 14875 7159 14881
rect 7101 14841 7113 14875
rect 7147 14872 7159 14875
rect 20533 14875 20591 14881
rect 20533 14872 20545 14875
rect 7147 14844 8156 14872
rect 7147 14841 7159 14844
rect 7101 14835 7159 14841
rect 5074 14804 5080 14816
rect 3344 14776 5080 14804
rect 5074 14764 5080 14776
rect 5132 14804 5138 14816
rect 5353 14807 5411 14813
rect 5353 14804 5365 14807
rect 5132 14776 5365 14804
rect 5132 14764 5138 14776
rect 5353 14773 5365 14776
rect 5399 14773 5411 14807
rect 5353 14767 5411 14773
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 8018 14804 8024 14816
rect 6512 14776 8024 14804
rect 6512 14764 6518 14776
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 8128 14804 8156 14844
rect 10428 14844 13400 14872
rect 10428 14804 10456 14844
rect 8128 14776 10456 14804
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 10873 14807 10931 14813
rect 10873 14804 10885 14807
rect 10652 14776 10885 14804
rect 10652 14764 10658 14776
rect 10873 14773 10885 14776
rect 10919 14773 10931 14807
rect 13262 14804 13268 14816
rect 13223 14776 13268 14804
rect 10873 14767 10931 14773
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 13372 14804 13400 14844
rect 15764 14844 20545 14872
rect 15764 14804 15792 14844
rect 20533 14841 20545 14844
rect 20579 14841 20591 14875
rect 20533 14835 20591 14841
rect 20993 14875 21051 14881
rect 20993 14841 21005 14875
rect 21039 14872 21051 14875
rect 26206 14872 26234 14980
rect 29181 14977 29193 14980
rect 29227 14977 29239 15011
rect 29181 14971 29239 14977
rect 29365 15011 29423 15017
rect 29365 14977 29377 15011
rect 29411 14977 29423 15011
rect 29365 14971 29423 14977
rect 29825 15011 29883 15017
rect 29825 14977 29837 15011
rect 29871 15008 29883 15011
rect 29914 15008 29920 15020
rect 29871 14980 29920 15008
rect 29871 14977 29883 14980
rect 29825 14971 29883 14977
rect 29380 14940 29408 14971
rect 29914 14968 29920 14980
rect 29972 14968 29978 15020
rect 30098 14940 30104 14952
rect 29380 14912 30104 14940
rect 30098 14900 30104 14912
rect 30156 14900 30162 14952
rect 29178 14872 29184 14884
rect 21039 14844 26234 14872
rect 29139 14844 29184 14872
rect 21039 14841 21051 14844
rect 20993 14835 21051 14841
rect 29178 14832 29184 14844
rect 29236 14832 29242 14884
rect 30006 14872 30012 14884
rect 29967 14844 30012 14872
rect 30006 14832 30012 14844
rect 30064 14832 30070 14884
rect 13372 14776 15792 14804
rect 15841 14807 15899 14813
rect 15841 14773 15853 14807
rect 15887 14804 15899 14807
rect 16206 14804 16212 14816
rect 15887 14776 16212 14804
rect 15887 14773 15899 14776
rect 15841 14767 15899 14773
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 16942 14764 16948 14816
rect 17000 14804 17006 14816
rect 17221 14807 17279 14813
rect 17221 14804 17233 14807
rect 17000 14776 17233 14804
rect 17000 14764 17006 14776
rect 17221 14773 17233 14776
rect 17267 14773 17279 14807
rect 17221 14767 17279 14773
rect 17310 14764 17316 14816
rect 17368 14804 17374 14816
rect 18598 14804 18604 14816
rect 17368 14776 18604 14804
rect 17368 14764 17374 14776
rect 18598 14764 18604 14776
rect 18656 14764 18662 14816
rect 18785 14807 18843 14813
rect 18785 14773 18797 14807
rect 18831 14804 18843 14807
rect 19334 14804 19340 14816
rect 18831 14776 19340 14804
rect 18831 14773 18843 14776
rect 18785 14767 18843 14773
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 1104 14714 30820 14736
rect 1104 14662 5915 14714
rect 5967 14662 5979 14714
rect 6031 14662 6043 14714
rect 6095 14662 6107 14714
rect 6159 14662 6171 14714
rect 6223 14662 15846 14714
rect 15898 14662 15910 14714
rect 15962 14662 15974 14714
rect 16026 14662 16038 14714
rect 16090 14662 16102 14714
rect 16154 14662 25776 14714
rect 25828 14662 25840 14714
rect 25892 14662 25904 14714
rect 25956 14662 25968 14714
rect 26020 14662 26032 14714
rect 26084 14662 30820 14714
rect 1104 14640 30820 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 2130 14600 2136 14612
rect 1627 14572 2136 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 2130 14560 2136 14572
rect 2188 14560 2194 14612
rect 5166 14600 5172 14612
rect 3068 14572 5172 14600
rect 2866 14532 2872 14544
rect 2792 14504 2872 14532
rect 2792 14473 2820 14504
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14433 2835 14467
rect 2777 14427 2835 14433
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 2498 14396 2504 14408
rect 2459 14368 2504 14396
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 2682 14396 2688 14408
rect 2643 14368 2688 14396
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14396 2927 14399
rect 2958 14396 2964 14408
rect 2915 14368 2964 14396
rect 2915 14365 2927 14368
rect 2869 14359 2927 14365
rect 2958 14356 2964 14368
rect 3016 14356 3022 14408
rect 3068 14405 3096 14572
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 6822 14600 6828 14612
rect 6288 14572 6828 14600
rect 5902 14464 5908 14476
rect 5863 14436 5908 14464
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14365 3111 14399
rect 3786 14396 3792 14408
rect 3747 14368 3792 14396
rect 3053 14359 3111 14365
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 5629 14399 5687 14405
rect 5629 14396 5641 14399
rect 5592 14368 5641 14396
rect 5592 14356 5598 14368
rect 5629 14365 5641 14368
rect 5675 14365 5687 14399
rect 5810 14396 5816 14408
rect 5771 14368 5816 14396
rect 5629 14359 5687 14365
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 5997 14399 6055 14405
rect 5997 14365 6009 14399
rect 6043 14365 6055 14399
rect 5997 14359 6055 14365
rect 6181 14399 6239 14405
rect 6181 14365 6193 14399
rect 6227 14396 6239 14399
rect 6288 14396 6316 14572
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7190 14560 7196 14612
rect 7248 14600 7254 14612
rect 7374 14600 7380 14612
rect 7248 14572 7380 14600
rect 7248 14560 7254 14572
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 8110 14600 8116 14612
rect 8071 14572 8116 14600
rect 8110 14560 8116 14572
rect 8168 14560 8174 14612
rect 9582 14600 9588 14612
rect 9543 14572 9588 14600
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 14461 14603 14519 14609
rect 9692 14572 14412 14600
rect 8018 14492 8024 14544
rect 8076 14532 8082 14544
rect 9692 14532 9720 14572
rect 12066 14532 12072 14544
rect 8076 14504 9720 14532
rect 9876 14504 12072 14532
rect 8076 14492 8082 14504
rect 6365 14467 6423 14473
rect 6365 14433 6377 14467
rect 6411 14464 6423 14467
rect 6914 14464 6920 14476
rect 6411 14436 6920 14464
rect 6411 14433 6423 14436
rect 6365 14427 6423 14433
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 7098 14424 7104 14476
rect 7156 14464 7162 14476
rect 7156 14436 7201 14464
rect 7156 14424 7162 14436
rect 8110 14424 8116 14476
rect 8168 14464 8174 14476
rect 8168 14436 9076 14464
rect 8168 14424 8174 14436
rect 6227 14368 6316 14396
rect 6227 14365 6239 14368
rect 6181 14359 6239 14365
rect 3237 14331 3295 14337
rect 3237 14297 3249 14331
rect 3283 14328 3295 14331
rect 4034 14331 4092 14337
rect 4034 14328 4046 14331
rect 3283 14300 4046 14328
rect 3283 14297 3295 14300
rect 3237 14291 3295 14297
rect 4034 14297 4046 14300
rect 4080 14297 4092 14331
rect 6012 14328 6040 14359
rect 6730 14356 6736 14408
rect 6788 14396 6794 14408
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 6788 14368 6837 14396
rect 6788 14356 6794 14368
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 7006 14396 7012 14408
rect 6967 14368 7012 14396
rect 6825 14359 6883 14365
rect 7006 14356 7012 14368
rect 7064 14356 7070 14408
rect 7190 14396 7196 14408
rect 7116 14368 7196 14396
rect 7116 14328 7144 14368
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 7374 14396 7380 14408
rect 7335 14368 7380 14396
rect 7374 14356 7380 14368
rect 7432 14356 7438 14408
rect 8938 14396 8944 14408
rect 8899 14368 8944 14396
rect 8938 14356 8944 14368
rect 8996 14356 9002 14408
rect 9048 14405 9076 14436
rect 9582 14424 9588 14476
rect 9640 14464 9646 14476
rect 9876 14464 9904 14504
rect 12066 14492 12072 14504
rect 12124 14492 12130 14544
rect 13354 14492 13360 14544
rect 13412 14532 13418 14544
rect 13541 14535 13599 14541
rect 13541 14532 13553 14535
rect 13412 14504 13553 14532
rect 13412 14492 13418 14504
rect 13541 14501 13553 14504
rect 13587 14501 13599 14535
rect 14384 14532 14412 14572
rect 14461 14569 14473 14603
rect 14507 14600 14519 14603
rect 14550 14600 14556 14612
rect 14507 14572 14556 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 16666 14560 16672 14612
rect 16724 14600 16730 14612
rect 18417 14603 18475 14609
rect 18417 14600 18429 14603
rect 16724 14572 18429 14600
rect 16724 14560 16730 14572
rect 18417 14569 18429 14572
rect 18463 14569 18475 14603
rect 18417 14563 18475 14569
rect 18598 14560 18604 14612
rect 18656 14600 18662 14612
rect 20714 14600 20720 14612
rect 18656 14572 20720 14600
rect 18656 14560 18662 14572
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 29914 14600 29920 14612
rect 29875 14572 29920 14600
rect 29914 14560 29920 14572
rect 29972 14560 29978 14612
rect 19889 14535 19947 14541
rect 19889 14532 19901 14535
rect 14384 14504 19901 14532
rect 13541 14495 13599 14501
rect 19889 14501 19901 14504
rect 19935 14501 19947 14535
rect 19889 14495 19947 14501
rect 20349 14535 20407 14541
rect 20349 14501 20361 14535
rect 20395 14532 20407 14535
rect 28994 14532 29000 14544
rect 20395 14504 29000 14532
rect 20395 14501 20407 14504
rect 20349 14495 20407 14501
rect 28994 14492 29000 14504
rect 29052 14492 29058 14544
rect 10594 14464 10600 14476
rect 9640 14436 9904 14464
rect 9968 14436 10600 14464
rect 9640 14424 9646 14436
rect 9034 14399 9092 14405
rect 9034 14365 9046 14399
rect 9080 14365 9092 14399
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 9034 14359 9092 14365
rect 9140 14368 9321 14396
rect 6012 14300 7144 14328
rect 8205 14331 8263 14337
rect 4034 14291 4092 14297
rect 8205 14297 8217 14331
rect 8251 14328 8263 14331
rect 8294 14328 8300 14340
rect 8251 14300 8300 14328
rect 8251 14297 8263 14300
rect 8205 14291 8263 14297
rect 8294 14288 8300 14300
rect 8352 14288 8358 14340
rect 8389 14331 8447 14337
rect 8389 14297 8401 14331
rect 8435 14297 8447 14331
rect 8389 14291 8447 14297
rect 7558 14260 7564 14272
rect 7519 14232 7564 14260
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 8404 14260 8432 14291
rect 8478 14288 8484 14340
rect 8536 14328 8542 14340
rect 9140 14328 9168 14368
rect 9309 14365 9321 14368
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 9398 14356 9404 14408
rect 9456 14405 9462 14408
rect 9456 14396 9464 14405
rect 9456 14368 9501 14396
rect 9456 14359 9464 14368
rect 9456 14356 9462 14359
rect 8536 14300 9168 14328
rect 9217 14331 9275 14337
rect 8536 14288 8542 14300
rect 9217 14297 9229 14331
rect 9263 14328 9275 14331
rect 9490 14328 9496 14340
rect 9263 14300 9496 14328
rect 9263 14297 9275 14300
rect 9217 14291 9275 14297
rect 9490 14288 9496 14300
rect 9548 14328 9554 14340
rect 9968 14328 9996 14436
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 12158 14464 12164 14476
rect 11756 14436 12164 14464
rect 11756 14424 11762 14436
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 14918 14464 14924 14476
rect 14879 14436 14924 14464
rect 14918 14424 14924 14436
rect 14976 14424 14982 14476
rect 16114 14464 16120 14476
rect 15028 14436 16120 14464
rect 10042 14356 10048 14408
rect 10100 14396 10106 14408
rect 10781 14399 10839 14405
rect 10781 14396 10793 14399
rect 10100 14368 10793 14396
rect 10100 14356 10106 14368
rect 10781 14365 10793 14368
rect 10827 14365 10839 14399
rect 10781 14359 10839 14365
rect 10870 14356 10876 14408
rect 10928 14396 10934 14408
rect 10965 14399 11023 14405
rect 10965 14396 10977 14399
rect 10928 14368 10977 14396
rect 10928 14356 10934 14368
rect 10965 14365 10977 14368
rect 11011 14365 11023 14399
rect 11514 14396 11520 14408
rect 11475 14368 11520 14396
rect 10965 14359 11023 14365
rect 11514 14356 11520 14368
rect 11572 14356 11578 14408
rect 12428 14399 12486 14405
rect 12428 14365 12440 14399
rect 12474 14396 12486 14399
rect 13262 14396 13268 14408
rect 12474 14368 13268 14396
rect 12474 14365 12486 14368
rect 12428 14359 12486 14365
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 14642 14396 14648 14408
rect 14603 14368 14648 14396
rect 14642 14356 14648 14368
rect 14700 14356 14706 14408
rect 14826 14396 14832 14408
rect 14787 14368 14832 14396
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 15028 14405 15056 14436
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 16298 14464 16304 14476
rect 16259 14436 16304 14464
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 16758 14464 16764 14476
rect 16500 14436 16764 14464
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14365 15071 14399
rect 15013 14359 15071 14365
rect 15194 14356 15200 14408
rect 15252 14396 15258 14408
rect 16209 14399 16267 14405
rect 15252 14368 15345 14396
rect 15252 14356 15258 14368
rect 16209 14365 16221 14399
rect 16255 14396 16267 14399
rect 16390 14396 16396 14408
rect 16255 14368 16396 14396
rect 16255 14365 16267 14368
rect 16209 14359 16267 14365
rect 16390 14356 16396 14368
rect 16448 14356 16454 14408
rect 16500 14405 16528 14436
rect 16758 14424 16764 14436
rect 16816 14424 16822 14476
rect 17218 14464 17224 14476
rect 17144 14436 17224 14464
rect 16485 14399 16543 14405
rect 16485 14365 16497 14399
rect 16531 14365 16543 14399
rect 16485 14359 16543 14365
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14396 16635 14399
rect 17144 14396 17172 14436
rect 17218 14424 17224 14436
rect 17276 14424 17282 14476
rect 17402 14464 17408 14476
rect 17363 14436 17408 14464
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 17865 14467 17923 14473
rect 17865 14433 17877 14467
rect 17911 14464 17923 14467
rect 29638 14464 29644 14476
rect 17911 14436 29644 14464
rect 17911 14433 17923 14436
rect 17865 14427 17923 14433
rect 29638 14424 29644 14436
rect 29696 14424 29702 14476
rect 17310 14396 17316 14408
rect 16623 14368 17172 14396
rect 17271 14368 17316 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 17586 14396 17592 14408
rect 17547 14368 17592 14396
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14396 17739 14399
rect 17954 14396 17960 14408
rect 17727 14368 17960 14396
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 18322 14396 18328 14408
rect 18283 14368 18328 14396
rect 18322 14356 18328 14368
rect 18380 14356 18386 14408
rect 19794 14396 19800 14408
rect 19755 14368 19800 14396
rect 19794 14356 19800 14368
rect 19852 14356 19858 14408
rect 20070 14396 20076 14408
rect 20031 14368 20076 14396
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14396 20223 14399
rect 20622 14396 20628 14408
rect 20211 14368 20628 14396
rect 20211 14365 20223 14368
rect 20165 14359 20223 14365
rect 20622 14356 20628 14368
rect 20680 14356 20686 14408
rect 20809 14399 20867 14405
rect 20809 14365 20821 14399
rect 20855 14396 20867 14399
rect 21174 14396 21180 14408
rect 20855 14368 21180 14396
rect 20855 14365 20867 14368
rect 20809 14359 20867 14365
rect 21174 14356 21180 14368
rect 21232 14356 21238 14408
rect 29917 14399 29975 14405
rect 29917 14396 29929 14399
rect 26206 14368 29929 14396
rect 10134 14328 10140 14340
rect 9548 14300 9996 14328
rect 10095 14300 10140 14328
rect 9548 14288 9554 14300
rect 10134 14288 10140 14300
rect 10192 14288 10198 14340
rect 10318 14328 10324 14340
rect 10279 14300 10324 14328
rect 10318 14288 10324 14300
rect 10376 14288 10382 14340
rect 13078 14288 13084 14340
rect 13136 14328 13142 14340
rect 15212 14328 15240 14356
rect 13136 14300 15240 14328
rect 16761 14331 16819 14337
rect 13136 14288 13142 14300
rect 16761 14297 16773 14331
rect 16807 14328 16819 14331
rect 26206 14328 26234 14368
rect 29917 14365 29929 14368
rect 29963 14365 29975 14399
rect 30098 14396 30104 14408
rect 30059 14368 30104 14396
rect 29917 14359 29975 14365
rect 30098 14356 30104 14368
rect 30156 14356 30162 14408
rect 16807 14300 26234 14328
rect 16807 14297 16819 14300
rect 16761 14291 16819 14297
rect 9674 14260 9680 14272
rect 8404 14232 9680 14260
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 10594 14220 10600 14272
rect 10652 14260 10658 14272
rect 10873 14263 10931 14269
rect 10873 14260 10885 14263
rect 10652 14232 10885 14260
rect 10652 14220 10658 14232
rect 10873 14229 10885 14232
rect 10919 14229 10931 14263
rect 10873 14223 10931 14229
rect 11701 14263 11759 14269
rect 11701 14229 11713 14263
rect 11747 14260 11759 14263
rect 12434 14260 12440 14272
rect 11747 14232 12440 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 16206 14220 16212 14272
rect 16264 14260 16270 14272
rect 18322 14260 18328 14272
rect 16264 14232 18328 14260
rect 16264 14220 16270 14232
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 20714 14220 20720 14272
rect 20772 14260 20778 14272
rect 21039 14263 21097 14269
rect 21039 14260 21051 14263
rect 20772 14232 21051 14260
rect 20772 14220 20778 14232
rect 21039 14229 21051 14232
rect 21085 14229 21097 14263
rect 21039 14223 21097 14229
rect 1104 14170 30820 14192
rect 1104 14118 10880 14170
rect 10932 14118 10944 14170
rect 10996 14118 11008 14170
rect 11060 14118 11072 14170
rect 11124 14118 11136 14170
rect 11188 14118 20811 14170
rect 20863 14118 20875 14170
rect 20927 14118 20939 14170
rect 20991 14118 21003 14170
rect 21055 14118 21067 14170
rect 21119 14118 30820 14170
rect 1104 14096 30820 14118
rect 1670 14016 1676 14068
rect 1728 14016 1734 14068
rect 1762 14016 1768 14068
rect 1820 14056 1826 14068
rect 2777 14059 2835 14065
rect 2777 14056 2789 14059
rect 1820 14028 2789 14056
rect 1820 14016 1826 14028
rect 2777 14025 2789 14028
rect 2823 14056 2835 14059
rect 5721 14059 5779 14065
rect 2823 14028 4936 14056
rect 2823 14025 2835 14028
rect 2777 14019 2835 14025
rect 1688 13988 1716 14016
rect 3786 13988 3792 14000
rect 1412 13960 3792 13988
rect 1412 13929 1440 13960
rect 3786 13948 3792 13960
rect 3844 13948 3850 14000
rect 1397 13923 1455 13929
rect 1397 13889 1409 13923
rect 1443 13889 1455 13923
rect 1397 13883 1455 13889
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1653 13923 1711 13929
rect 1653 13920 1665 13923
rect 1544 13892 1665 13920
rect 1544 13880 1550 13892
rect 1653 13889 1665 13892
rect 1699 13889 1711 13923
rect 1653 13883 1711 13889
rect 3050 13880 3056 13932
rect 3108 13920 3114 13932
rect 4908 13929 4936 14028
rect 5721 14025 5733 14059
rect 5767 14056 5779 14059
rect 5902 14056 5908 14068
rect 5767 14028 5908 14056
rect 5767 14025 5779 14028
rect 5721 14019 5779 14025
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 7101 14059 7159 14065
rect 7101 14025 7113 14059
rect 7147 14056 7159 14059
rect 11422 14056 11428 14068
rect 7147 14028 11428 14056
rect 7147 14025 7159 14028
rect 7101 14019 7159 14025
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 11701 14059 11759 14065
rect 11701 14056 11713 14059
rect 11572 14028 11713 14056
rect 11572 14016 11578 14028
rect 11701 14025 11713 14028
rect 11747 14025 11759 14059
rect 17586 14056 17592 14068
rect 11701 14019 11759 14025
rect 12406 14028 17592 14056
rect 6454 13948 6460 14000
rect 6512 13948 6518 14000
rect 7558 13948 7564 14000
rect 7616 13988 7622 14000
rect 12406 13988 12434 14028
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 18414 14016 18420 14068
rect 18472 14056 18478 14068
rect 19153 14059 19211 14065
rect 19153 14056 19165 14059
rect 18472 14028 19165 14056
rect 18472 14016 18478 14028
rect 19153 14025 19165 14028
rect 19199 14025 19211 14059
rect 19153 14019 19211 14025
rect 29822 14016 29828 14068
rect 29880 14056 29886 14068
rect 30009 14059 30067 14065
rect 30009 14056 30021 14059
rect 29880 14028 30021 14056
rect 29880 14016 29886 14028
rect 30009 14025 30021 14028
rect 30055 14025 30067 14059
rect 30009 14019 30067 14025
rect 12802 13988 12808 14000
rect 7616 13960 12434 13988
rect 12763 13960 12808 13988
rect 7616 13948 7622 13960
rect 12802 13948 12808 13960
rect 12860 13948 12866 14000
rect 13814 13948 13820 14000
rect 13872 13988 13878 14000
rect 14550 13988 14556 14000
rect 13872 13960 14556 13988
rect 13872 13948 13878 13960
rect 14550 13948 14556 13960
rect 14608 13948 14614 14000
rect 15470 13948 15476 14000
rect 15528 13988 15534 14000
rect 15565 13991 15623 13997
rect 15565 13988 15577 13991
rect 15528 13960 15577 13988
rect 15528 13948 15534 13960
rect 15565 13957 15577 13960
rect 15611 13957 15623 13991
rect 21174 13988 21180 14000
rect 15565 13951 15623 13957
rect 15672 13960 17632 13988
rect 3605 13923 3663 13929
rect 3605 13920 3617 13923
rect 3108 13892 3617 13920
rect 3108 13880 3114 13892
rect 3605 13889 3617 13892
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 4982 13880 4988 13932
rect 5040 13920 5046 13932
rect 5629 13923 5687 13929
rect 5040 13892 5085 13920
rect 5040 13880 5046 13892
rect 5629 13889 5641 13923
rect 5675 13920 5687 13923
rect 6353 13923 6411 13929
rect 5675 13892 6316 13920
rect 5675 13889 5687 13892
rect 5629 13883 5687 13889
rect 3329 13855 3387 13861
rect 3329 13821 3341 13855
rect 3375 13852 3387 13855
rect 3418 13852 3424 13864
rect 3375 13824 3424 13852
rect 3375 13821 3387 13824
rect 3329 13815 3387 13821
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 6288 13784 6316 13892
rect 6353 13889 6365 13923
rect 6399 13889 6411 13923
rect 6472 13920 6500 13948
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 6472 13892 6561 13920
rect 6353 13883 6411 13889
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6380 13852 6408 13883
rect 6638 13880 6644 13932
rect 6696 13920 6702 13932
rect 6696 13892 6741 13920
rect 6696 13880 6702 13892
rect 6822 13880 6828 13932
rect 6880 13920 6886 13932
rect 6917 13923 6975 13929
rect 6917 13920 6929 13923
rect 6880 13892 6929 13920
rect 6880 13880 6886 13892
rect 6917 13889 6929 13892
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 8297 13923 8355 13929
rect 8297 13889 8309 13923
rect 8343 13920 8355 13923
rect 8754 13920 8760 13932
rect 8343 13892 8760 13920
rect 8343 13889 8355 13892
rect 8297 13883 8355 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13920 8999 13923
rect 9674 13920 9680 13932
rect 8987 13892 9680 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 10042 13920 10048 13932
rect 10003 13892 10048 13920
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10502 13880 10508 13932
rect 10560 13920 10566 13932
rect 10597 13923 10655 13929
rect 10597 13920 10609 13923
rect 10560 13892 10609 13920
rect 10560 13880 10566 13892
rect 10597 13889 10609 13892
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12621 13923 12679 13929
rect 11931 13892 12434 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 6454 13852 6460 13864
rect 6380 13824 6460 13852
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 6733 13855 6791 13861
rect 6733 13821 6745 13855
rect 6779 13852 6791 13855
rect 7006 13852 7012 13864
rect 6779 13824 7012 13852
rect 6779 13821 6791 13824
rect 6733 13815 6791 13821
rect 6748 13784 6776 13815
rect 7006 13812 7012 13824
rect 7064 13852 7070 13864
rect 7558 13852 7564 13864
rect 7064 13824 7564 13852
rect 7064 13812 7070 13824
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 7834 13812 7840 13864
rect 7892 13852 7898 13864
rect 7892 13824 7972 13852
rect 7892 13812 7898 13824
rect 6288 13756 6776 13784
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 7374 13716 7380 13728
rect 4028 13688 7380 13716
rect 4028 13676 4034 13688
rect 7374 13676 7380 13688
rect 7432 13676 7438 13728
rect 7944 13716 7972 13824
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 8846 13852 8852 13864
rect 8444 13824 8852 13852
rect 8444 13812 8450 13824
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 9125 13855 9183 13861
rect 9125 13821 9137 13855
rect 9171 13852 9183 13855
rect 9582 13852 9588 13864
rect 9171 13824 9588 13852
rect 9171 13821 9183 13824
rect 9125 13815 9183 13821
rect 9582 13812 9588 13824
rect 9640 13852 9646 13864
rect 9950 13852 9956 13864
rect 9640 13824 9956 13852
rect 9640 13812 9646 13824
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 12066 13852 12072 13864
rect 12027 13824 12072 13852
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 12406 13852 12434 13892
rect 12621 13889 12633 13923
rect 12667 13920 12679 13923
rect 13078 13920 13084 13932
rect 12667 13892 13084 13920
rect 12667 13889 12679 13892
rect 12621 13883 12679 13889
rect 13078 13880 13084 13892
rect 13136 13880 13142 13932
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13920 13599 13923
rect 13722 13920 13728 13932
rect 13587 13892 13728 13920
rect 13587 13889 13599 13892
rect 13541 13883 13599 13889
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 15102 13920 15108 13932
rect 15063 13892 15108 13920
rect 15102 13880 15108 13892
rect 15160 13920 15166 13932
rect 15672 13920 15700 13960
rect 16850 13920 16856 13932
rect 15160 13892 15700 13920
rect 16811 13892 16856 13920
rect 15160 13880 15166 13892
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 17034 13880 17040 13932
rect 17092 13920 17098 13932
rect 17604 13929 17632 13960
rect 19720 13960 21180 13988
rect 17129 13923 17187 13929
rect 17129 13920 17141 13923
rect 17092 13892 17141 13920
rect 17092 13880 17098 13892
rect 17129 13889 17141 13892
rect 17175 13889 17187 13923
rect 17129 13883 17187 13889
rect 17589 13923 17647 13929
rect 17589 13889 17601 13923
rect 17635 13889 17647 13923
rect 17589 13883 17647 13889
rect 17773 13923 17831 13929
rect 17773 13889 17785 13923
rect 17819 13920 17831 13923
rect 18322 13920 18328 13932
rect 17819 13892 18328 13920
rect 17819 13889 17831 13892
rect 17773 13883 17831 13889
rect 18322 13880 18328 13892
rect 18380 13880 18386 13932
rect 18506 13880 18512 13932
rect 18564 13920 18570 13932
rect 18601 13923 18659 13929
rect 18601 13920 18613 13923
rect 18564 13892 18613 13920
rect 18564 13880 18570 13892
rect 18601 13889 18613 13892
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 19337 13923 19395 13929
rect 19337 13889 19349 13923
rect 19383 13920 19395 13923
rect 19720 13920 19748 13960
rect 21174 13948 21180 13960
rect 21232 13948 21238 14000
rect 19383 13892 19748 13920
rect 19383 13889 19395 13892
rect 19337 13883 19395 13889
rect 19794 13880 19800 13932
rect 19852 13920 19858 13932
rect 20257 13923 20315 13929
rect 20257 13920 20269 13923
rect 19852 13892 20269 13920
rect 19852 13880 19858 13892
rect 20257 13889 20269 13892
rect 20303 13920 20315 13923
rect 20346 13920 20352 13932
rect 20303 13892 20352 13920
rect 20303 13889 20315 13892
rect 20257 13883 20315 13889
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13889 20591 13923
rect 20533 13883 20591 13889
rect 20625 13923 20683 13929
rect 20625 13889 20637 13923
rect 20671 13920 20683 13923
rect 20714 13920 20720 13932
rect 20671 13892 20720 13920
rect 20671 13889 20683 13892
rect 20625 13883 20683 13889
rect 13354 13852 13360 13864
rect 12406 13824 13360 13852
rect 13354 13812 13360 13824
rect 13412 13812 13418 13864
rect 16574 13812 16580 13864
rect 16632 13852 16638 13864
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 16632 13824 16957 13852
rect 16632 13812 16638 13824
rect 16945 13821 16957 13824
rect 16991 13821 17003 13855
rect 16945 13815 17003 13821
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 20548 13852 20576 13883
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 29914 13920 29920 13932
rect 29875 13892 29920 13920
rect 29914 13880 29920 13892
rect 29972 13880 29978 13932
rect 30098 13920 30104 13932
rect 30059 13892 30104 13920
rect 30098 13880 30104 13892
rect 30156 13880 30162 13932
rect 17920 13824 20576 13852
rect 20809 13855 20867 13861
rect 17920 13812 17926 13824
rect 20809 13821 20821 13855
rect 20855 13852 20867 13855
rect 29270 13852 29276 13864
rect 20855 13824 29276 13852
rect 20855 13821 20867 13824
rect 20809 13815 20867 13821
rect 29270 13812 29276 13824
rect 29328 13812 29334 13864
rect 8018 13744 8024 13796
rect 8076 13784 8082 13796
rect 8113 13787 8171 13793
rect 8113 13784 8125 13787
rect 8076 13756 8125 13784
rect 8076 13744 8082 13756
rect 8113 13753 8125 13756
rect 8159 13753 8171 13787
rect 8113 13747 8171 13753
rect 8202 13744 8208 13796
rect 8260 13784 8266 13796
rect 15746 13784 15752 13796
rect 8260 13756 15752 13784
rect 8260 13744 8266 13756
rect 15746 13744 15752 13756
rect 15804 13744 15810 13796
rect 18414 13784 18420 13796
rect 17144 13756 18420 13784
rect 9861 13719 9919 13725
rect 9861 13716 9873 13719
rect 7944 13688 9873 13716
rect 9861 13685 9873 13688
rect 9907 13685 9919 13719
rect 9861 13679 9919 13685
rect 10781 13719 10839 13725
rect 10781 13685 10793 13719
rect 10827 13716 10839 13719
rect 11238 13716 11244 13728
rect 10827 13688 11244 13716
rect 10827 13685 10839 13688
rect 10781 13679 10839 13685
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 12802 13676 12808 13728
rect 12860 13716 12866 13728
rect 13449 13719 13507 13725
rect 13449 13716 13461 13719
rect 12860 13688 13461 13716
rect 12860 13676 12866 13688
rect 13449 13685 13461 13688
rect 13495 13685 13507 13719
rect 16666 13716 16672 13728
rect 16627 13688 16672 13716
rect 13449 13679 13507 13685
rect 16666 13676 16672 13688
rect 16724 13676 16730 13728
rect 17144 13725 17172 13756
rect 18414 13744 18420 13756
rect 18472 13744 18478 13796
rect 18598 13744 18604 13796
rect 18656 13784 18662 13796
rect 20349 13787 20407 13793
rect 20349 13784 20361 13787
rect 18656 13756 20361 13784
rect 18656 13744 18662 13756
rect 20349 13753 20361 13756
rect 20395 13753 20407 13787
rect 20349 13747 20407 13753
rect 17129 13719 17187 13725
rect 17129 13685 17141 13719
rect 17175 13685 17187 13719
rect 17129 13679 17187 13685
rect 17218 13676 17224 13728
rect 17276 13716 17282 13728
rect 17770 13716 17776 13728
rect 17276 13688 17776 13716
rect 17276 13676 17282 13688
rect 17770 13676 17776 13688
rect 17828 13716 17834 13728
rect 17865 13719 17923 13725
rect 17865 13716 17877 13719
rect 17828 13688 17877 13716
rect 17828 13676 17834 13688
rect 17865 13685 17877 13688
rect 17911 13685 17923 13719
rect 18506 13716 18512 13728
rect 18467 13688 18512 13716
rect 17865 13679 17923 13685
rect 18506 13676 18512 13688
rect 18564 13676 18570 13728
rect 1104 13626 30820 13648
rect 1104 13574 5915 13626
rect 5967 13574 5979 13626
rect 6031 13574 6043 13626
rect 6095 13574 6107 13626
rect 6159 13574 6171 13626
rect 6223 13574 15846 13626
rect 15898 13574 15910 13626
rect 15962 13574 15974 13626
rect 16026 13574 16038 13626
rect 16090 13574 16102 13626
rect 16154 13574 25776 13626
rect 25828 13574 25840 13626
rect 25892 13574 25904 13626
rect 25956 13574 25968 13626
rect 26020 13574 26032 13626
rect 26084 13574 30820 13626
rect 1104 13552 30820 13574
rect 4157 13515 4215 13521
rect 4157 13481 4169 13515
rect 4203 13512 4215 13515
rect 5350 13512 5356 13524
rect 4203 13484 5356 13512
rect 4203 13481 4215 13484
rect 4157 13475 4215 13481
rect 5350 13472 5356 13484
rect 5408 13512 5414 13524
rect 9306 13512 9312 13524
rect 5408 13484 9312 13512
rect 5408 13472 5414 13484
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 9582 13472 9588 13524
rect 9640 13512 9646 13524
rect 9677 13515 9735 13521
rect 9677 13512 9689 13515
rect 9640 13484 9689 13512
rect 9640 13472 9646 13484
rect 9677 13481 9689 13484
rect 9723 13481 9735 13515
rect 9677 13475 9735 13481
rect 9861 13515 9919 13521
rect 9861 13481 9873 13515
rect 9907 13512 9919 13515
rect 10042 13512 10048 13524
rect 9907 13484 10048 13512
rect 9907 13481 9919 13484
rect 9861 13475 9919 13481
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 11701 13515 11759 13521
rect 10152 13484 11275 13512
rect 6457 13447 6515 13453
rect 6457 13413 6469 13447
rect 6503 13444 6515 13447
rect 10152 13444 10180 13484
rect 6503 13416 10180 13444
rect 11247 13444 11275 13484
rect 11701 13481 11713 13515
rect 11747 13512 11759 13515
rect 12066 13512 12072 13524
rect 11747 13484 12072 13512
rect 11747 13481 11759 13484
rect 11701 13475 11759 13481
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 16298 13512 16304 13524
rect 12406 13484 16304 13512
rect 12406 13444 12434 13484
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 18233 13515 18291 13521
rect 18233 13512 18245 13515
rect 17552 13484 18245 13512
rect 17552 13472 17558 13484
rect 18233 13481 18245 13484
rect 18279 13512 18291 13515
rect 18506 13512 18512 13524
rect 18279 13484 18512 13512
rect 18279 13481 18291 13484
rect 18233 13475 18291 13481
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 19702 13512 19708 13524
rect 19615 13484 19708 13512
rect 19702 13472 19708 13484
rect 19760 13512 19766 13524
rect 20254 13512 20260 13524
rect 19760 13484 20260 13512
rect 19760 13472 19766 13484
rect 20254 13472 20260 13484
rect 20312 13472 20318 13524
rect 14458 13444 14464 13456
rect 11247 13416 12434 13444
rect 14419 13416 14464 13444
rect 6503 13413 6515 13416
rect 6457 13407 6515 13413
rect 14458 13404 14464 13416
rect 14516 13404 14522 13456
rect 15746 13444 15752 13456
rect 15707 13416 15752 13444
rect 15746 13404 15752 13416
rect 15804 13404 15810 13456
rect 19610 13444 19616 13456
rect 15856 13416 19616 13444
rect 2225 13379 2283 13385
rect 2225 13345 2237 13379
rect 2271 13376 2283 13379
rect 3234 13376 3240 13388
rect 2271 13348 3240 13376
rect 2271 13345 2283 13348
rect 2225 13339 2283 13345
rect 3234 13336 3240 13348
rect 3292 13376 3298 13388
rect 3970 13376 3976 13388
rect 3292 13348 3976 13376
rect 3292 13336 3298 13348
rect 3970 13336 3976 13348
rect 4028 13336 4034 13388
rect 5997 13379 6055 13385
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6638 13376 6644 13388
rect 6043 13348 6644 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 6638 13336 6644 13348
rect 6696 13376 6702 13388
rect 7193 13379 7251 13385
rect 7193 13376 7205 13379
rect 6696 13348 7205 13376
rect 6696 13336 6702 13348
rect 7193 13345 7205 13348
rect 7239 13345 7251 13379
rect 7193 13339 7251 13345
rect 7374 13336 7380 13388
rect 7432 13376 7438 13388
rect 9858 13376 9864 13388
rect 7432 13348 9864 13376
rect 7432 13336 7438 13348
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 13081 13379 13139 13385
rect 13081 13345 13093 13379
rect 13127 13376 13139 13379
rect 13814 13376 13820 13388
rect 13127 13348 13820 13376
rect 13127 13345 13139 13348
rect 13081 13339 13139 13345
rect 13814 13336 13820 13348
rect 13872 13376 13878 13388
rect 15856 13376 15884 13416
rect 19610 13404 19616 13416
rect 19668 13404 19674 13456
rect 13872 13348 15884 13376
rect 13872 13336 13878 13348
rect 16022 13336 16028 13388
rect 16080 13376 16086 13388
rect 20441 13379 20499 13385
rect 20441 13376 20453 13379
rect 16080 13348 20453 13376
rect 16080 13336 16086 13348
rect 20441 13345 20453 13348
rect 20487 13345 20499 13379
rect 20441 13339 20499 13345
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 2498 13308 2504 13320
rect 2459 13280 2504 13308
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 3510 13268 3516 13320
rect 3568 13308 3574 13320
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 3568 13280 4077 13308
rect 3568 13268 3574 13280
rect 4065 13277 4077 13280
rect 4111 13308 4123 13311
rect 4246 13308 4252 13320
rect 4111 13280 4252 13308
rect 4111 13277 4123 13280
rect 4065 13271 4123 13277
rect 4246 13268 4252 13280
rect 4304 13268 4310 13320
rect 5721 13311 5779 13317
rect 5721 13277 5733 13311
rect 5767 13277 5779 13311
rect 5902 13308 5908 13320
rect 5863 13280 5908 13308
rect 5721 13271 5779 13277
rect 5166 13240 5172 13252
rect 5127 13212 5172 13240
rect 5166 13200 5172 13212
rect 5224 13200 5230 13252
rect 5736 13240 5764 13271
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 6086 13268 6092 13320
rect 6144 13308 6150 13320
rect 6270 13308 6276 13320
rect 6144 13280 6189 13308
rect 6231 13280 6276 13308
rect 6144 13268 6150 13280
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13308 6975 13311
rect 8202 13308 8208 13320
rect 6963 13280 8208 13308
rect 6963 13277 6975 13280
rect 6917 13271 6975 13277
rect 7208 13252 7236 13280
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 8478 13308 8484 13320
rect 8435 13280 8484 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 10318 13308 10324 13320
rect 10279 13280 10324 13308
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 10594 13317 10600 13320
rect 10588 13308 10600 13317
rect 10555 13280 10600 13308
rect 10588 13271 10600 13280
rect 10594 13268 10600 13271
rect 10652 13268 10658 13320
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 14921 13311 14979 13317
rect 14921 13308 14933 13311
rect 11388 13280 14933 13308
rect 11388 13268 11394 13280
rect 14921 13277 14933 13280
rect 14967 13308 14979 13311
rect 15010 13308 15016 13320
rect 14967 13280 15016 13308
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 15289 13311 15347 13317
rect 15289 13277 15301 13311
rect 15335 13308 15347 13311
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 15335 13280 16129 13308
rect 15335 13277 15347 13280
rect 15289 13271 15347 13277
rect 16117 13277 16129 13280
rect 16163 13308 16175 13311
rect 16666 13308 16672 13320
rect 16163 13280 16672 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 17126 13308 17132 13320
rect 17087 13280 17132 13308
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 17221 13311 17279 13317
rect 17221 13277 17233 13311
rect 17267 13277 17279 13311
rect 17494 13308 17500 13320
rect 17455 13280 17500 13308
rect 17221 13271 17279 13277
rect 6362 13240 6368 13252
rect 5736 13212 6368 13240
rect 6362 13200 6368 13212
rect 6420 13200 6426 13252
rect 7190 13200 7196 13252
rect 7248 13200 7254 13252
rect 9490 13240 9496 13252
rect 9451 13212 9496 13240
rect 9490 13200 9496 13212
rect 9548 13200 9554 13252
rect 9582 13200 9588 13252
rect 9640 13240 9646 13252
rect 12802 13240 12808 13252
rect 9640 13212 12434 13240
rect 12763 13212 12808 13240
rect 9640 13200 9646 13212
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 2682 13172 2688 13184
rect 1627 13144 2688 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 3786 13132 3792 13184
rect 3844 13172 3850 13184
rect 5077 13175 5135 13181
rect 5077 13172 5089 13175
rect 3844 13144 5089 13172
rect 3844 13132 3850 13144
rect 5077 13141 5089 13144
rect 5123 13172 5135 13175
rect 7006 13172 7012 13184
rect 5123 13144 7012 13172
rect 5123 13141 5135 13144
rect 5077 13135 5135 13141
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 8297 13175 8355 13181
rect 8297 13141 8309 13175
rect 8343 13172 8355 13175
rect 8386 13172 8392 13184
rect 8343 13144 8392 13172
rect 8343 13141 8355 13144
rect 8297 13135 8355 13141
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 9703 13175 9761 13181
rect 9703 13141 9715 13175
rect 9749 13172 9761 13175
rect 9858 13172 9864 13184
rect 9749 13144 9864 13172
rect 9749 13141 9761 13144
rect 9703 13135 9761 13141
rect 9858 13132 9864 13144
rect 9916 13172 9922 13184
rect 10042 13172 10048 13184
rect 9916 13144 10048 13172
rect 9916 13132 9922 13144
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 12406 13172 12434 13212
rect 12802 13200 12808 13212
rect 12860 13200 12866 13252
rect 14274 13240 14280 13252
rect 14235 13212 14280 13240
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 14642 13200 14648 13252
rect 14700 13240 14706 13252
rect 15102 13240 15108 13252
rect 14700 13212 15108 13240
rect 14700 13200 14706 13212
rect 15102 13200 15108 13212
rect 15160 13200 15166 13252
rect 15933 13243 15991 13249
rect 15933 13209 15945 13243
rect 15979 13209 15991 13243
rect 15933 13203 15991 13209
rect 12618 13172 12624 13184
rect 12406 13144 12624 13172
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 15470 13132 15476 13184
rect 15528 13172 15534 13184
rect 15948 13172 15976 13203
rect 16574 13200 16580 13252
rect 16632 13240 16638 13252
rect 16945 13243 17003 13249
rect 16945 13240 16957 13243
rect 16632 13212 16957 13240
rect 16632 13200 16638 13212
rect 16945 13209 16957 13212
rect 16991 13209 17003 13243
rect 16945 13203 17003 13209
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 17236 13240 17264 13271
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13277 17831 13311
rect 18230 13308 18236 13320
rect 18191 13280 18236 13308
rect 17773 13271 17831 13277
rect 17092 13212 17264 13240
rect 17788 13240 17816 13271
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 18325 13311 18383 13317
rect 18325 13277 18337 13311
rect 18371 13277 18383 13311
rect 18325 13271 18383 13277
rect 18340 13240 18368 13271
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19797 13311 19855 13317
rect 19797 13308 19809 13311
rect 19484 13280 19809 13308
rect 19484 13268 19490 13280
rect 19797 13277 19809 13280
rect 19843 13308 19855 13311
rect 19886 13308 19892 13320
rect 19843 13280 19892 13308
rect 19843 13277 19855 13280
rect 19797 13271 19855 13277
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 20346 13308 20352 13320
rect 20307 13280 20352 13308
rect 20346 13268 20352 13280
rect 20404 13268 20410 13320
rect 20625 13311 20683 13317
rect 20625 13277 20637 13311
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 17788 13212 18368 13240
rect 17092 13200 17098 13212
rect 15528 13144 15976 13172
rect 15528 13132 15534 13144
rect 16850 13132 16856 13184
rect 16908 13172 16914 13184
rect 17310 13172 17316 13184
rect 16908 13144 17316 13172
rect 16908 13132 16914 13144
rect 17310 13132 17316 13144
rect 17368 13172 17374 13184
rect 17788 13172 17816 13212
rect 18966 13200 18972 13252
rect 19024 13240 19030 13252
rect 20640 13240 20668 13271
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 29825 13311 29883 13317
rect 20772 13280 20817 13308
rect 20772 13268 20778 13280
rect 29825 13277 29837 13311
rect 29871 13308 29883 13311
rect 30098 13308 30104 13320
rect 29871 13280 30104 13308
rect 29871 13277 29883 13280
rect 29825 13271 29883 13277
rect 30098 13268 30104 13280
rect 30156 13268 30162 13320
rect 19024 13212 20668 13240
rect 20901 13243 20959 13249
rect 19024 13200 19030 13212
rect 20901 13209 20913 13243
rect 20947 13240 20959 13243
rect 29914 13240 29920 13252
rect 20947 13212 29920 13240
rect 20947 13209 20959 13212
rect 20901 13203 20959 13209
rect 29914 13200 29920 13212
rect 29972 13200 29978 13252
rect 18598 13172 18604 13184
rect 17368 13144 17816 13172
rect 18559 13144 18604 13172
rect 17368 13132 17374 13144
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 30006 13172 30012 13184
rect 29967 13144 30012 13172
rect 30006 13132 30012 13144
rect 30064 13132 30070 13184
rect 1104 13082 30820 13104
rect 1104 13030 10880 13082
rect 10932 13030 10944 13082
rect 10996 13030 11008 13082
rect 11060 13030 11072 13082
rect 11124 13030 11136 13082
rect 11188 13030 20811 13082
rect 20863 13030 20875 13082
rect 20927 13030 20939 13082
rect 20991 13030 21003 13082
rect 21055 13030 21067 13082
rect 21119 13030 30820 13082
rect 1104 13008 30820 13030
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 5629 12971 5687 12977
rect 5629 12968 5641 12971
rect 5224 12940 5641 12968
rect 5224 12928 5230 12940
rect 5629 12937 5641 12940
rect 5675 12968 5687 12971
rect 10134 12968 10140 12980
rect 5675 12940 10140 12968
rect 5675 12937 5687 12940
rect 5629 12931 5687 12937
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 16022 12968 16028 12980
rect 10244 12940 16028 12968
rect 5721 12903 5779 12909
rect 5721 12869 5733 12903
rect 5767 12900 5779 12903
rect 8294 12900 8300 12912
rect 5767 12872 8300 12900
rect 5767 12869 5779 12872
rect 5721 12863 5779 12869
rect 8294 12860 8300 12872
rect 8352 12860 8358 12912
rect 10244 12900 10272 12940
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 16117 12971 16175 12977
rect 16117 12937 16129 12971
rect 16163 12937 16175 12971
rect 16117 12931 16175 12937
rect 18325 12971 18383 12977
rect 18325 12937 18337 12971
rect 18371 12968 18383 12971
rect 18414 12968 18420 12980
rect 18371 12940 18420 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 9416 12872 10272 12900
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12801 1455 12835
rect 1397 12795 1455 12801
rect 1412 12708 1440 12795
rect 2774 12792 2780 12844
rect 2832 12832 2838 12844
rect 3053 12835 3111 12841
rect 2832 12804 2877 12832
rect 2832 12792 2838 12804
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 3142 12832 3148 12844
rect 3099 12804 3148 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3694 12792 3700 12844
rect 3752 12832 3758 12844
rect 3861 12835 3919 12841
rect 3861 12832 3873 12835
rect 3752 12804 3873 12832
rect 3752 12792 3758 12804
rect 3861 12801 3873 12804
rect 3907 12801 3919 12835
rect 3861 12795 3919 12801
rect 5810 12792 5816 12844
rect 5868 12832 5874 12844
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 5868 12804 6377 12832
rect 5868 12792 5874 12804
rect 6365 12801 6377 12804
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 1394 12656 1400 12708
rect 1452 12656 1458 12708
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 2774 12628 2780 12640
rect 1627 12600 2780 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 2774 12588 2780 12600
rect 2832 12588 2838 12640
rect 3620 12628 3648 12727
rect 5626 12724 5632 12776
rect 5684 12764 5690 12776
rect 6564 12764 6592 12795
rect 6638 12792 6644 12844
rect 6696 12832 6702 12844
rect 6914 12832 6920 12844
rect 6696 12804 6741 12832
rect 6875 12804 6920 12832
rect 6696 12792 6702 12804
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12832 7159 12835
rect 9416 12832 9444 12872
rect 10502 12860 10508 12912
rect 10560 12900 10566 12912
rect 10597 12903 10655 12909
rect 10597 12900 10609 12903
rect 10560 12872 10609 12900
rect 10560 12860 10566 12872
rect 10597 12869 10609 12872
rect 10643 12869 10655 12903
rect 10597 12863 10655 12869
rect 12158 12860 12164 12912
rect 12216 12900 12222 12912
rect 13081 12903 13139 12909
rect 13081 12900 13093 12903
rect 12216 12872 13093 12900
rect 12216 12860 12222 12872
rect 13081 12869 13093 12872
rect 13127 12869 13139 12903
rect 13081 12863 13139 12869
rect 15289 12903 15347 12909
rect 15289 12869 15301 12903
rect 15335 12900 15347 12903
rect 15562 12900 15568 12912
rect 15335 12872 15568 12900
rect 15335 12869 15347 12872
rect 15289 12863 15347 12869
rect 15562 12860 15568 12872
rect 15620 12900 15626 12912
rect 16132 12900 16160 12931
rect 18230 12900 18236 12912
rect 15620 12872 15884 12900
rect 16132 12872 18236 12900
rect 15620 12860 15626 12872
rect 7147 12804 9444 12832
rect 9493 12835 9551 12841
rect 7147 12801 7159 12804
rect 7101 12795 7159 12801
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 9582 12832 9588 12844
rect 9539 12804 9588 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 5684 12736 6592 12764
rect 6733 12767 6791 12773
rect 5684 12724 5690 12736
rect 6733 12733 6745 12767
rect 6779 12764 6791 12767
rect 8018 12764 8024 12776
rect 6779 12736 8024 12764
rect 6779 12733 6791 12736
rect 6733 12727 6791 12733
rect 6086 12656 6092 12708
rect 6144 12696 6150 12708
rect 6748 12696 6776 12727
rect 8018 12724 8024 12736
rect 8076 12724 8082 12776
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12733 8539 12767
rect 8754 12764 8760 12776
rect 8667 12736 8760 12764
rect 8481 12727 8539 12733
rect 6144 12668 6776 12696
rect 6144 12656 6150 12668
rect 7558 12656 7564 12708
rect 7616 12696 7622 12708
rect 8496 12696 8524 12727
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 9398 12724 9404 12776
rect 9456 12764 9462 12776
rect 9508 12764 9536 12795
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12832 9735 12835
rect 9858 12832 9864 12844
rect 9723 12804 9864 12832
rect 9723 12801 9735 12804
rect 9677 12795 9735 12801
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 11790 12792 11796 12844
rect 11848 12830 11854 12844
rect 11885 12835 11943 12841
rect 11885 12830 11897 12835
rect 11848 12802 11897 12830
rect 11848 12792 11854 12802
rect 11885 12801 11897 12802
rect 11931 12801 11943 12835
rect 12066 12832 12072 12844
rect 12027 12804 12072 12832
rect 11885 12795 11943 12801
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12832 12495 12835
rect 12986 12832 12992 12844
rect 12483 12804 12992 12832
rect 12483 12801 12495 12804
rect 12437 12795 12495 12801
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12832 13323 12835
rect 14274 12832 14280 12844
rect 13311 12804 14280 12832
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 15010 12832 15016 12844
rect 14971 12804 15016 12832
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 15749 12835 15807 12841
rect 15749 12801 15761 12835
rect 15795 12801 15807 12835
rect 15749 12795 15807 12801
rect 9456 12736 9536 12764
rect 10781 12767 10839 12773
rect 9456 12724 9462 12736
rect 10781 12733 10793 12767
rect 10827 12764 10839 12767
rect 11974 12764 11980 12776
rect 10827 12736 11980 12764
rect 10827 12733 10839 12736
rect 10781 12727 10839 12733
rect 11974 12724 11980 12736
rect 12032 12764 12038 12776
rect 12161 12767 12219 12773
rect 12161 12764 12173 12767
rect 12032 12736 12173 12764
rect 12032 12724 12038 12736
rect 12161 12733 12173 12736
rect 12207 12733 12219 12767
rect 12161 12727 12219 12733
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12733 12311 12767
rect 12253 12727 12311 12733
rect 7616 12668 8524 12696
rect 8772 12696 8800 12724
rect 11330 12696 11336 12708
rect 8772 12668 11336 12696
rect 7616 12656 7622 12668
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 11882 12656 11888 12708
rect 11940 12696 11946 12708
rect 12268 12696 12296 12727
rect 11940 12668 12296 12696
rect 15764 12696 15792 12795
rect 15856 12764 15884 12872
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12832 15991 12835
rect 16206 12832 16212 12844
rect 15979 12804 16212 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 16206 12792 16212 12804
rect 16264 12792 16270 12844
rect 16868 12841 16896 12872
rect 18230 12860 18236 12872
rect 18288 12860 18294 12912
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12801 17095 12835
rect 17310 12832 17316 12844
rect 17271 12804 17316 12832
rect 17037 12795 17095 12801
rect 16482 12764 16488 12776
rect 15856 12736 16488 12764
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 16666 12764 16672 12776
rect 16627 12736 16672 12764
rect 16666 12724 16672 12736
rect 16724 12724 16730 12776
rect 17052 12764 17080 12795
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 18340 12764 18368 12931
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 30009 12971 30067 12977
rect 18748 12940 20300 12968
rect 18748 12928 18754 12940
rect 19334 12860 19340 12912
rect 19392 12900 19398 12912
rect 19438 12903 19496 12909
rect 19438 12900 19450 12903
rect 19392 12872 19450 12900
rect 19392 12860 19398 12872
rect 19438 12869 19450 12872
rect 19484 12869 19496 12903
rect 19438 12863 19496 12869
rect 19978 12860 19984 12912
rect 20036 12900 20042 12912
rect 20165 12903 20223 12909
rect 20165 12900 20177 12903
rect 20036 12872 20177 12900
rect 20036 12860 20042 12872
rect 20165 12869 20177 12872
rect 20211 12869 20223 12903
rect 20165 12863 20223 12869
rect 19610 12792 19616 12844
rect 19668 12832 19674 12844
rect 20272 12841 20300 12940
rect 30009 12937 30021 12971
rect 30055 12968 30067 12971
rect 30190 12968 30196 12980
rect 30055 12940 30196 12968
rect 30055 12937 30067 12940
rect 30009 12931 30067 12937
rect 30190 12928 30196 12940
rect 30248 12928 30254 12980
rect 19705 12835 19763 12841
rect 19705 12832 19717 12835
rect 19668 12804 19717 12832
rect 19668 12792 19674 12804
rect 19705 12801 19717 12804
rect 19751 12801 19763 12835
rect 19705 12795 19763 12801
rect 20257 12835 20315 12841
rect 20257 12801 20269 12835
rect 20303 12832 20315 12835
rect 21634 12832 21640 12844
rect 20303 12804 21640 12832
rect 20303 12801 20315 12804
rect 20257 12795 20315 12801
rect 21634 12792 21640 12804
rect 21692 12792 21698 12844
rect 29914 12832 29920 12844
rect 29875 12804 29920 12832
rect 29914 12792 29920 12804
rect 29972 12792 29978 12844
rect 30098 12832 30104 12844
rect 30059 12804 30104 12832
rect 30098 12792 30104 12804
rect 30156 12792 30162 12844
rect 17052 12736 18368 12764
rect 17034 12696 17040 12708
rect 15764 12668 17040 12696
rect 11940 12656 11946 12668
rect 17034 12656 17040 12668
rect 17092 12656 17098 12708
rect 3786 12628 3792 12640
rect 3620 12600 3792 12628
rect 3786 12588 3792 12600
rect 3844 12588 3850 12640
rect 4982 12628 4988 12640
rect 4943 12600 4988 12628
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 9309 12631 9367 12637
rect 9309 12597 9321 12631
rect 9355 12628 9367 12631
rect 9766 12628 9772 12640
rect 9355 12600 9772 12628
rect 9355 12597 9367 12600
rect 9309 12591 9367 12597
rect 9766 12588 9772 12600
rect 9824 12628 9830 12640
rect 10778 12628 10784 12640
rect 9824 12600 10784 12628
rect 9824 12588 9830 12600
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 12618 12628 12624 12640
rect 12579 12600 12624 12628
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 15470 12588 15476 12640
rect 15528 12628 15534 12640
rect 15749 12631 15807 12637
rect 15749 12628 15761 12631
rect 15528 12600 15761 12628
rect 15528 12588 15534 12600
rect 15749 12597 15761 12600
rect 15795 12597 15807 12631
rect 15749 12591 15807 12597
rect 16482 12588 16488 12640
rect 16540 12628 16546 12640
rect 18046 12628 18052 12640
rect 16540 12600 18052 12628
rect 16540 12588 16546 12600
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 1104 12538 30820 12560
rect 1104 12486 5915 12538
rect 5967 12486 5979 12538
rect 6031 12486 6043 12538
rect 6095 12486 6107 12538
rect 6159 12486 6171 12538
rect 6223 12486 15846 12538
rect 15898 12486 15910 12538
rect 15962 12486 15974 12538
rect 16026 12486 16038 12538
rect 16090 12486 16102 12538
rect 16154 12486 25776 12538
rect 25828 12486 25840 12538
rect 25892 12486 25904 12538
rect 25956 12486 25968 12538
rect 26020 12486 26032 12538
rect 26084 12486 30820 12538
rect 1104 12464 30820 12486
rect 5721 12427 5779 12433
rect 5721 12393 5733 12427
rect 5767 12424 5779 12427
rect 6270 12424 6276 12436
rect 5767 12396 6276 12424
rect 5767 12393 5779 12396
rect 5721 12387 5779 12393
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 6457 12427 6515 12433
rect 6457 12393 6469 12427
rect 6503 12424 6515 12427
rect 7098 12424 7104 12436
rect 6503 12396 7104 12424
rect 6503 12393 6515 12396
rect 6457 12387 6515 12393
rect 7098 12384 7104 12396
rect 7156 12424 7162 12436
rect 14185 12427 14243 12433
rect 7156 12396 12020 12424
rect 7156 12384 7162 12396
rect 3050 12316 3056 12368
rect 3108 12316 3114 12368
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12288 2927 12291
rect 3068 12288 3096 12316
rect 3786 12288 3792 12300
rect 2915 12260 3096 12288
rect 3747 12260 3792 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 3786 12248 3792 12260
rect 3844 12248 3850 12300
rect 7190 12288 7196 12300
rect 6564 12260 7196 12288
rect 1210 12180 1216 12232
rect 1268 12220 1274 12232
rect 1397 12223 1455 12229
rect 1397 12220 1409 12223
rect 1268 12192 1409 12220
rect 1268 12180 1274 12192
rect 1397 12189 1409 12192
rect 1443 12189 1455 12223
rect 2498 12220 2504 12232
rect 2459 12192 2504 12220
rect 1397 12183 1455 12189
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 2682 12220 2688 12232
rect 2643 12192 2688 12220
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12189 2835 12223
rect 2777 12183 2835 12189
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 2792 12152 2820 12183
rect 2866 12152 2872 12164
rect 2792 12124 2872 12152
rect 2866 12112 2872 12124
rect 2924 12112 2930 12164
rect 1581 12087 1639 12093
rect 1581 12053 1593 12087
rect 1627 12084 1639 12087
rect 2958 12084 2964 12096
rect 1627 12056 2964 12084
rect 1627 12053 1639 12056
rect 1581 12047 1639 12053
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 3068 12084 3096 12183
rect 5350 12180 5356 12232
rect 5408 12220 5414 12232
rect 6564 12229 6592 12260
rect 7190 12248 7196 12260
rect 7248 12288 7254 12300
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 7248 12260 7389 12288
rect 7248 12248 7254 12260
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 7377 12251 7435 12257
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12288 7527 12291
rect 7558 12288 7564 12300
rect 7515 12260 7564 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 8202 12248 8208 12300
rect 8260 12288 8266 12300
rect 8938 12288 8944 12300
rect 8260 12260 8944 12288
rect 8260 12248 8266 12260
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 11992 12288 12020 12396
rect 14185 12393 14197 12427
rect 14231 12424 14243 12427
rect 14274 12424 14280 12436
rect 14231 12396 14280 12424
rect 14231 12393 14243 12396
rect 14185 12387 14243 12393
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 16666 12424 16672 12436
rect 14568 12396 16672 12424
rect 12158 12316 12164 12368
rect 12216 12356 12222 12368
rect 14568 12356 14596 12396
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17865 12427 17923 12433
rect 17865 12424 17877 12427
rect 17000 12396 17877 12424
rect 17000 12384 17006 12396
rect 17865 12393 17877 12396
rect 17911 12393 17923 12427
rect 17865 12387 17923 12393
rect 18322 12356 18328 12368
rect 12216 12328 14596 12356
rect 15396 12328 18328 12356
rect 12216 12316 12222 12328
rect 15396 12288 15424 12328
rect 18322 12316 18328 12328
rect 18380 12356 18386 12368
rect 18417 12359 18475 12365
rect 18417 12356 18429 12359
rect 18380 12328 18429 12356
rect 18380 12316 18386 12328
rect 18417 12325 18429 12328
rect 18463 12325 18475 12359
rect 18417 12319 18475 12325
rect 11992 12260 15424 12288
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12288 15531 12291
rect 15654 12288 15660 12300
rect 15519 12260 15660 12288
rect 15519 12257 15531 12260
rect 15473 12251 15531 12257
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 18509 12291 18567 12297
rect 18509 12257 18521 12291
rect 18555 12288 18567 12291
rect 19334 12288 19340 12300
rect 18555 12260 19340 12288
rect 18555 12257 18567 12260
rect 18509 12251 18567 12257
rect 19334 12248 19340 12260
rect 19392 12248 19398 12300
rect 20533 12291 20591 12297
rect 20533 12257 20545 12291
rect 20579 12257 20591 12291
rect 20533 12251 20591 12257
rect 20993 12291 21051 12297
rect 20993 12257 21005 12291
rect 21039 12288 21051 12291
rect 29914 12288 29920 12300
rect 21039 12260 29920 12288
rect 21039 12257 21051 12260
rect 20993 12251 21051 12257
rect 5629 12223 5687 12229
rect 5629 12220 5641 12223
rect 5408 12192 5641 12220
rect 5408 12180 5414 12192
rect 5629 12189 5641 12192
rect 5675 12189 5687 12223
rect 5629 12183 5687 12189
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 7101 12223 7159 12229
rect 7101 12189 7113 12223
rect 7147 12189 7159 12223
rect 7101 12183 7159 12189
rect 7285 12223 7343 12229
rect 7285 12189 7297 12223
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 7653 12223 7711 12229
rect 7653 12189 7665 12223
rect 7699 12220 7711 12223
rect 7742 12220 7748 12232
rect 7699 12192 7748 12220
rect 7699 12189 7711 12192
rect 7653 12183 7711 12189
rect 3237 12155 3295 12161
rect 3237 12121 3249 12155
rect 3283 12152 3295 12155
rect 4034 12155 4092 12161
rect 4034 12152 4046 12155
rect 3283 12124 4046 12152
rect 3283 12121 3295 12124
rect 3237 12115 3295 12121
rect 4034 12121 4046 12124
rect 4080 12121 4092 12155
rect 4034 12115 4092 12121
rect 4890 12112 4896 12164
rect 4948 12152 4954 12164
rect 7116 12152 7144 12183
rect 4948 12124 7144 12152
rect 4948 12112 4954 12124
rect 5169 12087 5227 12093
rect 5169 12084 5181 12087
rect 3068 12056 5181 12084
rect 5169 12053 5181 12056
rect 5215 12084 5227 12087
rect 5626 12084 5632 12096
rect 5215 12056 5632 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5626 12044 5632 12056
rect 5684 12044 5690 12096
rect 7300 12084 7328 12183
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 10284 12192 10333 12220
rect 10284 12180 10290 12192
rect 10321 12189 10333 12192
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 10965 12223 11023 12229
rect 10965 12189 10977 12223
rect 11011 12220 11023 12223
rect 12250 12220 12256 12232
rect 11011 12192 12256 12220
rect 11011 12189 11023 12192
rect 10965 12183 11023 12189
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 12986 12180 12992 12232
rect 13044 12220 13050 12232
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 13044 12192 14841 12220
rect 13044 12180 13050 12192
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 15749 12223 15807 12229
rect 15749 12189 15761 12223
rect 15795 12220 15807 12223
rect 16298 12220 16304 12232
rect 15795 12192 16304 12220
rect 15795 12189 15807 12192
rect 15749 12183 15807 12189
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 16390 12180 16396 12232
rect 16448 12220 16454 12232
rect 17990 12223 18048 12229
rect 17990 12220 18002 12223
rect 16448 12192 18002 12220
rect 16448 12180 16454 12192
rect 17990 12189 18002 12192
rect 18036 12189 18048 12223
rect 17990 12183 18048 12189
rect 18598 12180 18604 12232
rect 18656 12220 18662 12232
rect 19058 12220 19064 12232
rect 18656 12192 19064 12220
rect 18656 12180 18662 12192
rect 19058 12180 19064 12192
rect 19116 12220 19122 12232
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 19116 12192 19441 12220
rect 19116 12180 19122 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19613 12223 19671 12229
rect 19613 12189 19625 12223
rect 19659 12220 19671 12223
rect 19702 12220 19708 12232
rect 19659 12192 19708 12220
rect 19659 12189 19671 12192
rect 19613 12183 19671 12189
rect 19702 12180 19708 12192
rect 19760 12180 19766 12232
rect 20346 12180 20352 12232
rect 20404 12220 20410 12232
rect 20441 12223 20499 12229
rect 20441 12220 20453 12223
rect 20404 12192 20453 12220
rect 20404 12180 20410 12192
rect 20441 12189 20453 12192
rect 20487 12189 20499 12223
rect 20441 12183 20499 12189
rect 7837 12155 7895 12161
rect 7837 12121 7849 12155
rect 7883 12152 7895 12155
rect 7883 12124 9352 12152
rect 7883 12121 7895 12124
rect 7837 12115 7895 12121
rect 8386 12084 8392 12096
rect 7300 12056 8392 12084
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 8941 12087 8999 12093
rect 8941 12053 8953 12087
rect 8987 12084 8999 12087
rect 9030 12084 9036 12096
rect 8987 12056 9036 12084
rect 8987 12053 8999 12056
rect 8941 12047 8999 12053
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 9324 12084 9352 12124
rect 9582 12112 9588 12164
rect 9640 12152 9646 12164
rect 11238 12161 11244 12164
rect 10054 12155 10112 12161
rect 10054 12152 10066 12155
rect 9640 12124 10066 12152
rect 9640 12112 9646 12124
rect 10054 12121 10066 12124
rect 10100 12121 10112 12155
rect 10054 12115 10112 12121
rect 11232 12115 11244 12161
rect 11296 12152 11302 12164
rect 11296 12124 11332 12152
rect 11238 12112 11244 12115
rect 11296 12112 11302 12124
rect 14182 12112 14188 12164
rect 14240 12152 14246 12164
rect 14277 12155 14335 12161
rect 14277 12152 14289 12155
rect 14240 12124 14289 12152
rect 14240 12112 14246 12124
rect 14277 12121 14289 12124
rect 14323 12121 14335 12155
rect 20548 12152 20576 12251
rect 29914 12248 29920 12260
rect 29972 12248 29978 12300
rect 20622 12180 20628 12232
rect 20680 12220 20686 12232
rect 20717 12223 20775 12229
rect 20717 12220 20729 12223
rect 20680 12192 20729 12220
rect 20680 12180 20686 12192
rect 20717 12189 20729 12192
rect 20763 12189 20775 12223
rect 20717 12183 20775 12189
rect 20806 12180 20812 12232
rect 20864 12220 20870 12232
rect 21450 12220 21456 12232
rect 20864 12192 20909 12220
rect 21411 12192 21456 12220
rect 20864 12180 20870 12192
rect 21450 12180 21456 12192
rect 21508 12180 21514 12232
rect 21634 12152 21640 12164
rect 14277 12115 14335 12121
rect 14384 12124 20576 12152
rect 21595 12124 21640 12152
rect 11330 12084 11336 12096
rect 9324 12056 11336 12084
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 12342 12084 12348 12096
rect 12303 12056 12348 12084
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 14384 12084 14412 12124
rect 21634 12112 21640 12124
rect 21692 12112 21698 12164
rect 12952 12056 14412 12084
rect 14921 12087 14979 12093
rect 12952 12044 12958 12056
rect 14921 12053 14933 12087
rect 14967 12084 14979 12087
rect 15654 12084 15660 12096
rect 14967 12056 15660 12084
rect 14967 12053 14979 12056
rect 14921 12047 14979 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 18046 12084 18052 12096
rect 18007 12056 18052 12084
rect 18046 12044 18052 12056
rect 18104 12044 18110 12096
rect 19797 12087 19855 12093
rect 19797 12053 19809 12087
rect 19843 12084 19855 12087
rect 19886 12084 19892 12096
rect 19843 12056 19892 12084
rect 19843 12053 19855 12056
rect 19797 12047 19855 12053
rect 19886 12044 19892 12056
rect 19944 12044 19950 12096
rect 21821 12087 21879 12093
rect 21821 12053 21833 12087
rect 21867 12084 21879 12087
rect 22186 12084 22192 12096
rect 21867 12056 22192 12084
rect 21867 12053 21879 12056
rect 21821 12047 21879 12053
rect 22186 12044 22192 12056
rect 22244 12044 22250 12096
rect 1104 11994 30820 12016
rect 1104 11942 10880 11994
rect 10932 11942 10944 11994
rect 10996 11942 11008 11994
rect 11060 11942 11072 11994
rect 11124 11942 11136 11994
rect 11188 11942 20811 11994
rect 20863 11942 20875 11994
rect 20927 11942 20939 11994
rect 20991 11942 21003 11994
rect 21055 11942 21067 11994
rect 21119 11942 30820 11994
rect 1104 11920 30820 11942
rect 3329 11883 3387 11889
rect 3329 11849 3341 11883
rect 3375 11880 3387 11883
rect 3694 11880 3700 11892
rect 3375 11852 3700 11880
rect 3375 11849 3387 11852
rect 3329 11843 3387 11849
rect 3694 11840 3700 11852
rect 3752 11840 3758 11892
rect 4798 11880 4804 11892
rect 4759 11852 4804 11880
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 6914 11880 6920 11892
rect 5767 11852 6920 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 8846 11880 8852 11892
rect 8807 11852 8852 11880
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 10965 11883 11023 11889
rect 8956 11852 9674 11880
rect 2498 11772 2504 11824
rect 2556 11812 2562 11824
rect 3786 11812 3792 11824
rect 2556 11784 3792 11812
rect 2556 11772 2562 11784
rect 1394 11744 1400 11756
rect 1355 11716 1400 11744
rect 1394 11704 1400 11716
rect 1452 11704 1458 11756
rect 2608 11753 2636 11784
rect 3786 11772 3792 11784
rect 3844 11772 3850 11824
rect 4614 11772 4620 11824
rect 4672 11812 4678 11824
rect 4709 11815 4767 11821
rect 4709 11812 4721 11815
rect 4672 11784 4721 11812
rect 4672 11772 4678 11784
rect 4709 11781 4721 11784
rect 4755 11781 4767 11815
rect 4816 11812 4844 11840
rect 8956 11812 8984 11852
rect 4816 11784 8984 11812
rect 9646 11812 9674 11852
rect 10965 11849 10977 11883
rect 11011 11880 11023 11883
rect 11238 11880 11244 11892
rect 11011 11852 11244 11880
rect 11011 11849 11023 11852
rect 10965 11843 11023 11849
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 12894 11880 12900 11892
rect 11388 11852 12900 11880
rect 11388 11840 11394 11852
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 12986 11840 12992 11892
rect 13044 11880 13050 11892
rect 13633 11883 13691 11889
rect 13633 11880 13645 11883
rect 13044 11852 13645 11880
rect 13044 11840 13050 11852
rect 13633 11849 13645 11852
rect 13679 11849 13691 11883
rect 13633 11843 13691 11849
rect 17402 11840 17408 11892
rect 17460 11880 17466 11892
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 17460 11852 17785 11880
rect 17460 11840 17466 11852
rect 17773 11849 17785 11852
rect 17819 11849 17831 11883
rect 17773 11843 17831 11849
rect 17957 11883 18015 11889
rect 17957 11849 17969 11883
rect 18003 11880 18015 11883
rect 18046 11880 18052 11892
rect 18003 11852 18052 11880
rect 18003 11849 18015 11852
rect 17957 11843 18015 11849
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 20622 11880 20628 11892
rect 20583 11852 20628 11880
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 9950 11812 9956 11824
rect 9646 11784 9956 11812
rect 4709 11775 4767 11781
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11713 2651 11747
rect 2593 11707 2651 11713
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 2961 11747 3019 11753
rect 2832 11716 2877 11744
rect 2832 11704 2838 11716
rect 2961 11713 2973 11747
rect 3007 11744 3019 11747
rect 3050 11744 3056 11756
rect 3007 11716 3056 11744
rect 3007 11713 3019 11716
rect 2961 11707 3019 11713
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11744 3203 11747
rect 4982 11744 4988 11756
rect 3191 11716 4988 11744
rect 3191 11713 3203 11716
rect 3145 11707 3203 11713
rect 4982 11704 4988 11716
rect 5040 11744 5046 11756
rect 5350 11744 5356 11756
rect 5040 11716 5356 11744
rect 5040 11704 5046 11716
rect 5350 11704 5356 11716
rect 5408 11704 5414 11756
rect 5626 11744 5632 11756
rect 5587 11716 5632 11744
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 7208 11753 7236 11784
rect 9950 11772 9956 11784
rect 10008 11812 10014 11824
rect 12342 11812 12348 11824
rect 10008 11784 10272 11812
rect 10008 11772 10014 11784
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11744 7527 11747
rect 7745 11747 7803 11753
rect 7515 11716 7697 11744
rect 7515 11713 7527 11716
rect 7469 11707 7527 11713
rect 2866 11676 2872 11688
rect 2779 11648 2872 11676
rect 2866 11636 2872 11648
rect 2924 11676 2930 11688
rect 4062 11676 4068 11688
rect 2924 11648 4068 11676
rect 2924 11636 2930 11648
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 2222 11568 2228 11620
rect 2280 11608 2286 11620
rect 7392 11608 7420 11707
rect 7558 11676 7564 11688
rect 7519 11648 7564 11676
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 2280 11580 7420 11608
rect 7669 11608 7697 11716
rect 7745 11713 7757 11747
rect 7791 11744 7803 11747
rect 8478 11744 8484 11756
rect 7791 11716 8484 11744
rect 7791 11713 7803 11716
rect 7745 11707 7803 11713
rect 8478 11704 8484 11716
rect 8536 11704 8542 11756
rect 8662 11744 8668 11756
rect 8623 11716 8668 11744
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 8987 11747 9045 11753
rect 8987 11744 8999 11747
rect 8904 11716 8999 11744
rect 8904 11704 8910 11716
rect 8987 11713 8999 11716
rect 9033 11713 9045 11747
rect 8987 11707 9045 11713
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 10244 11753 10272 11784
rect 10796 11784 12348 11812
rect 10229 11747 10287 11753
rect 9364 11716 9409 11744
rect 9364 11704 9370 11716
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 10410 11744 10416 11756
rect 10371 11716 10416 11744
rect 10229 11707 10287 11713
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 10502 11704 10508 11756
rect 10560 11744 10566 11756
rect 10796 11753 10824 11784
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 12520 11815 12578 11821
rect 12520 11781 12532 11815
rect 12566 11812 12578 11815
rect 12618 11812 12624 11824
rect 12566 11784 12624 11812
rect 12566 11781 12578 11784
rect 12520 11775 12578 11781
rect 12618 11772 12624 11784
rect 12676 11772 12682 11824
rect 14458 11812 14464 11824
rect 14108 11784 14464 11812
rect 14108 11756 14136 11784
rect 14458 11772 14464 11784
rect 14516 11772 14522 11824
rect 19058 11812 19064 11824
rect 19019 11784 19064 11812
rect 19058 11772 19064 11784
rect 19116 11772 19122 11824
rect 19245 11815 19303 11821
rect 19245 11781 19257 11815
rect 19291 11812 19303 11815
rect 19978 11812 19984 11824
rect 19291 11784 19984 11812
rect 19291 11781 19303 11784
rect 19245 11775 19303 11781
rect 19978 11772 19984 11784
rect 20036 11772 20042 11824
rect 10781 11747 10839 11753
rect 10560 11716 10605 11744
rect 10560 11704 10566 11716
rect 10781 11713 10793 11747
rect 10827 11713 10839 11747
rect 12250 11744 12256 11756
rect 12211 11716 12256 11744
rect 10781 11707 10839 11713
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 14090 11744 14096 11756
rect 14003 11716 14096 11744
rect 14090 11704 14096 11716
rect 14148 11704 14154 11756
rect 14366 11753 14372 11756
rect 14360 11707 14372 11753
rect 14424 11744 14430 11756
rect 14424 11716 14460 11744
rect 14366 11704 14372 11707
rect 14424 11704 14430 11716
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15344 11716 15945 11744
rect 15344 11704 15350 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16669 11747 16727 11753
rect 16669 11713 16681 11747
rect 16715 11713 16727 11747
rect 16669 11707 16727 11713
rect 10520 11676 10548 11704
rect 9508 11648 10548 11676
rect 10597 11679 10655 11685
rect 9508 11608 9536 11648
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 11882 11676 11888 11688
rect 10643 11648 11888 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 11882 11636 11888 11648
rect 11940 11636 11946 11688
rect 9858 11608 9864 11620
rect 7669 11580 9536 11608
rect 9646 11580 9864 11608
rect 2280 11568 2286 11580
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3970 11540 3976 11552
rect 3016 11512 3976 11540
rect 3016 11500 3022 11512
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 7282 11500 7288 11552
rect 7340 11540 7346 11552
rect 7929 11543 7987 11549
rect 7929 11540 7941 11543
rect 7340 11512 7941 11540
rect 7340 11500 7346 11512
rect 7929 11509 7941 11512
rect 7975 11509 7987 11543
rect 7929 11503 7987 11509
rect 9031 11500 9037 11552
rect 9089 11549 9095 11552
rect 9089 11543 9137 11549
rect 9089 11509 9091 11543
rect 9125 11509 9137 11543
rect 9089 11503 9137 11509
rect 9089 11500 9095 11503
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 9646 11540 9674 11580
rect 9858 11568 9864 11580
rect 9916 11608 9922 11620
rect 11238 11608 11244 11620
rect 9916 11580 11244 11608
rect 9916 11568 9922 11580
rect 11238 11568 11244 11580
rect 11296 11568 11302 11620
rect 9364 11512 9674 11540
rect 12268 11540 12296 11704
rect 16684 11676 16712 11707
rect 16942 11704 16948 11756
rect 17000 11744 17006 11756
rect 17898 11747 17956 11753
rect 17898 11744 17910 11747
rect 17000 11716 17910 11744
rect 17000 11704 17006 11716
rect 17898 11713 17910 11716
rect 17944 11713 17956 11747
rect 18322 11744 18328 11756
rect 18283 11716 18328 11744
rect 17898 11707 17956 11713
rect 18322 11704 18328 11716
rect 18380 11704 18386 11756
rect 19886 11744 19892 11756
rect 19847 11716 19892 11744
rect 19886 11704 19892 11716
rect 19944 11704 19950 11756
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11744 20131 11747
rect 20346 11744 20352 11756
rect 20119 11716 20352 11744
rect 20119 11713 20131 11716
rect 20073 11707 20131 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 22186 11744 22192 11756
rect 20496 11716 20541 11744
rect 22147 11716 22192 11744
rect 20496 11704 20502 11716
rect 22186 11704 22192 11716
rect 22244 11704 22250 11756
rect 18414 11676 18420 11688
rect 15488 11648 16712 11676
rect 18375 11648 18420 11676
rect 12434 11540 12440 11552
rect 12268 11512 12440 11540
rect 9364 11500 9370 11512
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15488 11549 15516 11648
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 20162 11676 20168 11688
rect 20123 11648 20168 11676
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 20254 11636 20260 11688
rect 20312 11676 20318 11688
rect 22465 11679 22523 11685
rect 20312 11648 20357 11676
rect 20312 11636 20318 11648
rect 22465 11645 22477 11679
rect 22511 11676 22523 11679
rect 29822 11676 29828 11688
rect 22511 11648 29828 11676
rect 22511 11645 22523 11648
rect 22465 11639 22523 11645
rect 29822 11636 29828 11648
rect 29880 11636 29886 11688
rect 16025 11611 16083 11617
rect 16025 11577 16037 11611
rect 16071 11608 16083 11611
rect 16850 11608 16856 11620
rect 16071 11580 16856 11608
rect 16071 11577 16083 11580
rect 16025 11571 16083 11577
rect 16850 11568 16856 11580
rect 16908 11568 16914 11620
rect 15473 11543 15531 11549
rect 15473 11540 15485 11543
rect 14884 11512 15485 11540
rect 14884 11500 14890 11512
rect 15473 11509 15485 11512
rect 15519 11509 15531 11543
rect 15473 11503 15531 11509
rect 16761 11543 16819 11549
rect 16761 11509 16773 11543
rect 16807 11540 16819 11543
rect 17310 11540 17316 11552
rect 16807 11512 17316 11540
rect 16807 11509 16819 11512
rect 16761 11503 16819 11509
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 19429 11543 19487 11549
rect 19429 11509 19441 11543
rect 19475 11540 19487 11543
rect 20622 11540 20628 11552
rect 19475 11512 20628 11540
rect 19475 11509 19487 11512
rect 19429 11503 19487 11509
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 1104 11450 30820 11472
rect 1104 11398 5915 11450
rect 5967 11398 5979 11450
rect 6031 11398 6043 11450
rect 6095 11398 6107 11450
rect 6159 11398 6171 11450
rect 6223 11398 15846 11450
rect 15898 11398 15910 11450
rect 15962 11398 15974 11450
rect 16026 11398 16038 11450
rect 16090 11398 16102 11450
rect 16154 11398 25776 11450
rect 25828 11398 25840 11450
rect 25892 11398 25904 11450
rect 25956 11398 25968 11450
rect 26020 11398 26032 11450
rect 26084 11398 30820 11450
rect 1104 11376 30820 11398
rect 8389 11339 8447 11345
rect 8389 11305 8401 11339
rect 8435 11336 8447 11339
rect 8478 11336 8484 11348
rect 8435 11308 8484 11336
rect 8435 11305 8447 11308
rect 8389 11299 8447 11305
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 17862 11336 17868 11348
rect 9508 11308 17724 11336
rect 17823 11308 17868 11336
rect 2777 11271 2835 11277
rect 2777 11237 2789 11271
rect 2823 11268 2835 11271
rect 2958 11268 2964 11280
rect 2823 11240 2964 11268
rect 2823 11237 2835 11240
rect 2777 11231 2835 11237
rect 2958 11228 2964 11240
rect 3016 11268 3022 11280
rect 3016 11240 4476 11268
rect 3016 11228 3022 11240
rect 4157 11203 4215 11209
rect 4157 11200 4169 11203
rect 2884 11172 4169 11200
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 2774 11132 2780 11144
rect 1443 11104 2780 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 2774 11092 2780 11104
rect 2832 11092 2838 11144
rect 1664 11067 1722 11073
rect 1664 11033 1676 11067
rect 1710 11064 1722 11067
rect 2130 11064 2136 11076
rect 1710 11036 2136 11064
rect 1710 11033 1722 11036
rect 1664 11027 1722 11033
rect 2130 11024 2136 11036
rect 2188 11024 2194 11076
rect 1762 10956 1768 11008
rect 1820 10996 1826 11008
rect 2038 10996 2044 11008
rect 1820 10968 2044 10996
rect 1820 10956 1826 10968
rect 2038 10956 2044 10968
rect 2096 10996 2102 11008
rect 2884 10996 2912 11172
rect 4157 11169 4169 11172
rect 4203 11169 4215 11203
rect 4157 11163 4215 11169
rect 3786 11132 3792 11144
rect 3747 11104 3792 11132
rect 3786 11092 3792 11104
rect 3844 11092 3850 11144
rect 3970 11132 3976 11144
rect 3931 11104 3976 11132
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4338 11132 4344 11144
rect 4120 11104 4165 11132
rect 4299 11104 4344 11132
rect 4120 11092 4126 11104
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 4448 11132 4476 11240
rect 8018 11228 8024 11280
rect 8076 11268 8082 11280
rect 9508 11268 9536 11308
rect 12986 11268 12992 11280
rect 8076 11240 9536 11268
rect 12820 11240 12992 11268
rect 8076 11228 8082 11240
rect 5442 11200 5448 11212
rect 5403 11172 5448 11200
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 7006 11200 7012 11212
rect 6967 11172 7012 11200
rect 7006 11160 7012 11172
rect 7064 11160 7070 11212
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11200 9183 11203
rect 9582 11200 9588 11212
rect 9171 11172 9588 11200
rect 9171 11169 9183 11172
rect 9125 11163 9183 11169
rect 9582 11160 9588 11172
rect 9640 11160 9646 11212
rect 11790 11160 11796 11212
rect 11848 11200 11854 11212
rect 12820 11200 12848 11240
rect 12986 11228 12992 11240
rect 13044 11228 13050 11280
rect 15473 11271 15531 11277
rect 15473 11237 15485 11271
rect 15519 11268 15531 11271
rect 16942 11268 16948 11280
rect 15519 11240 16948 11268
rect 15519 11237 15531 11240
rect 15473 11231 15531 11237
rect 11848 11172 12848 11200
rect 11848 11160 11854 11172
rect 7282 11141 7288 11144
rect 5537 11135 5595 11141
rect 5537 11132 5549 11135
rect 4448 11104 5549 11132
rect 5537 11101 5549 11104
rect 5583 11101 5595 11135
rect 5537 11095 5595 11101
rect 5665 11135 5723 11141
rect 5665 11101 5677 11135
rect 5711 11132 5723 11135
rect 7276 11132 7288 11141
rect 5711 11104 6316 11132
rect 7243 11104 7288 11132
rect 5711 11101 5723 11104
rect 5665 11095 5723 11101
rect 6288 11076 6316 11104
rect 7276 11095 7288 11104
rect 7282 11092 7288 11095
rect 7340 11092 7346 11144
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 9306 11132 9312 11144
rect 8904 11104 9312 11132
rect 8904 11092 8910 11104
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11132 9459 11135
rect 9766 11132 9772 11144
rect 9447 11104 9772 11132
rect 9447 11101 9459 11104
rect 9401 11095 9459 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11132 10195 11135
rect 10226 11132 10232 11144
rect 10183 11104 10232 11132
rect 10183 11101 10195 11104
rect 10137 11095 10195 11101
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 12158 11132 12164 11144
rect 10336 11104 12164 11132
rect 5166 11024 5172 11076
rect 5224 11064 5230 11076
rect 5261 11067 5319 11073
rect 5261 11064 5273 11067
rect 5224 11036 5273 11064
rect 5224 11024 5230 11036
rect 5261 11033 5273 11036
rect 5307 11033 5319 11067
rect 5261 11027 5319 11033
rect 5350 11024 5356 11076
rect 5408 11064 5414 11076
rect 5445 11067 5503 11073
rect 5445 11064 5457 11067
rect 5408 11036 5457 11064
rect 5408 11024 5414 11036
rect 5445 11033 5457 11036
rect 5491 11033 5503 11067
rect 5445 11027 5503 11033
rect 6270 11024 6276 11076
rect 6328 11064 6334 11076
rect 7190 11064 7196 11076
rect 6328 11036 7196 11064
rect 6328 11024 6334 11036
rect 7190 11024 7196 11036
rect 7248 11064 7254 11076
rect 10336 11064 10364 11104
rect 12158 11092 12164 11104
rect 12216 11092 12222 11144
rect 12820 11141 12848 11172
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11200 13231 11203
rect 13722 11200 13728 11212
rect 13219 11172 13728 11200
rect 13219 11169 13231 11172
rect 13173 11163 13231 11169
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 14090 11200 14096 11212
rect 14051 11172 14096 11200
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 12894 11092 12900 11144
rect 12952 11132 12958 11144
rect 12989 11135 13047 11141
rect 12989 11132 13001 11135
rect 12952 11104 13001 11132
rect 12952 11092 12958 11104
rect 12989 11101 13001 11104
rect 13035 11101 13047 11135
rect 12989 11095 13047 11101
rect 13081 11135 13139 11141
rect 13081 11101 13093 11135
rect 13127 11132 13139 11135
rect 13262 11132 13268 11144
rect 13127 11104 13268 11132
rect 13127 11101 13139 11104
rect 13081 11095 13139 11101
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 15488 11132 15516 11231
rect 16942 11228 16948 11240
rect 17000 11228 17006 11280
rect 17696 11268 17724 11308
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 18414 11336 18420 11348
rect 18375 11308 18420 11336
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 19889 11339 19947 11345
rect 19889 11305 19901 11339
rect 19935 11336 19947 11339
rect 20070 11336 20076 11348
rect 19935 11308 20076 11336
rect 19935 11305 19947 11308
rect 19889 11299 19947 11305
rect 20070 11296 20076 11308
rect 20128 11296 20134 11348
rect 20346 11296 20352 11348
rect 20404 11336 20410 11348
rect 21177 11339 21235 11345
rect 21177 11336 21189 11339
rect 20404 11308 21189 11336
rect 20404 11296 20410 11308
rect 21177 11305 21189 11308
rect 21223 11305 21235 11339
rect 21177 11299 21235 11305
rect 17696 11240 18460 11268
rect 15654 11160 15660 11212
rect 15712 11200 15718 11212
rect 16298 11200 16304 11212
rect 15712 11172 16160 11200
rect 16259 11172 16304 11200
rect 15712 11160 15718 11172
rect 13403 11104 15516 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 15746 11092 15752 11144
rect 15804 11132 15810 11144
rect 16132 11141 16160 11172
rect 16298 11160 16304 11172
rect 16356 11200 16362 11212
rect 17034 11200 17040 11212
rect 16356 11172 17040 11200
rect 16356 11160 16362 11172
rect 17034 11160 17040 11172
rect 17092 11160 17098 11212
rect 17497 11203 17555 11209
rect 17497 11169 17509 11203
rect 17543 11200 17555 11203
rect 18322 11200 18328 11212
rect 17543 11172 18328 11200
rect 17543 11169 17555 11172
rect 17497 11163 17555 11169
rect 18322 11160 18328 11172
rect 18380 11160 18386 11212
rect 18432 11200 18460 11240
rect 18432 11172 18644 11200
rect 15933 11135 15991 11141
rect 15933 11132 15945 11135
rect 15804 11104 15945 11132
rect 15804 11092 15810 11104
rect 15933 11101 15945 11104
rect 15979 11101 15991 11135
rect 15933 11095 15991 11101
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 16209 11135 16267 11141
rect 16209 11101 16221 11135
rect 16255 11101 16267 11135
rect 16482 11132 16488 11144
rect 16443 11104 16488 11132
rect 16209 11095 16267 11101
rect 7248 11036 10364 11064
rect 10404 11067 10462 11073
rect 7248 11024 7254 11036
rect 10404 11033 10416 11067
rect 10450 11064 10462 11067
rect 10686 11064 10692 11076
rect 10450 11036 10692 11064
rect 10450 11033 10462 11036
rect 10404 11027 10462 11033
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 13541 11067 13599 11073
rect 13541 11033 13553 11067
rect 13587 11064 13599 11067
rect 14338 11067 14396 11073
rect 14338 11064 14350 11067
rect 13587 11036 14350 11064
rect 13587 11033 13599 11036
rect 13541 11027 13599 11033
rect 14338 11033 14350 11036
rect 14384 11033 14396 11067
rect 14338 11027 14396 11033
rect 14550 11024 14556 11076
rect 14608 11064 14614 11076
rect 16224 11064 16252 11095
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11132 16727 11135
rect 16758 11132 16764 11144
rect 16715 11104 16764 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 17126 11132 17132 11144
rect 17087 11104 17132 11132
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 17310 11132 17316 11144
rect 17271 11104 17316 11132
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 17405 11135 17463 11141
rect 17405 11101 17417 11135
rect 17451 11101 17463 11135
rect 17405 11095 17463 11101
rect 17681 11135 17739 11141
rect 17681 11101 17693 11135
rect 17727 11132 17739 11135
rect 18046 11132 18052 11144
rect 17727 11104 18052 11132
rect 17727 11101 17739 11104
rect 17681 11095 17739 11101
rect 16942 11064 16948 11076
rect 14608 11036 16948 11064
rect 14608 11024 14614 11036
rect 16942 11024 16948 11036
rect 17000 11064 17006 11076
rect 17420 11064 17448 11095
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18506 11132 18512 11144
rect 18467 11104 18512 11132
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 17000 11036 17448 11064
rect 18616 11064 18644 11172
rect 20162 11160 20168 11212
rect 20220 11200 20226 11212
rect 20349 11203 20407 11209
rect 20349 11200 20361 11203
rect 20220 11172 20361 11200
rect 20220 11160 20226 11172
rect 20349 11169 20361 11172
rect 20395 11169 20407 11203
rect 20349 11163 20407 11169
rect 19518 11092 19524 11144
rect 19576 11132 19582 11144
rect 20073 11135 20131 11141
rect 20073 11132 20085 11135
rect 19576 11104 20085 11132
rect 19576 11092 19582 11104
rect 20073 11101 20085 11104
rect 20119 11101 20131 11135
rect 20254 11132 20260 11144
rect 20167 11104 20260 11132
rect 20073 11095 20131 11101
rect 20254 11092 20260 11104
rect 20312 11092 20318 11144
rect 20441 11135 20499 11141
rect 20441 11101 20453 11135
rect 20487 11101 20499 11135
rect 20622 11132 20628 11144
rect 20583 11104 20628 11132
rect 20441 11095 20499 11101
rect 20272 11064 20300 11092
rect 18616 11036 20300 11064
rect 20456 11064 20484 11095
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 21269 11135 21327 11141
rect 21269 11101 21281 11135
rect 21315 11132 21327 11135
rect 21358 11132 21364 11144
rect 21315 11104 21364 11132
rect 21315 11101 21327 11104
rect 21269 11095 21327 11101
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 29822 11132 29828 11144
rect 29783 11104 29828 11132
rect 29822 11092 29828 11104
rect 29880 11092 29886 11144
rect 20714 11064 20720 11076
rect 20456 11036 20720 11064
rect 17000 11024 17006 11036
rect 20714 11024 20720 11036
rect 20772 11024 20778 11076
rect 4522 10996 4528 11008
rect 2096 10968 2912 10996
rect 4483 10968 4528 10996
rect 2096 10956 2102 10968
rect 4522 10956 4528 10968
rect 4580 10956 4586 11008
rect 11514 10996 11520 11008
rect 11475 10968 11520 10996
rect 11514 10956 11520 10968
rect 11572 10956 11578 11008
rect 11606 10956 11612 11008
rect 11664 10996 11670 11008
rect 13814 10996 13820 11008
rect 11664 10968 13820 10996
rect 11664 10956 11670 10968
rect 13814 10956 13820 10968
rect 13872 10996 13878 11008
rect 15010 10996 15016 11008
rect 13872 10968 15016 10996
rect 13872 10956 13878 10968
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 30006 10996 30012 11008
rect 29967 10968 30012 10996
rect 30006 10956 30012 10968
rect 30064 10956 30070 11008
rect 1104 10906 30820 10928
rect 1104 10854 10880 10906
rect 10932 10854 10944 10906
rect 10996 10854 11008 10906
rect 11060 10854 11072 10906
rect 11124 10854 11136 10906
rect 11188 10854 20811 10906
rect 20863 10854 20875 10906
rect 20927 10854 20939 10906
rect 20991 10854 21003 10906
rect 21055 10854 21067 10906
rect 21119 10854 30820 10906
rect 1104 10832 30820 10854
rect 2958 10792 2964 10804
rect 1964 10764 2964 10792
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10625 1455 10659
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1397 10619 1455 10625
rect 1412 10588 1440 10619
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 1964 10665 1992 10764
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 5460 10764 5764 10792
rect 2130 10724 2136 10736
rect 2091 10696 2136 10724
rect 2130 10684 2136 10696
rect 2188 10684 2194 10736
rect 3044 10727 3102 10733
rect 3044 10693 3056 10727
rect 3090 10724 3102 10727
rect 4522 10724 4528 10736
rect 3090 10696 4528 10724
rect 3090 10693 3102 10696
rect 3044 10687 3102 10693
rect 4522 10684 4528 10696
rect 4580 10684 4586 10736
rect 5166 10684 5172 10736
rect 5224 10724 5230 10736
rect 5353 10727 5411 10733
rect 5353 10724 5365 10727
rect 5224 10696 5365 10724
rect 5224 10684 5230 10696
rect 5353 10693 5365 10696
rect 5399 10724 5411 10727
rect 5460 10724 5488 10764
rect 5399 10696 5488 10724
rect 5537 10727 5595 10733
rect 5399 10693 5411 10696
rect 5353 10687 5411 10693
rect 5537 10693 5549 10727
rect 5583 10693 5595 10727
rect 5537 10687 5595 10693
rect 5629 10727 5687 10733
rect 5629 10693 5641 10727
rect 5675 10693 5687 10727
rect 5736 10724 5764 10764
rect 6546 10752 6552 10804
rect 6604 10792 6610 10804
rect 6914 10792 6920 10804
rect 6604 10764 6920 10792
rect 6604 10752 6610 10764
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 10686 10792 10692 10804
rect 10647 10764 10692 10792
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 10778 10752 10784 10804
rect 10836 10792 10842 10804
rect 12710 10792 12716 10804
rect 10836 10764 12716 10792
rect 10836 10752 10842 10764
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 13725 10795 13783 10801
rect 13725 10761 13737 10795
rect 13771 10792 13783 10795
rect 14366 10792 14372 10804
rect 13771 10764 14372 10792
rect 13771 10761 13783 10764
rect 13725 10755 13783 10761
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 16574 10752 16580 10804
rect 16632 10752 16638 10804
rect 18046 10792 18052 10804
rect 18007 10764 18052 10792
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 20530 10792 20536 10804
rect 20491 10764 20536 10792
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 21085 10795 21143 10801
rect 21085 10792 21097 10795
rect 20772 10764 21097 10792
rect 20772 10752 20778 10764
rect 21085 10761 21097 10764
rect 21131 10761 21143 10795
rect 21085 10755 21143 10761
rect 6825 10727 6883 10733
rect 6825 10724 6837 10727
rect 5736 10696 6837 10724
rect 5629 10687 5687 10693
rect 6825 10693 6837 10696
rect 6871 10724 6883 10727
rect 11606 10724 11612 10736
rect 6871 10696 11612 10724
rect 6871 10693 6883 10696
rect 6825 10687 6883 10693
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 1949 10659 2007 10665
rect 1719 10628 1900 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 1486 10588 1492 10600
rect 1412 10560 1492 10588
rect 1486 10548 1492 10560
rect 1544 10548 1550 10600
rect 1762 10588 1768 10600
rect 1723 10560 1768 10588
rect 1762 10548 1768 10560
rect 1820 10548 1826 10600
rect 1872 10588 1900 10628
rect 1949 10625 1961 10659
rect 1995 10625 2007 10659
rect 2774 10656 2780 10668
rect 2687 10628 2780 10656
rect 1949 10619 2007 10625
rect 2774 10616 2780 10628
rect 2832 10656 2838 10668
rect 3878 10656 3884 10668
rect 2832 10628 3884 10656
rect 2832 10616 2838 10628
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 5552 10656 5580 10687
rect 5500 10628 5580 10656
rect 5500 10616 5506 10628
rect 2682 10588 2688 10600
rect 1872 10560 2688 10588
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 5353 10591 5411 10597
rect 5353 10588 5365 10591
rect 4948 10560 5365 10588
rect 4948 10548 4954 10560
rect 5353 10557 5365 10560
rect 5399 10557 5411 10591
rect 5353 10551 5411 10557
rect 4157 10523 4215 10529
rect 4157 10489 4169 10523
rect 4203 10520 4215 10523
rect 4338 10520 4344 10532
rect 4203 10492 4344 10520
rect 4203 10489 4215 10492
rect 4157 10483 4215 10489
rect 4338 10480 4344 10492
rect 4396 10520 4402 10532
rect 5649 10520 5677 10687
rect 11606 10684 11612 10696
rect 11664 10684 11670 10736
rect 12342 10684 12348 10736
rect 12400 10724 12406 10736
rect 15841 10727 15899 10733
rect 15841 10724 15853 10727
rect 12400 10696 15853 10724
rect 12400 10684 12406 10696
rect 15841 10693 15853 10696
rect 15887 10693 15899 10727
rect 16592 10724 16620 10752
rect 15841 10687 15899 10693
rect 16500 10696 16620 10724
rect 17405 10727 17463 10733
rect 5757 10659 5815 10665
rect 5757 10625 5769 10659
rect 5803 10656 5815 10659
rect 6270 10656 6276 10668
rect 5803 10628 6276 10656
rect 5803 10625 5815 10628
rect 5757 10619 5815 10625
rect 6270 10616 6276 10628
rect 6328 10656 6334 10668
rect 6421 10659 6479 10665
rect 6421 10656 6433 10659
rect 6328 10628 6433 10656
rect 6328 10616 6334 10628
rect 6421 10625 6433 10628
rect 6467 10625 6479 10659
rect 6546 10656 6552 10668
rect 6507 10628 6552 10656
rect 6421 10619 6479 10625
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 6696 10628 6741 10656
rect 6696 10616 6702 10628
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 8205 10659 8263 10665
rect 8205 10656 8217 10659
rect 8168 10628 8217 10656
rect 8168 10616 8174 10628
rect 8205 10625 8217 10628
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10656 8999 10659
rect 9858 10656 9864 10668
rect 8987 10628 9864 10656
rect 8987 10625 8999 10628
rect 8941 10619 8999 10625
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10134 10656 10140 10668
rect 10008 10628 10053 10656
rect 10095 10628 10140 10656
rect 10008 10616 10014 10628
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10656 10563 10659
rect 11422 10656 11428 10668
rect 10551 10628 11428 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 11422 10616 11428 10628
rect 11480 10616 11486 10668
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10625 11575 10659
rect 11698 10656 11704 10668
rect 11659 10628 11704 10656
rect 11517 10619 11575 10625
rect 10229 10591 10287 10597
rect 10229 10557 10241 10591
rect 10275 10557 10287 10591
rect 10229 10551 10287 10557
rect 10321 10591 10379 10597
rect 10321 10557 10333 10591
rect 10367 10588 10379 10591
rect 10367 10560 10640 10588
rect 10367 10557 10379 10560
rect 10321 10551 10379 10557
rect 4396 10492 5677 10520
rect 4396 10480 4402 10492
rect 5718 10480 5724 10532
rect 5776 10520 5782 10532
rect 6825 10523 6883 10529
rect 6825 10520 6837 10523
rect 5776 10492 6837 10520
rect 5776 10480 5782 10492
rect 6825 10489 6837 10492
rect 6871 10489 6883 10523
rect 6825 10483 6883 10489
rect 8294 10480 8300 10532
rect 8352 10520 8358 10532
rect 8757 10523 8815 10529
rect 8757 10520 8769 10523
rect 8352 10492 8769 10520
rect 8352 10480 8358 10492
rect 8757 10489 8769 10492
rect 8803 10489 8815 10523
rect 10244 10520 10272 10551
rect 10502 10520 10508 10532
rect 10244 10492 10508 10520
rect 8757 10483 8815 10489
rect 10502 10480 10508 10492
rect 10560 10480 10566 10532
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 6546 10452 6552 10464
rect 3568 10424 6552 10452
rect 3568 10412 3574 10424
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 7558 10412 7564 10464
rect 7616 10452 7622 10464
rect 8113 10455 8171 10461
rect 8113 10452 8125 10455
rect 7616 10424 8125 10452
rect 7616 10412 7622 10424
rect 8113 10421 8125 10424
rect 8159 10452 8171 10455
rect 10612 10452 10640 10560
rect 10962 10480 10968 10532
rect 11020 10520 11026 10532
rect 11532 10520 11560 10619
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 11793 10659 11851 10665
rect 11793 10625 11805 10659
rect 11839 10656 11851 10659
rect 11974 10656 11980 10668
rect 11839 10628 11980 10656
rect 11839 10625 11851 10628
rect 11793 10619 11851 10625
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 12069 10659 12127 10665
rect 12069 10625 12081 10659
rect 12115 10656 12127 10659
rect 12618 10656 12624 10668
rect 12115 10628 12624 10656
rect 12115 10625 12127 10628
rect 12069 10619 12127 10625
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 12986 10656 12992 10668
rect 12947 10628 12992 10656
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10656 13231 10659
rect 13446 10656 13452 10668
rect 13219 10628 13452 10656
rect 13219 10625 13231 10628
rect 13173 10619 13231 10625
rect 13446 10616 13452 10628
rect 13504 10616 13510 10668
rect 13541 10659 13599 10665
rect 13541 10625 13553 10659
rect 13587 10656 13599 10659
rect 14826 10656 14832 10668
rect 13587 10628 14832 10656
rect 13587 10625 13599 10628
rect 13541 10619 13599 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 15010 10656 15016 10668
rect 14971 10628 15016 10656
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10656 15255 10659
rect 15654 10656 15660 10668
rect 15243 10628 15660 10656
rect 15243 10625 15255 10628
rect 15197 10619 15255 10625
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 16061 10659 16119 10665
rect 16061 10625 16073 10659
rect 16107 10656 16119 10659
rect 16500 10656 16528 10696
rect 17405 10693 17417 10727
rect 17451 10724 17463 10727
rect 18966 10724 18972 10736
rect 17451 10696 18972 10724
rect 17451 10693 17463 10696
rect 17405 10687 17463 10693
rect 18966 10684 18972 10696
rect 19024 10684 19030 10736
rect 16107 10628 16528 10656
rect 16107 10625 16119 10628
rect 16061 10619 16119 10625
rect 11882 10588 11888 10600
rect 11843 10560 11888 10588
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 11992 10588 12020 10616
rect 13262 10588 13268 10600
rect 11992 10560 13268 10588
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10588 13415 10591
rect 13722 10588 13728 10600
rect 13403 10560 13728 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 15746 10588 15752 10600
rect 15707 10560 15752 10588
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 11020 10492 11560 10520
rect 11020 10480 11026 10492
rect 11900 10452 11928 10548
rect 12250 10452 12256 10464
rect 8159 10424 11928 10452
rect 12211 10424 12256 10452
rect 8159 10421 8171 10424
rect 8113 10415 8171 10421
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 15948 10452 15976 10619
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 16632 10628 16681 10656
rect 16632 10616 16638 10628
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16850 10656 16856 10668
rect 16811 10628 16856 10656
rect 16669 10619 16727 10625
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 16942 10616 16948 10668
rect 17000 10656 17006 10668
rect 17218 10656 17224 10668
rect 17000 10628 17045 10656
rect 17179 10628 17224 10656
rect 17000 10616 17006 10628
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 17954 10656 17960 10668
rect 17915 10628 17960 10656
rect 17954 10616 17960 10628
rect 18012 10616 18018 10668
rect 18874 10656 18880 10668
rect 18835 10628 18880 10656
rect 18874 10616 18880 10628
rect 18932 10616 18938 10668
rect 19797 10659 19855 10665
rect 19797 10625 19809 10659
rect 19843 10625 19855 10659
rect 19978 10656 19984 10668
rect 19939 10628 19984 10656
rect 19797 10619 19855 10625
rect 17034 10588 17040 10600
rect 16995 10560 17040 10588
rect 17034 10548 17040 10560
rect 17092 10548 17098 10600
rect 19337 10591 19395 10597
rect 19337 10557 19349 10591
rect 19383 10588 19395 10591
rect 19812 10588 19840 10619
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 20346 10656 20352 10668
rect 20307 10628 20352 10656
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10656 21235 10659
rect 21450 10656 21456 10668
rect 21223 10628 21456 10656
rect 21223 10625 21235 10628
rect 21177 10619 21235 10625
rect 21450 10616 21456 10628
rect 21508 10616 21514 10668
rect 20070 10588 20076 10600
rect 19383 10560 19840 10588
rect 19983 10560 20076 10588
rect 19383 10557 19395 10560
rect 19337 10551 19395 10557
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10588 20223 10591
rect 20254 10588 20260 10600
rect 20211 10560 20260 10588
rect 20211 10557 20223 10560
rect 20165 10551 20223 10557
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 17052 10520 17080 10548
rect 20088 10520 20116 10548
rect 17052 10492 20116 10520
rect 18598 10452 18604 10464
rect 15948 10424 18604 10452
rect 18598 10412 18604 10424
rect 18656 10412 18662 10464
rect 19058 10452 19064 10464
rect 19019 10424 19064 10452
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 1104 10362 30820 10384
rect 1104 10310 5915 10362
rect 5967 10310 5979 10362
rect 6031 10310 6043 10362
rect 6095 10310 6107 10362
rect 6159 10310 6171 10362
rect 6223 10310 15846 10362
rect 15898 10310 15910 10362
rect 15962 10310 15974 10362
rect 16026 10310 16038 10362
rect 16090 10310 16102 10362
rect 16154 10310 25776 10362
rect 25828 10310 25840 10362
rect 25892 10310 25904 10362
rect 25956 10310 25968 10362
rect 26020 10310 26032 10362
rect 26084 10310 30820 10362
rect 1104 10288 30820 10310
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 9217 10251 9275 10257
rect 9217 10248 9229 10251
rect 8628 10220 9229 10248
rect 8628 10208 8634 10220
rect 9217 10217 9229 10220
rect 9263 10217 9275 10251
rect 9217 10211 9275 10217
rect 10226 10208 10232 10260
rect 10284 10248 10290 10260
rect 10321 10251 10379 10257
rect 10321 10248 10333 10251
rect 10284 10220 10333 10248
rect 10284 10208 10290 10220
rect 10321 10217 10333 10220
rect 10367 10217 10379 10251
rect 10321 10211 10379 10217
rect 11514 10208 11520 10260
rect 11572 10248 11578 10260
rect 15746 10248 15752 10260
rect 11572 10220 15752 10248
rect 11572 10208 11578 10220
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 16209 10251 16267 10257
rect 16209 10217 16221 10251
rect 16255 10248 16267 10251
rect 17678 10248 17684 10260
rect 16255 10220 17684 10248
rect 16255 10217 16267 10220
rect 16209 10211 16267 10217
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 19978 10208 19984 10260
rect 20036 10248 20042 10260
rect 20441 10251 20499 10257
rect 20441 10248 20453 10251
rect 20036 10220 20453 10248
rect 20036 10208 20042 10220
rect 20441 10217 20453 10220
rect 20487 10217 20499 10251
rect 28718 10248 28724 10260
rect 20441 10211 20499 10217
rect 20548 10220 28724 10248
rect 1486 10140 1492 10192
rect 1544 10180 1550 10192
rect 2590 10180 2596 10192
rect 1544 10152 2596 10180
rect 1544 10140 1550 10152
rect 1688 10053 1716 10152
rect 2590 10140 2596 10152
rect 2648 10140 2654 10192
rect 2869 10183 2927 10189
rect 2869 10180 2881 10183
rect 2746 10152 2881 10180
rect 2746 10112 2774 10152
rect 2869 10149 2881 10152
rect 2915 10149 2927 10183
rect 2869 10143 2927 10149
rect 6270 10140 6276 10192
rect 6328 10180 6334 10192
rect 8754 10180 8760 10192
rect 6328 10152 8760 10180
rect 6328 10140 6334 10152
rect 8754 10140 8760 10152
rect 8812 10140 8818 10192
rect 9950 10140 9956 10192
rect 10008 10180 10014 10192
rect 10962 10180 10968 10192
rect 10008 10152 10968 10180
rect 10008 10140 10014 10152
rect 10962 10140 10968 10152
rect 11020 10140 11026 10192
rect 12618 10180 12624 10192
rect 12531 10152 12624 10180
rect 12618 10140 12624 10152
rect 12676 10180 12682 10192
rect 20548 10180 20576 10220
rect 28718 10208 28724 10220
rect 28776 10208 28782 10260
rect 12676 10152 17540 10180
rect 12676 10140 12682 10152
rect 6638 10112 6644 10124
rect 1872 10084 2774 10112
rect 5920 10084 6644 10112
rect 1872 10053 1900 10084
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 1943 10047 2001 10053
rect 1943 10013 1955 10047
rect 1989 10013 2001 10047
rect 1943 10007 2001 10013
rect 1958 9920 1986 10007
rect 2038 10004 2044 10056
rect 2096 10053 2102 10056
rect 2096 10047 2145 10053
rect 2096 10013 2099 10047
rect 2133 10013 2145 10047
rect 2096 10007 2145 10013
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 3050 10044 3056 10056
rect 2271 10016 2774 10044
rect 3011 10016 3056 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 2096 10004 2102 10007
rect 2746 9976 2774 10016
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 3881 10047 3939 10053
rect 3881 10013 3893 10047
rect 3927 10044 3939 10047
rect 5074 10044 5080 10056
rect 3927 10016 5080 10044
rect 3927 10013 3939 10016
rect 3881 10007 3939 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5920 10053 5948 10084
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 13722 10072 13728 10124
rect 13780 10112 13786 10124
rect 14461 10115 14519 10121
rect 14461 10112 14473 10115
rect 13780 10084 14473 10112
rect 13780 10072 13786 10084
rect 14461 10081 14473 10084
rect 14507 10081 14519 10115
rect 16390 10112 16396 10124
rect 14461 10075 14519 10081
rect 14660 10084 16396 10112
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 6089 10047 6147 10053
rect 6089 10044 6101 10047
rect 6052 10016 6101 10044
rect 6052 10004 6058 10016
rect 6089 10013 6101 10016
rect 6135 10013 6147 10047
rect 6089 10007 6147 10013
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 3510 9976 3516 9988
rect 2746 9948 3516 9976
rect 3510 9936 3516 9948
rect 3568 9936 3574 9988
rect 4148 9979 4206 9985
rect 4148 9945 4160 9979
rect 4194 9976 4206 9979
rect 4982 9976 4988 9988
rect 4194 9948 4988 9976
rect 4194 9945 4206 9948
rect 4148 9939 4206 9945
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 6196 9976 6224 10007
rect 6270 10004 6276 10056
rect 6328 10044 6334 10056
rect 6457 10047 6515 10053
rect 6328 10016 6373 10044
rect 6328 10004 6334 10016
rect 6457 10013 6469 10047
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 7190 10044 7196 10056
rect 7147 10016 7196 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 6472 9976 6500 10007
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 10778 10044 10784 10056
rect 7883 10016 10784 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10044 11299 10047
rect 12434 10044 12440 10056
rect 11287 10016 12440 10044
rect 11287 10013 11299 10016
rect 11241 10007 11299 10013
rect 12434 10004 12440 10016
rect 12492 10004 12498 10056
rect 12986 10004 12992 10056
rect 13044 10044 13050 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13044 10016 14105 10044
rect 13044 10004 13050 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14274 10044 14280 10056
rect 14235 10016 14280 10044
rect 14093 10007 14151 10013
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 14369 10047 14427 10053
rect 14369 10013 14381 10047
rect 14415 10044 14427 10047
rect 14550 10044 14556 10056
rect 14415 10016 14556 10044
rect 14415 10013 14427 10016
rect 14369 10007 14427 10013
rect 14550 10004 14556 10016
rect 14608 10004 14614 10056
rect 14660 10053 14688 10084
rect 16390 10072 16396 10084
rect 16448 10072 16454 10124
rect 16574 10112 16580 10124
rect 16535 10084 16580 10112
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 17126 10072 17132 10124
rect 17184 10112 17190 10124
rect 17405 10115 17463 10121
rect 17405 10112 17417 10115
rect 17184 10084 17417 10112
rect 17184 10072 17190 10084
rect 17405 10081 17417 10084
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 14645 10047 14703 10053
rect 14645 10013 14657 10047
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 15746 10004 15752 10056
rect 15804 10044 15810 10056
rect 16485 10047 16543 10053
rect 16485 10044 16497 10047
rect 15804 10016 16497 10044
rect 15804 10004 15810 10016
rect 16485 10013 16497 10016
rect 16531 10013 16543 10047
rect 16666 10044 16672 10056
rect 16724 10053 16730 10056
rect 16724 10047 16763 10053
rect 16615 10016 16672 10044
rect 16485 10007 16543 10013
rect 16666 10004 16672 10016
rect 16751 10044 16763 10047
rect 17277 10047 17335 10053
rect 17277 10044 17289 10047
rect 16751 10016 17289 10044
rect 16751 10013 16763 10016
rect 16724 10007 16763 10013
rect 17277 10013 17289 10016
rect 17323 10013 17335 10047
rect 17277 10007 17335 10013
rect 16724 10004 16730 10007
rect 5408 9948 6224 9976
rect 6288 9948 6500 9976
rect 5408 9936 5414 9948
rect 6288 9920 6316 9948
rect 6546 9936 6552 9988
rect 6604 9976 6610 9988
rect 6917 9979 6975 9985
rect 6917 9976 6929 9979
rect 6604 9948 6929 9976
rect 6604 9936 6610 9948
rect 6917 9945 6929 9948
rect 6963 9945 6975 9979
rect 6917 9939 6975 9945
rect 7006 9936 7012 9988
rect 7064 9976 7070 9988
rect 7653 9979 7711 9985
rect 7653 9976 7665 9979
rect 7064 9948 7665 9976
rect 7064 9936 7070 9948
rect 7653 9945 7665 9948
rect 7699 9945 7711 9979
rect 7653 9939 7711 9945
rect 9401 9979 9459 9985
rect 9401 9945 9413 9979
rect 9447 9945 9459 9979
rect 9401 9939 9459 9945
rect 1946 9868 1952 9920
rect 2004 9868 2010 9920
rect 2406 9908 2412 9920
rect 2367 9880 2412 9908
rect 2406 9868 2412 9880
rect 2464 9868 2470 9920
rect 5258 9908 5264 9920
rect 5219 9880 5264 9908
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 5718 9908 5724 9920
rect 5679 9880 5724 9908
rect 5718 9868 5724 9880
rect 5776 9868 5782 9920
rect 6270 9868 6276 9920
rect 6328 9868 6334 9920
rect 9416 9908 9444 9939
rect 9490 9936 9496 9988
rect 9548 9976 9554 9988
rect 9585 9979 9643 9985
rect 9585 9976 9597 9979
rect 9548 9948 9597 9976
rect 9548 9936 9554 9948
rect 9585 9945 9597 9948
rect 9631 9976 9643 9979
rect 10045 9979 10103 9985
rect 10045 9976 10057 9979
rect 9631 9948 10057 9976
rect 9631 9945 9643 9948
rect 9585 9939 9643 9945
rect 10045 9945 10057 9948
rect 10091 9945 10103 9979
rect 10226 9976 10232 9988
rect 10187 9948 10232 9976
rect 10045 9939 10103 9945
rect 10226 9936 10232 9948
rect 10284 9936 10290 9988
rect 11508 9979 11566 9985
rect 11508 9945 11520 9979
rect 11554 9976 11566 9979
rect 12250 9976 12256 9988
rect 11554 9948 12256 9976
rect 11554 9945 11566 9948
rect 11508 9939 11566 9945
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 13173 9979 13231 9985
rect 13173 9976 13185 9979
rect 12406 9948 13185 9976
rect 9950 9908 9956 9920
rect 9416 9880 9956 9908
rect 9950 9868 9956 9880
rect 10008 9868 10014 9920
rect 10686 9868 10692 9920
rect 10744 9908 10750 9920
rect 12406 9908 12434 9948
rect 13173 9945 13185 9948
rect 13219 9945 13231 9979
rect 13173 9939 13231 9945
rect 13357 9979 13415 9985
rect 13357 9945 13369 9979
rect 13403 9976 13415 9979
rect 14182 9976 14188 9988
rect 13403 9948 14188 9976
rect 13403 9945 13415 9948
rect 13357 9939 13415 9945
rect 14182 9936 14188 9948
rect 14240 9976 14246 9988
rect 15381 9979 15439 9985
rect 15381 9976 15393 9979
rect 14240 9948 15393 9976
rect 14240 9936 14246 9948
rect 15381 9945 15393 9948
rect 15427 9945 15439 9979
rect 15562 9976 15568 9988
rect 15523 9948 15568 9976
rect 15381 9939 15439 9945
rect 15562 9936 15568 9948
rect 15620 9936 15626 9988
rect 15654 9936 15660 9988
rect 15712 9976 15718 9988
rect 16209 9979 16267 9985
rect 16209 9976 16221 9979
rect 15712 9948 16221 9976
rect 15712 9936 15718 9948
rect 16209 9945 16221 9948
rect 16255 9976 16267 9979
rect 16301 9979 16359 9985
rect 16301 9976 16313 9979
rect 16255 9948 16313 9976
rect 16255 9945 16267 9948
rect 16209 9939 16267 9945
rect 16301 9945 16313 9948
rect 16347 9945 16359 9979
rect 16301 9939 16359 9945
rect 16577 9979 16635 9985
rect 16577 9945 16589 9979
rect 16623 9945 16635 9979
rect 17402 9976 17408 9988
rect 17363 9948 17408 9976
rect 16577 9939 16635 9945
rect 10744 9880 12434 9908
rect 10744 9868 10750 9880
rect 12618 9868 12624 9920
rect 12676 9908 12682 9920
rect 14642 9908 14648 9920
rect 12676 9880 14648 9908
rect 12676 9868 12682 9880
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 14826 9908 14832 9920
rect 14787 9880 14832 9908
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 16592 9908 16620 9939
rect 17402 9936 17408 9948
rect 17460 9936 17466 9988
rect 17512 9985 17540 10152
rect 18340 10152 20576 10180
rect 17678 10044 17684 10056
rect 17639 10016 17684 10044
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 18138 10004 18144 10056
rect 18196 10044 18202 10056
rect 18340 10053 18368 10152
rect 18509 10115 18567 10121
rect 18509 10081 18521 10115
rect 18555 10112 18567 10115
rect 18690 10112 18696 10124
rect 18555 10084 18696 10112
rect 18555 10081 18567 10084
rect 18509 10075 18567 10081
rect 18690 10072 18696 10084
rect 18748 10072 18754 10124
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 18196 10016 18337 10044
rect 18196 10004 18202 10016
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 18601 10047 18659 10053
rect 18601 10013 18613 10047
rect 18647 10044 18659 10047
rect 18874 10044 18880 10056
rect 18647 10016 18880 10044
rect 18647 10013 18659 10016
rect 18601 10007 18659 10013
rect 18874 10004 18880 10016
rect 18932 10044 18938 10056
rect 19242 10044 19248 10056
rect 18932 10016 19248 10044
rect 18932 10004 18938 10016
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 19886 10004 19892 10056
rect 19944 10044 19950 10056
rect 20349 10047 20407 10053
rect 20349 10044 20361 10047
rect 19944 10016 20361 10044
rect 19944 10004 19950 10016
rect 20349 10013 20361 10016
rect 20395 10013 20407 10047
rect 21266 10044 21272 10056
rect 21227 10016 21272 10044
rect 20349 10007 20407 10013
rect 21266 10004 21272 10016
rect 21324 10004 21330 10056
rect 17497 9979 17555 9985
rect 17497 9945 17509 9979
rect 17543 9945 17555 9979
rect 20714 9976 20720 9988
rect 17497 9939 17555 9945
rect 17972 9948 20720 9976
rect 17972 9908 18000 9948
rect 20714 9936 20720 9948
rect 20772 9936 20778 9988
rect 21174 9936 21180 9988
rect 21232 9976 21238 9988
rect 21514 9979 21572 9985
rect 21514 9976 21526 9979
rect 21232 9948 21526 9976
rect 21232 9936 21238 9948
rect 21514 9945 21526 9948
rect 21560 9945 21572 9979
rect 21514 9939 21572 9945
rect 18138 9908 18144 9920
rect 16592 9880 18000 9908
rect 18099 9880 18144 9908
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 20732 9908 20760 9936
rect 22649 9911 22707 9917
rect 22649 9908 22661 9911
rect 20732 9880 22661 9908
rect 22649 9877 22661 9880
rect 22695 9877 22707 9911
rect 22649 9871 22707 9877
rect 1104 9818 30820 9840
rect 1104 9766 10880 9818
rect 10932 9766 10944 9818
rect 10996 9766 11008 9818
rect 11060 9766 11072 9818
rect 11124 9766 11136 9818
rect 11188 9766 20811 9818
rect 20863 9766 20875 9818
rect 20927 9766 20939 9818
rect 20991 9766 21003 9818
rect 21055 9766 21067 9818
rect 21119 9766 30820 9818
rect 1104 9744 30820 9766
rect 3510 9704 3516 9716
rect 3471 9676 3516 9704
rect 3510 9664 3516 9676
rect 3568 9664 3574 9716
rect 13170 9664 13176 9716
rect 13228 9664 13234 9716
rect 13262 9664 13268 9716
rect 13320 9704 13326 9716
rect 13320 9676 15148 9704
rect 13320 9664 13326 9676
rect 2406 9645 2412 9648
rect 2400 9636 2412 9645
rect 2367 9608 2412 9636
rect 2400 9599 2412 9608
rect 2406 9596 2412 9599
rect 2464 9596 2470 9648
rect 3050 9596 3056 9648
rect 3108 9636 3114 9648
rect 6733 9639 6791 9645
rect 6733 9636 6745 9639
rect 3108 9608 6745 9636
rect 3108 9596 3114 9608
rect 6733 9605 6745 9608
rect 6779 9605 6791 9639
rect 6733 9599 6791 9605
rect 6825 9639 6883 9645
rect 6825 9605 6837 9639
rect 6871 9636 6883 9639
rect 7098 9636 7104 9648
rect 6871 9608 7104 9636
rect 6871 9605 6883 9608
rect 6825 9599 6883 9605
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 7653 9639 7711 9645
rect 7653 9605 7665 9639
rect 7699 9636 7711 9639
rect 8294 9636 8300 9648
rect 7699 9608 8300 9636
rect 7699 9605 7711 9608
rect 7653 9599 7711 9605
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 9858 9596 9864 9648
rect 9916 9636 9922 9648
rect 10686 9636 10692 9648
rect 9916 9608 10692 9636
rect 9916 9596 9922 9608
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 10873 9639 10931 9645
rect 10873 9605 10885 9639
rect 10919 9636 10931 9639
rect 13188 9636 13216 9664
rect 13722 9636 13728 9648
rect 10919 9608 13216 9636
rect 13372 9608 13728 9636
rect 10919 9605 10931 9608
rect 10873 9599 10931 9605
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 4062 9568 4068 9580
rect 4023 9540 4068 9568
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9568 4307 9571
rect 4522 9568 4528 9580
rect 4295 9540 4528 9568
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 5534 9568 5540 9580
rect 4663 9540 5540 9568
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 1670 9460 1676 9512
rect 1728 9500 1734 9512
rect 2133 9503 2191 9509
rect 2133 9500 2145 9503
rect 1728 9472 2145 9500
rect 1728 9460 1734 9472
rect 2133 9469 2145 9472
rect 2179 9469 2191 9503
rect 2133 9463 2191 9469
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 4356 9432 4384 9463
rect 4430 9460 4436 9512
rect 4488 9500 4494 9512
rect 5350 9500 5356 9512
rect 4488 9472 4533 9500
rect 4632 9472 5356 9500
rect 4488 9460 4494 9472
rect 4632 9432 4660 9472
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 5644 9500 5672 9531
rect 6546 9528 6552 9580
rect 6604 9577 6610 9580
rect 6604 9571 6663 9577
rect 6604 9537 6617 9571
rect 6651 9537 6663 9571
rect 7006 9568 7012 9580
rect 6967 9540 7012 9568
rect 6604 9531 6663 9537
rect 6604 9528 6610 9531
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 8110 9528 8116 9580
rect 8168 9568 8174 9580
rect 8168 9540 8616 9568
rect 8168 9528 8174 9540
rect 8202 9500 8208 9512
rect 5644 9472 7604 9500
rect 8163 9472 8208 9500
rect 4356 9404 4660 9432
rect 4706 9392 4712 9444
rect 4764 9432 4770 9444
rect 4764 9404 4936 9432
rect 4764 9392 4770 9404
rect 1486 9324 1492 9376
rect 1544 9364 1550 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 1544 9336 1593 9364
rect 1544 9324 1550 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 4798 9364 4804 9376
rect 4759 9336 4804 9364
rect 1581 9327 1639 9333
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 4908 9364 4936 9404
rect 5074 9392 5080 9444
rect 5132 9432 5138 9444
rect 5445 9435 5503 9441
rect 5445 9432 5457 9435
rect 5132 9404 5457 9432
rect 5132 9392 5138 9404
rect 5445 9401 5457 9404
rect 5491 9401 5503 9435
rect 5445 9395 5503 9401
rect 6730 9392 6736 9444
rect 6788 9432 6794 9444
rect 7009 9435 7067 9441
rect 7009 9432 7021 9435
rect 6788 9404 7021 9432
rect 6788 9392 6794 9404
rect 7009 9401 7021 9404
rect 7055 9401 7067 9435
rect 7009 9395 7067 9401
rect 7576 9376 7604 9472
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 8478 9500 8484 9512
rect 8439 9472 8484 9500
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 8588 9500 8616 9540
rect 10226 9528 10232 9580
rect 10284 9568 10290 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 10284 9540 11529 9568
rect 10284 9528 10290 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9568 12495 9571
rect 13372 9568 13400 9608
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 15120 9636 15148 9676
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 17313 9707 17371 9713
rect 17313 9704 17325 9707
rect 17276 9676 17325 9704
rect 17276 9664 17282 9676
rect 17313 9673 17325 9676
rect 17359 9673 17371 9707
rect 17313 9667 17371 9673
rect 17402 9664 17408 9716
rect 17460 9704 17466 9716
rect 19058 9704 19064 9716
rect 17460 9676 19064 9704
rect 17460 9664 17466 9676
rect 19058 9664 19064 9676
rect 19116 9664 19122 9716
rect 19242 9704 19248 9716
rect 19203 9676 19248 9704
rect 19242 9664 19248 9676
rect 19300 9664 19306 9716
rect 19797 9707 19855 9713
rect 19797 9673 19809 9707
rect 19843 9704 19855 9707
rect 20346 9704 20352 9716
rect 19843 9676 20352 9704
rect 19843 9673 19855 9676
rect 19797 9667 19855 9673
rect 20346 9664 20352 9676
rect 20404 9664 20410 9716
rect 16025 9639 16083 9645
rect 15120 9608 15424 9636
rect 12483 9540 13400 9568
rect 13449 9571 13507 9577
rect 12483 9537 12495 9540
rect 12437 9531 12495 9537
rect 13449 9537 13461 9571
rect 13495 9568 13507 9571
rect 13630 9568 13636 9580
rect 13495 9540 13636 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 14737 9571 14795 9577
rect 14737 9570 14749 9571
rect 14660 9568 14749 9570
rect 13740 9542 14749 9568
rect 13740 9540 14688 9542
rect 12161 9503 12219 9509
rect 12161 9500 12173 9503
rect 8588 9472 12173 9500
rect 12161 9469 12173 9472
rect 12207 9469 12219 9503
rect 12161 9463 12219 9469
rect 12986 9460 12992 9512
rect 13044 9500 13050 9512
rect 13740 9509 13768 9540
rect 14737 9537 14749 9542
rect 14783 9537 14795 9571
rect 14737 9531 14795 9537
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 13725 9503 13783 9509
rect 13725 9500 13737 9503
rect 13044 9472 13737 9500
rect 13044 9460 13050 9472
rect 13725 9469 13737 9472
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 13078 9392 13084 9444
rect 13136 9432 13142 9444
rect 14936 9432 14964 9531
rect 15102 9528 15108 9580
rect 15160 9568 15166 9580
rect 15286 9568 15292 9580
rect 15160 9540 15205 9568
rect 15247 9540 15292 9568
rect 15160 9528 15166 9540
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 15013 9503 15071 9509
rect 15013 9469 15025 9503
rect 15059 9500 15071 9503
rect 15396 9500 15424 9608
rect 16025 9605 16037 9639
rect 16071 9636 16083 9639
rect 16482 9636 16488 9648
rect 16071 9608 16488 9636
rect 16071 9605 16083 9608
rect 16025 9599 16083 9605
rect 16482 9596 16488 9608
rect 16540 9596 16546 9648
rect 18138 9645 18144 9648
rect 18132 9636 18144 9645
rect 18099 9608 18144 9636
rect 18132 9599 18144 9608
rect 18138 9596 18144 9599
rect 18196 9596 18202 9648
rect 15654 9528 15660 9580
rect 15712 9568 15718 9580
rect 15933 9571 15991 9577
rect 15933 9568 15945 9571
rect 15712 9540 15945 9568
rect 15712 9528 15718 9540
rect 15933 9537 15945 9540
rect 15979 9537 15991 9571
rect 17218 9568 17224 9580
rect 17179 9540 17224 9568
rect 15933 9531 15991 9537
rect 17218 9528 17224 9540
rect 17276 9528 17282 9580
rect 19705 9571 19763 9577
rect 19705 9568 19717 9571
rect 17328 9540 19717 9568
rect 15059 9472 15424 9500
rect 15059 9469 15071 9472
rect 15013 9463 15071 9469
rect 15746 9460 15752 9512
rect 15804 9500 15810 9512
rect 17328 9500 17356 9540
rect 19705 9537 19717 9540
rect 19751 9537 19763 9571
rect 19705 9531 19763 9537
rect 17862 9500 17868 9512
rect 15804 9472 17356 9500
rect 17823 9472 17868 9500
rect 15804 9460 15810 9472
rect 17862 9460 17868 9472
rect 17920 9460 17926 9512
rect 13136 9404 14964 9432
rect 13136 9392 13142 9404
rect 7374 9364 7380 9376
rect 4908 9336 7380 9364
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 7558 9364 7564 9376
rect 7519 9336 7564 9364
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 9582 9364 9588 9376
rect 9543 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 10008 9336 11621 9364
rect 10008 9324 10014 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 11609 9327 11667 9333
rect 13262 9324 13268 9376
rect 13320 9364 13326 9376
rect 15473 9367 15531 9373
rect 15473 9364 15485 9367
rect 13320 9336 15485 9364
rect 13320 9324 13326 9336
rect 15473 9333 15485 9336
rect 15519 9333 15531 9367
rect 15473 9327 15531 9333
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 19426 9364 19432 9376
rect 16356 9336 19432 9364
rect 16356 9324 16362 9336
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 20254 9324 20260 9376
rect 20312 9364 20318 9376
rect 21266 9364 21272 9376
rect 20312 9336 21272 9364
rect 20312 9324 20318 9336
rect 21266 9324 21272 9336
rect 21324 9364 21330 9376
rect 21542 9364 21548 9376
rect 21324 9336 21548 9364
rect 21324 9324 21330 9336
rect 21542 9324 21548 9336
rect 21600 9324 21606 9376
rect 1104 9274 30820 9296
rect 1104 9222 5915 9274
rect 5967 9222 5979 9274
rect 6031 9222 6043 9274
rect 6095 9222 6107 9274
rect 6159 9222 6171 9274
rect 6223 9222 15846 9274
rect 15898 9222 15910 9274
rect 15962 9222 15974 9274
rect 16026 9222 16038 9274
rect 16090 9222 16102 9274
rect 16154 9222 25776 9274
rect 25828 9222 25840 9274
rect 25892 9222 25904 9274
rect 25956 9222 25968 9274
rect 26020 9222 26032 9274
rect 26084 9222 30820 9274
rect 1104 9200 30820 9222
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 6457 9163 6515 9169
rect 3660 9132 6132 9160
rect 3660 9120 3666 9132
rect 2869 9027 2927 9033
rect 2869 8993 2881 9027
rect 2915 9024 2927 9027
rect 3234 9024 3240 9036
rect 2915 8996 3240 9024
rect 2915 8993 2927 8996
rect 2869 8987 2927 8993
rect 3234 8984 3240 8996
rect 3292 9024 3298 9036
rect 3786 9024 3792 9036
rect 3292 8996 3792 9024
rect 3292 8984 3298 8996
rect 3786 8984 3792 8996
rect 3844 8984 3850 9036
rect 5074 9024 5080 9036
rect 5035 8996 5080 9024
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 2590 8956 2596 8968
rect 2551 8928 2596 8956
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 4062 8956 4068 8968
rect 3975 8928 4068 8956
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 5344 8959 5402 8965
rect 5344 8925 5356 8959
rect 5390 8956 5402 8959
rect 5718 8956 5724 8968
rect 5390 8928 5724 8956
rect 5390 8925 5402 8928
rect 5344 8919 5402 8925
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 6104 8956 6132 9132
rect 6457 9129 6469 9163
rect 6503 9160 6515 9163
rect 6638 9160 6644 9172
rect 6503 9132 6644 9160
rect 6503 9129 6515 9132
rect 6457 9123 6515 9129
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 6880 9132 8432 9160
rect 6880 9120 6886 9132
rect 8404 9092 8432 9132
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 9677 9163 9735 9169
rect 9677 9160 9689 9163
rect 8536 9132 9689 9160
rect 8536 9120 8542 9132
rect 9677 9129 9689 9132
rect 9723 9129 9735 9163
rect 9677 9123 9735 9129
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 10192 9132 10241 9160
rect 10192 9120 10198 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 10229 9123 10287 9129
rect 13538 9120 13544 9172
rect 13596 9160 13602 9172
rect 17129 9163 17187 9169
rect 17129 9160 17141 9163
rect 13596 9132 17141 9160
rect 13596 9120 13602 9132
rect 17129 9129 17141 9132
rect 17175 9160 17187 9163
rect 17862 9160 17868 9172
rect 17175 9132 17868 9160
rect 17175 9129 17187 9132
rect 17129 9123 17187 9129
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 19797 9163 19855 9169
rect 19797 9129 19809 9163
rect 19843 9160 19855 9163
rect 20438 9160 20444 9172
rect 19843 9132 20444 9160
rect 19843 9129 19855 9132
rect 19797 9123 19855 9129
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 21085 9163 21143 9169
rect 21085 9129 21097 9163
rect 21131 9160 21143 9163
rect 21174 9160 21180 9172
rect 21131 9132 21180 9160
rect 21131 9129 21143 9132
rect 21085 9123 21143 9129
rect 21174 9120 21180 9132
rect 21232 9120 21238 9172
rect 11330 9092 11336 9104
rect 8404 9064 11336 9092
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 15565 9095 15623 9101
rect 15565 9061 15577 9095
rect 15611 9092 15623 9095
rect 16390 9092 16396 9104
rect 15611 9064 16396 9092
rect 15611 9061 15623 9064
rect 15565 9055 15623 9061
rect 16390 9052 16396 9064
rect 16448 9052 16454 9104
rect 17880 9092 17908 9120
rect 17880 9064 18175 9092
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 9024 9275 9027
rect 9766 9024 9772 9036
rect 9263 8996 9772 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 10873 9027 10931 9033
rect 10873 8993 10885 9027
rect 10919 9024 10931 9027
rect 11882 9024 11888 9036
rect 10919 8996 11888 9024
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 18147 9024 18175 9064
rect 18230 9052 18236 9104
rect 18288 9092 18294 9104
rect 18288 9064 20392 9092
rect 18288 9052 18294 9064
rect 20254 9024 20260 9036
rect 18147 8996 20260 9024
rect 20254 8984 20260 8996
rect 20312 8984 20318 9036
rect 20364 8968 20392 9064
rect 20625 9027 20683 9033
rect 20625 8993 20637 9027
rect 20671 9024 20683 9027
rect 21266 9024 21272 9036
rect 20671 8996 21272 9024
rect 20671 8993 20683 8996
rect 20625 8987 20683 8993
rect 21266 8984 21272 8996
rect 21324 8984 21330 9036
rect 21542 9024 21548 9036
rect 21503 8996 21548 9024
rect 21542 8984 21548 8996
rect 21600 8984 21606 9036
rect 8294 8956 8300 8968
rect 6104 8928 8156 8956
rect 8255 8928 8300 8956
rect 4080 8888 4108 8916
rect 6270 8888 6276 8900
rect 4080 8860 6276 8888
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 6380 8860 7236 8888
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 3602 8780 3608 8832
rect 3660 8820 3666 8832
rect 6380 8820 6408 8860
rect 3660 8792 6408 8820
rect 6917 8823 6975 8829
rect 3660 8780 3666 8792
rect 6917 8789 6929 8823
rect 6963 8820 6975 8823
rect 7098 8820 7104 8832
rect 6963 8792 7104 8820
rect 6963 8789 6975 8792
rect 6917 8783 6975 8789
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 7208 8820 7236 8860
rect 7282 8848 7288 8900
rect 7340 8888 7346 8900
rect 8030 8891 8088 8897
rect 8030 8888 8042 8891
rect 7340 8860 8042 8888
rect 7340 8848 7346 8860
rect 8030 8857 8042 8860
rect 8076 8857 8088 8891
rect 8128 8888 8156 8928
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 8386 8916 8392 8968
rect 8444 8956 8450 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8444 8928 8953 8956
rect 8444 8916 8450 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9306 8956 9312 8968
rect 9267 8928 9312 8956
rect 9125 8919 9183 8925
rect 9140 8888 9168 8919
rect 9306 8916 9312 8928
rect 9364 8916 9370 8968
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8956 9551 8959
rect 9582 8956 9588 8968
rect 9539 8928 9588 8956
rect 9539 8925 9551 8928
rect 9493 8919 9551 8925
rect 8128 8860 9168 8888
rect 9508 8888 9536 8919
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 10597 8959 10655 8965
rect 10597 8925 10609 8959
rect 10643 8956 10655 8959
rect 11422 8956 11428 8968
rect 10643 8928 11428 8956
rect 10643 8925 10655 8928
rect 10597 8919 10655 8925
rect 11422 8916 11428 8928
rect 11480 8916 11486 8968
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 11974 8956 11980 8968
rect 11655 8928 11980 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 13262 8916 13268 8968
rect 13320 8965 13326 8968
rect 13320 8956 13332 8965
rect 13538 8956 13544 8968
rect 13320 8928 13365 8956
rect 13499 8928 13544 8956
rect 13320 8919 13332 8928
rect 13320 8916 13326 8919
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 14185 8959 14243 8965
rect 14185 8925 14197 8959
rect 14231 8956 14243 8959
rect 14231 8928 15516 8956
rect 14231 8925 14243 8928
rect 14185 8919 14243 8925
rect 14090 8888 14096 8900
rect 9508 8860 14096 8888
rect 8030 8851 8088 8857
rect 14090 8848 14096 8860
rect 14148 8848 14154 8900
rect 14452 8891 14510 8897
rect 14452 8857 14464 8891
rect 14498 8888 14510 8891
rect 14826 8888 14832 8900
rect 14498 8860 14832 8888
rect 14498 8857 14510 8860
rect 14452 8851 14510 8857
rect 14826 8848 14832 8860
rect 14884 8848 14890 8900
rect 15488 8888 15516 8928
rect 15562 8916 15568 8968
rect 15620 8956 15626 8968
rect 16393 8959 16451 8965
rect 16393 8956 16405 8959
rect 15620 8928 16405 8956
rect 15620 8916 15626 8928
rect 16393 8925 16405 8928
rect 16439 8956 16451 8959
rect 17037 8959 17095 8965
rect 17037 8956 17049 8959
rect 16439 8928 17049 8956
rect 16439 8925 16451 8928
rect 16393 8919 16451 8925
rect 17037 8925 17049 8928
rect 17083 8925 17095 8959
rect 17770 8956 17776 8968
rect 17731 8928 17776 8956
rect 17037 8919 17095 8925
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 17957 8957 18015 8963
rect 17957 8956 17969 8957
rect 17880 8928 17969 8956
rect 15488 8860 16344 8888
rect 8110 8820 8116 8832
rect 7208 8792 8116 8820
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 10689 8823 10747 8829
rect 10689 8820 10701 8823
rect 10284 8792 10701 8820
rect 10284 8780 10290 8792
rect 10689 8789 10701 8792
rect 10735 8789 10747 8823
rect 11514 8820 11520 8832
rect 11475 8792 11520 8820
rect 10689 8783 10747 8789
rect 11514 8780 11520 8792
rect 11572 8780 11578 8832
rect 12158 8820 12164 8832
rect 12119 8792 12164 8820
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 12894 8780 12900 8832
rect 12952 8820 12958 8832
rect 15286 8820 15292 8832
rect 12952 8792 15292 8820
rect 12952 8780 12958 8792
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 16316 8829 16344 8860
rect 16301 8823 16359 8829
rect 16301 8789 16313 8823
rect 16347 8820 16359 8823
rect 16482 8820 16488 8832
rect 16347 8792 16488 8820
rect 16347 8789 16359 8792
rect 16301 8783 16359 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 17880 8820 17908 8928
rect 17957 8923 17969 8928
rect 18003 8923 18015 8957
rect 17957 8917 18015 8923
rect 18043 8959 18101 8965
rect 18043 8925 18055 8959
rect 18089 8925 18101 8959
rect 18043 8919 18101 8925
rect 18058 8888 18086 8919
rect 18138 8916 18144 8968
rect 18196 8965 18202 8968
rect 18196 8959 18245 8965
rect 18196 8925 18199 8959
rect 18233 8925 18245 8959
rect 18196 8919 18245 8925
rect 18196 8916 18202 8919
rect 18322 8916 18328 8968
rect 18380 8956 18386 8968
rect 19705 8959 19763 8965
rect 18380 8928 18425 8956
rect 18380 8916 18386 8928
rect 19705 8925 19717 8959
rect 19751 8925 19763 8959
rect 20346 8956 20352 8968
rect 20259 8928 20352 8956
rect 19705 8919 19763 8925
rect 18782 8888 18788 8900
rect 18058 8860 18788 8888
rect 18782 8848 18788 8860
rect 18840 8848 18846 8900
rect 18874 8848 18880 8900
rect 18932 8888 18938 8900
rect 19720 8888 19748 8919
rect 20346 8916 20352 8928
rect 20404 8916 20410 8968
rect 20530 8956 20536 8968
rect 20491 8928 20536 8956
rect 20530 8916 20536 8928
rect 20588 8916 20594 8968
rect 20714 8956 20720 8968
rect 20675 8928 20720 8956
rect 20714 8916 20720 8928
rect 20772 8916 20778 8968
rect 20898 8916 20904 8968
rect 20956 8956 20962 8968
rect 29822 8956 29828 8968
rect 20956 8928 21001 8956
rect 29783 8928 29828 8956
rect 20956 8916 20962 8928
rect 29822 8916 29828 8928
rect 29880 8916 29886 8968
rect 18932 8860 19748 8888
rect 18932 8848 18938 8860
rect 19794 8848 19800 8900
rect 19852 8888 19858 8900
rect 21634 8888 21640 8900
rect 19852 8860 21640 8888
rect 19852 8848 19858 8860
rect 21634 8848 21640 8860
rect 21692 8848 21698 8900
rect 21818 8897 21824 8900
rect 21812 8851 21824 8897
rect 21876 8888 21882 8900
rect 21876 8860 21912 8888
rect 21818 8848 21824 8851
rect 21876 8848 21882 8860
rect 18414 8820 18420 8832
rect 17880 8792 18420 8820
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 18509 8823 18567 8829
rect 18509 8789 18521 8823
rect 18555 8820 18567 8823
rect 18690 8820 18696 8832
rect 18555 8792 18696 8820
rect 18555 8789 18567 8792
rect 18509 8783 18567 8789
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 19058 8780 19064 8832
rect 19116 8820 19122 8832
rect 22002 8820 22008 8832
rect 19116 8792 22008 8820
rect 19116 8780 19122 8792
rect 22002 8780 22008 8792
rect 22060 8820 22066 8832
rect 22925 8823 22983 8829
rect 22925 8820 22937 8823
rect 22060 8792 22937 8820
rect 22060 8780 22066 8792
rect 22925 8789 22937 8792
rect 22971 8789 22983 8823
rect 30006 8820 30012 8832
rect 29967 8792 30012 8820
rect 22925 8783 22983 8789
rect 30006 8780 30012 8792
rect 30064 8780 30070 8832
rect 1104 8730 30820 8752
rect 1104 8678 10880 8730
rect 10932 8678 10944 8730
rect 10996 8678 11008 8730
rect 11060 8678 11072 8730
rect 11124 8678 11136 8730
rect 11188 8678 20811 8730
rect 20863 8678 20875 8730
rect 20927 8678 20939 8730
rect 20991 8678 21003 8730
rect 21055 8678 21067 8730
rect 21119 8678 30820 8730
rect 1104 8656 30820 8678
rect 3050 8616 3056 8628
rect 3011 8588 3056 8616
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 3602 8616 3608 8628
rect 3563 8588 3608 8616
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 3786 8576 3792 8628
rect 3844 8616 3850 8628
rect 3844 8588 5488 8616
rect 3844 8576 3850 8588
rect 5074 8548 5080 8560
rect 4264 8520 5080 8548
rect 1670 8480 1676 8492
rect 1631 8452 1676 8480
rect 1670 8440 1676 8452
rect 1728 8440 1734 8492
rect 1940 8483 1998 8489
rect 1940 8449 1952 8483
rect 1986 8480 1998 8483
rect 2222 8480 2228 8492
rect 1986 8452 2228 8480
rect 1986 8449 1998 8452
rect 1940 8443 1998 8449
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 3786 8480 3792 8492
rect 3747 8452 3792 8480
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4264 8489 4292 8520
rect 5074 8508 5080 8520
rect 5132 8508 5138 8560
rect 5460 8548 5488 8588
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 5629 8619 5687 8625
rect 5629 8616 5641 8619
rect 5592 8588 5641 8616
rect 5592 8576 5598 8588
rect 5629 8585 5641 8588
rect 5675 8585 5687 8619
rect 5629 8579 5687 8585
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 8352 8588 10793 8616
rect 8352 8576 8358 8588
rect 10781 8585 10793 8588
rect 10827 8585 10839 8619
rect 10781 8579 10839 8585
rect 11517 8619 11575 8625
rect 11517 8585 11529 8619
rect 11563 8616 11575 8619
rect 11698 8616 11704 8628
rect 11563 8588 11704 8616
rect 11563 8585 11575 8588
rect 11517 8579 11575 8585
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 12158 8576 12164 8628
rect 12216 8616 12222 8628
rect 12894 8616 12900 8628
rect 12216 8588 12900 8616
rect 12216 8576 12222 8588
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13004 8588 17172 8616
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 5460 8520 6377 8548
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 6365 8511 6423 8517
rect 6546 8508 6552 8560
rect 6604 8508 6610 8560
rect 7558 8508 7564 8560
rect 7616 8548 7622 8560
rect 10873 8551 10931 8557
rect 10873 8548 10885 8551
rect 7616 8520 10885 8548
rect 7616 8508 7622 8520
rect 10873 8517 10885 8520
rect 10919 8517 10931 8551
rect 10873 8511 10931 8517
rect 11330 8508 11336 8560
rect 11388 8548 11394 8560
rect 13004 8548 13032 8588
rect 13630 8548 13636 8560
rect 11388 8520 13032 8548
rect 13096 8520 13636 8548
rect 11388 8508 11394 8520
rect 4249 8483 4307 8489
rect 4249 8480 4261 8483
rect 4212 8452 4261 8480
rect 4212 8440 4218 8452
rect 4249 8449 4261 8452
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 4516 8483 4574 8489
rect 4516 8449 4528 8483
rect 4562 8480 4574 8483
rect 4798 8480 4804 8492
rect 4562 8452 4804 8480
rect 4562 8449 4574 8452
rect 4516 8443 4574 8449
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 6564 8480 6592 8508
rect 5644 8452 6592 8480
rect 5644 8424 5672 8452
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 8297 8483 8355 8489
rect 8297 8480 8309 8483
rect 6880 8452 8309 8480
rect 6880 8440 6886 8452
rect 8297 8449 8309 8452
rect 8343 8449 8355 8483
rect 9950 8480 9956 8492
rect 9911 8452 9956 8480
rect 8297 8443 8355 8449
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10686 8480 10692 8492
rect 10275 8452 10692 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12894 8480 12900 8492
rect 11931 8452 12900 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13096 8489 13124 8520
rect 13630 8508 13636 8520
rect 13688 8508 13694 8560
rect 14476 8520 17080 8548
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 13538 8440 13544 8492
rect 13596 8480 13602 8492
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 13596 8452 14381 8480
rect 13596 8440 13602 8452
rect 14369 8449 14381 8452
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 5626 8372 5632 8424
rect 5684 8372 5690 8424
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8412 6423 8415
rect 6457 8415 6515 8421
rect 6457 8412 6469 8415
rect 6411 8384 6469 8412
rect 6411 8381 6423 8384
rect 6365 8375 6423 8381
rect 6457 8381 6469 8384
rect 6503 8381 6515 8415
rect 6457 8375 6515 8381
rect 6546 8372 6552 8424
rect 6604 8412 6610 8424
rect 6733 8415 6791 8421
rect 6733 8412 6745 8415
rect 6604 8384 6745 8412
rect 6604 8372 6610 8384
rect 6733 8381 6745 8384
rect 6779 8381 6791 8415
rect 6733 8375 6791 8381
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 8444 8384 8585 8412
rect 8444 8372 8450 8384
rect 8573 8381 8585 8384
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 10137 8415 10195 8421
rect 9364 8384 9904 8412
rect 9364 8372 9370 8384
rect 9674 8304 9680 8356
rect 9732 8344 9738 8356
rect 9769 8347 9827 8353
rect 9769 8344 9781 8347
rect 9732 8316 9781 8344
rect 9732 8304 9738 8316
rect 9769 8313 9781 8316
rect 9815 8313 9827 8347
rect 9876 8344 9904 8384
rect 10137 8381 10149 8415
rect 10183 8412 10195 8415
rect 11974 8412 11980 8424
rect 10183 8384 11980 8412
rect 10183 8381 10195 8384
rect 10137 8375 10195 8381
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12069 8415 12127 8421
rect 12069 8381 12081 8415
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8412 13415 8415
rect 13998 8412 14004 8424
rect 13403 8384 14004 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 9876 8316 11836 8344
rect 9769 8307 9827 8313
rect 2406 8236 2412 8288
rect 2464 8276 2470 8288
rect 9398 8276 9404 8288
rect 2464 8248 9404 8276
rect 2464 8236 2470 8248
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 10134 8276 10140 8288
rect 10095 8248 10140 8276
rect 10134 8236 10140 8248
rect 10192 8236 10198 8288
rect 11808 8276 11836 8316
rect 11882 8304 11888 8356
rect 11940 8344 11946 8356
rect 12084 8344 12112 8375
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 14476 8412 14504 8520
rect 14642 8489 14648 8492
rect 14636 8443 14648 8489
rect 14700 8480 14706 8492
rect 14700 8452 14736 8480
rect 14642 8440 14648 8443
rect 14700 8440 14706 8452
rect 14384 8384 14504 8412
rect 17052 8412 17080 8520
rect 17144 8489 17172 8588
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 19794 8616 19800 8628
rect 18472 8588 19800 8616
rect 18472 8576 18478 8588
rect 19794 8576 19800 8588
rect 19852 8576 19858 8628
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 21818 8616 21824 8628
rect 20404 8588 21496 8616
rect 21779 8588 21824 8616
rect 20404 8576 20410 8588
rect 21358 8548 21364 8560
rect 20732 8520 21364 8548
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8480 17187 8483
rect 17310 8480 17316 8492
rect 17175 8452 17316 8480
rect 17175 8449 17187 8452
rect 17129 8443 17187 8449
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 17770 8480 17776 8492
rect 17451 8452 17776 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 17770 8440 17776 8452
rect 17828 8440 17834 8492
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 18417 8483 18475 8489
rect 18417 8480 18429 8483
rect 17920 8452 18429 8480
rect 17920 8440 17926 8452
rect 18417 8449 18429 8452
rect 18463 8449 18475 8483
rect 18690 8480 18696 8492
rect 18651 8452 18696 8480
rect 18417 8443 18475 8449
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 20732 8489 20760 8520
rect 21358 8508 21364 8520
rect 21416 8508 21422 8560
rect 21468 8548 21496 8588
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 29822 8576 29828 8628
rect 29880 8616 29886 8628
rect 30009 8619 30067 8625
rect 30009 8616 30021 8619
rect 29880 8588 30021 8616
rect 29880 8576 29886 8588
rect 30009 8585 30021 8588
rect 30055 8585 30067 8619
rect 30009 8579 30067 8585
rect 21468 8520 22600 8548
rect 20717 8483 20775 8489
rect 20717 8449 20729 8483
rect 20763 8449 20775 8483
rect 20717 8443 20775 8449
rect 21085 8483 21143 8489
rect 21085 8449 21097 8483
rect 21131 8480 21143 8483
rect 21174 8480 21180 8492
rect 21131 8452 21180 8480
rect 21131 8449 21143 8452
rect 21085 8443 21143 8449
rect 21174 8440 21180 8452
rect 21232 8440 21238 8492
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21468 8480 21496 8520
rect 22002 8480 22008 8492
rect 21315 8452 21496 8480
rect 21963 8452 22008 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 22186 8440 22192 8492
rect 22244 8480 22250 8492
rect 22370 8480 22376 8492
rect 22244 8452 22289 8480
rect 22331 8452 22376 8480
rect 22244 8440 22250 8452
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 22572 8489 22600 8520
rect 22557 8483 22615 8489
rect 22557 8449 22569 8483
rect 22603 8449 22615 8483
rect 29914 8480 29920 8492
rect 29875 8452 29920 8480
rect 22557 8443 22615 8449
rect 29914 8440 29920 8452
rect 29972 8440 29978 8492
rect 30098 8480 30104 8492
rect 30059 8452 30104 8480
rect 30098 8440 30104 8452
rect 30156 8440 30162 8492
rect 17052 8384 19380 8412
rect 14384 8344 14412 8384
rect 15746 8344 15752 8356
rect 11940 8316 12112 8344
rect 12176 8316 14412 8344
rect 15707 8316 15752 8344
rect 11940 8304 11946 8316
rect 12176 8276 12204 8316
rect 15746 8304 15752 8316
rect 15804 8304 15810 8356
rect 19352 8344 19380 8384
rect 19426 8372 19432 8424
rect 19484 8412 19490 8424
rect 20438 8412 20444 8424
rect 19484 8384 20444 8412
rect 19484 8372 19490 8384
rect 20438 8372 20444 8384
rect 20496 8412 20502 8424
rect 20901 8415 20959 8421
rect 20901 8412 20913 8415
rect 20496 8384 20913 8412
rect 20496 8372 20502 8384
rect 20901 8381 20913 8384
rect 20947 8381 20959 8415
rect 20901 8375 20959 8381
rect 20993 8415 21051 8421
rect 20993 8381 21005 8415
rect 21039 8381 21051 8415
rect 20993 8375 21051 8381
rect 22281 8415 22339 8421
rect 22281 8381 22293 8415
rect 22327 8381 22339 8415
rect 22281 8375 22339 8381
rect 20714 8344 20720 8356
rect 19352 8316 20720 8344
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 21008 8344 21036 8375
rect 21266 8344 21272 8356
rect 21008 8316 21272 8344
rect 21266 8304 21272 8316
rect 21324 8344 21330 8356
rect 22296 8344 22324 8375
rect 21324 8316 22324 8344
rect 21324 8304 21330 8316
rect 11808 8248 12204 8276
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 15764 8276 15792 8304
rect 20530 8276 20536 8288
rect 15344 8248 15792 8276
rect 20491 8248 20536 8276
rect 15344 8236 15350 8248
rect 20530 8236 20536 8248
rect 20588 8236 20594 8288
rect 20732 8276 20760 8304
rect 22186 8276 22192 8288
rect 20732 8248 22192 8276
rect 22186 8236 22192 8248
rect 22244 8236 22250 8288
rect 1104 8186 30820 8208
rect 1104 8134 5915 8186
rect 5967 8134 5979 8186
rect 6031 8134 6043 8186
rect 6095 8134 6107 8186
rect 6159 8134 6171 8186
rect 6223 8134 15846 8186
rect 15898 8134 15910 8186
rect 15962 8134 15974 8186
rect 16026 8134 16038 8186
rect 16090 8134 16102 8186
rect 16154 8134 25776 8186
rect 25828 8134 25840 8186
rect 25892 8134 25904 8186
rect 25956 8134 25968 8186
rect 26020 8134 26032 8186
rect 26084 8134 30820 8186
rect 1104 8112 30820 8134
rect 2222 8072 2228 8084
rect 2183 8044 2228 8072
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 5040 8044 5089 8072
rect 5040 8032 5046 8044
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 5077 8035 5135 8041
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 7282 8072 7288 8084
rect 6788 8044 7052 8072
rect 7243 8044 7288 8072
rect 6788 8032 6794 8044
rect 2038 7964 2044 8016
rect 2096 7964 2102 8016
rect 5442 7964 5448 8016
rect 5500 8004 5506 8016
rect 5810 8004 5816 8016
rect 5500 7976 5816 8004
rect 5500 7964 5506 7976
rect 5810 7964 5816 7976
rect 5868 8004 5874 8016
rect 7024 8004 7052 8044
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8041 9551 8075
rect 10042 8072 10048 8084
rect 10003 8044 10048 8072
rect 9493 8035 9551 8041
rect 9214 8004 9220 8016
rect 5868 7976 6960 8004
rect 7024 7976 9220 8004
rect 5868 7964 5874 7976
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7936 1915 7939
rect 2056 7936 2084 7964
rect 4062 7936 4068 7948
rect 1903 7908 2084 7936
rect 3975 7908 4068 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 4062 7896 4068 7908
rect 4120 7936 4126 7948
rect 4430 7936 4436 7948
rect 4120 7908 4436 7936
rect 4120 7896 4126 7908
rect 4430 7896 4436 7908
rect 4488 7936 4494 7948
rect 6932 7945 6960 7976
rect 9214 7964 9220 7976
rect 9272 7964 9278 8016
rect 9508 8004 9536 8035
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 10505 8075 10563 8081
rect 10505 8041 10517 8075
rect 10551 8072 10563 8075
rect 11974 8072 11980 8084
rect 10551 8044 11980 8072
rect 10551 8041 10563 8044
rect 10505 8035 10563 8041
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 12124 8044 12265 8072
rect 12124 8032 12130 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 12894 8072 12900 8084
rect 12855 8044 12900 8072
rect 12253 8035 12311 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 17405 8075 17463 8081
rect 17405 8072 17417 8075
rect 15396 8044 17417 8072
rect 10134 8004 10140 8016
rect 9508 7976 10140 8004
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 6917 7939 6975 7945
rect 4488 7908 5488 7936
rect 4488 7896 4494 7908
rect 5460 7880 5488 7908
rect 6917 7905 6929 7939
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 9401 7939 9459 7945
rect 9401 7905 9413 7939
rect 9447 7936 9459 7939
rect 11514 7936 11520 7948
rect 9447 7908 11520 7936
rect 9447 7905 9459 7908
rect 9401 7899 9459 7905
rect 11514 7896 11520 7908
rect 11572 7896 11578 7948
rect 11701 7939 11759 7945
rect 11701 7905 11713 7939
rect 11747 7936 11759 7939
rect 11882 7936 11888 7948
rect 11747 7908 11888 7936
rect 11747 7905 11759 7908
rect 11701 7899 11759 7905
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 14185 7939 14243 7945
rect 14185 7936 14197 7939
rect 12912 7908 14197 7936
rect 1489 7871 1547 7877
rect 1489 7837 1501 7871
rect 1535 7837 1547 7871
rect 1489 7831 1547 7837
rect 1504 7800 1532 7831
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 1673 7871 1731 7877
rect 1673 7868 1685 7871
rect 1636 7840 1685 7868
rect 1636 7828 1642 7840
rect 1673 7837 1685 7840
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7868 1823 7871
rect 1946 7868 1952 7880
rect 1811 7840 1952 7868
rect 1811 7837 1823 7840
rect 1765 7831 1823 7837
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 3050 7868 3056 7880
rect 2087 7840 3056 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 3786 7868 3792 7880
rect 3747 7840 3792 7868
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 5258 7868 5264 7880
rect 5219 7840 5264 7868
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5442 7868 5448 7880
rect 5403 7840 5448 7868
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7868 5871 7871
rect 6270 7868 6276 7880
rect 5859 7840 6276 7868
rect 5859 7837 5871 7840
rect 5813 7831 5871 7837
rect 2590 7800 2596 7812
rect 1504 7772 2596 7800
rect 1596 7744 1624 7772
rect 2590 7760 2596 7772
rect 2648 7760 2654 7812
rect 5074 7760 5080 7812
rect 5132 7800 5138 7812
rect 5350 7800 5356 7812
rect 5132 7772 5356 7800
rect 5132 7760 5138 7772
rect 5350 7760 5356 7772
rect 5408 7800 5414 7812
rect 5552 7800 5580 7831
rect 5408 7772 5580 7800
rect 5644 7800 5672 7831
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 6546 7868 6552 7880
rect 6507 7840 6552 7868
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 6730 7868 6736 7880
rect 6691 7840 6736 7868
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 7098 7868 7104 7880
rect 6880 7840 6925 7868
rect 7059 7840 7104 7868
rect 6880 7828 6886 7840
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 7926 7868 7932 7880
rect 7208 7840 7932 7868
rect 7208 7800 7236 7840
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7837 9551 7871
rect 10226 7868 10232 7880
rect 10187 7840 10232 7868
rect 9493 7831 9551 7837
rect 7834 7800 7840 7812
rect 5644 7772 7236 7800
rect 7795 7772 7840 7800
rect 5408 7760 5414 7772
rect 6748 7744 6776 7772
rect 7834 7760 7840 7772
rect 7892 7760 7898 7812
rect 8021 7803 8079 7809
rect 8021 7769 8033 7803
rect 8067 7800 8079 7803
rect 8478 7800 8484 7812
rect 8067 7772 8484 7800
rect 8067 7769 8079 7772
rect 8021 7763 8079 7769
rect 8478 7760 8484 7772
rect 8536 7760 8542 7812
rect 9508 7800 9536 7831
rect 10226 7828 10232 7840
rect 10284 7828 10290 7880
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 11532 7868 11560 7896
rect 12912 7877 12940 7908
rect 14185 7905 14197 7908
rect 14231 7905 14243 7939
rect 14185 7899 14243 7905
rect 14550 7896 14556 7948
rect 14608 7936 14614 7948
rect 15105 7939 15163 7945
rect 15105 7936 15117 7939
rect 14608 7908 15117 7936
rect 14608 7896 14614 7908
rect 15105 7905 15117 7908
rect 15151 7905 15163 7939
rect 15105 7899 15163 7905
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 10376 7840 10421 7868
rect 11532 7840 12725 7868
rect 10376 7828 10382 7840
rect 12713 7837 12725 7840
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7837 12955 7871
rect 14090 7868 14096 7880
rect 14051 7840 14096 7868
rect 12897 7831 12955 7837
rect 10505 7803 10563 7809
rect 10505 7800 10517 7803
rect 9508 7772 10517 7800
rect 10505 7769 10517 7772
rect 10551 7800 10563 7803
rect 10686 7800 10692 7812
rect 10551 7772 10692 7800
rect 10551 7769 10563 7772
rect 10505 7763 10563 7769
rect 10686 7760 10692 7772
rect 10744 7760 10750 7812
rect 11698 7760 11704 7812
rect 11756 7800 11762 7812
rect 12912 7800 12940 7831
rect 14090 7828 14096 7840
rect 14148 7828 14154 7880
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7868 14335 7871
rect 14366 7868 14372 7880
rect 14323 7840 14372 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 14366 7828 14372 7840
rect 14424 7828 14430 7880
rect 14826 7870 14832 7880
rect 14752 7868 14832 7870
rect 14660 7842 14832 7868
rect 14660 7840 14780 7842
rect 11756 7772 12940 7800
rect 11756 7760 11762 7772
rect 13998 7760 14004 7812
rect 14056 7800 14062 7812
rect 14660 7800 14688 7840
rect 14826 7828 14832 7842
rect 14884 7870 14890 7880
rect 15013 7871 15071 7877
rect 14884 7842 14975 7870
rect 14884 7828 14890 7842
rect 15013 7837 15025 7871
rect 15059 7837 15071 7871
rect 15194 7868 15200 7880
rect 15155 7840 15200 7868
rect 15013 7831 15071 7837
rect 14056 7772 14688 7800
rect 15028 7800 15056 7831
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 15396 7877 15424 8044
rect 17405 8041 17417 8044
rect 17451 8072 17463 8075
rect 18874 8072 18880 8084
rect 17451 8044 18880 8072
rect 17451 8041 17463 8044
rect 17405 8035 17463 8041
rect 18874 8032 18880 8044
rect 18932 8032 18938 8084
rect 21269 8075 21327 8081
rect 21269 8041 21281 8075
rect 21315 8072 21327 8075
rect 21358 8072 21364 8084
rect 21315 8044 21364 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 21358 8032 21364 8044
rect 21416 8032 21422 8084
rect 18509 8007 18567 8013
rect 18509 7973 18521 8007
rect 18555 8004 18567 8007
rect 19426 8004 19432 8016
rect 18555 7976 19432 8004
rect 18555 7973 18567 7976
rect 18509 7967 18567 7973
rect 19426 7964 19432 7976
rect 19484 7964 19490 8016
rect 15381 7871 15439 7877
rect 15381 7837 15393 7871
rect 15427 7837 15439 7871
rect 15381 7831 15439 7837
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7868 16083 7871
rect 16071 7840 16528 7868
rect 16071 7837 16083 7840
rect 16025 7831 16083 7837
rect 16500 7812 16528 7840
rect 19702 7828 19708 7880
rect 19760 7868 19766 7880
rect 19889 7871 19947 7877
rect 19889 7868 19901 7871
rect 19760 7840 19901 7868
rect 19760 7828 19766 7840
rect 19889 7837 19901 7840
rect 19935 7837 19947 7871
rect 19889 7831 19947 7837
rect 20156 7871 20214 7877
rect 20156 7837 20168 7871
rect 20202 7868 20214 7871
rect 20530 7868 20536 7880
rect 20202 7840 20536 7868
rect 20202 7837 20214 7840
rect 20156 7831 20214 7837
rect 20530 7828 20536 7840
rect 20588 7828 20594 7880
rect 15470 7800 15476 7812
rect 15028 7772 15476 7800
rect 14056 7760 14062 7772
rect 15470 7760 15476 7772
rect 15528 7760 15534 7812
rect 15565 7803 15623 7809
rect 15565 7769 15577 7803
rect 15611 7800 15623 7803
rect 16270 7803 16328 7809
rect 16270 7800 16282 7803
rect 15611 7772 16282 7800
rect 15611 7769 15623 7772
rect 15565 7763 15623 7769
rect 16270 7769 16282 7772
rect 16316 7769 16328 7803
rect 16270 7763 16328 7769
rect 16482 7760 16488 7812
rect 16540 7760 16546 7812
rect 18046 7760 18052 7812
rect 18104 7800 18110 7812
rect 18325 7803 18383 7809
rect 18325 7800 18337 7803
rect 18104 7772 18337 7800
rect 18104 7760 18110 7772
rect 18325 7769 18337 7772
rect 18371 7769 18383 7803
rect 18325 7763 18383 7769
rect 1578 7692 1584 7744
rect 1636 7692 1642 7744
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 6638 7732 6644 7744
rect 4856 7704 6644 7732
rect 4856 7692 4862 7704
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 6730 7692 6736 7744
rect 6788 7692 6794 7744
rect 7190 7692 7196 7744
rect 7248 7732 7254 7744
rect 9030 7732 9036 7744
rect 7248 7704 9036 7732
rect 7248 7692 7254 7704
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9125 7735 9183 7741
rect 9125 7701 9137 7735
rect 9171 7732 9183 7735
rect 9490 7732 9496 7744
rect 9171 7704 9496 7732
rect 9171 7701 9183 7704
rect 9125 7695 9183 7701
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 11790 7732 11796 7744
rect 10652 7704 11796 7732
rect 10652 7692 10658 7704
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 11940 7704 11985 7732
rect 11940 7692 11946 7704
rect 1104 7642 30820 7664
rect 1104 7590 10880 7642
rect 10932 7590 10944 7642
rect 10996 7590 11008 7642
rect 11060 7590 11072 7642
rect 11124 7590 11136 7642
rect 11188 7590 20811 7642
rect 20863 7590 20875 7642
rect 20927 7590 20939 7642
rect 20991 7590 21003 7642
rect 21055 7590 21067 7642
rect 21119 7590 30820 7642
rect 1104 7568 30820 7590
rect 2038 7488 2044 7540
rect 2096 7488 2102 7540
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7528 2283 7531
rect 4338 7528 4344 7540
rect 2271 7500 4344 7528
rect 2271 7497 2283 7500
rect 2225 7491 2283 7497
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 6457 7531 6515 7537
rect 6457 7528 6469 7531
rect 5644 7500 6469 7528
rect 1762 7420 1768 7472
rect 1820 7460 1826 7472
rect 2056 7460 2084 7488
rect 2777 7463 2835 7469
rect 2777 7460 2789 7463
rect 1820 7432 2789 7460
rect 1820 7420 1826 7432
rect 2777 7429 2789 7432
rect 2823 7429 2835 7463
rect 2777 7423 2835 7429
rect 2961 7463 3019 7469
rect 2961 7429 2973 7463
rect 3007 7460 3019 7463
rect 3786 7460 3792 7472
rect 3007 7432 3792 7460
rect 3007 7429 3019 7432
rect 2961 7423 3019 7429
rect 3786 7420 3792 7432
rect 3844 7460 3850 7472
rect 5644 7469 5672 7500
rect 6457 7497 6469 7500
rect 6503 7528 6515 7531
rect 7834 7528 7840 7540
rect 6503 7500 7840 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 10134 7528 10140 7540
rect 10095 7500 10140 7528
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 10318 7488 10324 7540
rect 10376 7528 10382 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 10376 7500 12173 7528
rect 10376 7488 10382 7500
rect 5629 7463 5687 7469
rect 5629 7460 5641 7463
rect 3844 7432 5641 7460
rect 3844 7420 3850 7432
rect 5629 7429 5641 7432
rect 5675 7429 5687 7463
rect 5810 7460 5816 7472
rect 5771 7432 5816 7460
rect 5629 7423 5687 7429
rect 5810 7420 5816 7432
rect 5868 7420 5874 7472
rect 7374 7460 7380 7472
rect 6564 7432 7380 7460
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 5166 7392 5172 7404
rect 4571 7364 5172 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 5166 7352 5172 7364
rect 5224 7392 5230 7404
rect 6564 7401 6592 7432
rect 7374 7420 7380 7432
rect 7432 7460 7438 7472
rect 9674 7460 9680 7472
rect 7432 7432 9680 7460
rect 7432 7420 7438 7432
rect 9674 7420 9680 7432
rect 9732 7420 9738 7472
rect 9950 7420 9956 7472
rect 10008 7460 10014 7472
rect 10520 7469 10548 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12161 7491 12219 7497
rect 14642 7488 14648 7540
rect 14700 7528 14706 7540
rect 14737 7531 14795 7537
rect 14737 7528 14749 7531
rect 14700 7500 14749 7528
rect 14700 7488 14706 7500
rect 14737 7497 14749 7500
rect 14783 7497 14795 7531
rect 14737 7491 14795 7497
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 17954 7528 17960 7540
rect 15252 7500 15608 7528
rect 17915 7500 17960 7528
rect 15252 7488 15258 7500
rect 10505 7463 10563 7469
rect 10008 7432 10456 7460
rect 10008 7420 10014 7432
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 5224 7364 6561 7392
rect 5224 7352 5230 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6696 7364 7021 7392
rect 6696 7352 6702 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7190 7392 7196 7404
rect 7151 7364 7196 7392
rect 7009 7355 7067 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 7561 7395 7619 7401
rect 7561 7392 7573 7395
rect 7524 7364 7573 7392
rect 7524 7352 7530 7364
rect 7561 7361 7573 7364
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 8481 7395 8539 7401
rect 8481 7392 8493 7395
rect 8444 7364 8493 7392
rect 8444 7352 8450 7364
rect 8481 7361 8493 7364
rect 8527 7361 8539 7395
rect 8662 7392 8668 7404
rect 8623 7364 8668 7392
rect 8481 7355 8539 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 9030 7392 9036 7404
rect 8991 7364 9036 7392
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10428 7392 10456 7432
rect 10505 7429 10517 7463
rect 10551 7429 10563 7463
rect 10505 7423 10563 7429
rect 11422 7420 11428 7472
rect 11480 7460 11486 7472
rect 11609 7463 11667 7469
rect 11609 7460 11621 7463
rect 11480 7432 11621 7460
rect 11480 7420 11486 7432
rect 11609 7429 11621 7432
rect 11655 7429 11667 7463
rect 15010 7460 15016 7472
rect 11609 7423 11667 7429
rect 14476 7432 15016 7460
rect 14476 7404 14504 7432
rect 15010 7420 15016 7432
rect 15068 7460 15074 7472
rect 15068 7432 15516 7460
rect 15068 7420 15074 7432
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 10428 7364 11529 7392
rect 10321 7355 10379 7361
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11698 7392 11704 7404
rect 11659 7364 11704 7392
rect 11517 7355 11575 7361
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7324 4307 7327
rect 4430 7324 4436 7336
rect 4295 7296 4436 7324
rect 4295 7293 4307 7296
rect 4249 7287 4307 7293
rect 4430 7284 4436 7296
rect 4488 7284 4494 7336
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 7285 7327 7343 7333
rect 7285 7324 7297 7327
rect 6880 7296 7297 7324
rect 6880 7284 6886 7296
rect 7285 7293 7297 7296
rect 7331 7293 7343 7327
rect 7285 7287 7343 7293
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 8757 7327 8815 7333
rect 7423 7296 8524 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 3510 7256 3516 7268
rect 1627 7228 3516 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 3510 7216 3516 7228
rect 3568 7216 3574 7268
rect 7300 7256 7328 7287
rect 8496 7268 8524 7296
rect 8757 7293 8769 7327
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 8849 7327 8907 7333
rect 8849 7293 8861 7327
rect 8895 7324 8907 7327
rect 9306 7324 9312 7336
rect 8895 7296 9312 7324
rect 8895 7293 8907 7296
rect 8849 7287 8907 7293
rect 7650 7256 7656 7268
rect 7300 7228 7656 7256
rect 7650 7216 7656 7228
rect 7708 7216 7714 7268
rect 8478 7216 8484 7268
rect 8536 7216 8542 7268
rect 8772 7256 8800 7287
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 10336 7324 10364 7355
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7392 12587 7395
rect 12894 7392 12900 7404
rect 12575 7364 12900 7392
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7361 13231 7395
rect 13998 7392 14004 7404
rect 13959 7364 14004 7392
rect 13173 7355 13231 7361
rect 10594 7324 10600 7336
rect 10336 7296 10600 7324
rect 10594 7284 10600 7296
rect 10652 7284 10658 7336
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 12492 7296 12537 7324
rect 12492 7284 12498 7296
rect 9766 7256 9772 7268
rect 8772 7228 9772 7256
rect 9766 7216 9772 7228
rect 9824 7256 9830 7268
rect 9950 7256 9956 7268
rect 9824 7228 9956 7256
rect 9824 7216 9830 7228
rect 9950 7216 9956 7228
rect 10008 7216 10014 7268
rect 13188 7256 13216 7355
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 14182 7392 14188 7404
rect 14143 7364 14188 7392
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7392 14335 7395
rect 14458 7392 14464 7404
rect 14323 7364 14464 7392
rect 14323 7361 14335 7364
rect 14277 7355 14335 7361
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 14553 7395 14611 7401
rect 14553 7361 14565 7395
rect 14599 7361 14611 7395
rect 14553 7355 14611 7361
rect 13449 7327 13507 7333
rect 13449 7293 13461 7327
rect 13495 7324 13507 7327
rect 13538 7324 13544 7336
rect 13495 7296 13544 7324
rect 13495 7293 13507 7296
rect 13449 7287 13507 7293
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7293 14427 7327
rect 14568 7324 14596 7355
rect 14826 7352 14832 7404
rect 14884 7392 14890 7404
rect 15194 7392 15200 7404
rect 14884 7364 15200 7392
rect 14884 7352 14890 7364
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 15378 7392 15384 7404
rect 15339 7364 15384 7392
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 15488 7401 15516 7432
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15286 7324 15292 7336
rect 14568 7296 15292 7324
rect 14369 7287 14427 7293
rect 12544 7228 13216 7256
rect 14384 7256 14412 7287
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 15580 7333 15608 7500
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 18598 7488 18604 7540
rect 18656 7528 18662 7540
rect 23201 7531 23259 7537
rect 23201 7528 23213 7531
rect 18656 7500 23213 7528
rect 18656 7488 18662 7500
rect 17310 7460 17316 7472
rect 17271 7432 17316 7460
rect 17310 7420 17316 7432
rect 17368 7420 17374 7472
rect 18046 7420 18052 7472
rect 18104 7460 18110 7472
rect 19981 7463 20039 7469
rect 19981 7460 19993 7463
rect 18104 7432 19993 7460
rect 18104 7420 18110 7432
rect 19981 7429 19993 7432
rect 20027 7429 20039 7463
rect 19981 7423 20039 7429
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7392 15807 7395
rect 16942 7392 16948 7404
rect 15795 7364 16948 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 18230 7352 18236 7404
rect 18288 7392 18294 7404
rect 19070 7395 19128 7401
rect 19070 7392 19082 7395
rect 18288 7364 19082 7392
rect 18288 7352 18294 7364
rect 19070 7361 19082 7364
rect 19116 7361 19128 7395
rect 19070 7355 19128 7361
rect 20346 7352 20352 7404
rect 20404 7392 20410 7404
rect 20533 7395 20591 7401
rect 20533 7392 20545 7395
rect 20404 7364 20545 7392
rect 20404 7352 20410 7364
rect 20533 7361 20545 7364
rect 20579 7361 20591 7395
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 20533 7355 20591 7361
rect 20640 7364 20729 7392
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7324 15623 7327
rect 19337 7327 19395 7333
rect 15611 7296 16896 7324
rect 15611 7293 15623 7296
rect 15565 7287 15623 7293
rect 15102 7256 15108 7268
rect 14384 7228 15108 7256
rect 12544 7200 12572 7228
rect 15102 7216 15108 7228
rect 15160 7216 15166 7268
rect 16868 7200 16896 7296
rect 19337 7293 19349 7327
rect 19383 7324 19395 7327
rect 19702 7324 19708 7336
rect 19383 7296 19708 7324
rect 19383 7293 19395 7296
rect 19337 7287 19395 7293
rect 19702 7284 19708 7296
rect 19760 7284 19766 7336
rect 17494 7256 17500 7268
rect 17455 7228 17500 7256
rect 17494 7216 17500 7228
rect 17552 7216 17558 7268
rect 20640 7256 20668 7364
rect 20717 7361 20729 7364
rect 20763 7361 20775 7395
rect 20898 7392 20904 7404
rect 20859 7364 20904 7392
rect 20717 7355 20775 7361
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 21100 7401 21128 7500
rect 23201 7497 23213 7500
rect 23247 7497 23259 7531
rect 23201 7491 23259 7497
rect 21269 7463 21327 7469
rect 21269 7429 21281 7463
rect 21315 7460 21327 7463
rect 22066 7463 22124 7469
rect 22066 7460 22078 7463
rect 21315 7432 22078 7460
rect 21315 7429 21327 7432
rect 21269 7423 21327 7429
rect 22066 7429 22078 7432
rect 22112 7429 22124 7463
rect 22066 7423 22124 7429
rect 21085 7395 21143 7401
rect 21085 7361 21097 7395
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 21634 7352 21640 7404
rect 21692 7392 21698 7404
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 21692 7364 21833 7392
rect 21692 7352 21698 7364
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 29546 7352 29552 7404
rect 29604 7392 29610 7404
rect 29825 7395 29883 7401
rect 29825 7392 29837 7395
rect 29604 7364 29837 7392
rect 29604 7352 29610 7364
rect 29825 7361 29837 7364
rect 29871 7361 29883 7395
rect 29825 7355 29883 7361
rect 20806 7324 20812 7336
rect 20767 7296 20812 7324
rect 20806 7284 20812 7296
rect 20864 7284 20870 7336
rect 20640 7228 21864 7256
rect 7742 7188 7748 7200
rect 7703 7160 7748 7188
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 9214 7188 9220 7200
rect 9175 7160 9220 7188
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 12526 7188 12532 7200
rect 12487 7160 12532 7188
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12986 7188 12992 7200
rect 12947 7160 12992 7188
rect 12986 7148 12992 7160
rect 13044 7148 13050 7200
rect 13357 7191 13415 7197
rect 13357 7157 13369 7191
rect 13403 7188 13415 7191
rect 13630 7188 13636 7200
rect 13403 7160 13636 7188
rect 13403 7157 13415 7160
rect 13357 7151 13415 7157
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 15933 7191 15991 7197
rect 15933 7188 15945 7191
rect 15804 7160 15945 7188
rect 15804 7148 15810 7160
rect 15933 7157 15945 7160
rect 15979 7157 15991 7191
rect 15933 7151 15991 7157
rect 16850 7148 16856 7200
rect 16908 7188 16914 7200
rect 17586 7188 17592 7200
rect 16908 7160 17592 7188
rect 16908 7148 16914 7160
rect 17586 7148 17592 7160
rect 17644 7188 17650 7200
rect 19889 7191 19947 7197
rect 19889 7188 19901 7191
rect 17644 7160 19901 7188
rect 17644 7148 17650 7160
rect 19889 7157 19901 7160
rect 19935 7157 19947 7191
rect 19889 7151 19947 7157
rect 20806 7148 20812 7200
rect 20864 7188 20870 7200
rect 21266 7188 21272 7200
rect 20864 7160 21272 7188
rect 20864 7148 20870 7160
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 21836 7188 21864 7228
rect 22094 7188 22100 7200
rect 21836 7160 22100 7188
rect 22094 7148 22100 7160
rect 22152 7148 22158 7200
rect 30006 7188 30012 7200
rect 29967 7160 30012 7188
rect 30006 7148 30012 7160
rect 30064 7148 30070 7200
rect 1104 7098 30820 7120
rect 1104 7046 5915 7098
rect 5967 7046 5979 7098
rect 6031 7046 6043 7098
rect 6095 7046 6107 7098
rect 6159 7046 6171 7098
rect 6223 7046 15846 7098
rect 15898 7046 15910 7098
rect 15962 7046 15974 7098
rect 16026 7046 16038 7098
rect 16090 7046 16102 7098
rect 16154 7046 25776 7098
rect 25828 7046 25840 7098
rect 25892 7046 25904 7098
rect 25956 7046 25968 7098
rect 26020 7046 26032 7098
rect 26084 7046 30820 7098
rect 1104 7024 30820 7046
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 6549 6987 6607 6993
rect 6549 6984 6561 6987
rect 6420 6956 6561 6984
rect 6420 6944 6426 6956
rect 6549 6953 6561 6956
rect 6595 6953 6607 6987
rect 6549 6947 6607 6953
rect 7009 6987 7067 6993
rect 7009 6953 7021 6987
rect 7055 6984 7067 6987
rect 7466 6984 7472 6996
rect 7055 6956 7472 6984
rect 7055 6953 7067 6956
rect 7009 6947 7067 6953
rect 5258 6916 5264 6928
rect 3988 6888 5264 6916
rect 1762 6848 1768 6860
rect 1723 6820 1768 6848
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1412 6644 1440 6743
rect 1486 6740 1492 6792
rect 1544 6780 1550 6792
rect 1581 6783 1639 6789
rect 1581 6780 1593 6783
rect 1544 6752 1593 6780
rect 1544 6740 1550 6752
rect 1581 6749 1593 6752
rect 1627 6749 1639 6783
rect 1581 6743 1639 6749
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1854 6780 1860 6792
rect 1719 6752 1860 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 1854 6740 1860 6752
rect 1912 6740 1918 6792
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 2774 6780 2780 6792
rect 2639 6752 2780 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 1964 6712 1992 6743
rect 2774 6740 2780 6752
rect 2832 6740 2838 6792
rect 3988 6789 4016 6888
rect 5258 6876 5264 6888
rect 5316 6876 5322 6928
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 6730 6848 6736 6860
rect 5500 6820 6736 6848
rect 5500 6808 5506 6820
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 4120 6752 4169 6780
rect 4120 6740 4126 6752
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 2866 6712 2872 6724
rect 1964 6684 2872 6712
rect 2866 6672 2872 6684
rect 2924 6672 2930 6724
rect 4264 6712 4292 6743
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 4525 6783 4583 6789
rect 4396 6752 4441 6780
rect 4396 6740 4402 6752
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 4571 6752 5304 6780
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 5166 6712 5172 6724
rect 4264 6684 4384 6712
rect 5127 6684 5172 6712
rect 4356 6656 4384 6684
rect 5166 6672 5172 6684
rect 5224 6672 5230 6724
rect 1578 6644 1584 6656
rect 1412 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6644 1642 6656
rect 1946 6644 1952 6656
rect 1636 6616 1952 6644
rect 1636 6604 1642 6616
rect 1946 6604 1952 6616
rect 2004 6604 2010 6656
rect 2130 6644 2136 6656
rect 2091 6616 2136 6644
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 2777 6647 2835 6653
rect 2777 6613 2789 6647
rect 2823 6644 2835 6647
rect 3694 6644 3700 6656
rect 2823 6616 3700 6644
rect 2823 6613 2835 6616
rect 2777 6607 2835 6613
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 3789 6647 3847 6653
rect 3789 6613 3801 6647
rect 3835 6644 3847 6647
rect 3878 6644 3884 6656
rect 3835 6616 3884 6644
rect 3835 6613 3847 6616
rect 3789 6607 3847 6613
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 4338 6604 4344 6656
rect 4396 6604 4402 6656
rect 5074 6644 5080 6656
rect 5035 6616 5080 6644
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 5276 6644 5304 6752
rect 5350 6740 5356 6792
rect 5408 6780 5414 6792
rect 5626 6780 5632 6792
rect 5408 6752 5632 6780
rect 5408 6740 5414 6752
rect 5626 6740 5632 6752
rect 5684 6780 5690 6792
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 5684 6752 5733 6780
rect 5684 6740 5690 6752
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 5810 6740 5816 6792
rect 5868 6780 5874 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5868 6752 6009 6780
rect 5868 6740 5874 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 6914 6780 6920 6792
rect 6595 6752 6920 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 5442 6672 5448 6724
rect 5500 6712 5506 6724
rect 5902 6712 5908 6724
rect 5500 6684 5908 6712
rect 5500 6672 5506 6684
rect 5902 6672 5908 6684
rect 5960 6672 5966 6724
rect 6380 6712 6408 6743
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7024 6712 7052 6947
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 11701 6987 11759 6993
rect 7708 6956 8432 6984
rect 7708 6944 7714 6956
rect 8404 6916 8432 6956
rect 11701 6953 11713 6987
rect 11747 6984 11759 6987
rect 11882 6984 11888 6996
rect 11747 6956 11888 6984
rect 11747 6953 11759 6956
rect 11701 6947 11759 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 18414 6984 18420 6996
rect 12406 6956 18420 6984
rect 12406 6916 12434 6956
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 12802 6916 12808 6928
rect 8404 6888 12434 6916
rect 12763 6888 12808 6916
rect 12802 6876 12808 6888
rect 12860 6876 12866 6928
rect 13998 6876 14004 6928
rect 14056 6916 14062 6928
rect 18049 6919 18107 6925
rect 18049 6916 18061 6919
rect 14056 6888 18061 6916
rect 14056 6876 14062 6888
rect 18049 6885 18061 6888
rect 18095 6916 18107 6919
rect 18782 6916 18788 6928
rect 18095 6888 18788 6916
rect 18095 6885 18107 6888
rect 18049 6879 18107 6885
rect 18782 6876 18788 6888
rect 18840 6876 18846 6928
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 12069 6851 12127 6857
rect 9732 6820 11008 6848
rect 9732 6808 9738 6820
rect 7742 6740 7748 6792
rect 7800 6780 7806 6792
rect 8122 6783 8180 6789
rect 8122 6780 8134 6783
rect 7800 6752 8134 6780
rect 7800 6740 7806 6752
rect 8122 6749 8134 6752
rect 8168 6749 8180 6783
rect 8122 6743 8180 6749
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 8352 6752 8401 6780
rect 8352 6740 8358 6752
rect 8389 6749 8401 6752
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 9950 6740 9956 6792
rect 10008 6780 10014 6792
rect 10980 6789 11008 6820
rect 12069 6817 12081 6851
rect 12115 6848 12127 6851
rect 13449 6851 13507 6857
rect 12115 6820 13308 6848
rect 12115 6817 12127 6820
rect 12069 6811 12127 6817
rect 10045 6783 10103 6789
rect 10045 6780 10057 6783
rect 10008 6752 10057 6780
rect 10008 6740 10014 6752
rect 10045 6749 10057 6752
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6780 10379 6783
rect 10965 6783 11023 6789
rect 10367 6752 10916 6780
rect 10367 6749 10379 6752
rect 10321 6743 10379 6749
rect 6380 6684 7052 6712
rect 6270 6644 6276 6656
rect 5276 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 6362 6604 6368 6656
rect 6420 6644 6426 6656
rect 6638 6644 6644 6656
rect 6420 6616 6644 6644
rect 6420 6604 6426 6616
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 10888 6653 10916 6752
rect 10965 6749 10977 6783
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11422 6740 11428 6792
rect 11480 6780 11486 6792
rect 11790 6780 11796 6792
rect 11480 6752 11796 6780
rect 11480 6740 11486 6752
rect 11790 6740 11796 6752
rect 11848 6780 11854 6792
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 11848 6752 11897 6780
rect 11848 6740 11854 6752
rect 11885 6749 11897 6752
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6780 12219 6783
rect 12710 6780 12716 6792
rect 12207 6752 12716 6780
rect 12207 6749 12219 6752
rect 12161 6743 12219 6749
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 12986 6740 12992 6792
rect 13044 6780 13050 6792
rect 13173 6783 13231 6789
rect 13173 6780 13185 6783
rect 13044 6752 13185 6780
rect 13044 6740 13050 6752
rect 13173 6749 13185 6752
rect 13219 6749 13231 6783
rect 13280 6780 13308 6820
rect 13449 6817 13461 6851
rect 13495 6848 13507 6851
rect 13722 6848 13728 6860
rect 13495 6820 13728 6848
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 15010 6848 15016 6860
rect 14971 6820 15016 6848
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15562 6848 15568 6860
rect 15252 6820 15568 6848
rect 15252 6808 15258 6820
rect 15562 6808 15568 6820
rect 15620 6848 15626 6860
rect 16850 6848 16856 6860
rect 15620 6820 16528 6848
rect 16811 6820 16856 6848
rect 15620 6808 15626 6820
rect 13630 6780 13636 6792
rect 13280 6752 13636 6780
rect 13173 6743 13231 6749
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 15286 6780 15292 6792
rect 14476 6752 15292 6780
rect 12526 6672 12532 6724
rect 12584 6712 12590 6724
rect 13265 6715 13323 6721
rect 13265 6712 13277 6715
rect 12584 6684 13277 6712
rect 12584 6672 12590 6684
rect 13265 6681 13277 6684
rect 13311 6681 13323 6715
rect 13265 6675 13323 6681
rect 10873 6647 10931 6653
rect 10873 6613 10885 6647
rect 10919 6644 10931 6647
rect 14476 6644 14504 6752
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 16500 6789 16528 6820
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 16942 6808 16948 6860
rect 17000 6848 17006 6860
rect 19518 6848 19524 6860
rect 17000 6820 17448 6848
rect 19479 6820 19524 6848
rect 17000 6808 17006 6820
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6749 15991 6783
rect 15933 6743 15991 6749
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6749 16543 6783
rect 16666 6780 16672 6792
rect 16627 6752 16672 6780
rect 16485 6743 16543 6749
rect 14826 6672 14832 6724
rect 14884 6712 14890 6724
rect 15948 6712 15976 6743
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 16770 6783 16828 6789
rect 16770 6749 16782 6783
rect 16816 6780 16828 6783
rect 16816 6752 16988 6780
rect 16816 6749 16828 6752
rect 16770 6743 16828 6749
rect 14884 6684 15976 6712
rect 16960 6712 16988 6752
rect 17034 6740 17040 6792
rect 17092 6780 17098 6792
rect 17218 6780 17224 6792
rect 17092 6752 17224 6780
rect 17092 6740 17098 6752
rect 17218 6740 17224 6752
rect 17276 6740 17282 6792
rect 17420 6780 17448 6820
rect 19518 6808 19524 6820
rect 19576 6808 19582 6860
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 17420 6752 19441 6780
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 20073 6783 20131 6789
rect 20073 6749 20085 6783
rect 20119 6780 20131 6783
rect 21266 6780 21272 6792
rect 20119 6752 21272 6780
rect 20119 6749 20131 6752
rect 20073 6743 20131 6749
rect 21266 6740 21272 6752
rect 21324 6780 21330 6792
rect 21634 6780 21640 6792
rect 21324 6752 21640 6780
rect 21324 6740 21330 6752
rect 21634 6740 21640 6752
rect 21692 6740 21698 6792
rect 17770 6712 17776 6724
rect 16960 6684 17776 6712
rect 14884 6672 14890 6684
rect 17770 6672 17776 6684
rect 17828 6672 17834 6724
rect 17865 6715 17923 6721
rect 17865 6681 17877 6715
rect 17911 6712 17923 6715
rect 18046 6712 18052 6724
rect 17911 6684 18052 6712
rect 17911 6681 17923 6684
rect 17865 6675 17923 6681
rect 18046 6672 18052 6684
rect 18104 6672 18110 6724
rect 20340 6715 20398 6721
rect 20340 6681 20352 6715
rect 20386 6712 20398 6715
rect 20714 6712 20720 6724
rect 20386 6684 20720 6712
rect 20386 6681 20398 6684
rect 20340 6675 20398 6681
rect 20714 6672 20720 6684
rect 20772 6672 20778 6724
rect 10919 6616 14504 6644
rect 10919 6613 10931 6616
rect 10873 6607 10931 6613
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 15749 6647 15807 6653
rect 15749 6644 15761 6647
rect 14608 6616 15761 6644
rect 14608 6604 14614 6616
rect 15749 6613 15761 6616
rect 15795 6613 15807 6647
rect 17218 6644 17224 6656
rect 17179 6616 17224 6644
rect 15749 6607 15807 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 21450 6644 21456 6656
rect 21411 6616 21456 6644
rect 21450 6604 21456 6616
rect 21508 6604 21514 6656
rect 1104 6554 30820 6576
rect 1104 6502 10880 6554
rect 10932 6502 10944 6554
rect 10996 6502 11008 6554
rect 11060 6502 11072 6554
rect 11124 6502 11136 6554
rect 11188 6502 20811 6554
rect 20863 6502 20875 6554
rect 20927 6502 20939 6554
rect 20991 6502 21003 6554
rect 21055 6502 21067 6554
rect 21119 6502 30820 6554
rect 1104 6480 30820 6502
rect 1670 6400 1676 6452
rect 1728 6400 1734 6452
rect 2866 6440 2872 6452
rect 2779 6412 2872 6440
rect 2866 6400 2872 6412
rect 2924 6440 2930 6452
rect 7006 6440 7012 6452
rect 2924 6412 7012 6440
rect 2924 6400 2930 6412
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 8941 6443 8999 6449
rect 8941 6409 8953 6443
rect 8987 6440 8999 6443
rect 9030 6440 9036 6452
rect 8987 6412 9036 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 9030 6400 9036 6412
rect 9088 6440 9094 6452
rect 9677 6443 9735 6449
rect 9677 6440 9689 6443
rect 9088 6412 9689 6440
rect 9088 6400 9094 6412
rect 9677 6409 9689 6412
rect 9723 6409 9735 6443
rect 30098 6440 30104 6452
rect 9677 6403 9735 6409
rect 10336 6412 30104 6440
rect 1489 6307 1547 6313
rect 1489 6273 1501 6307
rect 1535 6304 1547 6307
rect 1688 6304 1716 6400
rect 1756 6375 1814 6381
rect 1756 6341 1768 6375
rect 1802 6372 1814 6375
rect 2130 6372 2136 6384
rect 1802 6344 2136 6372
rect 1802 6341 1814 6344
rect 1756 6335 1814 6341
rect 2130 6332 2136 6344
rect 2188 6332 2194 6384
rect 3694 6332 3700 6384
rect 3752 6372 3758 6384
rect 8294 6372 8300 6384
rect 3752 6344 6500 6372
rect 3752 6332 3758 6344
rect 1535 6276 1716 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 2038 6264 2044 6316
rect 2096 6304 2102 6316
rect 3329 6307 3387 6313
rect 3329 6304 3341 6307
rect 2096 6276 3341 6304
rect 2096 6264 2102 6276
rect 3329 6273 3341 6276
rect 3375 6273 3387 6307
rect 3510 6304 3516 6316
rect 3471 6276 3516 6304
rect 3329 6267 3387 6273
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 3786 6264 3792 6316
rect 3844 6304 3850 6316
rect 3881 6307 3939 6313
rect 3881 6304 3893 6307
rect 3844 6276 3893 6304
rect 3844 6264 3850 6276
rect 3881 6273 3893 6276
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6273 5135 6307
rect 5258 6304 5264 6316
rect 5219 6276 5264 6304
rect 5077 6267 5135 6273
rect 3605 6239 3663 6245
rect 3605 6236 3617 6239
rect 2746 6208 3617 6236
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 2746 6100 2774 6208
rect 3605 6205 3617 6208
rect 3651 6205 3663 6239
rect 3605 6199 3663 6205
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6236 3755 6239
rect 4062 6236 4068 6248
rect 3743 6208 4068 6236
rect 3743 6205 3755 6208
rect 3697 6199 3755 6205
rect 3620 6168 3648 6199
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 5092 6236 5120 6267
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 5626 6304 5632 6316
rect 5587 6276 5632 6304
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 6086 6304 6092 6316
rect 5859 6276 6092 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6328 6276 6377 6304
rect 6328 6264 6334 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6472 6304 6500 6344
rect 7576 6344 8300 6372
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6472 6276 6561 6304
rect 6365 6267 6423 6273
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6730 6304 6736 6316
rect 6691 6276 6736 6304
rect 6549 6267 6607 6273
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 7576 6313 7604 6344
rect 8294 6332 8300 6344
rect 8352 6332 8358 6384
rect 10336 6372 10364 6412
rect 30098 6400 30104 6412
rect 30156 6400 30162 6452
rect 9508 6344 10364 6372
rect 10413 6375 10471 6381
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 7828 6307 7886 6313
rect 7828 6273 7840 6307
rect 7874 6304 7886 6307
rect 9214 6304 9220 6316
rect 7874 6276 9220 6304
rect 7874 6273 7886 6276
rect 7828 6267 7886 6273
rect 5350 6236 5356 6248
rect 5092 6208 5356 6236
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 5460 6208 6653 6236
rect 4338 6168 4344 6180
rect 3620 6140 4344 6168
rect 4338 6128 4344 6140
rect 4396 6128 4402 6180
rect 5074 6128 5080 6180
rect 5132 6168 5138 6180
rect 5460 6168 5488 6208
rect 6641 6205 6653 6208
rect 6687 6205 6699 6239
rect 6641 6199 6699 6205
rect 5132 6140 5488 6168
rect 5629 6171 5687 6177
rect 5132 6128 5138 6140
rect 5629 6137 5641 6171
rect 5675 6168 5687 6171
rect 5718 6168 5724 6180
rect 5675 6140 5724 6168
rect 5675 6137 5687 6140
rect 5629 6131 5687 6137
rect 5718 6128 5724 6140
rect 5776 6128 5782 6180
rect 5902 6128 5908 6180
rect 5960 6168 5966 6180
rect 6932 6168 6960 6267
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 9508 6177 9536 6344
rect 10413 6341 10425 6375
rect 10459 6372 10471 6375
rect 10594 6372 10600 6384
rect 10459 6344 10600 6372
rect 10459 6341 10471 6344
rect 10413 6335 10471 6341
rect 10594 6332 10600 6344
rect 10652 6332 10658 6384
rect 10778 6372 10784 6384
rect 10739 6344 10784 6372
rect 10778 6332 10784 6344
rect 10836 6332 10842 6384
rect 10962 6332 10968 6384
rect 11020 6372 11026 6384
rect 12618 6372 12624 6384
rect 11020 6344 12624 6372
rect 11020 6332 11026 6344
rect 12618 6332 12624 6344
rect 12676 6332 12682 6384
rect 12802 6332 12808 6384
rect 12860 6372 12866 6384
rect 13538 6372 13544 6384
rect 12860 6344 13544 6372
rect 12860 6332 12866 6344
rect 13538 6332 13544 6344
rect 13596 6372 13602 6384
rect 16482 6372 16488 6384
rect 13596 6344 13768 6372
rect 13596 6332 13602 6344
rect 10042 6304 10048 6316
rect 10003 6276 10048 6304
rect 10042 6264 10048 6276
rect 10100 6264 10106 6316
rect 10502 6304 10508 6316
rect 10463 6276 10508 6304
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 13740 6313 13768 6344
rect 14292 6344 16488 6372
rect 14292 6313 14320 6344
rect 16482 6332 16488 6344
rect 16540 6372 16546 6384
rect 19702 6372 19708 6384
rect 16540 6344 19708 6372
rect 16540 6332 16546 6344
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 13265 6307 13323 6313
rect 13265 6304 13277 6307
rect 12483 6276 13277 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 13265 6273 13277 6276
rect 13311 6273 13323 6307
rect 13265 6267 13323 6273
rect 13449 6307 13507 6313
rect 13449 6273 13461 6307
rect 13495 6273 13507 6307
rect 13449 6267 13507 6273
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 14544 6307 14602 6313
rect 14544 6273 14556 6307
rect 14590 6304 14602 6307
rect 14918 6304 14924 6316
rect 14590 6276 14924 6304
rect 14590 6273 14602 6276
rect 14544 6267 14602 6273
rect 10968 6248 11020 6254
rect 11974 6196 11980 6248
rect 12032 6236 12038 6248
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 12032 6208 12173 6236
rect 12032 6196 12038 6208
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 12342 6236 12348 6248
rect 12255 6208 12348 6236
rect 12161 6199 12219 6205
rect 10968 6190 11020 6196
rect 5960 6140 6960 6168
rect 9493 6171 9551 6177
rect 5960 6128 5966 6140
rect 9493 6137 9505 6171
rect 9539 6137 9551 6171
rect 12176 6168 12204 6199
rect 12342 6196 12348 6208
rect 12400 6236 12406 6248
rect 12618 6236 12624 6248
rect 12400 6208 12624 6236
rect 12400 6196 12406 6208
rect 12618 6196 12624 6208
rect 12676 6236 12682 6248
rect 13464 6236 13492 6267
rect 14918 6264 14924 6276
rect 14976 6264 14982 6316
rect 17218 6264 17224 6316
rect 17276 6304 17282 6316
rect 18064 6313 18092 6344
rect 19702 6332 19708 6344
rect 19760 6332 19766 6384
rect 17782 6307 17840 6313
rect 17782 6304 17794 6307
rect 17276 6276 17794 6304
rect 17276 6264 17282 6276
rect 17782 6273 17794 6276
rect 17828 6273 17840 6307
rect 17782 6267 17840 6273
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6273 18107 6307
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 18049 6267 18107 6273
rect 18156 6276 18705 6304
rect 12676 6208 13492 6236
rect 12676 6196 12682 6208
rect 12434 6168 12440 6180
rect 12176 6140 12440 6168
rect 9493 6131 9551 6137
rect 12434 6128 12440 6140
rect 12492 6128 12498 6180
rect 12805 6171 12863 6177
rect 12805 6137 12817 6171
rect 12851 6168 12863 6171
rect 13078 6168 13084 6180
rect 12851 6140 13084 6168
rect 12851 6137 12863 6140
rect 12805 6131 12863 6137
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 15654 6168 15660 6180
rect 15615 6140 15660 6168
rect 15654 6128 15660 6140
rect 15712 6128 15718 6180
rect 16669 6171 16727 6177
rect 16669 6137 16681 6171
rect 16715 6168 16727 6171
rect 17034 6168 17040 6180
rect 16715 6140 17040 6168
rect 16715 6137 16727 6140
rect 16669 6131 16727 6137
rect 17034 6128 17040 6140
rect 17092 6128 17098 6180
rect 4062 6100 4068 6112
rect 1912 6072 2774 6100
rect 4023 6072 4068 6100
rect 1912 6060 1918 6072
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4430 6060 4436 6112
rect 4488 6100 4494 6112
rect 7101 6103 7159 6109
rect 7101 6100 7113 6103
rect 4488 6072 7113 6100
rect 4488 6060 4494 6072
rect 7101 6069 7113 6072
rect 7147 6069 7159 6103
rect 13630 6100 13636 6112
rect 13591 6072 13636 6100
rect 7101 6063 7159 6069
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 15286 6060 15292 6112
rect 15344 6100 15350 6112
rect 18156 6100 18184 6276
rect 18693 6273 18705 6276
rect 18739 6304 18751 6307
rect 19426 6304 19432 6316
rect 18739 6276 19432 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 19426 6264 19432 6276
rect 19484 6304 19490 6316
rect 19613 6307 19671 6313
rect 19613 6304 19625 6307
rect 19484 6276 19625 6304
rect 19484 6264 19490 6276
rect 19613 6273 19625 6276
rect 19659 6273 19671 6307
rect 19613 6267 19671 6273
rect 19889 6307 19947 6313
rect 19889 6273 19901 6307
rect 19935 6304 19947 6307
rect 20254 6304 20260 6316
rect 19935 6276 20260 6304
rect 19935 6273 19947 6276
rect 19889 6267 19947 6273
rect 20254 6264 20260 6276
rect 20312 6304 20318 6316
rect 20622 6304 20628 6316
rect 20312 6276 20628 6304
rect 20312 6264 20318 6276
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 18414 6196 18420 6248
rect 18472 6236 18478 6248
rect 18509 6239 18567 6245
rect 18509 6236 18521 6239
rect 18472 6208 18521 6236
rect 18472 6196 18478 6208
rect 18509 6205 18521 6208
rect 18555 6205 18567 6239
rect 18509 6199 18567 6205
rect 15344 6072 18184 6100
rect 15344 6060 15350 6072
rect 1104 6010 30820 6032
rect 1104 5958 5915 6010
rect 5967 5958 5979 6010
rect 6031 5958 6043 6010
rect 6095 5958 6107 6010
rect 6159 5958 6171 6010
rect 6223 5958 15846 6010
rect 15898 5958 15910 6010
rect 15962 5958 15974 6010
rect 16026 5958 16038 6010
rect 16090 5958 16102 6010
rect 16154 5958 25776 6010
rect 25828 5958 25840 6010
rect 25892 5958 25904 6010
rect 25956 5958 25968 6010
rect 26020 5958 26032 6010
rect 26084 5958 30820 6010
rect 1104 5936 30820 5958
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 3786 5896 3792 5908
rect 3283 5868 3792 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 3786 5856 3792 5868
rect 3844 5896 3850 5908
rect 3844 5868 6316 5896
rect 3844 5856 3850 5868
rect 5537 5831 5595 5837
rect 5537 5797 5549 5831
rect 5583 5828 5595 5831
rect 5810 5828 5816 5840
rect 5583 5800 5816 5828
rect 5583 5797 5595 5800
rect 5537 5791 5595 5797
rect 5810 5788 5816 5800
rect 5868 5788 5874 5840
rect 1670 5720 1676 5772
rect 1728 5760 1734 5772
rect 1857 5763 1915 5769
rect 1857 5760 1869 5763
rect 1728 5732 1869 5760
rect 1728 5720 1734 5732
rect 1857 5729 1869 5732
rect 1903 5729 1915 5763
rect 4154 5760 4160 5772
rect 4115 5732 4160 5760
rect 1857 5723 1915 5729
rect 1872 5692 1900 5723
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 4172 5692 4200 5720
rect 4430 5701 4436 5704
rect 4424 5692 4436 5701
rect 1872 5664 4200 5692
rect 4391 5664 4436 5692
rect 4424 5655 4436 5664
rect 4430 5652 4436 5655
rect 4488 5652 4494 5704
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 5994 5692 6000 5704
rect 5408 5664 6000 5692
rect 5408 5652 5414 5664
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 6288 5701 6316 5868
rect 9306 5856 9312 5908
rect 9364 5896 9370 5908
rect 9401 5899 9459 5905
rect 9401 5896 9413 5899
rect 9364 5868 9413 5896
rect 9364 5856 9370 5868
rect 9401 5865 9413 5868
rect 9447 5865 9459 5899
rect 9401 5859 9459 5865
rect 10410 5856 10416 5908
rect 10468 5896 10474 5908
rect 10781 5899 10839 5905
rect 10781 5896 10793 5899
rect 10468 5868 10793 5896
rect 10468 5856 10474 5868
rect 10781 5865 10793 5868
rect 10827 5865 10839 5899
rect 13446 5896 13452 5908
rect 13407 5868 13452 5896
rect 10781 5859 10839 5865
rect 13446 5856 13452 5868
rect 13504 5856 13510 5908
rect 16942 5896 16948 5908
rect 15580 5868 16804 5896
rect 16903 5868 16948 5896
rect 6454 5828 6460 5840
rect 6415 5800 6460 5828
rect 6454 5788 6460 5800
rect 6512 5788 6518 5840
rect 8478 5788 8484 5840
rect 8536 5828 8542 5840
rect 15580 5828 15608 5868
rect 8536 5800 15608 5828
rect 16776 5828 16804 5868
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 18046 5896 18052 5908
rect 17696 5868 18052 5896
rect 17696 5828 17724 5868
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 18230 5896 18236 5908
rect 18191 5868 18236 5896
rect 18230 5856 18236 5868
rect 18288 5856 18294 5908
rect 20714 5896 20720 5908
rect 20675 5868 20720 5896
rect 20714 5856 20720 5868
rect 20772 5856 20778 5908
rect 16776 5800 17724 5828
rect 8536 5788 8542 5800
rect 6914 5760 6920 5772
rect 6840 5732 6920 5760
rect 6840 5701 6868 5732
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 9508 5701 9536 5800
rect 17770 5788 17776 5840
rect 17828 5828 17834 5840
rect 19245 5831 19303 5837
rect 19245 5828 19257 5831
rect 17828 5800 19257 5828
rect 17828 5788 17834 5800
rect 19245 5797 19257 5800
rect 19291 5828 19303 5831
rect 19978 5828 19984 5840
rect 19291 5800 19984 5828
rect 19291 5797 19303 5800
rect 19245 5791 19303 5797
rect 19978 5788 19984 5800
rect 20036 5788 20042 5840
rect 11425 5763 11483 5769
rect 11425 5729 11437 5763
rect 11471 5760 11483 5763
rect 12434 5760 12440 5772
rect 11471 5732 12440 5760
rect 11471 5729 11483 5732
rect 11425 5723 11483 5729
rect 12434 5720 12440 5732
rect 12492 5760 12498 5772
rect 12805 5763 12863 5769
rect 12805 5760 12817 5763
rect 12492 5732 12817 5760
rect 12492 5720 12498 5732
rect 12805 5729 12817 5732
rect 12851 5729 12863 5763
rect 12805 5723 12863 5729
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5661 9551 5695
rect 9493 5655 9551 5661
rect 2124 5627 2182 5633
rect 2124 5593 2136 5627
rect 2170 5624 2182 5627
rect 4062 5624 4068 5636
rect 2170 5596 4068 5624
rect 2170 5593 2182 5596
rect 2124 5587 2182 5593
rect 4062 5584 4068 5596
rect 4120 5584 4126 5636
rect 6656 5624 6684 5655
rect 11238 5652 11244 5704
rect 11296 5692 11302 5704
rect 11790 5692 11796 5704
rect 11296 5664 11796 5692
rect 11296 5652 11302 5664
rect 11790 5652 11796 5664
rect 11848 5692 11854 5704
rect 11977 5695 12035 5701
rect 11977 5692 11989 5695
rect 11848 5664 11989 5692
rect 11848 5652 11854 5664
rect 11977 5661 11989 5664
rect 12023 5661 12035 5695
rect 12820 5692 12848 5723
rect 12894 5720 12900 5772
rect 12952 5760 12958 5772
rect 12989 5763 13047 5769
rect 12989 5760 13001 5763
rect 12952 5732 13001 5760
rect 12952 5720 12958 5732
rect 12989 5729 13001 5732
rect 13035 5729 13047 5763
rect 12989 5723 13047 5729
rect 13630 5720 13636 5772
rect 13688 5760 13694 5772
rect 14369 5763 14427 5769
rect 14369 5760 14381 5763
rect 13688 5732 14381 5760
rect 13688 5720 13694 5732
rect 14369 5729 14381 5732
rect 14415 5729 14427 5763
rect 14369 5723 14427 5729
rect 17586 5720 17592 5772
rect 17644 5760 17650 5772
rect 17865 5763 17923 5769
rect 17865 5760 17877 5763
rect 17644 5732 17877 5760
rect 17644 5720 17650 5732
rect 17865 5729 17877 5732
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 17954 5720 17960 5772
rect 18012 5720 18018 5772
rect 20254 5760 20260 5772
rect 20215 5732 20260 5760
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 20349 5763 20407 5769
rect 20349 5729 20361 5763
rect 20395 5760 20407 5763
rect 20438 5760 20444 5772
rect 20395 5732 20444 5760
rect 20395 5729 20407 5732
rect 20349 5723 20407 5729
rect 20438 5720 20444 5732
rect 20496 5720 20502 5772
rect 13538 5692 13544 5704
rect 12820 5664 13544 5692
rect 11977 5655 12035 5661
rect 13538 5652 13544 5664
rect 13596 5692 13602 5704
rect 13722 5692 13728 5704
rect 13596 5664 13728 5692
rect 13596 5652 13602 5664
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 14090 5692 14096 5704
rect 14051 5664 14096 5692
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 15565 5695 15623 5701
rect 15565 5661 15577 5695
rect 15611 5692 15623 5695
rect 16390 5692 16396 5704
rect 15611 5664 16396 5692
rect 15611 5661 15623 5664
rect 15565 5655 15623 5661
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5661 17739 5695
rect 17681 5655 17739 5661
rect 6914 5624 6920 5636
rect 6656 5596 6920 5624
rect 6914 5584 6920 5596
rect 6972 5584 6978 5636
rect 11149 5627 11207 5633
rect 11149 5593 11161 5627
rect 11195 5624 11207 5627
rect 11514 5624 11520 5636
rect 11195 5596 11520 5624
rect 11195 5593 11207 5596
rect 11149 5587 11207 5593
rect 11514 5584 11520 5596
rect 11572 5584 11578 5636
rect 12069 5627 12127 5633
rect 12069 5593 12081 5627
rect 12115 5624 12127 5627
rect 13354 5624 13360 5636
rect 12115 5596 13360 5624
rect 12115 5593 12127 5596
rect 12069 5587 12127 5593
rect 13354 5584 13360 5596
rect 13412 5584 13418 5636
rect 15746 5584 15752 5636
rect 15804 5633 15810 5636
rect 15804 5627 15868 5633
rect 15804 5593 15822 5627
rect 15856 5593 15868 5627
rect 17696 5624 17724 5655
rect 17770 5652 17776 5704
rect 17828 5692 17834 5704
rect 17972 5692 18000 5720
rect 18049 5695 18107 5701
rect 18049 5692 18061 5695
rect 17828 5664 17873 5692
rect 17972 5664 18061 5692
rect 17828 5652 17834 5664
rect 18049 5661 18061 5664
rect 18095 5661 18107 5695
rect 19426 5692 19432 5704
rect 19387 5664 19432 5692
rect 18049 5655 18107 5661
rect 19426 5652 19432 5664
rect 19484 5652 19490 5704
rect 19794 5652 19800 5704
rect 19852 5692 19858 5704
rect 19981 5695 20039 5701
rect 19981 5692 19993 5695
rect 19852 5664 19993 5692
rect 19852 5652 19858 5664
rect 19981 5661 19993 5664
rect 20027 5661 20039 5695
rect 19981 5655 20039 5661
rect 20165 5695 20223 5701
rect 20165 5661 20177 5695
rect 20211 5661 20223 5695
rect 20165 5655 20223 5661
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5692 20591 5695
rect 21450 5692 21456 5704
rect 20579 5664 21456 5692
rect 20579 5661 20591 5664
rect 20533 5655 20591 5661
rect 17954 5624 17960 5636
rect 17696 5596 17960 5624
rect 15804 5587 15868 5593
rect 15804 5584 15810 5587
rect 17954 5584 17960 5596
rect 18012 5584 18018 5636
rect 20180 5624 20208 5655
rect 21450 5652 21456 5664
rect 21508 5652 21514 5704
rect 20438 5624 20444 5636
rect 20180 5596 20444 5624
rect 20438 5584 20444 5596
rect 20496 5584 20502 5636
rect 2498 5516 2504 5568
rect 2556 5556 2562 5568
rect 9122 5556 9128 5568
rect 2556 5528 9128 5556
rect 2556 5516 2562 5528
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 11238 5556 11244 5568
rect 11199 5528 11244 5556
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 13078 5516 13084 5568
rect 13136 5556 13142 5568
rect 13136 5528 13181 5556
rect 13136 5516 13142 5528
rect 1104 5466 30820 5488
rect 1104 5414 10880 5466
rect 10932 5414 10944 5466
rect 10996 5414 11008 5466
rect 11060 5414 11072 5466
rect 11124 5414 11136 5466
rect 11188 5414 20811 5466
rect 20863 5414 20875 5466
rect 20927 5414 20939 5466
rect 20991 5414 21003 5466
rect 21055 5414 21067 5466
rect 21119 5414 30820 5466
rect 1104 5392 30820 5414
rect 4985 5355 5043 5361
rect 2746 5324 4292 5352
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 2746 5216 2774 5324
rect 4154 5284 4160 5296
rect 3620 5256 4160 5284
rect 3620 5225 3648 5256
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 4264 5284 4292 5324
rect 4985 5321 4997 5355
rect 5031 5352 5043 5355
rect 5258 5352 5264 5364
rect 5031 5324 5264 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 6362 5352 6368 5364
rect 5368 5324 6368 5352
rect 5368 5284 5396 5324
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 7006 5352 7012 5364
rect 6932 5324 7012 5352
rect 6822 5284 6828 5296
rect 4264 5256 5396 5284
rect 6380 5256 6828 5284
rect 3878 5225 3884 5228
rect 1719 5188 2774 5216
rect 3605 5219 3663 5225
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 3605 5185 3617 5219
rect 3651 5185 3663 5219
rect 3872 5216 3884 5225
rect 3839 5188 3884 5216
rect 3605 5179 3663 5185
rect 3872 5179 3884 5188
rect 3878 5176 3884 5179
rect 3936 5176 3942 5228
rect 6380 5225 6408 5256
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 6932 5225 6960 5324
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 11514 5352 11520 5364
rect 11475 5324 11520 5352
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 13078 5312 13084 5364
rect 13136 5352 13142 5364
rect 13265 5355 13323 5361
rect 13265 5352 13277 5355
rect 13136 5324 13277 5352
rect 13136 5312 13142 5324
rect 13265 5321 13277 5324
rect 13311 5321 13323 5355
rect 14918 5352 14924 5364
rect 14879 5324 14924 5352
rect 13265 5315 13323 5321
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 19886 5352 19892 5364
rect 19847 5324 19892 5352
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 9674 5284 9680 5296
rect 8772 5256 9680 5284
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6512 5188 6561 5216
rect 6512 5176 6518 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5185 6975 5219
rect 6917 5179 6975 5185
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 8386 5216 8392 5228
rect 8347 5188 8392 5216
rect 7009 5179 7067 5185
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 7024 5148 7052 5179
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 8570 5216 8576 5228
rect 8531 5188 8576 5216
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 8772 5225 8800 5256
rect 9674 5244 9680 5256
rect 9732 5284 9738 5296
rect 10594 5284 10600 5296
rect 9732 5256 10600 5284
rect 9732 5244 9738 5256
rect 10594 5244 10600 5256
rect 10652 5284 10658 5296
rect 13998 5284 14004 5296
rect 10652 5256 14004 5284
rect 10652 5244 10658 5256
rect 13998 5244 14004 5256
rect 14056 5244 14062 5296
rect 15746 5284 15752 5296
rect 15120 5256 15752 5284
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 8941 5219 8999 5225
rect 8941 5185 8953 5219
rect 8987 5216 8999 5219
rect 10042 5216 10048 5228
rect 8987 5188 10048 5216
rect 8987 5185 8999 5188
rect 8941 5179 8999 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 6052 5120 7052 5148
rect 8665 5151 8723 5157
rect 6052 5108 6058 5120
rect 8665 5117 8677 5151
rect 8711 5148 8723 5151
rect 9950 5148 9956 5160
rect 8711 5120 9956 5148
rect 8711 5117 8723 5120
rect 8665 5111 8723 5117
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 10796 5148 10824 5179
rect 11238 5176 11244 5228
rect 11296 5216 11302 5228
rect 11698 5216 11704 5228
rect 11296 5188 11704 5216
rect 11296 5176 11302 5188
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 12894 5176 12900 5228
rect 12952 5216 12958 5228
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 12952 5188 13093 5216
rect 12952 5176 12958 5188
rect 13081 5185 13093 5188
rect 13127 5185 13139 5219
rect 13906 5216 13912 5228
rect 13867 5188 13912 5216
rect 13081 5179 13139 5185
rect 11514 5148 11520 5160
rect 10796 5120 11520 5148
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5148 12035 5151
rect 12802 5148 12808 5160
rect 12023 5120 12808 5148
rect 12023 5117 12035 5120
rect 11977 5111 12035 5117
rect 12802 5108 12808 5120
rect 12860 5108 12866 5160
rect 5534 5040 5540 5092
rect 5592 5080 5598 5092
rect 6365 5083 6423 5089
rect 6365 5080 6377 5083
rect 5592 5052 6377 5080
rect 5592 5040 5598 5052
rect 6365 5049 6377 5052
rect 6411 5049 6423 5083
rect 6365 5043 6423 5049
rect 10965 5083 11023 5089
rect 10965 5049 10977 5083
rect 11011 5080 11023 5083
rect 12526 5080 12532 5092
rect 11011 5052 12532 5080
rect 11011 5049 11023 5052
rect 10965 5043 11023 5049
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 13096 5080 13124 5179
rect 13906 5176 13912 5188
rect 13964 5176 13970 5228
rect 15120 5225 15148 5256
rect 15746 5244 15752 5256
rect 15804 5244 15810 5296
rect 15105 5219 15163 5225
rect 15105 5185 15117 5219
rect 15151 5185 15163 5219
rect 15381 5219 15439 5225
rect 15381 5216 15393 5219
rect 15105 5179 15163 5185
rect 15212 5188 15393 5216
rect 15010 5108 15016 5160
rect 15068 5148 15074 5160
rect 15212 5148 15240 5188
rect 15381 5185 15393 5188
rect 15427 5185 15439 5219
rect 15381 5179 15439 5185
rect 15473 5219 15531 5225
rect 15473 5185 15485 5219
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 15068 5120 15240 5148
rect 15289 5151 15347 5157
rect 15068 5108 15074 5120
rect 15289 5117 15301 5151
rect 15335 5117 15347 5151
rect 15488 5148 15516 5179
rect 15562 5176 15568 5228
rect 15620 5216 15626 5228
rect 15657 5219 15715 5225
rect 15657 5216 15669 5219
rect 15620 5188 15669 5216
rect 15620 5176 15626 5188
rect 15657 5185 15669 5188
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 16298 5176 16304 5228
rect 16356 5216 16362 5228
rect 16853 5219 16911 5225
rect 16853 5216 16865 5219
rect 16356 5188 16865 5216
rect 16356 5176 16362 5188
rect 16853 5185 16865 5188
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5216 18107 5219
rect 18138 5216 18144 5228
rect 18095 5188 18144 5216
rect 18095 5185 18107 5188
rect 18049 5179 18107 5185
rect 18138 5176 18144 5188
rect 18196 5176 18202 5228
rect 20622 5176 20628 5228
rect 20680 5216 20686 5228
rect 21002 5219 21060 5225
rect 21002 5216 21014 5219
rect 20680 5188 21014 5216
rect 20680 5176 20686 5188
rect 21002 5185 21014 5188
rect 21048 5185 21060 5219
rect 21266 5216 21272 5228
rect 21227 5188 21272 5216
rect 21002 5179 21060 5185
rect 21266 5176 21272 5188
rect 21324 5176 21330 5228
rect 29730 5176 29736 5228
rect 29788 5216 29794 5228
rect 29825 5219 29883 5225
rect 29825 5216 29837 5219
rect 29788 5188 29837 5216
rect 29788 5176 29794 5188
rect 29825 5185 29837 5188
rect 29871 5185 29883 5219
rect 29825 5179 29883 5185
rect 16574 5148 16580 5160
rect 15488 5120 16580 5148
rect 15289 5111 15347 5117
rect 13725 5083 13783 5089
rect 13725 5080 13737 5083
rect 13096 5052 13737 5080
rect 13725 5049 13737 5052
rect 13771 5049 13783 5083
rect 15304 5080 15332 5111
rect 16574 5108 16580 5120
rect 16632 5108 16638 5160
rect 17773 5151 17831 5157
rect 17773 5117 17785 5151
rect 17819 5148 17831 5151
rect 18230 5148 18236 5160
rect 17819 5120 18236 5148
rect 17819 5117 17831 5120
rect 17773 5111 17831 5117
rect 18230 5108 18236 5120
rect 18288 5148 18294 5160
rect 18966 5148 18972 5160
rect 18288 5120 18972 5148
rect 18288 5108 18294 5120
rect 18966 5108 18972 5120
rect 19024 5108 19030 5160
rect 17586 5080 17592 5092
rect 15304 5052 17592 5080
rect 13725 5043 13783 5049
rect 17586 5040 17592 5052
rect 17644 5040 17650 5092
rect 9122 5012 9128 5024
rect 9083 4984 9128 5012
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 11885 5015 11943 5021
rect 11885 4981 11897 5015
rect 11931 5012 11943 5015
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 11931 4984 12909 5012
rect 11931 4981 11943 4984
rect 11885 4975 11943 4981
rect 12897 4981 12909 4984
rect 12943 5012 12955 5015
rect 13630 5012 13636 5024
rect 12943 4984 13636 5012
rect 12943 4981 12955 4984
rect 12897 4975 12955 4981
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 15102 4972 15108 5024
rect 15160 5012 15166 5024
rect 16669 5015 16727 5021
rect 16669 5012 16681 5015
rect 15160 4984 16681 5012
rect 15160 4972 15166 4984
rect 16669 4981 16681 4984
rect 16715 4981 16727 5015
rect 16669 4975 16727 4981
rect 17865 5015 17923 5021
rect 17865 4981 17877 5015
rect 17911 5012 17923 5015
rect 18046 5012 18052 5024
rect 17911 4984 18052 5012
rect 17911 4981 17923 4984
rect 17865 4975 17923 4981
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 30006 5012 30012 5024
rect 29967 4984 30012 5012
rect 30006 4972 30012 4984
rect 30064 4972 30070 5024
rect 1104 4922 30820 4944
rect 1104 4870 5915 4922
rect 5967 4870 5979 4922
rect 6031 4870 6043 4922
rect 6095 4870 6107 4922
rect 6159 4870 6171 4922
rect 6223 4870 15846 4922
rect 15898 4870 15910 4922
rect 15962 4870 15974 4922
rect 16026 4870 16038 4922
rect 16090 4870 16102 4922
rect 16154 4870 25776 4922
rect 25828 4870 25840 4922
rect 25892 4870 25904 4922
rect 25956 4870 25968 4922
rect 26020 4870 26032 4922
rect 26084 4870 30820 4922
rect 1104 4848 30820 4870
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 6454 4808 6460 4820
rect 5224 4780 6460 4808
rect 5224 4768 5230 4780
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 6549 4811 6607 4817
rect 6549 4777 6561 4811
rect 6595 4808 6607 4811
rect 6914 4808 6920 4820
rect 6595 4780 6920 4808
rect 6595 4777 6607 4780
rect 6549 4771 6607 4777
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 9858 4808 9864 4820
rect 7024 4780 9864 4808
rect 5902 4700 5908 4752
rect 5960 4740 5966 4752
rect 7024 4740 7052 4780
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 10686 4768 10692 4820
rect 10744 4808 10750 4820
rect 11241 4811 11299 4817
rect 11241 4808 11253 4811
rect 10744 4780 11253 4808
rect 10744 4768 10750 4780
rect 11241 4777 11253 4780
rect 11287 4777 11299 4811
rect 11241 4771 11299 4777
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 14182 4808 14188 4820
rect 14139 4780 14188 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4808 15347 4811
rect 15378 4808 15384 4820
rect 15335 4780 15384 4808
rect 15335 4777 15347 4780
rect 15289 4771 15347 4777
rect 15378 4768 15384 4780
rect 15436 4768 15442 4820
rect 18690 4808 18696 4820
rect 18064 4780 18696 4808
rect 18064 4752 18092 4780
rect 18690 4768 18696 4780
rect 18748 4768 18754 4820
rect 19334 4808 19340 4820
rect 19295 4780 19340 4808
rect 19334 4768 19340 4780
rect 19392 4768 19398 4820
rect 20254 4808 20260 4820
rect 19444 4780 20260 4808
rect 5960 4712 7052 4740
rect 12437 4743 12495 4749
rect 5960 4700 5966 4712
rect 12437 4709 12449 4743
rect 12483 4709 12495 4743
rect 18046 4740 18052 4752
rect 12437 4703 12495 4709
rect 14108 4712 18052 4740
rect 1210 4632 1216 4684
rect 1268 4672 1274 4684
rect 1397 4675 1455 4681
rect 1397 4672 1409 4675
rect 1268 4644 1409 4672
rect 1268 4632 1274 4644
rect 1397 4641 1409 4644
rect 1443 4641 1455 4675
rect 1397 4635 1455 4641
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4672 1731 4675
rect 4614 4672 4620 4684
rect 1719 4644 4620 4672
rect 1719 4641 1731 4644
rect 1673 4635 1731 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 5442 4632 5448 4684
rect 5500 4672 5506 4684
rect 5721 4675 5779 4681
rect 5721 4672 5733 4675
rect 5500 4644 5733 4672
rect 5500 4632 5506 4644
rect 5721 4641 5733 4644
rect 5767 4672 5779 4675
rect 6638 4672 6644 4684
rect 5767 4644 6644 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 7929 4675 7987 4681
rect 7929 4641 7941 4675
rect 7975 4672 7987 4675
rect 8294 4672 8300 4684
rect 7975 4644 8300 4672
rect 7975 4641 7987 4644
rect 7929 4635 7987 4641
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 9309 4675 9367 4681
rect 9309 4641 9321 4675
rect 9355 4672 9367 4675
rect 9674 4672 9680 4684
rect 9355 4644 9680 4672
rect 9355 4641 9367 4644
rect 9309 4635 9367 4641
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4604 5595 4607
rect 5626 4604 5632 4616
rect 5583 4576 5632 4604
rect 5583 4573 5595 4576
rect 5537 4567 5595 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 5828 4536 5856 4567
rect 5902 4564 5908 4616
rect 5960 4604 5966 4616
rect 6089 4607 6147 4613
rect 5960 4576 6005 4604
rect 5960 4564 5966 4576
rect 6089 4573 6101 4607
rect 6135 4604 6147 4607
rect 6362 4604 6368 4616
rect 6135 4576 6368 4604
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 6362 4564 6368 4576
rect 6420 4604 6426 4616
rect 6546 4604 6552 4616
rect 6420 4576 6552 4604
rect 6420 4564 6426 4576
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8444 4576 8953 4604
rect 8444 4564 8450 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 6730 4536 6736 4548
rect 5828 4508 6736 4536
rect 6730 4496 6736 4508
rect 6788 4496 6794 4548
rect 7098 4496 7104 4548
rect 7156 4536 7162 4548
rect 7662 4539 7720 4545
rect 7662 4536 7674 4539
rect 7156 4508 7674 4536
rect 7156 4496 7162 4508
rect 7662 4505 7674 4508
rect 7708 4505 7720 4539
rect 8956 4536 8984 4567
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 9088 4576 9137 4604
rect 9088 4564 9094 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9493 4607 9551 4613
rect 9263 4576 9444 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 9306 4536 9312 4548
rect 8956 4508 9312 4536
rect 7662 4499 7720 4505
rect 9306 4496 9312 4508
rect 9364 4496 9370 4548
rect 9416 4536 9444 4576
rect 9493 4573 9505 4607
rect 9539 4604 9551 4607
rect 9766 4604 9772 4616
rect 9539 4576 9772 4604
rect 9539 4573 9551 4576
rect 9493 4567 9551 4573
rect 9766 4564 9772 4576
rect 9824 4604 9830 4616
rect 10502 4604 10508 4616
rect 9824 4576 10508 4604
rect 9824 4564 9830 4576
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 10689 4607 10747 4613
rect 10689 4573 10701 4607
rect 10735 4604 10747 4607
rect 12452 4604 12480 4703
rect 14108 4684 14136 4712
rect 18046 4700 18052 4712
rect 18104 4700 18110 4752
rect 19444 4740 19472 4780
rect 20254 4768 20260 4780
rect 20312 4768 20318 4820
rect 20622 4808 20628 4820
rect 20583 4780 20628 4808
rect 20622 4768 20628 4780
rect 20680 4768 20686 4820
rect 18340 4712 19472 4740
rect 13078 4672 13084 4684
rect 12544 4644 13084 4672
rect 12544 4613 12572 4644
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13541 4675 13599 4681
rect 13541 4641 13553 4675
rect 13587 4672 13599 4675
rect 14090 4672 14096 4684
rect 13587 4644 14096 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 14550 4672 14556 4684
rect 14511 4644 14556 4672
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 15841 4675 15899 4681
rect 15841 4672 15853 4675
rect 14783 4644 15853 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 15841 4641 15853 4644
rect 15887 4641 15899 4675
rect 15841 4635 15899 4641
rect 10735 4576 12480 4604
rect 12529 4607 12587 4613
rect 10735 4573 10747 4576
rect 10689 4567 10747 4573
rect 9416 4508 9812 4536
rect 5353 4471 5411 4477
rect 5353 4437 5365 4471
rect 5399 4468 5411 4471
rect 5534 4468 5540 4480
rect 5399 4440 5540 4468
rect 5399 4437 5411 4440
rect 5353 4431 5411 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 9674 4468 9680 4480
rect 9635 4440 9680 4468
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 9784 4468 9812 4508
rect 9858 4496 9864 4548
rect 9916 4536 9922 4548
rect 10612 4536 10640 4567
rect 9916 4508 10640 4536
rect 11425 4539 11483 4545
rect 9916 4496 9922 4508
rect 11425 4505 11437 4539
rect 11471 4505 11483 4539
rect 11606 4536 11612 4548
rect 11567 4508 11612 4536
rect 11425 4499 11483 4505
rect 9950 4468 9956 4480
rect 9784 4440 9956 4468
rect 9950 4428 9956 4440
rect 10008 4468 10014 4480
rect 10410 4468 10416 4480
rect 10008 4440 10416 4468
rect 10008 4428 10014 4440
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 11440 4468 11468 4499
rect 11606 4496 11612 4508
rect 11664 4496 11670 4548
rect 11882 4496 11888 4548
rect 11940 4536 11946 4548
rect 12253 4539 12311 4545
rect 12253 4536 12265 4539
rect 11940 4508 12265 4536
rect 11940 4496 11946 4508
rect 12253 4505 12265 4508
rect 12299 4505 12311 4539
rect 12360 4536 12388 4576
rect 12529 4573 12541 4607
rect 12575 4573 12587 4607
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 12529 4567 12587 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13630 4564 13636 4616
rect 13688 4604 13694 4616
rect 14752 4604 14780 4635
rect 13688 4576 14780 4604
rect 15856 4604 15884 4635
rect 15930 4632 15936 4684
rect 15988 4672 15994 4684
rect 16853 4675 16911 4681
rect 16853 4672 16865 4675
rect 15988 4644 16865 4672
rect 15988 4632 15994 4644
rect 16853 4641 16865 4644
rect 16899 4641 16911 4675
rect 16853 4635 16911 4641
rect 17770 4632 17776 4684
rect 17828 4672 17834 4684
rect 18340 4681 18368 4712
rect 19886 4700 19892 4752
rect 19944 4700 19950 4752
rect 18233 4675 18291 4681
rect 18233 4672 18245 4675
rect 17828 4644 18245 4672
rect 17828 4632 17834 4644
rect 18233 4641 18245 4644
rect 18279 4641 18291 4675
rect 18233 4635 18291 4641
rect 18325 4675 18383 4681
rect 18325 4641 18337 4675
rect 18371 4641 18383 4675
rect 19904 4672 19932 4700
rect 18325 4635 18383 4641
rect 18616 4644 19564 4672
rect 19904 4644 20484 4672
rect 16390 4604 16396 4616
rect 15856 4576 16396 4604
rect 13688 4564 13694 4576
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 16669 4607 16727 4613
rect 16669 4573 16681 4607
rect 16715 4604 16727 4607
rect 16758 4604 16764 4616
rect 16715 4576 16764 4604
rect 16715 4573 16727 4576
rect 16669 4567 16727 4573
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4573 17003 4607
rect 16945 4567 17003 4573
rect 12434 4536 12440 4548
rect 12360 4508 12440 4536
rect 12253 4499 12311 4505
rect 12434 4496 12440 4508
rect 12492 4496 12498 4548
rect 14461 4539 14519 4545
rect 14461 4505 14473 4539
rect 14507 4536 14519 4539
rect 15010 4536 15016 4548
rect 14507 4508 15016 4536
rect 14507 4505 14519 4508
rect 14461 4499 14519 4505
rect 15010 4496 15016 4508
rect 15068 4496 15074 4548
rect 16022 4496 16028 4548
rect 16080 4536 16086 4548
rect 16960 4536 16988 4567
rect 17494 4564 17500 4616
rect 17552 4604 17558 4616
rect 17957 4607 18015 4613
rect 17957 4604 17969 4607
rect 17552 4576 17969 4604
rect 17552 4564 17558 4576
rect 17957 4573 17969 4576
rect 18003 4573 18015 4607
rect 17957 4567 18015 4573
rect 16080 4508 16988 4536
rect 16080 4496 16086 4508
rect 12066 4468 12072 4480
rect 11440 4440 12072 4468
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 12526 4468 12532 4480
rect 12487 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 15562 4428 15568 4480
rect 15620 4468 15626 4480
rect 15657 4471 15715 4477
rect 15657 4468 15669 4471
rect 15620 4440 15669 4468
rect 15620 4428 15626 4440
rect 15657 4437 15669 4440
rect 15703 4437 15715 4471
rect 15657 4431 15715 4437
rect 15746 4428 15752 4480
rect 15804 4468 15810 4480
rect 16482 4468 16488 4480
rect 15804 4440 15849 4468
rect 16443 4440 16488 4468
rect 15804 4428 15810 4440
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 17972 4468 18000 4567
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 18141 4607 18199 4613
rect 18141 4604 18153 4607
rect 18104 4576 18153 4604
rect 18104 4564 18110 4576
rect 18141 4573 18153 4576
rect 18187 4573 18199 4607
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 18141 4567 18199 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 18616 4468 18644 4644
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19392 4576 19441 4604
rect 19392 4564 19398 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19536 4604 19564 4644
rect 19794 4604 19800 4616
rect 19536 4576 19800 4604
rect 19429 4567 19487 4573
rect 19794 4564 19800 4576
rect 19852 4604 19858 4616
rect 19889 4607 19947 4613
rect 19889 4604 19901 4607
rect 19852 4576 19901 4604
rect 19852 4564 19858 4576
rect 19889 4573 19901 4576
rect 19935 4573 19947 4607
rect 20070 4604 20076 4616
rect 20031 4576 20076 4604
rect 19889 4567 19947 4573
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20165 4607 20223 4613
rect 20165 4573 20177 4607
rect 20211 4573 20223 4607
rect 20165 4567 20223 4573
rect 18693 4539 18751 4545
rect 18693 4505 18705 4539
rect 18739 4536 18751 4539
rect 18739 4508 19472 4536
rect 18739 4505 18751 4508
rect 18693 4499 18751 4505
rect 19444 4480 19472 4508
rect 19978 4496 19984 4548
rect 20036 4536 20042 4548
rect 20180 4536 20208 4567
rect 20254 4564 20260 4616
rect 20312 4604 20318 4616
rect 20456 4613 20484 4644
rect 20441 4607 20499 4613
rect 20312 4576 20357 4604
rect 20312 4564 20318 4576
rect 20441 4573 20453 4607
rect 20487 4573 20499 4607
rect 20441 4567 20499 4573
rect 30101 4607 30159 4613
rect 30101 4573 30113 4607
rect 30147 4604 30159 4607
rect 30929 4607 30987 4613
rect 30929 4604 30941 4607
rect 30147 4576 30941 4604
rect 30147 4573 30159 4576
rect 30101 4567 30159 4573
rect 30929 4573 30941 4576
rect 30975 4573 30987 4607
rect 30929 4567 30987 4573
rect 20036 4508 20208 4536
rect 20272 4536 20300 4564
rect 20530 4536 20536 4548
rect 20272 4508 20536 4536
rect 20036 4496 20042 4508
rect 20530 4496 20536 4508
rect 20588 4496 20594 4548
rect 17972 4440 18644 4468
rect 19426 4428 19432 4480
rect 19484 4428 19490 4480
rect 29638 4428 29644 4480
rect 29696 4468 29702 4480
rect 29917 4471 29975 4477
rect 29917 4468 29929 4471
rect 29696 4440 29929 4468
rect 29696 4428 29702 4440
rect 29917 4437 29929 4440
rect 29963 4437 29975 4471
rect 29917 4431 29975 4437
rect 1104 4378 30820 4400
rect 1104 4326 10880 4378
rect 10932 4326 10944 4378
rect 10996 4326 11008 4378
rect 11060 4326 11072 4378
rect 11124 4326 11136 4378
rect 11188 4326 20811 4378
rect 20863 4326 20875 4378
rect 20927 4326 20939 4378
rect 20991 4326 21003 4378
rect 21055 4326 21067 4378
rect 21119 4326 30820 4378
rect 1104 4304 30820 4326
rect 5902 4264 5908 4276
rect 5184 4236 5908 4264
rect 1854 4196 1860 4208
rect 1815 4168 1860 4196
rect 1854 4156 1860 4168
rect 1912 4156 1918 4208
rect 5184 4196 5212 4236
rect 5902 4224 5908 4236
rect 5960 4224 5966 4276
rect 6730 4224 6736 4276
rect 6788 4224 6794 4276
rect 7098 4264 7104 4276
rect 7059 4236 7104 4264
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 9677 4267 9735 4273
rect 9677 4233 9689 4267
rect 9723 4264 9735 4267
rect 10042 4264 10048 4276
rect 9723 4236 10048 4264
rect 9723 4233 9735 4236
rect 9677 4227 9735 4233
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 15562 4264 15568 4276
rect 15523 4236 15568 4264
rect 15562 4224 15568 4236
rect 15620 4224 15626 4276
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 16669 4267 16727 4273
rect 16669 4264 16681 4267
rect 16632 4236 16681 4264
rect 16632 4224 16638 4236
rect 16669 4233 16681 4236
rect 16715 4233 16727 4267
rect 16669 4227 16727 4233
rect 18325 4267 18383 4273
rect 18325 4233 18337 4267
rect 18371 4264 18383 4267
rect 18506 4264 18512 4276
rect 18371 4236 18512 4264
rect 18371 4233 18383 4236
rect 18325 4227 18383 4233
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 6748 4196 6776 4224
rect 3528 4168 3740 4196
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 2832 4100 2877 4128
rect 2832 4088 2838 4100
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3528 4128 3556 4168
rect 3200 4100 3556 4128
rect 3605 4131 3663 4137
rect 3200 4088 3206 4100
rect 3605 4097 3617 4131
rect 3651 4097 3663 4131
rect 3712 4128 3740 4168
rect 5092 4168 5212 4196
rect 6656 4168 6776 4196
rect 8564 4199 8622 4205
rect 5092 4128 5120 4168
rect 3712 4100 5120 4128
rect 3605 4091 3663 4097
rect 2590 4020 2596 4072
rect 2648 4060 2654 4072
rect 3620 4060 3648 4091
rect 5166 4088 5172 4140
rect 5224 4128 5230 4140
rect 5350 4128 5356 4140
rect 5224 4100 5269 4128
rect 5311 4100 5356 4128
rect 5224 4088 5230 4100
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4097 5595 4131
rect 5537 4091 5595 4097
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 6362 4128 6368 4140
rect 5767 4100 6368 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 2648 4032 3648 4060
rect 2648 4020 2654 4032
rect 5074 4020 5080 4072
rect 5132 4060 5138 4072
rect 5445 4063 5503 4069
rect 5132 4032 5304 4060
rect 5132 4020 5138 4032
rect 3050 3992 3056 4004
rect 3011 3964 3056 3992
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 3789 3995 3847 4001
rect 3789 3961 3801 3995
rect 3835 3992 3847 3995
rect 5276 3992 5304 4032
rect 5445 4029 5457 4063
rect 5491 4029 5503 4063
rect 5552 4060 5580 4091
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 6546 4128 6552 4140
rect 6507 4100 6552 4128
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 6656 4137 6684 4168
rect 8564 4165 8576 4199
rect 8610 4196 8622 4199
rect 9122 4196 9128 4208
rect 8610 4168 9128 4196
rect 8610 4165 8622 4168
rect 8564 4159 8622 4165
rect 9122 4156 9128 4168
rect 9180 4156 9186 4208
rect 13354 4156 13360 4208
rect 13412 4196 13418 4208
rect 17034 4196 17040 4208
rect 13412 4168 13952 4196
rect 16995 4168 17040 4196
rect 13412 4156 13418 4168
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 6914 4128 6920 4140
rect 6788 4100 6833 4128
rect 6875 4100 6920 4128
rect 6788 4088 6794 4100
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 8294 4128 8300 4140
rect 8255 4100 8300 4128
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 9858 4128 9864 4140
rect 8404 4100 9864 4128
rect 5810 4060 5816 4072
rect 5552 4032 5816 4060
rect 5445 4023 5503 4029
rect 5460 3992 5488 4023
rect 5810 4020 5816 4032
rect 5868 4060 5874 4072
rect 7558 4060 7564 4072
rect 5868 4032 7564 4060
rect 5868 4020 5874 4032
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 8404 4060 8432 4100
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 8312 4032 8432 4060
rect 8312 3992 8340 4032
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 10152 4060 10180 4091
rect 9364 4032 10180 4060
rect 9364 4020 9370 4032
rect 3835 3964 5120 3992
rect 5276 3964 5488 3992
rect 6656 3964 8340 3992
rect 3835 3961 3847 3964
rect 3789 3955 3847 3961
rect 2133 3927 2191 3933
rect 2133 3893 2145 3927
rect 2179 3924 2191 3927
rect 4798 3924 4804 3936
rect 2179 3896 4804 3924
rect 2179 3893 2191 3896
rect 2133 3887 2191 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5092 3924 5120 3964
rect 6656 3924 6684 3964
rect 5092 3896 6684 3924
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 10336 3924 10364 4091
rect 10410 4088 10416 4140
rect 10468 4128 10474 4140
rect 10689 4131 10747 4137
rect 10468 4100 10513 4128
rect 10468 4088 10474 4100
rect 10689 4097 10701 4131
rect 10735 4128 10747 4131
rect 10778 4128 10784 4140
rect 10735 4100 10784 4128
rect 10735 4097 10747 4100
rect 10689 4091 10747 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4128 12035 4131
rect 12066 4128 12072 4140
rect 12023 4100 12072 4128
rect 12023 4097 12035 4100
rect 11977 4091 12035 4097
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12526 4088 12532 4140
rect 12584 4128 12590 4140
rect 13722 4128 13728 4140
rect 12584 4100 13728 4128
rect 12584 4088 12590 4100
rect 13722 4088 13728 4100
rect 13780 4128 13786 4140
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13780 4100 13829 4128
rect 13780 4088 13786 4100
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 13924 4128 13952 4168
rect 17034 4156 17040 4168
rect 17092 4156 17098 4208
rect 19334 4156 19340 4208
rect 19392 4196 19398 4208
rect 19392 4168 20484 4196
rect 19392 4156 19398 4168
rect 14277 4131 14335 4137
rect 14277 4128 14289 4131
rect 13924 4100 14289 4128
rect 13817 4091 13875 4097
rect 14277 4097 14289 4100
rect 14323 4097 14335 4131
rect 14277 4091 14335 4097
rect 15378 4088 15384 4140
rect 15436 4128 15442 4140
rect 15746 4128 15752 4140
rect 15436 4100 15752 4128
rect 15436 4088 15442 4100
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 15930 4128 15936 4140
rect 15891 4100 15936 4128
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 16022 4088 16028 4140
rect 16080 4128 16086 4140
rect 17129 4131 17187 4137
rect 16080 4100 16125 4128
rect 16080 4088 16086 4100
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17310 4128 17316 4140
rect 17175 4100 17316 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 19426 4088 19432 4140
rect 19484 4137 19490 4140
rect 19484 4128 19496 4137
rect 19702 4128 19708 4140
rect 19484 4100 19529 4128
rect 19663 4100 19708 4128
rect 19484 4091 19496 4100
rect 19484 4088 19490 4091
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 19794 4088 19800 4140
rect 19852 4128 19858 4140
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 19852 4100 20177 4128
rect 19852 4088 19858 4100
rect 20165 4097 20177 4100
rect 20211 4097 20223 4131
rect 20346 4128 20352 4140
rect 20307 4100 20352 4128
rect 20165 4091 20223 4097
rect 20346 4088 20352 4100
rect 20404 4088 20410 4140
rect 20456 4128 20484 4168
rect 20717 4131 20775 4137
rect 20717 4128 20729 4131
rect 20456 4100 20729 4128
rect 20717 4097 20729 4100
rect 20763 4097 20775 4131
rect 20717 4091 20775 4097
rect 21358 4088 21364 4140
rect 21416 4128 21422 4140
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 21416 4100 22017 4128
rect 21416 4088 21422 4100
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 29273 4131 29331 4137
rect 29273 4097 29285 4131
rect 29319 4097 29331 4131
rect 30098 4128 30104 4140
rect 30059 4100 30104 4128
rect 29273 4091 29331 4097
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4060 10563 4063
rect 10594 4060 10600 4072
rect 10551 4032 10600 4060
rect 10551 4029 10563 4032
rect 10505 4023 10563 4029
rect 10594 4020 10600 4032
rect 10652 4020 10658 4072
rect 11882 4060 11888 4072
rect 11843 4032 11888 4060
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 12158 4020 12164 4072
rect 12216 4060 12222 4072
rect 12618 4060 12624 4072
rect 12216 4032 12624 4060
rect 12216 4020 12222 4032
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 12802 4020 12808 4072
rect 12860 4060 12866 4072
rect 13541 4063 13599 4069
rect 13541 4060 13553 4063
rect 12860 4032 13553 4060
rect 12860 4020 12866 4032
rect 13541 4029 13553 4032
rect 13587 4029 13599 4063
rect 13541 4023 13599 4029
rect 14553 4063 14611 4069
rect 14553 4029 14565 4063
rect 14599 4060 14611 4063
rect 15286 4060 15292 4072
rect 14599 4032 15292 4060
rect 14599 4029 14611 4032
rect 14553 4023 14611 4029
rect 15286 4020 15292 4032
rect 15344 4060 15350 4072
rect 15948 4060 15976 4088
rect 15344 4032 15976 4060
rect 15344 4020 15350 4032
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 17218 4060 17224 4072
rect 16448 4032 17224 4060
rect 16448 4020 16454 4032
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 19978 4020 19984 4072
rect 20036 4060 20042 4072
rect 20441 4063 20499 4069
rect 20441 4060 20453 4063
rect 20036 4032 20453 4060
rect 20036 4020 20042 4032
rect 20441 4029 20453 4032
rect 20487 4029 20499 4063
rect 20441 4023 20499 4029
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 29288 4060 29316 4091
rect 30098 4088 30104 4100
rect 30156 4088 30162 4140
rect 31570 4060 31576 4072
rect 20588 4032 20633 4060
rect 29288 4032 31576 4060
rect 20588 4020 20594 4032
rect 31570 4020 31576 4032
rect 31628 4020 31634 4072
rect 11609 3995 11667 4001
rect 11609 3961 11621 3995
rect 11655 3992 11667 3995
rect 11790 3992 11796 4004
rect 11655 3964 11796 3992
rect 11655 3961 11667 3964
rect 11609 3955 11667 3961
rect 11790 3952 11796 3964
rect 11848 3952 11854 4004
rect 12526 3952 12532 4004
rect 12584 3992 12590 4004
rect 13906 3992 13912 4004
rect 12584 3964 13912 3992
rect 12584 3952 12590 3964
rect 13906 3952 13912 3964
rect 13964 3952 13970 4004
rect 14182 3952 14188 4004
rect 14240 3992 14246 4004
rect 16298 3992 16304 4004
rect 14240 3964 16304 3992
rect 14240 3952 14246 3964
rect 16298 3952 16304 3964
rect 16356 3952 16362 4004
rect 20070 3952 20076 4004
rect 20128 3992 20134 4004
rect 20622 3992 20628 4004
rect 20128 3964 20628 3992
rect 20128 3952 20134 3964
rect 20622 3952 20628 3964
rect 20680 3992 20686 4004
rect 21450 3992 21456 4004
rect 20680 3964 21456 3992
rect 20680 3952 20686 3964
rect 21450 3952 21456 3964
rect 21508 3992 21514 4004
rect 21821 3995 21879 4001
rect 21821 3992 21833 3995
rect 21508 3964 21833 3992
rect 21508 3952 21514 3964
rect 21821 3961 21833 3964
rect 21867 3961 21879 3995
rect 21821 3955 21879 3961
rect 10870 3924 10876 3936
rect 6788 3896 10364 3924
rect 10831 3896 10876 3924
rect 6788 3884 6794 3896
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 11977 3927 12035 3933
rect 11977 3893 11989 3927
rect 12023 3924 12035 3927
rect 12434 3924 12440 3936
rect 12023 3896 12440 3924
rect 12023 3893 12035 3896
rect 11977 3887 12035 3893
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 20898 3924 20904 3936
rect 20859 3896 20904 3924
rect 20898 3884 20904 3896
rect 20956 3884 20962 3936
rect 21174 3884 21180 3936
rect 21232 3924 21238 3936
rect 21542 3924 21548 3936
rect 21232 3896 21548 3924
rect 21232 3884 21238 3896
rect 21542 3884 21548 3896
rect 21600 3884 21606 3936
rect 29457 3927 29515 3933
rect 29457 3893 29469 3927
rect 29503 3924 29515 3927
rect 29546 3924 29552 3936
rect 29503 3896 29552 3924
rect 29503 3893 29515 3896
rect 29457 3887 29515 3893
rect 29546 3884 29552 3896
rect 29604 3884 29610 3936
rect 29917 3927 29975 3933
rect 29917 3893 29929 3927
rect 29963 3924 29975 3927
rect 30006 3924 30012 3936
rect 29963 3896 30012 3924
rect 29963 3893 29975 3896
rect 29917 3887 29975 3893
rect 30006 3884 30012 3896
rect 30064 3884 30070 3936
rect 1104 3834 30820 3856
rect 1104 3782 5915 3834
rect 5967 3782 5979 3834
rect 6031 3782 6043 3834
rect 6095 3782 6107 3834
rect 6159 3782 6171 3834
rect 6223 3782 15846 3834
rect 15898 3782 15910 3834
rect 15962 3782 15974 3834
rect 16026 3782 16038 3834
rect 16090 3782 16102 3834
rect 16154 3782 25776 3834
rect 25828 3782 25840 3834
rect 25892 3782 25904 3834
rect 25956 3782 25968 3834
rect 26020 3782 26032 3834
rect 26084 3782 30820 3834
rect 1104 3760 30820 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 2314 3720 2320 3732
rect 1627 3692 2320 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 2464 3692 2509 3720
rect 2464 3680 2470 3692
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4433 3723 4491 3729
rect 4433 3720 4445 3723
rect 4304 3692 4445 3720
rect 4304 3680 4310 3692
rect 4433 3689 4445 3692
rect 4479 3689 4491 3723
rect 4433 3683 4491 3689
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 6641 3723 6699 3729
rect 6641 3720 6653 3723
rect 5684 3692 6653 3720
rect 5684 3680 5690 3692
rect 6641 3689 6653 3692
rect 6687 3689 6699 3723
rect 6641 3683 6699 3689
rect 10134 3680 10140 3732
rect 10192 3720 10198 3732
rect 10778 3720 10784 3732
rect 10192 3692 10640 3720
rect 10739 3692 10784 3720
rect 10192 3680 10198 3692
rect 6546 3612 6552 3664
rect 6604 3652 6610 3664
rect 6822 3652 6828 3664
rect 6604 3624 6828 3652
rect 6604 3612 6610 3624
rect 6822 3612 6828 3624
rect 6880 3652 6886 3664
rect 8938 3652 8944 3664
rect 6880 3624 8944 3652
rect 6880 3612 6886 3624
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 4212 3556 5273 3584
rect 4212 3544 4218 3556
rect 5261 3553 5273 3556
rect 5307 3553 5319 3587
rect 5261 3547 5319 3553
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 9214 3584 9220 3596
rect 8352 3556 9220 3584
rect 8352 3544 8358 3556
rect 9214 3544 9220 3556
rect 9272 3584 9278 3596
rect 9401 3587 9459 3593
rect 9401 3584 9413 3587
rect 9272 3556 9413 3584
rect 9272 3544 9278 3556
rect 9401 3553 9413 3556
rect 9447 3553 9459 3587
rect 10612 3584 10640 3692
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 11425 3723 11483 3729
rect 11425 3689 11437 3723
rect 11471 3720 11483 3723
rect 12434 3720 12440 3732
rect 11471 3692 12440 3720
rect 11471 3689 11483 3692
rect 11425 3683 11483 3689
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 13173 3723 13231 3729
rect 13173 3689 13185 3723
rect 13219 3720 13231 3723
rect 13630 3720 13636 3732
rect 13219 3692 13636 3720
rect 13219 3689 13231 3692
rect 13173 3683 13231 3689
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 15470 3680 15476 3732
rect 15528 3720 15534 3732
rect 15565 3723 15623 3729
rect 15565 3720 15577 3723
rect 15528 3692 15577 3720
rect 15528 3680 15534 3692
rect 15565 3689 15577 3692
rect 15611 3689 15623 3723
rect 15565 3683 15623 3689
rect 16666 3680 16672 3732
rect 16724 3720 16730 3732
rect 16761 3723 16819 3729
rect 16761 3720 16773 3723
rect 16724 3692 16773 3720
rect 16724 3680 16730 3692
rect 16761 3689 16773 3692
rect 16807 3689 16819 3723
rect 17954 3720 17960 3732
rect 17915 3692 17960 3720
rect 16761 3683 16819 3689
rect 17954 3680 17960 3692
rect 18012 3680 18018 3732
rect 19245 3723 19303 3729
rect 19245 3689 19257 3723
rect 19291 3720 19303 3723
rect 19334 3720 19340 3732
rect 19291 3692 19340 3720
rect 19291 3689 19303 3692
rect 19245 3683 19303 3689
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 20438 3680 20444 3732
rect 20496 3720 20502 3732
rect 21269 3723 21327 3729
rect 21269 3720 21281 3723
rect 20496 3692 21281 3720
rect 20496 3680 20502 3692
rect 21269 3689 21281 3692
rect 21315 3689 21327 3723
rect 21269 3683 21327 3689
rect 11609 3655 11667 3661
rect 11609 3621 11621 3655
rect 11655 3652 11667 3655
rect 16206 3652 16212 3664
rect 11655 3624 12434 3652
rect 11655 3621 11667 3624
rect 11609 3615 11667 3621
rect 10778 3584 10784 3596
rect 10612 3556 10784 3584
rect 9401 3547 9459 3553
rect 10778 3544 10784 3556
rect 10836 3584 10842 3596
rect 12406 3584 12434 3624
rect 14384 3624 16212 3652
rect 13170 3584 13176 3596
rect 10836 3556 11284 3584
rect 12406 3556 13176 3584
rect 10836 3544 10842 3556
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 2498 3516 2504 3528
rect 2459 3488 2504 3516
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 5534 3525 5540 3528
rect 5528 3516 5540 3525
rect 5495 3488 5540 3516
rect 5528 3479 5540 3488
rect 5534 3476 5540 3479
rect 5592 3476 5598 3528
rect 9668 3519 9726 3525
rect 9668 3485 9680 3519
rect 9714 3516 9726 3519
rect 10870 3516 10876 3528
rect 9714 3488 10876 3516
rect 9714 3485 9726 3488
rect 9668 3479 9726 3485
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 11256 3525 11284 3556
rect 13170 3544 13176 3556
rect 13228 3544 13234 3596
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 14384 3593 14412 3624
rect 16206 3612 16212 3624
rect 16264 3612 16270 3664
rect 21284 3652 21312 3683
rect 21542 3680 21548 3732
rect 21600 3720 21606 3732
rect 22833 3723 22891 3729
rect 22833 3720 22845 3723
rect 21600 3692 22845 3720
rect 21600 3680 21606 3692
rect 22833 3689 22845 3692
rect 22879 3689 22891 3723
rect 22833 3683 22891 3689
rect 22922 3652 22928 3664
rect 21284 3624 22928 3652
rect 22922 3612 22928 3624
rect 22980 3612 22986 3664
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 13780 3556 14105 3584
rect 13780 3544 13786 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 14369 3587 14427 3593
rect 14369 3553 14381 3587
rect 14415 3553 14427 3587
rect 14369 3547 14427 3553
rect 16117 3587 16175 3593
rect 16117 3553 16129 3587
rect 16163 3584 16175 3587
rect 17218 3584 17224 3596
rect 16163 3556 17224 3584
rect 16163 3553 16175 3556
rect 16117 3547 16175 3553
rect 17218 3544 17224 3556
rect 17276 3584 17282 3596
rect 17405 3587 17463 3593
rect 17405 3584 17417 3587
rect 17276 3556 17417 3584
rect 17276 3544 17282 3556
rect 17405 3553 17417 3556
rect 17451 3584 17463 3587
rect 18506 3584 18512 3596
rect 17451 3556 18512 3584
rect 17451 3553 17463 3556
rect 17405 3547 17463 3553
rect 18506 3544 18512 3556
rect 18564 3544 18570 3596
rect 20625 3587 20683 3593
rect 20625 3553 20637 3587
rect 20671 3584 20683 3587
rect 21174 3584 21180 3596
rect 20671 3556 21180 3584
rect 20671 3553 20683 3556
rect 20625 3547 20683 3553
rect 21174 3544 21180 3556
rect 21232 3544 21238 3596
rect 21450 3584 21456 3596
rect 21411 3556 21456 3584
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 11241 3519 11299 3525
rect 11241 3485 11253 3519
rect 11287 3485 11299 3519
rect 11241 3479 11299 3485
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 11882 3516 11888 3528
rect 11379 3488 11888 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 2685 3451 2743 3457
rect 2685 3417 2697 3451
rect 2731 3448 2743 3451
rect 2866 3448 2872 3460
rect 2731 3420 2872 3448
rect 2731 3417 2743 3420
rect 2685 3411 2743 3417
rect 2866 3408 2872 3420
rect 2924 3408 2930 3460
rect 4246 3408 4252 3460
rect 4304 3448 4310 3460
rect 4341 3451 4399 3457
rect 4341 3448 4353 3451
rect 4304 3420 4353 3448
rect 4304 3408 4310 3420
rect 4341 3417 4353 3420
rect 4387 3417 4399 3451
rect 4341 3411 4399 3417
rect 9582 3408 9588 3460
rect 9640 3448 9646 3460
rect 11348 3448 11376 3479
rect 11882 3476 11888 3488
rect 11940 3516 11946 3528
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 11940 3488 12081 3516
rect 11940 3476 11946 3488
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 12492 3488 12541 3516
rect 12492 3476 12498 3488
rect 12529 3485 12541 3488
rect 12575 3485 12587 3519
rect 12529 3479 12587 3485
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3516 12955 3519
rect 12986 3516 12992 3528
rect 12943 3488 12992 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 16482 3516 16488 3528
rect 15979 3488 16488 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 20369 3519 20427 3525
rect 20369 3485 20381 3519
rect 20415 3516 20427 3519
rect 20898 3516 20904 3528
rect 20415 3488 20904 3516
rect 20415 3485 20427 3488
rect 20369 3479 20427 3485
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 21140 3488 21281 3516
rect 21140 3476 21146 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 22373 3519 22431 3525
rect 22373 3516 22385 3519
rect 21269 3479 21327 3485
rect 21376 3488 22385 3516
rect 9640 3420 11376 3448
rect 9640 3408 9646 3420
rect 11514 3408 11520 3460
rect 11572 3448 11578 3460
rect 13262 3448 13268 3460
rect 11572 3420 13268 3448
rect 11572 3408 11578 3420
rect 13262 3408 13268 3420
rect 13320 3408 13326 3460
rect 16025 3451 16083 3457
rect 16025 3417 16037 3451
rect 16071 3448 16083 3451
rect 16758 3448 16764 3460
rect 16071 3420 16764 3448
rect 16071 3417 16083 3420
rect 16025 3411 16083 3417
rect 16758 3408 16764 3420
rect 16816 3408 16822 3460
rect 17954 3408 17960 3460
rect 18012 3448 18018 3460
rect 18417 3451 18475 3457
rect 18417 3448 18429 3451
rect 18012 3420 18429 3448
rect 18012 3408 18018 3420
rect 18417 3417 18429 3420
rect 18463 3448 18475 3451
rect 19242 3448 19248 3460
rect 18463 3420 19248 3448
rect 18463 3417 18475 3420
rect 18417 3411 18475 3417
rect 19242 3408 19248 3420
rect 19300 3408 19306 3460
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 21376 3448 21404 3488
rect 22373 3485 22385 3488
rect 22419 3485 22431 3519
rect 22373 3479 22431 3485
rect 22462 3476 22468 3528
rect 22520 3516 22526 3528
rect 23017 3519 23075 3525
rect 23017 3516 23029 3519
rect 22520 3488 23029 3516
rect 22520 3476 22526 3488
rect 23017 3485 23029 3488
rect 23063 3485 23075 3519
rect 23017 3479 23075 3485
rect 27890 3476 27896 3528
rect 27948 3516 27954 3528
rect 28077 3519 28135 3525
rect 28077 3516 28089 3519
rect 27948 3488 28089 3516
rect 27948 3476 27954 3488
rect 28077 3485 28089 3488
rect 28123 3485 28135 3519
rect 28077 3479 28135 3485
rect 28534 3476 28540 3528
rect 28592 3516 28598 3528
rect 28813 3519 28871 3525
rect 28813 3516 28825 3519
rect 28592 3488 28825 3516
rect 28592 3476 28598 3488
rect 28813 3485 28825 3488
rect 28859 3485 28871 3519
rect 28813 3479 28871 3485
rect 29270 3476 29276 3528
rect 29328 3516 29334 3528
rect 29733 3519 29791 3525
rect 29733 3516 29745 3519
rect 29328 3488 29745 3516
rect 29328 3476 29334 3488
rect 29733 3485 29745 3488
rect 29779 3485 29791 3519
rect 29733 3479 29791 3485
rect 19484 3420 21404 3448
rect 21729 3451 21787 3457
rect 19484 3408 19490 3420
rect 21729 3417 21741 3451
rect 21775 3448 21787 3451
rect 21818 3448 21824 3460
rect 21775 3420 21824 3448
rect 21775 3417 21787 3420
rect 21729 3411 21787 3417
rect 21818 3408 21824 3420
rect 21876 3408 21882 3460
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 12158 3380 12164 3392
rect 8168 3352 12164 3380
rect 8168 3340 8174 3352
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 17126 3380 17132 3392
rect 17087 3352 17132 3380
rect 17126 3340 17132 3352
rect 17184 3340 17190 3392
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 18322 3380 18328 3392
rect 17276 3352 17321 3380
rect 18283 3352 18328 3380
rect 17276 3340 17282 3352
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 21085 3383 21143 3389
rect 21085 3380 21097 3383
rect 20772 3352 21097 3380
rect 20772 3340 20778 3352
rect 21085 3349 21097 3352
rect 21131 3349 21143 3383
rect 21085 3343 21143 3349
rect 21266 3340 21272 3392
rect 21324 3380 21330 3392
rect 22189 3383 22247 3389
rect 22189 3380 22201 3383
rect 21324 3352 22201 3380
rect 21324 3340 21330 3352
rect 22189 3349 22201 3352
rect 22235 3349 22247 3383
rect 22189 3343 22247 3349
rect 27798 3340 27804 3392
rect 27856 3380 27862 3392
rect 27893 3383 27951 3389
rect 27893 3380 27905 3383
rect 27856 3352 27905 3380
rect 27856 3340 27862 3352
rect 27893 3349 27905 3352
rect 27939 3349 27951 3383
rect 27893 3343 27951 3349
rect 27982 3340 27988 3392
rect 28040 3380 28046 3392
rect 28629 3383 28687 3389
rect 28629 3380 28641 3383
rect 28040 3352 28641 3380
rect 28040 3340 28046 3352
rect 28629 3349 28641 3352
rect 28675 3349 28687 3383
rect 28629 3343 28687 3349
rect 29549 3383 29607 3389
rect 29549 3349 29561 3383
rect 29595 3380 29607 3383
rect 29914 3380 29920 3392
rect 29595 3352 29920 3380
rect 29595 3349 29607 3352
rect 29549 3343 29607 3349
rect 29914 3340 29920 3352
rect 29972 3340 29978 3392
rect 1104 3290 30820 3312
rect 1104 3238 10880 3290
rect 10932 3238 10944 3290
rect 10996 3238 11008 3290
rect 11060 3238 11072 3290
rect 11124 3238 11136 3290
rect 11188 3238 20811 3290
rect 20863 3238 20875 3290
rect 20927 3238 20939 3290
rect 20991 3238 21003 3290
rect 21055 3238 21067 3290
rect 21119 3238 30820 3290
rect 1104 3216 30820 3238
rect 3789 3179 3847 3185
rect 3789 3145 3801 3179
rect 3835 3176 3847 3179
rect 8665 3179 8723 3185
rect 3835 3148 8616 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 1857 3111 1915 3117
rect 1857 3077 1869 3111
rect 1903 3108 1915 3111
rect 2958 3108 2964 3120
rect 1903 3080 2964 3108
rect 1903 3077 1915 3080
rect 1857 3071 1915 3077
rect 2958 3068 2964 3080
rect 3016 3068 3022 3120
rect 3142 3108 3148 3120
rect 3103 3080 3148 3108
rect 3142 3068 3148 3080
rect 3200 3068 3206 3120
rect 4700 3111 4758 3117
rect 4700 3077 4712 3111
rect 4746 3108 4758 3111
rect 4982 3108 4988 3120
rect 4746 3080 4988 3108
rect 4746 3077 4758 3080
rect 4700 3071 4758 3077
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 2832 3012 2877 3040
rect 2832 3000 2838 3012
rect 3418 3000 3424 3052
rect 3476 3040 3482 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3476 3012 3617 3040
rect 3476 3000 3482 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4212 3012 4445 3040
rect 4212 3000 4218 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 5224 3012 5764 3040
rect 5224 3000 5230 3012
rect 5736 2904 5764 3012
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 6512 3012 6561 3040
rect 6512 3000 6518 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 8588 3049 8616 3148
rect 8665 3145 8677 3179
rect 8711 3176 8723 3179
rect 9582 3176 9588 3188
rect 8711 3148 9588 3176
rect 8711 3145 8723 3148
rect 8665 3139 8723 3145
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 9824 3148 10609 3176
rect 9824 3136 9830 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 11517 3179 11575 3185
rect 11517 3145 11529 3179
rect 11563 3176 11575 3179
rect 11606 3176 11612 3188
rect 11563 3148 11612 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 14274 3136 14280 3188
rect 14332 3176 14338 3188
rect 14461 3179 14519 3185
rect 14461 3176 14473 3179
rect 14332 3148 14473 3176
rect 14332 3136 14338 3148
rect 14461 3145 14473 3148
rect 14507 3145 14519 3179
rect 14461 3139 14519 3145
rect 15841 3179 15899 3185
rect 15841 3145 15853 3179
rect 15887 3176 15899 3179
rect 15933 3179 15991 3185
rect 15933 3176 15945 3179
rect 15887 3148 15945 3176
rect 15887 3145 15899 3148
rect 15841 3139 15899 3145
rect 15933 3145 15945 3148
rect 15979 3176 15991 3179
rect 16758 3176 16764 3188
rect 15979 3148 16764 3176
rect 15979 3145 15991 3148
rect 15933 3139 15991 3145
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 16853 3179 16911 3185
rect 16853 3145 16865 3179
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 17773 3179 17831 3185
rect 17773 3145 17785 3179
rect 17819 3176 17831 3179
rect 18046 3176 18052 3188
rect 17819 3148 18052 3176
rect 17819 3145 17831 3148
rect 17773 3139 17831 3145
rect 9484 3111 9542 3117
rect 9484 3077 9496 3111
rect 9530 3108 9542 3111
rect 9674 3108 9680 3120
rect 9530 3080 9680 3108
rect 9530 3077 9542 3080
rect 9484 3071 9542 3077
rect 9674 3068 9680 3080
rect 9732 3068 9738 3120
rect 10778 3068 10784 3120
rect 10836 3108 10842 3120
rect 11977 3111 12035 3117
rect 10836 3080 11836 3108
rect 10836 3068 10842 3080
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 7248 3012 7297 3040
rect 7248 3000 7254 3012
rect 7285 3009 7297 3012
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3009 7987 3043
rect 7929 3003 7987 3009
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3009 8631 3043
rect 9214 3040 9220 3052
rect 9175 3012 9220 3040
rect 8573 3003 8631 3009
rect 7944 2972 7972 3003
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 11698 3040 11704 3052
rect 9324 3012 11560 3040
rect 11659 3012 11704 3040
rect 9324 2972 9352 3012
rect 7944 2944 9352 2972
rect 11532 2972 11560 3012
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 11808 3040 11836 3080
rect 11977 3077 11989 3111
rect 12023 3108 12035 3111
rect 16868 3108 16896 3139
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 18141 3179 18199 3185
rect 18141 3145 18153 3179
rect 18187 3176 18199 3179
rect 18230 3176 18236 3188
rect 18187 3148 18236 3176
rect 18187 3145 18199 3148
rect 18141 3139 18199 3145
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 18322 3136 18328 3188
rect 18380 3176 18386 3188
rect 19429 3179 19487 3185
rect 19429 3176 19441 3179
rect 18380 3148 19441 3176
rect 18380 3136 18386 3148
rect 19429 3145 19441 3148
rect 19475 3145 19487 3179
rect 21266 3176 21272 3188
rect 19429 3139 19487 3145
rect 19536 3148 21272 3176
rect 12023 3080 16896 3108
rect 17313 3111 17371 3117
rect 12023 3077 12035 3080
rect 11977 3071 12035 3077
rect 17313 3077 17325 3111
rect 17359 3108 17371 3111
rect 17954 3108 17960 3120
rect 17359 3080 17960 3108
rect 17359 3077 17371 3080
rect 17313 3071 17371 3077
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 19536 3108 19564 3148
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 22094 3136 22100 3188
rect 22152 3176 22158 3188
rect 23569 3179 23627 3185
rect 23569 3176 23581 3179
rect 22152 3148 23581 3176
rect 22152 3136 22158 3148
rect 23569 3145 23581 3148
rect 23615 3145 23627 3179
rect 23569 3139 23627 3145
rect 27341 3179 27399 3185
rect 27341 3145 27353 3179
rect 27387 3176 27399 3179
rect 29365 3179 29423 3185
rect 29365 3176 29377 3179
rect 27387 3148 28304 3176
rect 27387 3145 27399 3148
rect 27341 3139 27399 3145
rect 18248 3080 19564 3108
rect 12529 3043 12587 3049
rect 12529 3040 12541 3043
rect 11808 3012 12541 3040
rect 12529 3009 12541 3012
rect 12575 3009 12587 3043
rect 12986 3040 12992 3052
rect 12947 3012 12992 3040
rect 12529 3003 12587 3009
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 13078 3000 13084 3052
rect 13136 3040 13142 3052
rect 14090 3040 14096 3052
rect 13136 3012 13181 3040
rect 14051 3012 14096 3040
rect 13136 3000 13142 3012
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 15102 3040 15108 3052
rect 14608 3012 15108 3040
rect 14608 3000 14614 3012
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 15378 3040 15384 3052
rect 15339 3012 15384 3040
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3040 16175 3043
rect 16390 3040 16396 3052
rect 16163 3012 16396 3040
rect 16163 3009 16175 3012
rect 16117 3003 16175 3009
rect 16390 3000 16396 3012
rect 16448 3000 16454 3052
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 17218 3040 17224 3052
rect 17083 3012 17224 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 18138 3000 18144 3052
rect 18196 3040 18202 3052
rect 18248 3049 18276 3080
rect 20346 3068 20352 3120
rect 20404 3108 20410 3120
rect 20441 3111 20499 3117
rect 20441 3108 20453 3111
rect 20404 3080 20453 3108
rect 20404 3068 20410 3080
rect 20441 3077 20453 3080
rect 20487 3108 20499 3111
rect 21818 3108 21824 3120
rect 20487 3080 21824 3108
rect 20487 3077 20499 3080
rect 20441 3071 20499 3077
rect 21818 3068 21824 3080
rect 21876 3068 21882 3120
rect 22370 3108 22376 3120
rect 22020 3080 22376 3108
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 18196 3012 18245 3040
rect 18196 3000 18202 3012
rect 18233 3009 18245 3012
rect 18279 3009 18291 3043
rect 19242 3040 19248 3052
rect 19203 3012 19248 3040
rect 18233 3003 18291 3009
rect 11790 2972 11796 2984
rect 11532 2944 11796 2972
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 11885 2975 11943 2981
rect 11885 2941 11897 2975
rect 11931 2972 11943 2975
rect 11931 2944 13400 2972
rect 11931 2941 11943 2944
rect 11885 2935 11943 2941
rect 5813 2907 5871 2913
rect 5813 2904 5825 2907
rect 5736 2876 5825 2904
rect 5813 2873 5825 2876
rect 5859 2873 5871 2907
rect 6730 2904 6736 2916
rect 6691 2876 6736 2904
rect 5813 2867 5871 2873
rect 6730 2864 6736 2876
rect 6788 2864 6794 2916
rect 7469 2907 7527 2913
rect 7469 2873 7481 2907
rect 7515 2904 7527 2907
rect 9030 2904 9036 2916
rect 7515 2876 9036 2904
rect 7515 2873 7527 2876
rect 7469 2867 7527 2873
rect 9030 2864 9036 2876
rect 9088 2864 9094 2916
rect 13372 2904 13400 2944
rect 13630 2932 13636 2984
rect 13688 2972 13694 2984
rect 13817 2975 13875 2981
rect 13817 2972 13829 2975
rect 13688 2944 13829 2972
rect 13688 2932 13694 2944
rect 13817 2941 13829 2944
rect 13863 2941 13875 2975
rect 13817 2935 13875 2941
rect 13998 2932 14004 2984
rect 14056 2972 14062 2984
rect 15194 2972 15200 2984
rect 14056 2944 15200 2972
rect 14056 2932 14062 2944
rect 15194 2932 15200 2944
rect 15252 2932 15258 2984
rect 15289 2975 15347 2981
rect 15289 2941 15301 2975
rect 15335 2972 15347 2975
rect 15841 2975 15899 2981
rect 15841 2972 15853 2975
rect 15335 2944 15853 2972
rect 15335 2941 15347 2944
rect 15289 2935 15347 2941
rect 15841 2941 15853 2944
rect 15887 2941 15899 2975
rect 15841 2935 15899 2941
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2972 17187 2975
rect 18248 2972 18276 3003
rect 19242 3000 19248 3012
rect 19300 3040 19306 3052
rect 20257 3043 20315 3049
rect 20257 3040 20269 3043
rect 19300 3012 20269 3040
rect 19300 3000 19306 3012
rect 20257 3009 20269 3012
rect 20303 3009 20315 3043
rect 20622 3040 20628 3052
rect 20583 3012 20628 3040
rect 20257 3003 20315 3009
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 20717 3043 20775 3049
rect 20717 3009 20729 3043
rect 20763 3040 20775 3043
rect 21174 3040 21180 3052
rect 20763 3012 21180 3040
rect 20763 3009 20775 3012
rect 20717 3003 20775 3009
rect 21174 3000 21180 3012
rect 21232 3000 21238 3052
rect 21910 3040 21916 3052
rect 21284 3012 21916 3040
rect 17175 2944 18276 2972
rect 18325 2975 18383 2981
rect 17175 2941 17187 2944
rect 17129 2935 17187 2941
rect 18325 2941 18337 2975
rect 18371 2972 18383 2975
rect 18506 2972 18512 2984
rect 18371 2944 18512 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 18506 2932 18512 2944
rect 18564 2932 18570 2984
rect 18966 2972 18972 2984
rect 18927 2944 18972 2972
rect 18966 2932 18972 2944
rect 19024 2932 19030 2984
rect 21284 2972 21312 3012
rect 21910 3000 21916 3012
rect 21968 3000 21974 3052
rect 22020 3049 22048 3080
rect 22370 3068 22376 3080
rect 22428 3108 22434 3120
rect 25038 3108 25044 3120
rect 22428 3080 25044 3108
rect 22428 3068 22434 3080
rect 25038 3068 25044 3080
rect 25096 3068 25102 3120
rect 27801 3111 27859 3117
rect 27801 3077 27813 3111
rect 27847 3108 27859 3111
rect 27982 3108 27988 3120
rect 27847 3080 27988 3108
rect 27847 3077 27859 3080
rect 27801 3071 27859 3077
rect 27982 3068 27988 3080
rect 28040 3068 28046 3120
rect 28276 3117 28304 3148
rect 28460 3148 29377 3176
rect 28460 3117 28488 3148
rect 29365 3145 29377 3148
rect 29411 3145 29423 3179
rect 29365 3139 29423 3145
rect 28261 3111 28319 3117
rect 28261 3077 28273 3111
rect 28307 3077 28319 3111
rect 28261 3071 28319 3077
rect 28445 3111 28503 3117
rect 28445 3077 28457 3111
rect 28491 3077 28503 3111
rect 28445 3071 28503 3077
rect 22005 3043 22063 3049
rect 22005 3009 22017 3043
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 22094 3000 22100 3052
rect 22152 3040 22158 3052
rect 22465 3043 22523 3049
rect 22152 3012 22197 3040
rect 22152 3000 22158 3012
rect 22465 3009 22477 3043
rect 22511 3040 22523 3043
rect 22554 3040 22560 3052
rect 22511 3012 22560 3040
rect 22511 3009 22523 3012
rect 22465 3003 22523 3009
rect 22554 3000 22560 3012
rect 22612 3000 22618 3052
rect 23109 3043 23167 3049
rect 23109 3009 23121 3043
rect 23155 3009 23167 3043
rect 23109 3003 23167 3009
rect 19306 2944 21312 2972
rect 14921 2907 14979 2913
rect 14921 2904 14933 2907
rect 10152 2876 11744 2904
rect 13372 2876 14933 2904
rect 2133 2839 2191 2845
rect 2133 2805 2145 2839
rect 2179 2836 2191 2839
rect 7098 2836 7104 2848
rect 2179 2808 7104 2836
rect 2179 2805 2191 2808
rect 2133 2799 2191 2805
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 8110 2836 8116 2848
rect 8071 2808 8116 2836
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 8754 2796 8760 2848
rect 8812 2836 8818 2848
rect 10152 2836 10180 2876
rect 11716 2845 11744 2876
rect 14921 2873 14933 2876
rect 14967 2873 14979 2907
rect 19306 2904 19334 2944
rect 21726 2932 21732 2984
rect 21784 2972 21790 2984
rect 23124 2972 23152 3003
rect 23198 3000 23204 3052
rect 23256 3040 23262 3052
rect 23753 3043 23811 3049
rect 23753 3040 23765 3043
rect 23256 3012 23765 3040
rect 23256 3000 23262 3012
rect 23753 3009 23765 3012
rect 23799 3009 23811 3043
rect 23753 3003 23811 3009
rect 27154 3000 27160 3052
rect 27212 3040 27218 3052
rect 27525 3043 27583 3049
rect 27525 3040 27537 3043
rect 27212 3012 27537 3040
rect 27212 3000 27218 3012
rect 27525 3009 27537 3012
rect 27571 3009 27583 3043
rect 29546 3040 29552 3052
rect 29507 3012 29552 3040
rect 27525 3003 27583 3009
rect 29546 3000 29552 3012
rect 29604 3000 29610 3052
rect 29914 3040 29920 3052
rect 29875 3012 29920 3040
rect 29914 3000 29920 3012
rect 29972 3000 29978 3052
rect 30006 3000 30012 3052
rect 30064 3040 30070 3052
rect 30064 3012 30109 3040
rect 30064 3000 30070 3012
rect 27614 2972 27620 2984
rect 21784 2944 23152 2972
rect 27575 2944 27620 2972
rect 21784 2932 21790 2944
rect 27614 2932 27620 2944
rect 27672 2932 27678 2984
rect 14921 2867 14979 2873
rect 15028 2876 19334 2904
rect 20257 2907 20315 2913
rect 8812 2808 10180 2836
rect 11701 2839 11759 2845
rect 8812 2796 8818 2808
rect 11701 2805 11713 2839
rect 11747 2805 11759 2839
rect 11701 2799 11759 2805
rect 12986 2796 12992 2848
rect 13044 2836 13050 2848
rect 15028 2836 15056 2876
rect 20257 2873 20269 2907
rect 20303 2904 20315 2907
rect 22002 2904 22008 2916
rect 20303 2876 22008 2904
rect 20303 2873 20315 2876
rect 20257 2867 20315 2873
rect 22002 2864 22008 2876
rect 22060 2864 22066 2916
rect 24394 2904 24400 2916
rect 22296 2876 24400 2904
rect 22296 2848 22324 2876
rect 24394 2864 24400 2876
rect 24452 2864 24458 2916
rect 15194 2836 15200 2848
rect 13044 2808 15056 2836
rect 15155 2808 15200 2836
rect 13044 2796 13050 2808
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 17310 2836 17316 2848
rect 17271 2808 17316 2836
rect 17310 2796 17316 2808
rect 17368 2836 17374 2848
rect 17678 2836 17684 2848
rect 17368 2808 17684 2836
rect 17368 2796 17374 2808
rect 17678 2796 17684 2808
rect 17736 2796 17742 2848
rect 18138 2796 18144 2848
rect 18196 2836 18202 2848
rect 18690 2836 18696 2848
rect 18196 2808 18696 2836
rect 18196 2796 18202 2808
rect 18690 2796 18696 2808
rect 18748 2836 18754 2848
rect 19061 2839 19119 2845
rect 19061 2836 19073 2839
rect 18748 2808 19073 2836
rect 18748 2796 18754 2808
rect 19061 2805 19073 2808
rect 19107 2805 19119 2839
rect 20438 2836 20444 2848
rect 20399 2808 20444 2836
rect 19061 2799 19119 2805
rect 20438 2796 20444 2808
rect 20496 2796 20502 2848
rect 20901 2839 20959 2845
rect 20901 2805 20913 2839
rect 20947 2836 20959 2839
rect 21082 2836 21088 2848
rect 20947 2808 21088 2836
rect 20947 2805 20959 2808
rect 20901 2799 20959 2805
rect 21082 2796 21088 2808
rect 21140 2796 21146 2848
rect 21174 2796 21180 2848
rect 21232 2836 21238 2848
rect 21821 2839 21879 2845
rect 21821 2836 21833 2839
rect 21232 2808 21833 2836
rect 21232 2796 21238 2808
rect 21821 2805 21833 2808
rect 21867 2805 21879 2839
rect 22278 2836 22284 2848
rect 22239 2808 22284 2836
rect 21821 2799 21879 2805
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 22922 2836 22928 2848
rect 22883 2808 22928 2836
rect 22922 2796 22928 2808
rect 22980 2796 22986 2848
rect 27798 2836 27804 2848
rect 27759 2808 27804 2836
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 28626 2836 28632 2848
rect 28587 2808 28632 2836
rect 28626 2796 28632 2808
rect 28684 2796 28690 2848
rect 29638 2836 29644 2848
rect 29599 2808 29644 2836
rect 29638 2796 29644 2808
rect 29696 2796 29702 2848
rect 30834 2796 30840 2848
rect 30892 2836 30898 2848
rect 30929 2839 30987 2845
rect 30929 2836 30941 2839
rect 30892 2808 30941 2836
rect 30892 2796 30898 2808
rect 30929 2805 30941 2808
rect 30975 2805 30987 2839
rect 30929 2799 30987 2805
rect 1104 2746 30820 2768
rect 1104 2694 5915 2746
rect 5967 2694 5979 2746
rect 6031 2694 6043 2746
rect 6095 2694 6107 2746
rect 6159 2694 6171 2746
rect 6223 2694 15846 2746
rect 15898 2694 15910 2746
rect 15962 2694 15974 2746
rect 16026 2694 16038 2746
rect 16090 2694 16102 2746
rect 16154 2694 25776 2746
rect 25828 2694 25840 2746
rect 25892 2694 25904 2746
rect 25956 2694 25968 2746
rect 26020 2694 26032 2746
rect 26084 2694 30820 2746
rect 1104 2672 30820 2694
rect 2866 2632 2872 2644
rect 2827 2604 2872 2632
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 4433 2635 4491 2641
rect 4433 2601 4445 2635
rect 4479 2632 4491 2635
rect 6822 2632 6828 2644
rect 4479 2604 6828 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 7653 2635 7711 2641
rect 7653 2601 7665 2635
rect 7699 2632 7711 2635
rect 8754 2632 8760 2644
rect 7699 2604 8760 2632
rect 7699 2601 7711 2604
rect 7653 2595 7711 2601
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 11698 2632 11704 2644
rect 9171 2604 11704 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 14090 2632 14096 2644
rect 14051 2604 14096 2632
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 15010 2632 15016 2644
rect 14971 2604 15016 2632
rect 15010 2592 15016 2604
rect 15068 2592 15074 2644
rect 15378 2592 15384 2644
rect 15436 2632 15442 2644
rect 15933 2635 15991 2641
rect 15933 2632 15945 2635
rect 15436 2604 15945 2632
rect 15436 2592 15442 2604
rect 15933 2601 15945 2604
rect 15979 2601 15991 2635
rect 15933 2595 15991 2601
rect 17126 2592 17132 2644
rect 17184 2632 17190 2644
rect 17589 2635 17647 2641
rect 17589 2632 17601 2635
rect 17184 2604 17601 2632
rect 17184 2592 17190 2604
rect 17589 2601 17601 2604
rect 17635 2601 17647 2635
rect 17589 2595 17647 2601
rect 17678 2592 17684 2644
rect 17736 2632 17742 2644
rect 18509 2635 18567 2641
rect 18509 2632 18521 2635
rect 17736 2604 18521 2632
rect 17736 2592 17742 2604
rect 18509 2601 18521 2604
rect 18555 2601 18567 2635
rect 18509 2595 18567 2601
rect 20441 2635 20499 2641
rect 20441 2601 20453 2635
rect 20487 2632 20499 2635
rect 20714 2632 20720 2644
rect 20487 2604 20720 2632
rect 20487 2601 20499 2604
rect 20441 2595 20499 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 21082 2632 21088 2644
rect 21043 2604 21088 2632
rect 21082 2592 21088 2604
rect 21140 2592 21146 2644
rect 21910 2632 21916 2644
rect 21871 2604 21916 2632
rect 21910 2592 21916 2604
rect 21968 2592 21974 2644
rect 22554 2592 22560 2644
rect 22612 2632 22618 2644
rect 25685 2635 25743 2641
rect 25685 2632 25697 2635
rect 22612 2604 25697 2632
rect 22612 2592 22618 2604
rect 25685 2601 25697 2604
rect 25731 2601 25743 2635
rect 27154 2632 27160 2644
rect 27115 2604 27160 2632
rect 25685 2595 25743 2601
rect 27154 2592 27160 2604
rect 27212 2592 27218 2644
rect 27614 2632 27620 2644
rect 27575 2604 27620 2632
rect 27614 2592 27620 2604
rect 27672 2592 27678 2644
rect 30006 2632 30012 2644
rect 29967 2604 30012 2632
rect 30006 2592 30012 2604
rect 30064 2592 30070 2644
rect 6549 2567 6607 2573
rect 6549 2533 6561 2567
rect 6595 2564 6607 2567
rect 8570 2564 8576 2576
rect 6595 2536 8576 2564
rect 6595 2533 6607 2536
rect 6549 2527 6607 2533
rect 8570 2524 8576 2536
rect 8628 2524 8634 2576
rect 11422 2564 11428 2576
rect 9784 2536 11428 2564
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2496 2283 2499
rect 2498 2496 2504 2508
rect 2271 2468 2504 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 8389 2499 8447 2505
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 9784 2496 9812 2536
rect 11422 2524 11428 2536
rect 11480 2524 11486 2576
rect 14461 2567 14519 2573
rect 14461 2533 14473 2567
rect 14507 2564 14519 2567
rect 15286 2564 15292 2576
rect 14507 2536 15292 2564
rect 14507 2533 14519 2536
rect 14461 2527 14519 2533
rect 15286 2524 15292 2536
rect 15344 2564 15350 2576
rect 16761 2567 16819 2573
rect 16761 2564 16773 2567
rect 15344 2536 16773 2564
rect 15344 2524 15350 2536
rect 16761 2533 16773 2536
rect 16807 2533 16819 2567
rect 16761 2527 16819 2533
rect 17218 2524 17224 2576
rect 17276 2564 17282 2576
rect 19245 2567 19303 2573
rect 19245 2564 19257 2567
rect 17276 2536 19257 2564
rect 17276 2524 17282 2536
rect 8435 2468 9812 2496
rect 9861 2499 9919 2505
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 9950 2496 9956 2508
rect 9907 2468 9956 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 9950 2456 9956 2468
rect 10008 2456 10014 2508
rect 11793 2499 11851 2505
rect 11793 2465 11805 2499
rect 11839 2496 11851 2499
rect 11974 2496 11980 2508
rect 11839 2468 11980 2496
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 14553 2499 14611 2505
rect 14553 2465 14565 2499
rect 14599 2496 14611 2499
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 14599 2468 15485 2496
rect 14599 2465 14611 2468
rect 14553 2459 14611 2465
rect 15473 2465 15485 2468
rect 15519 2496 15531 2499
rect 16206 2496 16212 2508
rect 15519 2468 16212 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 16206 2456 16212 2468
rect 16264 2496 16270 2508
rect 16669 2499 16727 2505
rect 16669 2496 16681 2499
rect 16264 2468 16681 2496
rect 16264 2456 16270 2468
rect 16669 2465 16681 2468
rect 16715 2465 16727 2499
rect 16669 2459 16727 2465
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 17092 2468 17141 2496
rect 17092 2456 17098 2468
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 1854 2388 1860 2440
rect 1912 2428 1918 2440
rect 1949 2431 2007 2437
rect 1949 2428 1961 2431
rect 1912 2400 1961 2428
rect 1912 2388 1918 2400
rect 1949 2397 1961 2400
rect 1995 2397 2007 2431
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 1949 2391 2007 2397
rect 2056 2400 3065 2428
rect 382 2320 388 2372
rect 440 2360 446 2372
rect 2056 2360 2084 2400
rect 3053 2397 3065 2400
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 4890 2388 4896 2440
rect 4948 2428 4954 2440
rect 4985 2431 5043 2437
rect 4985 2428 4997 2431
rect 4948 2400 4997 2428
rect 4948 2388 4954 2400
rect 4985 2397 4997 2400
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 440 2332 2084 2360
rect 440 2320 446 2332
rect 2774 2320 2780 2372
rect 2832 2360 2838 2372
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 2832 2332 4169 2360
rect 2832 2320 2838 2332
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 5276 2360 5304 2391
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5776 2400 6377 2428
rect 5776 2388 5782 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7926 2428 7932 2440
rect 7515 2400 7932 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 8662 2428 8668 2440
rect 8036 2400 8668 2428
rect 8036 2360 8064 2400
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8812 2400 8953 2428
rect 8812 2388 8818 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9490 2388 9496 2440
rect 9548 2428 9554 2440
rect 9585 2431 9643 2437
rect 9585 2428 9597 2431
rect 9548 2400 9597 2428
rect 9548 2388 9554 2400
rect 9585 2397 9597 2400
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 10284 2400 11529 2428
rect 10284 2388 10290 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2428 13415 2431
rect 13722 2428 13728 2440
rect 13403 2400 13728 2428
rect 13403 2397 13415 2400
rect 13357 2391 13415 2397
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14056 2400 14289 2428
rect 14056 2388 14062 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 15102 2388 15108 2440
rect 15160 2428 15166 2440
rect 15197 2431 15255 2437
rect 15197 2428 15209 2431
rect 15160 2400 15209 2428
rect 15160 2388 15166 2400
rect 15197 2397 15209 2400
rect 15243 2397 15255 2431
rect 15197 2391 15255 2397
rect 15286 2388 15292 2440
rect 15344 2428 15350 2440
rect 15381 2431 15439 2437
rect 15381 2428 15393 2431
rect 15344 2400 15393 2428
rect 15344 2388 15350 2400
rect 15381 2397 15393 2400
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 15620 2400 16129 2428
rect 15620 2388 15626 2400
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2428 17003 2431
rect 17678 2428 17684 2440
rect 16991 2400 17684 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 17788 2437 17816 2536
rect 19245 2533 19257 2536
rect 19291 2533 19303 2567
rect 19245 2527 19303 2533
rect 20254 2524 20260 2576
rect 20312 2564 20318 2576
rect 24394 2564 24400 2576
rect 20312 2536 23520 2564
rect 24355 2536 24400 2564
rect 20312 2524 20318 2536
rect 17862 2456 17868 2508
rect 17920 2496 17926 2508
rect 20349 2499 20407 2505
rect 17920 2468 19472 2496
rect 17920 2456 17926 2468
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2397 17831 2431
rect 17954 2428 17960 2440
rect 17915 2400 17960 2428
rect 17773 2391 17831 2397
rect 17954 2388 17960 2400
rect 18012 2388 18018 2440
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2397 18107 2431
rect 18690 2428 18696 2440
rect 18651 2400 18696 2428
rect 18049 2391 18107 2397
rect 5276 2332 8064 2360
rect 8205 2363 8263 2369
rect 4157 2323 4215 2329
rect 8205 2329 8217 2363
rect 8251 2360 8263 2363
rect 9398 2360 9404 2372
rect 8251 2332 9404 2360
rect 8251 2329 8263 2332
rect 8205 2323 8263 2329
rect 9398 2320 9404 2332
rect 9456 2320 9462 2372
rect 13541 2363 13599 2369
rect 13541 2329 13553 2363
rect 13587 2360 13599 2363
rect 14366 2360 14372 2372
rect 13587 2332 14372 2360
rect 13587 2329 13599 2332
rect 13541 2323 13599 2329
rect 14366 2320 14372 2332
rect 14424 2360 14430 2372
rect 18064 2360 18092 2391
rect 18690 2388 18696 2400
rect 18748 2388 18754 2440
rect 19444 2437 19472 2468
rect 20349 2465 20361 2499
rect 20395 2496 20407 2499
rect 21174 2496 21180 2508
rect 20395 2468 21180 2496
rect 20395 2465 20407 2468
rect 20349 2459 20407 2465
rect 21174 2456 21180 2468
rect 21232 2456 21238 2508
rect 21818 2456 21824 2508
rect 21876 2496 21882 2508
rect 23290 2496 23296 2508
rect 21876 2468 23296 2496
rect 21876 2456 21882 2468
rect 23290 2456 23296 2468
rect 23348 2456 23354 2508
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 20441 2431 20499 2437
rect 20441 2397 20453 2431
rect 20487 2428 20499 2431
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 20487 2400 21281 2428
rect 20487 2397 20499 2400
rect 20441 2391 20499 2397
rect 21269 2397 21281 2400
rect 21315 2428 21327 2431
rect 21315 2400 22232 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 18966 2360 18972 2372
rect 14424 2332 18972 2360
rect 14424 2320 14430 2332
rect 18966 2320 18972 2332
rect 19024 2320 19030 2372
rect 22204 2369 22232 2400
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 22646 2428 22652 2440
rect 22336 2400 22652 2428
rect 22336 2388 22342 2400
rect 22646 2388 22652 2400
rect 22704 2388 22710 2440
rect 22830 2428 22836 2440
rect 22791 2400 22836 2428
rect 22830 2388 22836 2400
rect 22888 2388 22894 2440
rect 23492 2437 23520 2536
rect 24394 2524 24400 2536
rect 24452 2524 24458 2576
rect 25038 2564 25044 2576
rect 24999 2536 25044 2564
rect 25038 2524 25044 2536
rect 25096 2524 25102 2576
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 23934 2388 23940 2440
rect 23992 2428 23998 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23992 2400 24593 2428
rect 23992 2388 23998 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 24762 2388 24768 2440
rect 24820 2428 24826 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 24820 2400 25237 2428
rect 24820 2388 24826 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 25498 2388 25504 2440
rect 25556 2428 25562 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 25556 2400 25881 2428
rect 25556 2388 25562 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 26234 2388 26240 2440
rect 26292 2428 26298 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26292 2400 26985 2428
rect 26292 2388 26298 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27120 2400 27813 2428
rect 27120 2388 27126 2400
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 28718 2428 28724 2440
rect 28679 2400 28724 2428
rect 27801 2391 27859 2397
rect 28718 2388 28724 2400
rect 28776 2388 28782 2440
rect 29086 2388 29092 2440
rect 29144 2428 29150 2440
rect 29825 2431 29883 2437
rect 29825 2428 29837 2431
rect 29144 2400 29837 2428
rect 29144 2388 29150 2400
rect 29825 2397 29837 2400
rect 29871 2397 29883 2431
rect 29825 2391 29883 2397
rect 22005 2363 22063 2369
rect 22005 2329 22017 2363
rect 22051 2329 22063 2363
rect 22005 2323 22063 2329
rect 22189 2363 22247 2369
rect 22189 2329 22201 2363
rect 22235 2360 22247 2363
rect 28626 2360 28632 2372
rect 22235 2332 28632 2360
rect 22235 2329 22247 2332
rect 22189 2323 22247 2329
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 16850 2292 16856 2304
rect 12124 2264 16856 2292
rect 12124 2252 12130 2264
rect 16850 2252 16856 2264
rect 16908 2252 16914 2304
rect 18322 2252 18328 2304
rect 18380 2292 18386 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 18380 2264 20085 2292
rect 18380 2252 18386 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 20162 2252 20168 2304
rect 20220 2292 20226 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20220 2264 20913 2292
rect 20220 2252 20226 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 22020 2292 22048 2323
rect 28626 2320 28632 2332
rect 28684 2320 28690 2372
rect 22554 2292 22560 2304
rect 22020 2264 22560 2292
rect 20901 2255 20959 2261
rect 22554 2252 22560 2264
rect 22612 2252 22618 2304
rect 22646 2252 22652 2304
rect 22704 2292 22710 2304
rect 23290 2292 23296 2304
rect 22704 2264 22749 2292
rect 23251 2264 23296 2292
rect 22704 2252 22710 2264
rect 23290 2252 23296 2264
rect 23348 2252 23354 2304
rect 28902 2292 28908 2304
rect 28863 2264 28908 2292
rect 28902 2252 28908 2264
rect 28960 2252 28966 2304
rect 1104 2202 30820 2224
rect 1104 2150 10880 2202
rect 10932 2150 10944 2202
rect 10996 2150 11008 2202
rect 11060 2150 11072 2202
rect 11124 2150 11136 2202
rect 11188 2150 20811 2202
rect 20863 2150 20875 2202
rect 20927 2150 20939 2202
rect 20991 2150 21003 2202
rect 21055 2150 21067 2202
rect 21119 2150 30820 2202
rect 1104 2128 30820 2150
rect 16850 2048 16856 2100
rect 16908 2088 16914 2100
rect 18322 2088 18328 2100
rect 16908 2060 18328 2088
rect 16908 2048 16914 2060
rect 18322 2048 18328 2060
rect 18380 2048 18386 2100
rect 18598 2048 18604 2100
rect 18656 2088 18662 2100
rect 22830 2088 22836 2100
rect 18656 2060 22836 2088
rect 18656 2048 18662 2060
rect 22830 2048 22836 2060
rect 22888 2048 22894 2100
rect 13078 1912 13084 1964
rect 13136 1952 13142 1964
rect 20162 1952 20168 1964
rect 13136 1924 20168 1952
rect 13136 1912 13142 1924
rect 20162 1912 20168 1924
rect 20220 1912 20226 1964
rect 9398 1368 9404 1420
rect 9456 1408 9462 1420
rect 11054 1408 11060 1420
rect 9456 1380 11060 1408
rect 9456 1368 9462 1380
rect 11054 1368 11060 1380
rect 11112 1368 11118 1420
rect 17126 1368 17132 1420
rect 17184 1408 17190 1420
rect 18690 1408 18696 1420
rect 17184 1380 18696 1408
rect 17184 1368 17190 1380
rect 18690 1368 18696 1380
rect 18748 1368 18754 1420
<< via1 >>
rect 10880 45670 10932 45722
rect 10944 45670 10996 45722
rect 11008 45670 11060 45722
rect 11072 45670 11124 45722
rect 11136 45670 11188 45722
rect 20811 45670 20863 45722
rect 20875 45670 20927 45722
rect 20939 45670 20991 45722
rect 21003 45670 21055 45722
rect 21067 45670 21119 45722
rect 1676 45475 1728 45484
rect 1676 45441 1685 45475
rect 1685 45441 1719 45475
rect 1719 45441 1728 45475
rect 1676 45432 1728 45441
rect 4528 45432 4580 45484
rect 4896 45432 4948 45484
rect 5448 45432 5500 45484
rect 6460 45475 6512 45484
rect 6460 45441 6469 45475
rect 6469 45441 6503 45475
rect 6503 45441 6512 45475
rect 6460 45432 6512 45441
rect 7288 45475 7340 45484
rect 7288 45441 7297 45475
rect 7297 45441 7331 45475
rect 7331 45441 7340 45475
rect 7288 45432 7340 45441
rect 30104 45475 30156 45484
rect 30104 45441 30113 45475
rect 30113 45441 30147 45475
rect 30147 45441 30156 45475
rect 30104 45432 30156 45441
rect 2228 45339 2280 45348
rect 2228 45305 2237 45339
rect 2237 45305 2271 45339
rect 2271 45305 2280 45339
rect 2228 45296 2280 45305
rect 2964 45339 3016 45348
rect 2964 45305 2973 45339
rect 2973 45305 3007 45339
rect 3007 45305 3016 45339
rect 2964 45296 3016 45305
rect 2780 45228 2832 45280
rect 3792 45271 3844 45280
rect 3792 45237 3801 45271
rect 3801 45237 3835 45271
rect 3835 45237 3844 45271
rect 3792 45228 3844 45237
rect 4436 45271 4488 45280
rect 4436 45237 4445 45271
rect 4445 45237 4479 45271
rect 4479 45237 4488 45271
rect 4436 45228 4488 45237
rect 6736 45228 6788 45280
rect 29000 45228 29052 45280
rect 5915 45126 5967 45178
rect 5979 45126 6031 45178
rect 6043 45126 6095 45178
rect 6107 45126 6159 45178
rect 6171 45126 6223 45178
rect 15846 45126 15898 45178
rect 15910 45126 15962 45178
rect 15974 45126 16026 45178
rect 16038 45126 16090 45178
rect 16102 45126 16154 45178
rect 25776 45126 25828 45178
rect 25840 45126 25892 45178
rect 25904 45126 25956 45178
rect 25968 45126 26020 45178
rect 26032 45126 26084 45178
rect 2872 45024 2924 45076
rect 4252 45024 4304 45076
rect 7288 45024 7340 45076
rect 7380 44956 7432 45008
rect 4436 44888 4488 44940
rect 2412 44863 2464 44872
rect 2412 44829 2421 44863
rect 2421 44829 2455 44863
rect 2455 44829 2464 44863
rect 2412 44820 2464 44829
rect 3148 44820 3200 44872
rect 4068 44863 4120 44872
rect 4068 44829 4077 44863
rect 4077 44829 4111 44863
rect 4111 44829 4120 44863
rect 4068 44820 4120 44829
rect 5356 44820 5408 44872
rect 5724 44863 5776 44872
rect 5724 44829 5733 44863
rect 5733 44829 5767 44863
rect 5767 44829 5776 44863
rect 5724 44820 5776 44829
rect 6644 44820 6696 44872
rect 7196 44863 7248 44872
rect 7196 44829 7205 44863
rect 7205 44829 7239 44863
rect 7239 44829 7248 44863
rect 7196 44820 7248 44829
rect 1492 44727 1544 44736
rect 1492 44693 1501 44727
rect 1501 44693 1535 44727
rect 1535 44693 1544 44727
rect 1492 44684 1544 44693
rect 2872 44727 2924 44736
rect 2872 44693 2881 44727
rect 2881 44693 2915 44727
rect 2915 44693 2924 44727
rect 2872 44684 2924 44693
rect 4252 44727 4304 44736
rect 4252 44693 4261 44727
rect 4261 44693 4295 44727
rect 4295 44693 4304 44727
rect 4252 44684 4304 44693
rect 5540 44684 5592 44736
rect 5816 44684 5868 44736
rect 6828 44727 6880 44736
rect 6828 44693 6837 44727
rect 6837 44693 6871 44727
rect 6871 44693 6880 44727
rect 6828 44684 6880 44693
rect 7472 44820 7524 44872
rect 8208 44863 8260 44872
rect 8208 44829 8217 44863
rect 8217 44829 8251 44863
rect 8251 44829 8260 44863
rect 8208 44820 8260 44829
rect 30012 44820 30064 44872
rect 7656 44684 7708 44736
rect 8024 44727 8076 44736
rect 8024 44693 8033 44727
rect 8033 44693 8067 44727
rect 8067 44693 8076 44727
rect 8024 44684 8076 44693
rect 29920 44727 29972 44736
rect 29920 44693 29929 44727
rect 29929 44693 29963 44727
rect 29963 44693 29972 44727
rect 29920 44684 29972 44693
rect 10880 44582 10932 44634
rect 10944 44582 10996 44634
rect 11008 44582 11060 44634
rect 11072 44582 11124 44634
rect 11136 44582 11188 44634
rect 20811 44582 20863 44634
rect 20875 44582 20927 44634
rect 20939 44582 20991 44634
rect 21003 44582 21055 44634
rect 21067 44582 21119 44634
rect 4436 44523 4488 44532
rect 4436 44489 4445 44523
rect 4445 44489 4479 44523
rect 4479 44489 4488 44523
rect 4436 44480 4488 44489
rect 4896 44523 4948 44532
rect 4896 44489 4905 44523
rect 4905 44489 4939 44523
rect 4939 44489 4948 44523
rect 4896 44480 4948 44489
rect 6644 44480 6696 44532
rect 3792 44412 3844 44464
rect 2320 44387 2372 44396
rect 2320 44353 2329 44387
rect 2329 44353 2363 44387
rect 2363 44353 2372 44387
rect 2320 44344 2372 44353
rect 2964 44387 3016 44396
rect 2964 44353 2973 44387
rect 2973 44353 3007 44387
rect 3007 44353 3016 44387
rect 2964 44344 3016 44353
rect 6828 44412 6880 44464
rect 7196 44412 7248 44464
rect 6736 44387 6788 44396
rect 6736 44353 6745 44387
rect 6745 44353 6779 44387
rect 6779 44353 6788 44387
rect 6736 44344 6788 44353
rect 1492 44183 1544 44192
rect 1492 44149 1501 44183
rect 1501 44149 1535 44183
rect 1535 44149 1544 44183
rect 1492 44140 1544 44149
rect 1768 44140 1820 44192
rect 3056 44140 3108 44192
rect 4252 44183 4304 44192
rect 4252 44149 4261 44183
rect 4261 44149 4295 44183
rect 4295 44149 4304 44183
rect 4252 44140 4304 44149
rect 5356 44208 5408 44260
rect 8852 44276 8904 44328
rect 9864 44344 9916 44396
rect 9496 44276 9548 44328
rect 20076 44344 20128 44396
rect 9956 44208 10008 44260
rect 5264 44140 5316 44192
rect 8576 44183 8628 44192
rect 8576 44149 8585 44183
rect 8585 44149 8619 44183
rect 8619 44149 8628 44183
rect 8576 44140 8628 44149
rect 5915 44038 5967 44090
rect 5979 44038 6031 44090
rect 6043 44038 6095 44090
rect 6107 44038 6159 44090
rect 6171 44038 6223 44090
rect 15846 44038 15898 44090
rect 15910 44038 15962 44090
rect 15974 44038 16026 44090
rect 16038 44038 16090 44090
rect 16102 44038 16154 44090
rect 25776 44038 25828 44090
rect 25840 44038 25892 44090
rect 25904 44038 25956 44090
rect 25968 44038 26020 44090
rect 26032 44038 26084 44090
rect 4068 43936 4120 43988
rect 4988 43936 5040 43988
rect 5264 43979 5316 43988
rect 5264 43945 5273 43979
rect 5273 43945 5307 43979
rect 5307 43945 5316 43979
rect 5264 43936 5316 43945
rect 5448 43979 5500 43988
rect 5448 43945 5457 43979
rect 5457 43945 5491 43979
rect 5491 43945 5500 43979
rect 5448 43936 5500 43945
rect 7656 43936 7708 43988
rect 8852 43936 8904 43988
rect 20076 43979 20128 43988
rect 20076 43945 20085 43979
rect 20085 43945 20119 43979
rect 20119 43945 20128 43979
rect 20076 43936 20128 43945
rect 3332 43868 3384 43920
rect 2872 43800 2924 43852
rect 2596 43732 2648 43784
rect 5816 43800 5868 43852
rect 3976 43775 4028 43784
rect 3976 43741 3985 43775
rect 3985 43741 4019 43775
rect 4019 43741 4028 43775
rect 3976 43732 4028 43741
rect 5356 43732 5408 43784
rect 10416 43732 10468 43784
rect 20168 43732 20220 43784
rect 29000 43800 29052 43852
rect 29920 43732 29972 43784
rect 6644 43664 6696 43716
rect 8116 43664 8168 43716
rect 9772 43664 9824 43716
rect 1492 43639 1544 43648
rect 1492 43605 1501 43639
rect 1501 43605 1535 43639
rect 1535 43605 1544 43639
rect 1492 43596 1544 43605
rect 2504 43596 2556 43648
rect 3792 43639 3844 43648
rect 3792 43605 3801 43639
rect 3801 43605 3835 43639
rect 3835 43605 3844 43639
rect 3792 43596 3844 43605
rect 6828 43596 6880 43648
rect 8024 43596 8076 43648
rect 10880 43494 10932 43546
rect 10944 43494 10996 43546
rect 11008 43494 11060 43546
rect 11072 43494 11124 43546
rect 11136 43494 11188 43546
rect 20811 43494 20863 43546
rect 20875 43494 20927 43546
rect 20939 43494 20991 43546
rect 21003 43494 21055 43546
rect 21067 43494 21119 43546
rect 5724 43392 5776 43444
rect 8116 43435 8168 43444
rect 8116 43401 8125 43435
rect 8125 43401 8159 43435
rect 8159 43401 8168 43435
rect 8116 43392 8168 43401
rect 9956 43435 10008 43444
rect 9956 43401 9965 43435
rect 9965 43401 9999 43435
rect 9999 43401 10008 43435
rect 9956 43392 10008 43401
rect 10416 43435 10468 43444
rect 10416 43401 10425 43435
rect 10425 43401 10459 43435
rect 10459 43401 10468 43435
rect 10416 43392 10468 43401
rect 5540 43324 5592 43376
rect 8024 43324 8076 43376
rect 8576 43324 8628 43376
rect 1860 43256 1912 43308
rect 2780 43299 2832 43308
rect 2780 43265 2789 43299
rect 2789 43265 2823 43299
rect 2823 43265 2832 43299
rect 3608 43299 3660 43308
rect 2780 43256 2832 43265
rect 3608 43265 3617 43299
rect 3617 43265 3651 43299
rect 3651 43265 3660 43299
rect 3608 43256 3660 43265
rect 3884 43256 3936 43308
rect 4344 43256 4396 43308
rect 5724 43256 5776 43308
rect 7380 43299 7432 43308
rect 7380 43265 7389 43299
rect 7389 43265 7423 43299
rect 7423 43265 7432 43299
rect 7380 43256 7432 43265
rect 7012 43188 7064 43240
rect 7656 43231 7708 43240
rect 7656 43197 7665 43231
rect 7665 43197 7699 43231
rect 7699 43197 7708 43231
rect 7656 43188 7708 43197
rect 9128 43256 9180 43308
rect 30104 43299 30156 43308
rect 30104 43265 30113 43299
rect 30113 43265 30147 43299
rect 30147 43265 30156 43299
rect 30104 43256 30156 43265
rect 6460 43120 6512 43172
rect 7196 43120 7248 43172
rect 8024 43188 8076 43240
rect 8576 43231 8628 43240
rect 8576 43197 8585 43231
rect 8585 43197 8619 43231
rect 8619 43197 8628 43231
rect 8576 43188 8628 43197
rect 1400 43052 1452 43104
rect 2136 43095 2188 43104
rect 2136 43061 2145 43095
rect 2145 43061 2179 43095
rect 2179 43061 2188 43095
rect 2136 43052 2188 43061
rect 2964 43095 3016 43104
rect 2964 43061 2973 43095
rect 2973 43061 3007 43095
rect 3007 43061 3016 43095
rect 2964 43052 3016 43061
rect 3424 43095 3476 43104
rect 3424 43061 3433 43095
rect 3433 43061 3467 43095
rect 3467 43061 3476 43095
rect 3424 43052 3476 43061
rect 3516 43052 3568 43104
rect 29920 43095 29972 43104
rect 29920 43061 29929 43095
rect 29929 43061 29963 43095
rect 29963 43061 29972 43095
rect 29920 43052 29972 43061
rect 5915 42950 5967 43002
rect 5979 42950 6031 43002
rect 6043 42950 6095 43002
rect 6107 42950 6159 43002
rect 6171 42950 6223 43002
rect 15846 42950 15898 43002
rect 15910 42950 15962 43002
rect 15974 42950 16026 43002
rect 16038 42950 16090 43002
rect 16102 42950 16154 43002
rect 25776 42950 25828 43002
rect 25840 42950 25892 43002
rect 25904 42950 25956 43002
rect 25968 42950 26020 43002
rect 26032 42950 26084 43002
rect 2504 42891 2556 42900
rect 2504 42857 2513 42891
rect 2513 42857 2547 42891
rect 2547 42857 2556 42891
rect 2504 42848 2556 42857
rect 5264 42848 5316 42900
rect 6644 42891 6696 42900
rect 6644 42857 6653 42891
rect 6653 42857 6687 42891
rect 6687 42857 6696 42891
rect 6644 42848 6696 42857
rect 8576 42848 8628 42900
rect 3792 42712 3844 42764
rect 7196 42780 7248 42832
rect 8024 42780 8076 42832
rect 9772 42780 9824 42832
rect 9864 42712 9916 42764
rect 2228 42644 2280 42696
rect 3700 42644 3752 42696
rect 5080 42687 5132 42696
rect 5080 42653 5089 42687
rect 5089 42653 5123 42687
rect 5123 42653 5132 42687
rect 5080 42644 5132 42653
rect 5724 42644 5776 42696
rect 6828 42687 6880 42696
rect 6828 42653 6837 42687
rect 6837 42653 6871 42687
rect 6871 42653 6880 42687
rect 6828 42644 6880 42653
rect 6736 42576 6788 42628
rect 7012 42576 7064 42628
rect 7380 42687 7432 42696
rect 7380 42653 7389 42687
rect 7389 42653 7423 42687
rect 7423 42653 7432 42687
rect 7380 42644 7432 42653
rect 9128 42687 9180 42696
rect 7656 42576 7708 42628
rect 1492 42551 1544 42560
rect 1492 42517 1501 42551
rect 1501 42517 1535 42551
rect 1535 42517 1544 42551
rect 1492 42508 1544 42517
rect 3148 42508 3200 42560
rect 3792 42551 3844 42560
rect 3792 42517 3801 42551
rect 3801 42517 3835 42551
rect 3835 42517 3844 42551
rect 3792 42508 3844 42517
rect 4528 42551 4580 42560
rect 4528 42517 4537 42551
rect 4537 42517 4571 42551
rect 4571 42517 4580 42551
rect 4528 42508 4580 42517
rect 4712 42551 4764 42560
rect 4712 42517 4721 42551
rect 4721 42517 4755 42551
rect 4755 42517 4764 42551
rect 4712 42508 4764 42517
rect 6552 42508 6604 42560
rect 9128 42653 9137 42687
rect 9137 42653 9171 42687
rect 9171 42653 9180 42687
rect 9128 42644 9180 42653
rect 29920 42644 29972 42696
rect 20168 42576 20220 42628
rect 10232 42508 10284 42560
rect 10880 42406 10932 42458
rect 10944 42406 10996 42458
rect 11008 42406 11060 42458
rect 11072 42406 11124 42458
rect 11136 42406 11188 42458
rect 20811 42406 20863 42458
rect 20875 42406 20927 42458
rect 20939 42406 20991 42458
rect 21003 42406 21055 42458
rect 21067 42406 21119 42458
rect 3056 42304 3108 42356
rect 3700 42347 3752 42356
rect 3700 42313 3709 42347
rect 3709 42313 3743 42347
rect 3743 42313 3752 42347
rect 3700 42304 3752 42313
rect 2228 42032 2280 42084
rect 3240 42168 3292 42220
rect 5724 42168 5776 42220
rect 6460 42168 6512 42220
rect 7288 42304 7340 42356
rect 7748 42168 7800 42220
rect 2688 42100 2740 42152
rect 5080 42100 5132 42152
rect 7012 42143 7064 42152
rect 7012 42109 7021 42143
rect 7021 42109 7055 42143
rect 7055 42109 7064 42143
rect 7012 42100 7064 42109
rect 7196 42100 7248 42152
rect 1400 41964 1452 42016
rect 2504 42007 2556 42016
rect 2504 41973 2513 42007
rect 2513 41973 2547 42007
rect 2547 41973 2556 42007
rect 2504 41964 2556 41973
rect 4344 41964 4396 42016
rect 4896 42007 4948 42016
rect 4896 41973 4905 42007
rect 4905 41973 4939 42007
rect 4939 41973 4948 42007
rect 4896 41964 4948 41973
rect 21916 42168 21968 42220
rect 6920 41964 6972 42016
rect 7472 42007 7524 42016
rect 7472 41973 7481 42007
rect 7481 41973 7515 42007
rect 7515 41973 7524 42007
rect 7472 41964 7524 41973
rect 8392 41964 8444 42016
rect 5915 41862 5967 41914
rect 5979 41862 6031 41914
rect 6043 41862 6095 41914
rect 6107 41862 6159 41914
rect 6171 41862 6223 41914
rect 15846 41862 15898 41914
rect 15910 41862 15962 41914
rect 15974 41862 16026 41914
rect 16038 41862 16090 41914
rect 16102 41862 16154 41914
rect 25776 41862 25828 41914
rect 25840 41862 25892 41914
rect 25904 41862 25956 41914
rect 25968 41862 26020 41914
rect 26032 41862 26084 41914
rect 2504 41803 2556 41812
rect 2504 41769 2513 41803
rect 2513 41769 2547 41803
rect 2547 41769 2556 41803
rect 2504 41760 2556 41769
rect 3976 41760 4028 41812
rect 4712 41760 4764 41812
rect 7748 41760 7800 41812
rect 3516 41624 3568 41676
rect 3792 41667 3844 41676
rect 3792 41633 3801 41667
rect 3801 41633 3835 41667
rect 3835 41633 3844 41667
rect 3792 41624 3844 41633
rect 5080 41624 5132 41676
rect 8392 41667 8444 41676
rect 8392 41633 8401 41667
rect 8401 41633 8435 41667
rect 8435 41633 8444 41667
rect 8392 41624 8444 41633
rect 2228 41556 2280 41608
rect 2688 41556 2740 41608
rect 5632 41599 5684 41608
rect 4068 41531 4120 41540
rect 4068 41497 4102 41531
rect 4102 41497 4120 41531
rect 5632 41565 5641 41599
rect 5641 41565 5675 41599
rect 5675 41565 5684 41599
rect 5632 41556 5684 41565
rect 6552 41556 6604 41608
rect 4068 41488 4120 41497
rect 6276 41488 6328 41540
rect 7472 41488 7524 41540
rect 1308 41420 1360 41472
rect 3792 41420 3844 41472
rect 7656 41420 7708 41472
rect 10232 41488 10284 41540
rect 8944 41463 8996 41472
rect 8944 41429 8953 41463
rect 8953 41429 8987 41463
rect 8987 41429 8996 41463
rect 8944 41420 8996 41429
rect 10880 41318 10932 41370
rect 10944 41318 10996 41370
rect 11008 41318 11060 41370
rect 11072 41318 11124 41370
rect 11136 41318 11188 41370
rect 20811 41318 20863 41370
rect 20875 41318 20927 41370
rect 20939 41318 20991 41370
rect 21003 41318 21055 41370
rect 21067 41318 21119 41370
rect 3884 41216 3936 41268
rect 4068 41216 4120 41268
rect 6736 41259 6788 41268
rect 6736 41225 6745 41259
rect 6745 41225 6779 41259
rect 6779 41225 6788 41259
rect 6736 41216 6788 41225
rect 7012 41216 7064 41268
rect 2136 41080 2188 41132
rect 2412 40876 2464 40928
rect 3700 41080 3752 41132
rect 3792 41123 3844 41132
rect 3792 41089 3812 41123
rect 3812 41089 3844 41123
rect 3792 41080 3844 41089
rect 4344 41080 4396 41132
rect 7104 41080 7156 41132
rect 8944 41080 8996 41132
rect 16212 41080 16264 41132
rect 16856 41080 16908 41132
rect 30104 41123 30156 41132
rect 30104 41089 30113 41123
rect 30113 41089 30147 41123
rect 30147 41089 30156 41123
rect 30104 41080 30156 41089
rect 3516 41055 3568 41064
rect 3516 41021 3525 41055
rect 3525 41021 3559 41055
rect 3559 41021 3568 41055
rect 3516 41012 3568 41021
rect 4160 41012 4212 41064
rect 5816 41055 5868 41064
rect 5816 41021 5825 41055
rect 5825 41021 5859 41055
rect 5859 41021 5868 41055
rect 5816 41012 5868 41021
rect 8484 41012 8536 41064
rect 4528 40944 4580 40996
rect 4436 40919 4488 40928
rect 4436 40885 4445 40919
rect 4445 40885 4479 40919
rect 4479 40885 4488 40919
rect 4436 40876 4488 40885
rect 5172 40876 5224 40928
rect 16764 40919 16816 40928
rect 16764 40885 16773 40919
rect 16773 40885 16807 40919
rect 16807 40885 16816 40919
rect 16764 40876 16816 40885
rect 29920 40919 29972 40928
rect 29920 40885 29929 40919
rect 29929 40885 29963 40919
rect 29963 40885 29972 40919
rect 29920 40876 29972 40885
rect 5915 40774 5967 40826
rect 5979 40774 6031 40826
rect 6043 40774 6095 40826
rect 6107 40774 6159 40826
rect 6171 40774 6223 40826
rect 15846 40774 15898 40826
rect 15910 40774 15962 40826
rect 15974 40774 16026 40826
rect 16038 40774 16090 40826
rect 16102 40774 16154 40826
rect 25776 40774 25828 40826
rect 25840 40774 25892 40826
rect 25904 40774 25956 40826
rect 25968 40774 26020 40826
rect 26032 40774 26084 40826
rect 2412 40672 2464 40724
rect 2872 40672 2924 40724
rect 4344 40715 4396 40724
rect 4344 40681 4353 40715
rect 4353 40681 4387 40715
rect 4387 40681 4396 40715
rect 4344 40672 4396 40681
rect 2228 40604 2280 40656
rect 3700 40604 3752 40656
rect 8024 40604 8076 40656
rect 4804 40579 4856 40588
rect 4804 40545 4813 40579
rect 4813 40545 4847 40579
rect 4847 40545 4856 40579
rect 4804 40536 4856 40545
rect 5632 40536 5684 40588
rect 7196 40579 7248 40588
rect 1768 40468 1820 40520
rect 4436 40468 4488 40520
rect 4712 40511 4764 40520
rect 4712 40477 4721 40511
rect 4721 40477 4755 40511
rect 4755 40477 4764 40511
rect 4712 40468 4764 40477
rect 5172 40468 5224 40520
rect 5356 40468 5408 40520
rect 6276 40468 6328 40520
rect 7196 40545 7205 40579
rect 7205 40545 7239 40579
rect 7239 40545 7248 40579
rect 7196 40536 7248 40545
rect 15108 40579 15160 40588
rect 15108 40545 15117 40579
rect 15117 40545 15151 40579
rect 15151 40545 15160 40579
rect 15108 40536 15160 40545
rect 16304 40536 16356 40588
rect 6552 40468 6604 40520
rect 7012 40468 7064 40520
rect 8300 40468 8352 40520
rect 9128 40511 9180 40520
rect 9128 40477 9137 40511
rect 9137 40477 9171 40511
rect 9171 40477 9180 40511
rect 9128 40468 9180 40477
rect 9588 40511 9640 40520
rect 9588 40477 9597 40511
rect 9597 40477 9631 40511
rect 9631 40477 9640 40511
rect 9588 40468 9640 40477
rect 12164 40468 12216 40520
rect 12992 40511 13044 40520
rect 12992 40477 13001 40511
rect 13001 40477 13035 40511
rect 13035 40477 13044 40511
rect 12992 40468 13044 40477
rect 14464 40511 14516 40520
rect 14464 40477 14473 40511
rect 14473 40477 14507 40511
rect 14507 40477 14516 40511
rect 14464 40468 14516 40477
rect 14648 40511 14700 40520
rect 14648 40477 14657 40511
rect 14657 40477 14691 40511
rect 14691 40477 14700 40511
rect 14648 40468 14700 40477
rect 15476 40511 15528 40520
rect 15476 40477 15510 40511
rect 15510 40477 15528 40511
rect 15476 40468 15528 40477
rect 9036 40400 9088 40452
rect 1492 40375 1544 40384
rect 1492 40341 1501 40375
rect 1501 40341 1535 40375
rect 1535 40341 1544 40375
rect 1492 40332 1544 40341
rect 8944 40375 8996 40384
rect 8944 40341 8953 40375
rect 8953 40341 8987 40375
rect 8987 40341 8996 40375
rect 8944 40332 8996 40341
rect 10416 40332 10468 40384
rect 12532 40375 12584 40384
rect 12532 40341 12541 40375
rect 12541 40341 12575 40375
rect 12575 40341 12584 40375
rect 12532 40332 12584 40341
rect 13544 40332 13596 40384
rect 15200 40332 15252 40384
rect 15752 40332 15804 40384
rect 17408 40468 17460 40520
rect 16580 40400 16632 40452
rect 17592 40443 17644 40452
rect 17592 40409 17601 40443
rect 17601 40409 17635 40443
rect 17635 40409 17644 40443
rect 17592 40400 17644 40409
rect 17040 40332 17092 40384
rect 17132 40375 17184 40384
rect 17132 40341 17141 40375
rect 17141 40341 17175 40375
rect 17175 40341 17184 40375
rect 17132 40332 17184 40341
rect 10880 40230 10932 40282
rect 10944 40230 10996 40282
rect 11008 40230 11060 40282
rect 11072 40230 11124 40282
rect 11136 40230 11188 40282
rect 20811 40230 20863 40282
rect 20875 40230 20927 40282
rect 20939 40230 20991 40282
rect 21003 40230 21055 40282
rect 21067 40230 21119 40282
rect 3424 40128 3476 40180
rect 3976 40128 4028 40180
rect 5816 40128 5868 40180
rect 4896 40060 4948 40112
rect 3056 39992 3108 40044
rect 3792 39992 3844 40044
rect 5632 40035 5684 40044
rect 5632 40001 5641 40035
rect 5641 40001 5675 40035
rect 5675 40001 5684 40035
rect 5632 39992 5684 40001
rect 6460 39992 6512 40044
rect 6736 40060 6788 40112
rect 9588 40128 9640 40180
rect 12164 40171 12216 40180
rect 12164 40137 12173 40171
rect 12173 40137 12207 40171
rect 12207 40137 12216 40171
rect 12164 40128 12216 40137
rect 13176 40128 13228 40180
rect 15200 40128 15252 40180
rect 17868 40128 17920 40180
rect 7104 40035 7156 40044
rect 7104 40001 7113 40035
rect 7113 40001 7147 40035
rect 7147 40001 7156 40035
rect 7104 39992 7156 40001
rect 6644 39967 6696 39976
rect 1400 39788 1452 39840
rect 6644 39933 6653 39967
rect 6653 39933 6687 39967
rect 6687 39933 6696 39967
rect 6644 39924 6696 39933
rect 7012 39924 7064 39976
rect 8300 40060 8352 40112
rect 8944 40060 8996 40112
rect 9036 40060 9088 40112
rect 9496 40060 9548 40112
rect 9864 40060 9916 40112
rect 9680 39992 9732 40044
rect 10416 40035 10468 40044
rect 10416 40001 10425 40035
rect 10425 40001 10459 40035
rect 10459 40001 10468 40035
rect 10416 39992 10468 40001
rect 12532 39992 12584 40044
rect 8760 39924 8812 39976
rect 16764 39992 16816 40044
rect 16856 40035 16908 40044
rect 16856 40001 16865 40035
rect 16865 40001 16899 40035
rect 16899 40001 16908 40035
rect 16856 39992 16908 40001
rect 17592 40035 17644 40044
rect 17592 40001 17601 40035
rect 17601 40001 17635 40035
rect 17635 40001 17644 40035
rect 17592 39992 17644 40001
rect 19340 39992 19392 40044
rect 22100 39992 22152 40044
rect 4344 39856 4396 39908
rect 7656 39856 7708 39908
rect 12624 39856 12676 39908
rect 13268 39899 13320 39908
rect 13268 39865 13277 39899
rect 13277 39865 13311 39899
rect 13311 39865 13320 39899
rect 13268 39856 13320 39865
rect 13636 39967 13688 39976
rect 13636 39933 13670 39967
rect 13670 39933 13688 39967
rect 13820 39967 13872 39976
rect 13636 39924 13688 39933
rect 13820 39933 13829 39967
rect 13829 39933 13863 39967
rect 13863 39933 13872 39967
rect 13820 39924 13872 39933
rect 15200 39967 15252 39976
rect 15200 39933 15209 39967
rect 15209 39933 15243 39967
rect 15243 39933 15252 39967
rect 15200 39924 15252 39933
rect 16304 39924 16356 39976
rect 17408 39924 17460 39976
rect 18052 39924 18104 39976
rect 21824 39967 21876 39976
rect 21824 39933 21833 39967
rect 21833 39933 21867 39967
rect 21867 39933 21876 39967
rect 21824 39924 21876 39933
rect 29920 39924 29972 39976
rect 16856 39856 16908 39908
rect 5816 39831 5868 39840
rect 5816 39797 5825 39831
rect 5825 39797 5859 39831
rect 5859 39797 5868 39831
rect 5816 39788 5868 39797
rect 8576 39831 8628 39840
rect 8576 39797 8585 39831
rect 8585 39797 8619 39831
rect 8619 39797 8628 39831
rect 8576 39788 8628 39797
rect 9496 39788 9548 39840
rect 13360 39788 13412 39840
rect 15476 39788 15528 39840
rect 17776 39788 17828 39840
rect 18972 39831 19024 39840
rect 18972 39797 18981 39831
rect 18981 39797 19015 39831
rect 19015 39797 19024 39831
rect 18972 39788 19024 39797
rect 5915 39686 5967 39738
rect 5979 39686 6031 39738
rect 6043 39686 6095 39738
rect 6107 39686 6159 39738
rect 6171 39686 6223 39738
rect 15846 39686 15898 39738
rect 15910 39686 15962 39738
rect 15974 39686 16026 39738
rect 16038 39686 16090 39738
rect 16102 39686 16154 39738
rect 25776 39686 25828 39738
rect 25840 39686 25892 39738
rect 25904 39686 25956 39738
rect 25968 39686 26020 39738
rect 26032 39686 26084 39738
rect 2136 39516 2188 39568
rect 2412 39584 2464 39636
rect 3056 39627 3108 39636
rect 3056 39593 3065 39627
rect 3065 39593 3099 39627
rect 3099 39593 3108 39627
rect 3056 39584 3108 39593
rect 3792 39627 3844 39636
rect 3792 39593 3801 39627
rect 3801 39593 3835 39627
rect 3835 39593 3844 39627
rect 3792 39584 3844 39593
rect 5632 39584 5684 39636
rect 2412 39448 2464 39500
rect 4160 39491 4212 39500
rect 4160 39457 4169 39491
rect 4169 39457 4203 39491
rect 4203 39457 4212 39491
rect 4160 39448 4212 39457
rect 4712 39448 4764 39500
rect 3240 39423 3292 39432
rect 3240 39389 3249 39423
rect 3249 39389 3283 39423
rect 3283 39389 3292 39423
rect 3240 39380 3292 39389
rect 3976 39423 4028 39432
rect 3976 39389 3985 39423
rect 3985 39389 4019 39423
rect 4019 39389 4028 39423
rect 3976 39380 4028 39389
rect 4252 39423 4304 39432
rect 4252 39389 4258 39423
rect 4258 39389 4292 39423
rect 4292 39389 4304 39423
rect 4252 39380 4304 39389
rect 4344 39423 4396 39432
rect 4344 39389 4353 39423
rect 4353 39389 4387 39423
rect 4387 39389 4396 39423
rect 4344 39380 4396 39389
rect 4528 39423 4580 39432
rect 4528 39389 4537 39423
rect 4537 39389 4571 39423
rect 4571 39389 4580 39423
rect 4528 39380 4580 39389
rect 5080 39380 5132 39432
rect 5724 39380 5776 39432
rect 9036 39584 9088 39636
rect 12992 39627 13044 39636
rect 12992 39593 13001 39627
rect 13001 39593 13035 39627
rect 13035 39593 13044 39627
rect 12992 39584 13044 39593
rect 7012 39448 7064 39500
rect 8576 39448 8628 39500
rect 13268 39516 13320 39568
rect 15660 39584 15712 39636
rect 16856 39584 16908 39636
rect 18052 39584 18104 39636
rect 18788 39516 18840 39568
rect 14648 39491 14700 39500
rect 14648 39457 14657 39491
rect 14657 39457 14691 39491
rect 14691 39457 14700 39491
rect 14648 39448 14700 39457
rect 6644 39423 6696 39432
rect 6644 39389 6653 39423
rect 6653 39389 6687 39423
rect 6687 39389 6696 39423
rect 6920 39423 6972 39432
rect 6644 39380 6696 39389
rect 6920 39389 6929 39423
rect 6929 39389 6963 39423
rect 6963 39389 6972 39423
rect 6920 39380 6972 39389
rect 6460 39312 6512 39364
rect 6828 39312 6880 39364
rect 8116 39380 8168 39432
rect 13728 39380 13780 39432
rect 14464 39423 14516 39432
rect 14464 39389 14473 39423
rect 14473 39389 14507 39423
rect 14507 39389 14516 39423
rect 15476 39491 15528 39500
rect 15476 39457 15510 39491
rect 15510 39457 15528 39491
rect 15476 39448 15528 39457
rect 16304 39448 16356 39500
rect 16856 39491 16908 39500
rect 16856 39457 16865 39491
rect 16865 39457 16899 39491
rect 16899 39457 16908 39491
rect 16856 39448 16908 39457
rect 17040 39491 17092 39500
rect 17040 39457 17049 39491
rect 17049 39457 17083 39491
rect 17083 39457 17092 39491
rect 17040 39448 17092 39457
rect 18144 39423 18196 39432
rect 14464 39380 14516 39389
rect 18144 39389 18153 39423
rect 18153 39389 18187 39423
rect 18187 39389 18196 39423
rect 18144 39380 18196 39389
rect 19432 39380 19484 39432
rect 30104 39423 30156 39432
rect 30104 39389 30113 39423
rect 30113 39389 30147 39423
rect 30147 39389 30156 39423
rect 30104 39380 30156 39389
rect 6644 39244 6696 39296
rect 8484 39312 8536 39364
rect 9312 39355 9364 39364
rect 9312 39321 9346 39355
rect 9346 39321 9364 39355
rect 12624 39355 12676 39364
rect 9312 39312 9364 39321
rect 12624 39321 12633 39355
rect 12633 39321 12667 39355
rect 12667 39321 12676 39355
rect 12624 39312 12676 39321
rect 7104 39287 7156 39296
rect 7104 39253 7113 39287
rect 7113 39253 7147 39287
rect 7147 39253 7156 39287
rect 7104 39244 7156 39253
rect 8208 39287 8260 39296
rect 8208 39253 8217 39287
rect 8217 39253 8251 39287
rect 8251 39253 8260 39287
rect 8208 39244 8260 39253
rect 9128 39244 9180 39296
rect 17868 39312 17920 39364
rect 19616 39355 19668 39364
rect 19616 39321 19625 39355
rect 19625 39321 19659 39355
rect 19659 39321 19668 39355
rect 19616 39312 19668 39321
rect 14832 39244 14884 39296
rect 17684 39244 17736 39296
rect 20260 39244 20312 39296
rect 29920 39287 29972 39296
rect 29920 39253 29929 39287
rect 29929 39253 29963 39287
rect 29963 39253 29972 39287
rect 29920 39244 29972 39253
rect 10880 39142 10932 39194
rect 10944 39142 10996 39194
rect 11008 39142 11060 39194
rect 11072 39142 11124 39194
rect 11136 39142 11188 39194
rect 20811 39142 20863 39194
rect 20875 39142 20927 39194
rect 20939 39142 20991 39194
rect 21003 39142 21055 39194
rect 21067 39142 21119 39194
rect 3608 39040 3660 39092
rect 5724 39040 5776 39092
rect 6920 39040 6972 39092
rect 9312 39083 9364 39092
rect 9312 39049 9321 39083
rect 9321 39049 9355 39083
rect 9355 39049 9364 39083
rect 9312 39040 9364 39049
rect 15200 39040 15252 39092
rect 16212 39040 16264 39092
rect 17408 39040 17460 39092
rect 17684 39083 17736 39092
rect 17684 39049 17693 39083
rect 17693 39049 17727 39083
rect 17727 39049 17736 39083
rect 17684 39040 17736 39049
rect 17776 39083 17828 39092
rect 17776 39049 17785 39083
rect 17785 39049 17819 39083
rect 17819 39049 17828 39083
rect 18788 39083 18840 39092
rect 17776 39040 17828 39049
rect 18788 39049 18797 39083
rect 18797 39049 18831 39083
rect 18831 39049 18840 39083
rect 18788 39040 18840 39049
rect 18972 39040 19024 39092
rect 19616 39040 19668 39092
rect 21916 39083 21968 39092
rect 21916 39049 21925 39083
rect 21925 39049 21959 39083
rect 21959 39049 21968 39083
rect 21916 39040 21968 39049
rect 2504 38972 2556 39024
rect 1860 38904 1912 38956
rect 2136 38904 2188 38956
rect 2780 38904 2832 38956
rect 3056 38904 3108 38956
rect 3516 38904 3568 38956
rect 3976 38947 4028 38956
rect 3976 38913 3985 38947
rect 3985 38913 4019 38947
rect 4019 38913 4028 38947
rect 3976 38904 4028 38913
rect 8024 38972 8076 39024
rect 5632 38947 5684 38956
rect 5632 38913 5641 38947
rect 5641 38913 5675 38947
rect 5675 38913 5684 38947
rect 5632 38904 5684 38913
rect 5816 38904 5868 38956
rect 7104 38904 7156 38956
rect 8576 38947 8628 38956
rect 8576 38913 8585 38947
rect 8585 38913 8619 38947
rect 8619 38913 8628 38947
rect 8576 38904 8628 38913
rect 8760 38947 8812 38956
rect 8760 38913 8769 38947
rect 8769 38913 8803 38947
rect 8803 38913 8812 38947
rect 8760 38904 8812 38913
rect 9128 38947 9180 38956
rect 9128 38913 9137 38947
rect 9137 38913 9171 38947
rect 9171 38913 9180 38947
rect 9128 38904 9180 38913
rect 11428 38904 11480 38956
rect 12532 38947 12584 38956
rect 12532 38913 12541 38947
rect 12541 38913 12575 38947
rect 12575 38913 12584 38947
rect 12532 38904 12584 38913
rect 13452 38947 13504 38956
rect 13452 38913 13461 38947
rect 13461 38913 13495 38947
rect 13495 38913 13504 38947
rect 13452 38904 13504 38913
rect 14832 38904 14884 38956
rect 16580 38972 16632 39024
rect 15660 38904 15712 38956
rect 17132 38904 17184 38956
rect 20076 38947 20128 38956
rect 20076 38913 20085 38947
rect 20085 38913 20119 38947
rect 20119 38913 20128 38947
rect 20076 38904 20128 38913
rect 22100 38947 22152 38956
rect 22100 38913 22109 38947
rect 22109 38913 22143 38947
rect 22143 38913 22152 38947
rect 22100 38904 22152 38913
rect 2780 38768 2832 38820
rect 2412 38743 2464 38752
rect 2412 38709 2421 38743
rect 2421 38709 2455 38743
rect 2455 38709 2464 38743
rect 2412 38700 2464 38709
rect 2872 38700 2924 38752
rect 4160 38743 4212 38752
rect 4160 38709 4169 38743
rect 4169 38709 4203 38743
rect 4203 38709 4212 38743
rect 4160 38700 4212 38709
rect 6736 38700 6788 38752
rect 9312 38836 9364 38888
rect 12624 38836 12676 38888
rect 13268 38836 13320 38888
rect 13544 38879 13596 38888
rect 13544 38845 13578 38879
rect 13578 38845 13596 38879
rect 13544 38836 13596 38845
rect 13912 38836 13964 38888
rect 16304 38836 16356 38888
rect 17960 38879 18012 38888
rect 17960 38845 17969 38879
rect 17969 38845 18003 38879
rect 18003 38845 18012 38879
rect 17960 38836 18012 38845
rect 29920 38836 29972 38888
rect 13176 38811 13228 38820
rect 13176 38777 13185 38811
rect 13185 38777 13219 38811
rect 13219 38777 13228 38811
rect 13176 38768 13228 38777
rect 9220 38700 9272 38752
rect 10600 38700 10652 38752
rect 16764 38700 16816 38752
rect 19156 38700 19208 38752
rect 21364 38700 21416 38752
rect 5915 38598 5967 38650
rect 5979 38598 6031 38650
rect 6043 38598 6095 38650
rect 6107 38598 6159 38650
rect 6171 38598 6223 38650
rect 15846 38598 15898 38650
rect 15910 38598 15962 38650
rect 15974 38598 16026 38650
rect 16038 38598 16090 38650
rect 16102 38598 16154 38650
rect 25776 38598 25828 38650
rect 25840 38598 25892 38650
rect 25904 38598 25956 38650
rect 25968 38598 26020 38650
rect 26032 38598 26084 38650
rect 2412 38496 2464 38548
rect 2596 38496 2648 38548
rect 4252 38496 4304 38548
rect 8300 38496 8352 38548
rect 9680 38539 9732 38548
rect 9680 38505 9689 38539
rect 9689 38505 9723 38539
rect 9723 38505 9732 38539
rect 9680 38496 9732 38505
rect 13728 38496 13780 38548
rect 18144 38496 18196 38548
rect 19340 38496 19392 38548
rect 20076 38539 20128 38548
rect 20076 38505 20085 38539
rect 20085 38505 20119 38539
rect 20119 38505 20128 38539
rect 20076 38496 20128 38505
rect 2136 38428 2188 38480
rect 9128 38428 9180 38480
rect 13268 38428 13320 38480
rect 13360 38428 13412 38480
rect 2504 38360 2556 38412
rect 2964 38335 3016 38344
rect 2964 38301 2973 38335
rect 2973 38301 3007 38335
rect 3007 38301 3016 38335
rect 2964 38292 3016 38301
rect 4712 38360 4764 38412
rect 6736 38403 6788 38412
rect 6736 38369 6745 38403
rect 6745 38369 6779 38403
rect 6779 38369 6788 38403
rect 6736 38360 6788 38369
rect 9220 38403 9272 38412
rect 9220 38369 9229 38403
rect 9229 38369 9263 38403
rect 9263 38369 9272 38403
rect 9220 38360 9272 38369
rect 14372 38360 14424 38412
rect 4252 38335 4304 38344
rect 4252 38301 4261 38335
rect 4261 38301 4295 38335
rect 4295 38301 4304 38335
rect 4252 38292 4304 38301
rect 3148 38199 3200 38208
rect 3148 38165 3157 38199
rect 3157 38165 3191 38199
rect 3191 38165 3200 38199
rect 3148 38156 3200 38165
rect 3792 38199 3844 38208
rect 3792 38165 3801 38199
rect 3801 38165 3835 38199
rect 3835 38165 3844 38199
rect 3792 38156 3844 38165
rect 4620 38292 4672 38344
rect 4896 38224 4948 38276
rect 8024 38292 8076 38344
rect 8576 38292 8628 38344
rect 5632 38224 5684 38276
rect 9036 38292 9088 38344
rect 9312 38335 9364 38344
rect 9312 38301 9321 38335
rect 9321 38301 9355 38335
rect 9355 38301 9364 38335
rect 9312 38292 9364 38301
rect 9496 38335 9548 38344
rect 9496 38301 9505 38335
rect 9505 38301 9539 38335
rect 9539 38301 9548 38335
rect 9496 38292 9548 38301
rect 10416 38335 10468 38344
rect 10416 38301 10425 38335
rect 10425 38301 10459 38335
rect 10459 38301 10468 38335
rect 10416 38292 10468 38301
rect 4528 38156 4580 38208
rect 7564 38156 7616 38208
rect 9680 38224 9732 38276
rect 9312 38156 9364 38208
rect 12716 38292 12768 38344
rect 13360 38335 13412 38344
rect 13360 38301 13369 38335
rect 13369 38301 13403 38335
rect 13403 38301 13412 38335
rect 13360 38292 13412 38301
rect 14280 38335 14332 38344
rect 14280 38301 14289 38335
rect 14289 38301 14323 38335
rect 14323 38301 14332 38335
rect 14280 38292 14332 38301
rect 14924 38335 14976 38344
rect 13544 38224 13596 38276
rect 11520 38156 11572 38208
rect 13268 38156 13320 38208
rect 14924 38301 14933 38335
rect 14933 38301 14967 38335
rect 14967 38301 14976 38335
rect 14924 38292 14976 38301
rect 15108 38335 15160 38344
rect 15108 38301 15117 38335
rect 15117 38301 15151 38335
rect 15151 38301 15160 38335
rect 15108 38292 15160 38301
rect 17776 38292 17828 38344
rect 18788 38292 18840 38344
rect 20260 38335 20312 38344
rect 20260 38301 20269 38335
rect 20269 38301 20303 38335
rect 20303 38301 20312 38335
rect 20260 38292 20312 38301
rect 19432 38267 19484 38276
rect 19432 38233 19441 38267
rect 19441 38233 19475 38267
rect 19475 38233 19484 38267
rect 19432 38224 19484 38233
rect 10880 38054 10932 38106
rect 10944 38054 10996 38106
rect 11008 38054 11060 38106
rect 11072 38054 11124 38106
rect 11136 38054 11188 38106
rect 20811 38054 20863 38106
rect 20875 38054 20927 38106
rect 20939 38054 20991 38106
rect 21003 38054 21055 38106
rect 21067 38054 21119 38106
rect 2504 37952 2556 38004
rect 3792 37884 3844 37936
rect 4160 37859 4212 37868
rect 4160 37825 4169 37859
rect 4169 37825 4203 37859
rect 4203 37825 4212 37859
rect 4160 37816 4212 37825
rect 4436 37859 4488 37868
rect 4436 37825 4470 37859
rect 4470 37825 4488 37859
rect 4436 37816 4488 37825
rect 6368 37816 6420 37868
rect 7012 37884 7064 37936
rect 3700 37791 3752 37800
rect 3700 37757 3709 37791
rect 3709 37757 3743 37791
rect 3743 37757 3752 37791
rect 3700 37748 3752 37757
rect 6644 37748 6696 37800
rect 7104 37859 7156 37868
rect 7104 37825 7113 37859
rect 7113 37825 7147 37859
rect 7147 37825 7156 37859
rect 7748 37859 7800 37868
rect 7104 37816 7156 37825
rect 7748 37825 7757 37859
rect 7757 37825 7791 37859
rect 7791 37825 7800 37859
rect 7748 37816 7800 37825
rect 5632 37680 5684 37732
rect 7932 37748 7984 37800
rect 8208 37859 8260 37868
rect 8208 37825 8217 37859
rect 8217 37825 8251 37859
rect 8251 37825 8260 37859
rect 8208 37816 8260 37825
rect 8944 37816 8996 37868
rect 10140 37816 10192 37868
rect 10324 37884 10376 37936
rect 11244 37884 11296 37936
rect 11520 37859 11572 37868
rect 9772 37748 9824 37800
rect 10508 37748 10560 37800
rect 1492 37655 1544 37664
rect 1492 37621 1501 37655
rect 1501 37621 1535 37655
rect 1535 37621 1544 37655
rect 1492 37612 1544 37621
rect 5540 37655 5592 37664
rect 5540 37621 5549 37655
rect 5549 37621 5583 37655
rect 5583 37621 5592 37655
rect 5540 37612 5592 37621
rect 6368 37655 6420 37664
rect 6368 37621 6377 37655
rect 6377 37621 6411 37655
rect 6411 37621 6420 37655
rect 6368 37612 6420 37621
rect 9588 37655 9640 37664
rect 9588 37621 9597 37655
rect 9597 37621 9631 37655
rect 9631 37621 9640 37655
rect 9588 37612 9640 37621
rect 10048 37680 10100 37732
rect 11520 37825 11529 37859
rect 11529 37825 11563 37859
rect 11563 37825 11572 37859
rect 11520 37816 11572 37825
rect 14280 37952 14332 38004
rect 14464 37952 14516 38004
rect 16212 37952 16264 38004
rect 12992 37748 13044 37800
rect 13360 37791 13412 37800
rect 13360 37757 13369 37791
rect 13369 37757 13403 37791
rect 13403 37757 13412 37791
rect 13360 37748 13412 37757
rect 13820 37816 13872 37868
rect 14188 37816 14240 37868
rect 14372 37859 14424 37868
rect 14372 37825 14381 37859
rect 14381 37825 14415 37859
rect 14415 37825 14424 37859
rect 14372 37816 14424 37825
rect 19432 37884 19484 37936
rect 17684 37859 17736 37868
rect 17684 37825 17693 37859
rect 17693 37825 17727 37859
rect 17727 37825 17736 37859
rect 17684 37816 17736 37825
rect 14004 37748 14056 37800
rect 15108 37791 15160 37800
rect 15108 37757 15117 37791
rect 15117 37757 15151 37791
rect 15151 37757 15160 37791
rect 15108 37748 15160 37757
rect 10876 37612 10928 37664
rect 14924 37680 14976 37732
rect 12440 37612 12492 37664
rect 12900 37655 12952 37664
rect 12900 37621 12909 37655
rect 12909 37621 12943 37655
rect 12943 37621 12952 37655
rect 12900 37612 12952 37621
rect 13728 37612 13780 37664
rect 18512 37655 18564 37664
rect 18512 37621 18521 37655
rect 18521 37621 18555 37655
rect 18555 37621 18564 37655
rect 18512 37612 18564 37621
rect 5915 37510 5967 37562
rect 5979 37510 6031 37562
rect 6043 37510 6095 37562
rect 6107 37510 6159 37562
rect 6171 37510 6223 37562
rect 15846 37510 15898 37562
rect 15910 37510 15962 37562
rect 15974 37510 16026 37562
rect 16038 37510 16090 37562
rect 16102 37510 16154 37562
rect 25776 37510 25828 37562
rect 25840 37510 25892 37562
rect 25904 37510 25956 37562
rect 25968 37510 26020 37562
rect 26032 37510 26084 37562
rect 2412 37408 2464 37460
rect 6460 37408 6512 37460
rect 8944 37451 8996 37460
rect 8944 37417 8953 37451
rect 8953 37417 8987 37451
rect 8987 37417 8996 37451
rect 8944 37408 8996 37417
rect 12716 37451 12768 37460
rect 12716 37417 12725 37451
rect 12725 37417 12759 37451
rect 12759 37417 12768 37451
rect 12716 37408 12768 37417
rect 13820 37408 13872 37460
rect 14004 37408 14056 37460
rect 20352 37408 20404 37460
rect 1952 37247 2004 37256
rect 1952 37213 1961 37247
rect 1961 37213 1995 37247
rect 1995 37213 2004 37247
rect 1952 37204 2004 37213
rect 3240 37204 3292 37256
rect 3792 37204 3844 37256
rect 3332 37136 3384 37188
rect 4620 37272 4672 37324
rect 4804 37272 4856 37324
rect 5632 37315 5684 37324
rect 5632 37281 5641 37315
rect 5641 37281 5675 37315
rect 5675 37281 5684 37315
rect 5632 37272 5684 37281
rect 5816 37272 5868 37324
rect 9588 37340 9640 37392
rect 15200 37340 15252 37392
rect 9220 37272 9272 37324
rect 15384 37272 15436 37324
rect 15660 37272 15712 37324
rect 16120 37315 16172 37324
rect 16120 37281 16154 37315
rect 16154 37281 16172 37315
rect 16304 37315 16356 37324
rect 16120 37272 16172 37281
rect 16304 37281 16313 37315
rect 16313 37281 16347 37315
rect 16347 37281 16356 37315
rect 17960 37315 18012 37324
rect 16304 37272 16356 37281
rect 17960 37281 17969 37315
rect 17969 37281 18003 37315
rect 18003 37281 18012 37315
rect 17960 37272 18012 37281
rect 5724 37204 5776 37256
rect 6368 37247 6420 37256
rect 6368 37213 6402 37247
rect 6402 37213 6420 37247
rect 6368 37204 6420 37213
rect 8300 37204 8352 37256
rect 9128 37247 9180 37256
rect 9128 37213 9137 37247
rect 9137 37213 9171 37247
rect 9171 37213 9180 37247
rect 9128 37204 9180 37213
rect 9312 37247 9364 37256
rect 9312 37213 9321 37247
rect 9321 37213 9355 37247
rect 9355 37213 9364 37247
rect 9312 37204 9364 37213
rect 7748 37136 7800 37188
rect 7932 37136 7984 37188
rect 9680 37247 9732 37256
rect 9680 37213 9689 37247
rect 9689 37213 9723 37247
rect 9723 37213 9732 37247
rect 10600 37247 10652 37256
rect 9680 37204 9732 37213
rect 10600 37213 10609 37247
rect 10609 37213 10643 37247
rect 10643 37213 10652 37247
rect 10600 37204 10652 37213
rect 10876 37247 10928 37256
rect 10876 37213 10910 37247
rect 10910 37213 10928 37247
rect 10876 37204 10928 37213
rect 12992 37247 13044 37256
rect 12992 37213 13001 37247
rect 13001 37213 13035 37247
rect 13035 37213 13044 37247
rect 12992 37204 13044 37213
rect 13084 37247 13136 37256
rect 13084 37213 13093 37247
rect 13093 37213 13127 37247
rect 13127 37213 13136 37247
rect 14096 37247 14148 37256
rect 13084 37204 13136 37213
rect 14096 37213 14105 37247
rect 14105 37213 14139 37247
rect 14139 37213 14148 37247
rect 14096 37204 14148 37213
rect 11336 37136 11388 37188
rect 13728 37136 13780 37188
rect 14924 37204 14976 37256
rect 15292 37247 15344 37256
rect 15292 37213 15301 37247
rect 15301 37213 15335 37247
rect 15335 37213 15344 37247
rect 15292 37204 15344 37213
rect 17684 37204 17736 37256
rect 18512 37204 18564 37256
rect 18788 37204 18840 37256
rect 30104 37247 30156 37256
rect 30104 37213 30113 37247
rect 30113 37213 30147 37247
rect 30147 37213 30156 37247
rect 30104 37204 30156 37213
rect 15200 37136 15252 37188
rect 2964 37068 3016 37120
rect 3148 37111 3200 37120
rect 3148 37077 3157 37111
rect 3157 37077 3191 37111
rect 3191 37077 3200 37111
rect 3148 37068 3200 37077
rect 3424 37068 3476 37120
rect 4620 37068 4672 37120
rect 4988 37068 5040 37120
rect 7288 37068 7340 37120
rect 8116 37068 8168 37120
rect 8300 37068 8352 37120
rect 10048 37068 10100 37120
rect 14096 37068 14148 37120
rect 14832 37068 14884 37120
rect 16948 37111 17000 37120
rect 16948 37077 16957 37111
rect 16957 37077 16991 37111
rect 16991 37077 17000 37111
rect 16948 37068 17000 37077
rect 18144 37068 18196 37120
rect 19248 37111 19300 37120
rect 19248 37077 19257 37111
rect 19257 37077 19291 37111
rect 19291 37077 19300 37111
rect 19248 37068 19300 37077
rect 29920 37111 29972 37120
rect 29920 37077 29929 37111
rect 29929 37077 29963 37111
rect 29963 37077 29972 37111
rect 29920 37068 29972 37077
rect 10880 36966 10932 37018
rect 10944 36966 10996 37018
rect 11008 36966 11060 37018
rect 11072 36966 11124 37018
rect 11136 36966 11188 37018
rect 20811 36966 20863 37018
rect 20875 36966 20927 37018
rect 20939 36966 20991 37018
rect 21003 36966 21055 37018
rect 21067 36966 21119 37018
rect 1952 36864 2004 36916
rect 3056 36864 3108 36916
rect 3700 36864 3752 36916
rect 3792 36864 3844 36916
rect 11244 36864 11296 36916
rect 11428 36864 11480 36916
rect 14924 36907 14976 36916
rect 14924 36873 14933 36907
rect 14933 36873 14967 36907
rect 14967 36873 14976 36907
rect 14924 36864 14976 36873
rect 16948 36864 17000 36916
rect 17684 36864 17736 36916
rect 18788 36907 18840 36916
rect 18788 36873 18797 36907
rect 18797 36873 18831 36907
rect 18831 36873 18840 36907
rect 18788 36864 18840 36873
rect 1768 36728 1820 36780
rect 2136 36728 2188 36780
rect 3424 36771 3476 36780
rect 3424 36737 3433 36771
rect 3433 36737 3467 36771
rect 3467 36737 3476 36771
rect 3424 36728 3476 36737
rect 4436 36796 4488 36848
rect 5540 36796 5592 36848
rect 4620 36771 4672 36780
rect 4620 36737 4629 36771
rect 4629 36737 4663 36771
rect 4663 36737 4672 36771
rect 4620 36728 4672 36737
rect 4804 36771 4856 36780
rect 4804 36737 4813 36771
rect 4813 36737 4847 36771
rect 4847 36737 4856 36771
rect 5632 36771 5684 36780
rect 4804 36728 4856 36737
rect 5632 36737 5641 36771
rect 5641 36737 5675 36771
rect 5675 36737 5684 36771
rect 5632 36728 5684 36737
rect 7472 36728 7524 36780
rect 8116 36728 8168 36780
rect 10140 36771 10192 36780
rect 10140 36737 10149 36771
rect 10149 36737 10183 36771
rect 10183 36737 10192 36771
rect 10140 36728 10192 36737
rect 10324 36771 10376 36780
rect 10324 36737 10333 36771
rect 10333 36737 10367 36771
rect 10367 36737 10376 36771
rect 10324 36728 10376 36737
rect 10508 36771 10560 36780
rect 10508 36737 10517 36771
rect 10517 36737 10551 36771
rect 10551 36737 10560 36771
rect 10508 36728 10560 36737
rect 12900 36796 12952 36848
rect 10784 36728 10836 36780
rect 12440 36771 12492 36780
rect 12440 36737 12449 36771
rect 12449 36737 12483 36771
rect 12483 36737 12492 36771
rect 12440 36728 12492 36737
rect 13084 36728 13136 36780
rect 13728 36728 13780 36780
rect 13820 36771 13872 36780
rect 13820 36737 13829 36771
rect 13829 36737 13863 36771
rect 13863 36737 13872 36771
rect 13820 36728 13872 36737
rect 4528 36703 4580 36712
rect 4528 36669 4537 36703
rect 4537 36669 4571 36703
rect 4571 36669 4580 36703
rect 4528 36660 4580 36669
rect 4712 36592 4764 36644
rect 2412 36567 2464 36576
rect 2412 36533 2421 36567
rect 2421 36533 2455 36567
rect 2455 36533 2464 36567
rect 2412 36524 2464 36533
rect 2964 36524 3016 36576
rect 9496 36660 9548 36712
rect 9772 36660 9824 36712
rect 11888 36660 11940 36712
rect 14188 36771 14240 36780
rect 14188 36737 14197 36771
rect 14197 36737 14231 36771
rect 14231 36737 14240 36771
rect 14188 36728 14240 36737
rect 14924 36728 14976 36780
rect 19340 36796 19392 36848
rect 20168 36796 20220 36848
rect 19248 36771 19300 36780
rect 15292 36660 15344 36712
rect 16580 36660 16632 36712
rect 16856 36660 16908 36712
rect 17132 36703 17184 36712
rect 17132 36669 17141 36703
rect 17141 36669 17175 36703
rect 17175 36669 17184 36703
rect 17132 36660 17184 36669
rect 7564 36592 7616 36644
rect 8024 36592 8076 36644
rect 19248 36737 19257 36771
rect 19257 36737 19291 36771
rect 19291 36737 19300 36771
rect 19248 36728 19300 36737
rect 19524 36771 19576 36780
rect 19524 36737 19558 36771
rect 19558 36737 19576 36771
rect 22100 36771 22152 36780
rect 19524 36728 19576 36737
rect 22100 36737 22109 36771
rect 22109 36737 22143 36771
rect 22143 36737 22152 36771
rect 22100 36728 22152 36737
rect 29920 36660 29972 36712
rect 7196 36567 7248 36576
rect 7196 36533 7205 36567
rect 7205 36533 7239 36567
rect 7239 36533 7248 36567
rect 7196 36524 7248 36533
rect 7748 36524 7800 36576
rect 10416 36524 10468 36576
rect 10784 36524 10836 36576
rect 11336 36524 11388 36576
rect 13544 36524 13596 36576
rect 13728 36524 13780 36576
rect 20628 36567 20680 36576
rect 20628 36533 20637 36567
rect 20637 36533 20671 36567
rect 20671 36533 20680 36567
rect 20628 36524 20680 36533
rect 21272 36524 21324 36576
rect 5915 36422 5967 36474
rect 5979 36422 6031 36474
rect 6043 36422 6095 36474
rect 6107 36422 6159 36474
rect 6171 36422 6223 36474
rect 15846 36422 15898 36474
rect 15910 36422 15962 36474
rect 15974 36422 16026 36474
rect 16038 36422 16090 36474
rect 16102 36422 16154 36474
rect 25776 36422 25828 36474
rect 25840 36422 25892 36474
rect 25904 36422 25956 36474
rect 25968 36422 26020 36474
rect 26032 36422 26084 36474
rect 3976 36363 4028 36372
rect 3976 36329 3985 36363
rect 3985 36329 4019 36363
rect 4019 36329 4028 36363
rect 3976 36320 4028 36329
rect 5724 36320 5776 36372
rect 7196 36363 7248 36372
rect 7196 36329 7205 36363
rect 7205 36329 7239 36363
rect 7239 36329 7248 36363
rect 7196 36320 7248 36329
rect 9312 36320 9364 36372
rect 1768 36252 1820 36304
rect 2320 36252 2372 36304
rect 2872 36184 2924 36236
rect 2964 36116 3016 36168
rect 3792 36159 3844 36168
rect 3792 36125 3801 36159
rect 3801 36125 3835 36159
rect 3835 36125 3844 36159
rect 3792 36116 3844 36125
rect 3976 36116 4028 36168
rect 5540 36116 5592 36168
rect 6552 36116 6604 36168
rect 9680 36252 9732 36304
rect 10048 36184 10100 36236
rect 15200 36252 15252 36304
rect 17132 36320 17184 36372
rect 12900 36184 12952 36236
rect 15292 36227 15344 36236
rect 8116 36159 8168 36168
rect 8116 36125 8125 36159
rect 8125 36125 8159 36159
rect 8159 36125 8168 36159
rect 8116 36116 8168 36125
rect 8484 36116 8536 36168
rect 10324 36116 10376 36168
rect 13084 36116 13136 36168
rect 15292 36193 15301 36227
rect 15301 36193 15335 36227
rect 15335 36193 15344 36227
rect 15292 36184 15344 36193
rect 15752 36227 15804 36236
rect 15752 36193 15761 36227
rect 15761 36193 15795 36227
rect 15795 36193 15804 36227
rect 15752 36184 15804 36193
rect 21548 36252 21600 36304
rect 16120 36227 16172 36236
rect 16120 36193 16154 36227
rect 16154 36193 16172 36227
rect 16120 36184 16172 36193
rect 13268 36159 13320 36168
rect 13268 36125 13277 36159
rect 13277 36125 13311 36159
rect 13311 36125 13320 36159
rect 13268 36116 13320 36125
rect 15200 36116 15252 36168
rect 16304 36159 16356 36168
rect 16304 36125 16313 36159
rect 16313 36125 16347 36159
rect 16347 36125 16356 36159
rect 16304 36116 16356 36125
rect 19340 36184 19392 36236
rect 19800 36184 19852 36236
rect 20260 36227 20312 36236
rect 20260 36193 20269 36227
rect 20269 36193 20303 36227
rect 20303 36193 20312 36227
rect 20260 36184 20312 36193
rect 1492 36023 1544 36032
rect 1492 35989 1501 36023
rect 1501 35989 1535 36023
rect 1535 35989 1544 36023
rect 1492 35980 1544 35989
rect 2228 36023 2280 36032
rect 2228 35989 2237 36023
rect 2237 35989 2271 36023
rect 2271 35989 2280 36023
rect 2228 35980 2280 35989
rect 2872 36023 2924 36032
rect 2872 35989 2881 36023
rect 2881 35989 2915 36023
rect 2915 35989 2924 36023
rect 2872 35980 2924 35989
rect 3148 35980 3200 36032
rect 7196 35980 7248 36032
rect 7932 36023 7984 36032
rect 7932 35989 7941 36023
rect 7941 35989 7975 36023
rect 7975 35989 7984 36023
rect 7932 35980 7984 35989
rect 10692 36048 10744 36100
rect 10600 35980 10652 36032
rect 12624 36023 12676 36032
rect 12624 35989 12633 36023
rect 12633 35989 12667 36023
rect 12667 35989 12676 36023
rect 12624 35980 12676 35989
rect 13360 36048 13412 36100
rect 13176 35980 13228 36032
rect 16580 35980 16632 36032
rect 20628 36116 20680 36168
rect 21180 36116 21232 36168
rect 18512 36048 18564 36100
rect 19432 36048 19484 36100
rect 18236 36023 18288 36032
rect 18236 35989 18245 36023
rect 18245 35989 18279 36023
rect 18279 35989 18288 36023
rect 18236 35980 18288 35989
rect 19616 36023 19668 36032
rect 19616 35989 19625 36023
rect 19625 35989 19659 36023
rect 19659 35989 19668 36023
rect 19616 35980 19668 35989
rect 20260 35980 20312 36032
rect 10880 35878 10932 35930
rect 10944 35878 10996 35930
rect 11008 35878 11060 35930
rect 11072 35878 11124 35930
rect 11136 35878 11188 35930
rect 20811 35878 20863 35930
rect 20875 35878 20927 35930
rect 20939 35878 20991 35930
rect 21003 35878 21055 35930
rect 21067 35878 21119 35930
rect 5540 35819 5592 35828
rect 1952 35640 2004 35692
rect 3240 35708 3292 35760
rect 5540 35785 5549 35819
rect 5549 35785 5583 35819
rect 5583 35785 5592 35819
rect 5540 35776 5592 35785
rect 7472 35776 7524 35828
rect 8208 35776 8260 35828
rect 9404 35776 9456 35828
rect 10692 35819 10744 35828
rect 9128 35708 9180 35760
rect 5540 35640 5592 35692
rect 7932 35640 7984 35692
rect 8392 35640 8444 35692
rect 10048 35640 10100 35692
rect 10416 35708 10468 35760
rect 10692 35785 10701 35819
rect 10701 35785 10735 35819
rect 10735 35785 10744 35819
rect 10692 35776 10744 35785
rect 10232 35683 10284 35692
rect 10232 35649 10241 35683
rect 10241 35649 10275 35683
rect 10275 35649 10284 35683
rect 10600 35708 10652 35760
rect 10232 35640 10284 35649
rect 11980 35640 12032 35692
rect 13268 35776 13320 35828
rect 19432 35776 19484 35828
rect 20260 35776 20312 35828
rect 20720 35776 20772 35828
rect 21180 35776 21232 35828
rect 15752 35708 15804 35760
rect 12808 35683 12860 35692
rect 12808 35649 12815 35683
rect 12815 35649 12860 35683
rect 12808 35640 12860 35649
rect 2228 35479 2280 35488
rect 2228 35445 2237 35479
rect 2237 35445 2271 35479
rect 2271 35445 2280 35479
rect 2228 35436 2280 35445
rect 3792 35436 3844 35488
rect 4896 35436 4948 35488
rect 6276 35436 6328 35488
rect 10508 35504 10560 35556
rect 8484 35436 8536 35488
rect 10140 35436 10192 35488
rect 12900 35504 12952 35556
rect 12716 35436 12768 35488
rect 13084 35683 13136 35692
rect 13084 35649 13098 35683
rect 13098 35649 13132 35683
rect 13132 35649 13136 35683
rect 13084 35640 13136 35649
rect 16580 35640 16632 35692
rect 18236 35640 18288 35692
rect 18420 35683 18472 35692
rect 18420 35649 18454 35683
rect 18454 35649 18472 35683
rect 20260 35683 20312 35692
rect 18420 35640 18472 35649
rect 20260 35649 20269 35683
rect 20269 35649 20303 35683
rect 20303 35649 20312 35683
rect 20260 35640 20312 35649
rect 20628 35640 20680 35692
rect 16672 35572 16724 35624
rect 16948 35615 17000 35624
rect 16948 35581 16957 35615
rect 16957 35581 16991 35615
rect 16991 35581 17000 35615
rect 16948 35572 17000 35581
rect 14372 35436 14424 35488
rect 17316 35436 17368 35488
rect 5915 35334 5967 35386
rect 5979 35334 6031 35386
rect 6043 35334 6095 35386
rect 6107 35334 6159 35386
rect 6171 35334 6223 35386
rect 15846 35334 15898 35386
rect 15910 35334 15962 35386
rect 15974 35334 16026 35386
rect 16038 35334 16090 35386
rect 16102 35334 16154 35386
rect 25776 35334 25828 35386
rect 25840 35334 25892 35386
rect 25904 35334 25956 35386
rect 25968 35334 26020 35386
rect 26032 35334 26084 35386
rect 2228 35275 2280 35284
rect 2228 35241 2237 35275
rect 2237 35241 2271 35275
rect 2271 35241 2280 35275
rect 2228 35232 2280 35241
rect 3516 35232 3568 35284
rect 5632 35232 5684 35284
rect 8024 35232 8076 35284
rect 8392 35275 8444 35284
rect 8392 35241 8401 35275
rect 8401 35241 8435 35275
rect 8435 35241 8444 35275
rect 8392 35232 8444 35241
rect 10324 35232 10376 35284
rect 12900 35232 12952 35284
rect 16580 35275 16632 35284
rect 1952 35164 2004 35216
rect 3792 35139 3844 35148
rect 3792 35105 3801 35139
rect 3801 35105 3835 35139
rect 3835 35105 3844 35139
rect 3792 35096 3844 35105
rect 8300 35164 8352 35216
rect 8852 35164 8904 35216
rect 15200 35164 15252 35216
rect 16580 35241 16589 35275
rect 16589 35241 16623 35275
rect 16623 35241 16632 35275
rect 16580 35232 16632 35241
rect 20720 35232 20772 35284
rect 2780 35028 2832 35080
rect 4436 35028 4488 35080
rect 6644 35071 6696 35080
rect 6644 35037 6653 35071
rect 6653 35037 6687 35071
rect 6687 35037 6696 35071
rect 7656 35071 7708 35080
rect 6644 35028 6696 35037
rect 7656 35037 7665 35071
rect 7665 35037 7699 35071
rect 7699 35037 7708 35071
rect 7656 35028 7708 35037
rect 9956 35096 10008 35148
rect 10508 35096 10560 35148
rect 15384 35139 15436 35148
rect 15384 35105 15393 35139
rect 15393 35105 15427 35139
rect 15427 35105 15436 35139
rect 15384 35096 15436 35105
rect 17224 35164 17276 35216
rect 16304 35096 16356 35148
rect 17316 35139 17368 35148
rect 17316 35105 17325 35139
rect 17325 35105 17359 35139
rect 17359 35105 17368 35139
rect 17316 35096 17368 35105
rect 4068 35003 4120 35012
rect 4068 34969 4102 35003
rect 4102 34969 4120 35003
rect 4068 34960 4120 34969
rect 3056 34935 3108 34944
rect 3056 34901 3065 34935
rect 3065 34901 3099 34935
rect 3099 34901 3108 34935
rect 3056 34892 3108 34901
rect 3792 34892 3844 34944
rect 7932 34960 7984 35012
rect 8208 35071 8260 35080
rect 8208 35037 8234 35071
rect 8234 35037 8260 35071
rect 8208 35028 8260 35037
rect 8760 35028 8812 35080
rect 10784 35071 10836 35080
rect 10784 35037 10793 35071
rect 10793 35037 10827 35071
rect 10827 35037 10836 35071
rect 10784 35028 10836 35037
rect 11612 35028 11664 35080
rect 14648 35028 14700 35080
rect 12072 34960 12124 35012
rect 8668 34892 8720 34944
rect 13728 34960 13780 35012
rect 14464 34960 14516 35012
rect 15660 35071 15712 35080
rect 15660 35037 15669 35071
rect 15669 35037 15703 35071
rect 15703 35037 15712 35071
rect 15936 35071 15988 35080
rect 15660 35028 15712 35037
rect 15936 35037 15945 35071
rect 15945 35037 15979 35071
rect 15979 35037 15988 35071
rect 15936 35028 15988 35037
rect 18512 34960 18564 35012
rect 20444 35028 20496 35080
rect 22192 35028 22244 35080
rect 30104 35071 30156 35080
rect 20628 34960 20680 35012
rect 14648 34892 14700 34944
rect 14924 34892 14976 34944
rect 15660 34892 15712 34944
rect 17408 34935 17460 34944
rect 17408 34901 17417 34935
rect 17417 34901 17451 34935
rect 17451 34901 17460 34935
rect 17408 34892 17460 34901
rect 18328 34892 18380 34944
rect 18604 34935 18656 34944
rect 18604 34901 18613 34935
rect 18613 34901 18647 34935
rect 18647 34901 18656 34935
rect 18604 34892 18656 34901
rect 19984 34892 20036 34944
rect 21916 34935 21968 34944
rect 21916 34901 21925 34935
rect 21925 34901 21959 34935
rect 21959 34901 21968 34935
rect 21916 34892 21968 34901
rect 30104 35037 30113 35071
rect 30113 35037 30147 35071
rect 30147 35037 30156 35071
rect 30104 35028 30156 35037
rect 10880 34790 10932 34842
rect 10944 34790 10996 34842
rect 11008 34790 11060 34842
rect 11072 34790 11124 34842
rect 11136 34790 11188 34842
rect 20811 34790 20863 34842
rect 20875 34790 20927 34842
rect 20939 34790 20991 34842
rect 21003 34790 21055 34842
rect 21067 34790 21119 34842
rect 1860 34688 1912 34740
rect 4068 34688 4120 34740
rect 4436 34731 4488 34740
rect 4436 34697 4445 34731
rect 4445 34697 4479 34731
rect 4479 34697 4488 34731
rect 4436 34688 4488 34697
rect 5816 34688 5868 34740
rect 6828 34688 6880 34740
rect 4712 34620 4764 34672
rect 1952 34552 2004 34604
rect 3424 34595 3476 34604
rect 3424 34561 3433 34595
rect 3433 34561 3467 34595
rect 3467 34561 3476 34595
rect 3424 34552 3476 34561
rect 3516 34595 3568 34604
rect 3516 34561 3525 34595
rect 3525 34561 3559 34595
rect 3559 34561 3568 34595
rect 3516 34552 3568 34561
rect 3792 34595 3844 34604
rect 3792 34561 3801 34595
rect 3801 34561 3835 34595
rect 3835 34561 3844 34595
rect 3792 34552 3844 34561
rect 5724 34552 5776 34604
rect 6276 34552 6328 34604
rect 7840 34688 7892 34740
rect 8760 34731 8812 34740
rect 8760 34697 8769 34731
rect 8769 34697 8803 34731
rect 8803 34697 8812 34731
rect 8760 34688 8812 34697
rect 13360 34688 13412 34740
rect 16948 34688 17000 34740
rect 17408 34688 17460 34740
rect 12624 34663 12676 34672
rect 12624 34629 12658 34663
rect 12658 34629 12676 34663
rect 12624 34620 12676 34629
rect 8024 34552 8076 34604
rect 8668 34595 8720 34604
rect 8668 34561 8677 34595
rect 8677 34561 8711 34595
rect 8711 34561 8720 34595
rect 8668 34552 8720 34561
rect 3608 34527 3660 34536
rect 3608 34493 3617 34527
rect 3617 34493 3651 34527
rect 3651 34493 3660 34527
rect 3608 34484 3660 34493
rect 4528 34484 4580 34536
rect 7656 34484 7708 34536
rect 8484 34484 8536 34536
rect 8944 34552 8996 34604
rect 11704 34552 11756 34604
rect 13084 34552 13136 34604
rect 14464 34595 14516 34604
rect 14464 34561 14473 34595
rect 14473 34561 14507 34595
rect 14507 34561 14516 34595
rect 14464 34552 14516 34561
rect 15292 34595 15344 34604
rect 18604 34620 18656 34672
rect 19156 34688 19208 34740
rect 20352 34688 20404 34740
rect 20720 34731 20772 34740
rect 20720 34697 20729 34731
rect 20729 34697 20763 34731
rect 20763 34697 20772 34731
rect 20720 34688 20772 34697
rect 21180 34688 21232 34740
rect 20444 34620 20496 34672
rect 20628 34663 20680 34672
rect 20628 34629 20637 34663
rect 20637 34629 20671 34663
rect 20671 34629 20680 34663
rect 20628 34620 20680 34629
rect 15292 34561 15326 34595
rect 15326 34561 15344 34595
rect 15292 34552 15344 34561
rect 18052 34552 18104 34604
rect 19616 34552 19668 34604
rect 20996 34595 21048 34604
rect 20996 34561 21005 34595
rect 21005 34561 21039 34595
rect 21039 34561 21048 34595
rect 20996 34552 21048 34561
rect 9864 34527 9916 34536
rect 9864 34493 9873 34527
rect 9873 34493 9907 34527
rect 9907 34493 9916 34527
rect 9864 34484 9916 34493
rect 10140 34527 10192 34536
rect 10140 34493 10149 34527
rect 10149 34493 10183 34527
rect 10183 34493 10192 34527
rect 10140 34484 10192 34493
rect 10416 34484 10468 34536
rect 11612 34484 11664 34536
rect 14188 34484 14240 34536
rect 14648 34484 14700 34536
rect 15660 34484 15712 34536
rect 15844 34484 15896 34536
rect 17500 34527 17552 34536
rect 17500 34493 17509 34527
rect 17509 34493 17543 34527
rect 17543 34493 17552 34527
rect 17500 34484 17552 34493
rect 20076 34484 20128 34536
rect 2228 34391 2280 34400
rect 2228 34357 2237 34391
rect 2237 34357 2271 34391
rect 2271 34357 2280 34391
rect 2228 34348 2280 34357
rect 7656 34391 7708 34400
rect 7656 34357 7665 34391
rect 7665 34357 7699 34391
rect 7699 34357 7708 34391
rect 7656 34348 7708 34357
rect 9036 34348 9088 34400
rect 15016 34416 15068 34468
rect 19340 34391 19392 34400
rect 19340 34357 19349 34391
rect 19349 34357 19383 34391
rect 19383 34357 19392 34391
rect 19340 34348 19392 34357
rect 19892 34391 19944 34400
rect 19892 34357 19901 34391
rect 19901 34357 19935 34391
rect 19935 34357 19944 34391
rect 19892 34348 19944 34357
rect 21916 34348 21968 34400
rect 5915 34246 5967 34298
rect 5979 34246 6031 34298
rect 6043 34246 6095 34298
rect 6107 34246 6159 34298
rect 6171 34246 6223 34298
rect 15846 34246 15898 34298
rect 15910 34246 15962 34298
rect 15974 34246 16026 34298
rect 16038 34246 16090 34298
rect 16102 34246 16154 34298
rect 25776 34246 25828 34298
rect 25840 34246 25892 34298
rect 25904 34246 25956 34298
rect 25968 34246 26020 34298
rect 26032 34246 26084 34298
rect 2228 34187 2280 34196
rect 2228 34153 2237 34187
rect 2237 34153 2271 34187
rect 2271 34153 2280 34187
rect 2228 34144 2280 34153
rect 3976 34144 4028 34196
rect 5724 34144 5776 34196
rect 8116 34144 8168 34196
rect 1952 34076 2004 34128
rect 3148 33983 3200 33992
rect 3148 33949 3157 33983
rect 3157 33949 3191 33983
rect 3191 33949 3200 33983
rect 3148 33940 3200 33949
rect 3792 33983 3844 33992
rect 3792 33949 3801 33983
rect 3801 33949 3835 33983
rect 3835 33949 3844 33983
rect 3792 33940 3844 33949
rect 4436 33940 4488 33992
rect 7932 34008 7984 34060
rect 5816 33983 5868 33992
rect 5816 33949 5825 33983
rect 5825 33949 5859 33983
rect 5859 33949 5868 33983
rect 5816 33940 5868 33949
rect 2964 33847 3016 33856
rect 2964 33813 2973 33847
rect 2973 33813 3007 33847
rect 3007 33813 3016 33847
rect 2964 33804 3016 33813
rect 3884 33872 3936 33924
rect 4160 33872 4212 33924
rect 6184 33983 6236 33992
rect 6184 33949 6193 33983
rect 6193 33949 6227 33983
rect 6227 33949 6236 33983
rect 6368 33983 6420 33992
rect 6184 33940 6236 33949
rect 6368 33949 6377 33983
rect 6377 33949 6411 33983
rect 6411 33949 6420 33983
rect 6368 33940 6420 33949
rect 6736 33940 6788 33992
rect 7012 33983 7064 33992
rect 7012 33949 7021 33983
rect 7021 33949 7055 33983
rect 7055 33949 7064 33983
rect 7012 33940 7064 33949
rect 8116 33983 8168 33992
rect 8116 33949 8125 33983
rect 8125 33949 8159 33983
rect 8159 33949 8168 33983
rect 8116 33940 8168 33949
rect 8944 34144 8996 34196
rect 9864 34144 9916 34196
rect 18052 34187 18104 34196
rect 8300 34076 8352 34128
rect 9772 34076 9824 34128
rect 8944 34008 8996 34060
rect 15200 34076 15252 34128
rect 15752 34076 15804 34128
rect 18052 34153 18061 34187
rect 18061 34153 18095 34187
rect 18095 34153 18104 34187
rect 18052 34144 18104 34153
rect 20076 34144 20128 34196
rect 20812 34076 20864 34128
rect 22008 34076 22060 34128
rect 8484 33940 8536 33992
rect 9312 33983 9364 33992
rect 9312 33949 9321 33983
rect 9321 33949 9355 33983
rect 9355 33949 9364 33983
rect 9312 33940 9364 33949
rect 19984 34051 20036 34060
rect 19984 34017 19993 34051
rect 19993 34017 20027 34051
rect 20027 34017 20036 34051
rect 19984 34008 20036 34017
rect 8300 33872 8352 33924
rect 11520 33940 11572 33992
rect 11980 33940 12032 33992
rect 9588 33872 9640 33924
rect 10416 33872 10468 33924
rect 11244 33872 11296 33924
rect 11428 33872 11480 33924
rect 14004 33872 14056 33924
rect 14372 33915 14424 33924
rect 14372 33881 14406 33915
rect 14406 33881 14424 33915
rect 14372 33872 14424 33881
rect 14556 33872 14608 33924
rect 18604 33940 18656 33992
rect 19432 33940 19484 33992
rect 19616 33940 19668 33992
rect 19800 33940 19852 33992
rect 20168 34008 20220 34060
rect 20352 33940 20404 33992
rect 18236 33872 18288 33924
rect 5172 33847 5224 33856
rect 5172 33813 5181 33847
rect 5181 33813 5215 33847
rect 5215 33813 5224 33847
rect 5172 33804 5224 33813
rect 7288 33804 7340 33856
rect 8116 33804 8168 33856
rect 9036 33804 9088 33856
rect 9496 33847 9548 33856
rect 9496 33813 9505 33847
rect 9505 33813 9539 33847
rect 9539 33813 9548 33847
rect 9496 33804 9548 33813
rect 10324 33804 10376 33856
rect 10784 33804 10836 33856
rect 15384 33804 15436 33856
rect 19064 33804 19116 33856
rect 20076 33804 20128 33856
rect 20812 33940 20864 33992
rect 20996 33940 21048 33992
rect 21732 33983 21784 33992
rect 20720 33872 20772 33924
rect 21732 33949 21741 33983
rect 21741 33949 21775 33983
rect 21775 33949 21784 33983
rect 21732 33940 21784 33949
rect 21180 33804 21232 33856
rect 22376 33804 22428 33856
rect 10880 33702 10932 33754
rect 10944 33702 10996 33754
rect 11008 33702 11060 33754
rect 11072 33702 11124 33754
rect 11136 33702 11188 33754
rect 20811 33702 20863 33754
rect 20875 33702 20927 33754
rect 20939 33702 20991 33754
rect 21003 33702 21055 33754
rect 21067 33702 21119 33754
rect 3792 33600 3844 33652
rect 5540 33643 5592 33652
rect 5540 33609 5549 33643
rect 5549 33609 5583 33643
rect 5583 33609 5592 33643
rect 5540 33600 5592 33609
rect 8392 33600 8444 33652
rect 2872 33532 2924 33584
rect 3240 33507 3292 33516
rect 3240 33473 3249 33507
rect 3249 33473 3283 33507
rect 3283 33473 3292 33507
rect 3240 33464 3292 33473
rect 3884 33464 3936 33516
rect 5172 33532 5224 33584
rect 4344 33507 4396 33516
rect 4344 33473 4353 33507
rect 4353 33473 4387 33507
rect 4387 33473 4396 33507
rect 4344 33464 4396 33473
rect 4528 33507 4580 33516
rect 4528 33473 4537 33507
rect 4537 33473 4571 33507
rect 4571 33473 4580 33507
rect 4528 33464 4580 33473
rect 6276 33464 6328 33516
rect 7012 33532 7064 33584
rect 7656 33532 7708 33584
rect 9312 33532 9364 33584
rect 9496 33532 9548 33584
rect 11520 33600 11572 33652
rect 12072 33643 12124 33652
rect 12072 33609 12081 33643
rect 12081 33609 12115 33643
rect 12115 33609 12124 33643
rect 12072 33600 12124 33609
rect 3608 33396 3660 33448
rect 4160 33439 4212 33448
rect 4160 33405 4169 33439
rect 4169 33405 4203 33439
rect 4203 33405 4212 33439
rect 4160 33396 4212 33405
rect 3516 33328 3568 33380
rect 4344 33328 4396 33380
rect 8208 33464 8260 33516
rect 8392 33439 8444 33448
rect 8392 33405 8401 33439
rect 8401 33405 8435 33439
rect 8435 33405 8444 33439
rect 8392 33396 8444 33405
rect 8576 33464 8628 33516
rect 9772 33507 9824 33516
rect 9772 33473 9781 33507
rect 9781 33473 9815 33507
rect 9815 33473 9824 33507
rect 9772 33464 9824 33473
rect 9956 33507 10008 33516
rect 9956 33473 9965 33507
rect 9965 33473 9999 33507
rect 9999 33473 10008 33507
rect 9956 33464 10008 33473
rect 10140 33507 10192 33516
rect 10140 33473 10149 33507
rect 10149 33473 10183 33507
rect 10183 33473 10192 33507
rect 10140 33464 10192 33473
rect 10416 33464 10468 33516
rect 11428 33532 11480 33584
rect 11704 33464 11756 33516
rect 11888 33507 11940 33516
rect 11888 33473 11897 33507
rect 11897 33473 11931 33507
rect 11931 33473 11940 33507
rect 11888 33464 11940 33473
rect 12072 33507 12124 33516
rect 12072 33473 12081 33507
rect 12081 33473 12115 33507
rect 12115 33473 12124 33507
rect 12072 33464 12124 33473
rect 8944 33396 8996 33448
rect 10048 33439 10100 33448
rect 10048 33405 10057 33439
rect 10057 33405 10091 33439
rect 10091 33405 10100 33439
rect 10048 33396 10100 33405
rect 14004 33532 14056 33584
rect 14280 33507 14332 33516
rect 14280 33473 14298 33507
rect 14298 33473 14332 33507
rect 14280 33464 14332 33473
rect 14556 33507 14608 33516
rect 14556 33473 14565 33507
rect 14565 33473 14599 33507
rect 14599 33473 14608 33507
rect 14556 33464 14608 33473
rect 12808 33396 12860 33448
rect 8760 33328 8812 33380
rect 15384 33464 15436 33516
rect 18420 33600 18472 33652
rect 18604 33600 18656 33652
rect 19156 33600 19208 33652
rect 21732 33600 21784 33652
rect 18236 33507 18288 33516
rect 18236 33473 18245 33507
rect 18245 33473 18279 33507
rect 18279 33473 18288 33507
rect 18236 33464 18288 33473
rect 19340 33532 19392 33584
rect 19708 33532 19760 33584
rect 19064 33507 19116 33516
rect 19064 33473 19070 33507
rect 19070 33473 19104 33507
rect 19104 33473 19116 33507
rect 19064 33464 19116 33473
rect 19432 33507 19484 33516
rect 19432 33473 19441 33507
rect 19441 33473 19475 33507
rect 19475 33473 19484 33507
rect 19432 33464 19484 33473
rect 19892 33464 19944 33516
rect 20352 33464 20404 33516
rect 22376 33507 22428 33516
rect 20536 33396 20588 33448
rect 22376 33473 22385 33507
rect 22385 33473 22419 33507
rect 22419 33473 22428 33507
rect 22376 33464 22428 33473
rect 30104 33507 30156 33516
rect 30104 33473 30113 33507
rect 30113 33473 30147 33507
rect 30147 33473 30156 33507
rect 30104 33464 30156 33473
rect 20812 33439 20864 33448
rect 20812 33405 20821 33439
rect 20821 33405 20855 33439
rect 20855 33405 20864 33439
rect 20812 33396 20864 33405
rect 21180 33396 21232 33448
rect 21272 33328 21324 33380
rect 1492 33303 1544 33312
rect 1492 33269 1501 33303
rect 1501 33269 1535 33303
rect 1535 33269 1544 33303
rect 1492 33260 1544 33269
rect 6736 33260 6788 33312
rect 7104 33303 7156 33312
rect 7104 33269 7113 33303
rect 7113 33269 7147 33303
rect 7147 33269 7156 33303
rect 7104 33260 7156 33269
rect 7932 33303 7984 33312
rect 7932 33269 7941 33303
rect 7941 33269 7975 33303
rect 7975 33269 7984 33303
rect 7932 33260 7984 33269
rect 10692 33260 10744 33312
rect 11336 33260 11388 33312
rect 13820 33260 13872 33312
rect 14372 33260 14424 33312
rect 16856 33303 16908 33312
rect 16856 33269 16865 33303
rect 16865 33269 16899 33303
rect 16899 33269 16908 33303
rect 16856 33260 16908 33269
rect 16948 33260 17000 33312
rect 21824 33260 21876 33312
rect 22560 33303 22612 33312
rect 22560 33269 22569 33303
rect 22569 33269 22603 33303
rect 22603 33269 22612 33303
rect 22560 33260 22612 33269
rect 29920 33303 29972 33312
rect 29920 33269 29929 33303
rect 29929 33269 29963 33303
rect 29963 33269 29972 33303
rect 29920 33260 29972 33269
rect 5915 33158 5967 33210
rect 5979 33158 6031 33210
rect 6043 33158 6095 33210
rect 6107 33158 6159 33210
rect 6171 33158 6223 33210
rect 15846 33158 15898 33210
rect 15910 33158 15962 33210
rect 15974 33158 16026 33210
rect 16038 33158 16090 33210
rect 16102 33158 16154 33210
rect 25776 33158 25828 33210
rect 25840 33158 25892 33210
rect 25904 33158 25956 33210
rect 25968 33158 26020 33210
rect 26032 33158 26084 33210
rect 4712 33099 4764 33108
rect 4712 33065 4721 33099
rect 4721 33065 4755 33099
rect 4755 33065 4764 33099
rect 4712 33056 4764 33065
rect 4620 32988 4672 33040
rect 6368 32988 6420 33040
rect 8300 33056 8352 33108
rect 10048 33056 10100 33108
rect 11244 33056 11296 33108
rect 9956 32988 10008 33040
rect 6828 32920 6880 32972
rect 9680 32920 9732 32972
rect 15384 33056 15436 33108
rect 15476 33056 15528 33108
rect 19616 33056 19668 33108
rect 20352 33099 20404 33108
rect 20352 33065 20361 33099
rect 20361 33065 20395 33099
rect 20395 33065 20404 33099
rect 20352 33056 20404 33065
rect 20720 33099 20772 33108
rect 20720 33065 20729 33099
rect 20729 33065 20763 33099
rect 20763 33065 20772 33099
rect 20720 33056 20772 33065
rect 16856 32920 16908 32972
rect 20444 32963 20496 32972
rect 20444 32929 20453 32963
rect 20453 32929 20487 32963
rect 20487 32929 20496 32963
rect 20444 32920 20496 32929
rect 1400 32895 1452 32904
rect 1400 32861 1409 32895
rect 1409 32861 1443 32895
rect 1443 32861 1452 32895
rect 1400 32852 1452 32861
rect 2320 32895 2372 32904
rect 2320 32861 2329 32895
rect 2329 32861 2363 32895
rect 2363 32861 2372 32895
rect 2320 32852 2372 32861
rect 3240 32852 3292 32904
rect 4068 32895 4120 32904
rect 4068 32861 4077 32895
rect 4077 32861 4111 32895
rect 4111 32861 4120 32895
rect 4068 32852 4120 32861
rect 4896 32895 4948 32904
rect 4896 32861 4905 32895
rect 4905 32861 4939 32895
rect 4939 32861 4948 32895
rect 4896 32852 4948 32861
rect 5724 32784 5776 32836
rect 6920 32852 6972 32904
rect 7288 32895 7340 32904
rect 7288 32861 7322 32895
rect 7322 32861 7340 32895
rect 7288 32852 7340 32861
rect 9312 32852 9364 32904
rect 9588 32852 9640 32904
rect 9956 32895 10008 32904
rect 9956 32861 9965 32895
rect 9965 32861 9999 32895
rect 9999 32861 10008 32895
rect 9956 32852 10008 32861
rect 10324 32895 10376 32904
rect 10324 32861 10333 32895
rect 10333 32861 10367 32895
rect 10367 32861 10376 32895
rect 10324 32852 10376 32861
rect 11612 32895 11664 32904
rect 7104 32784 7156 32836
rect 11612 32861 11621 32895
rect 11621 32861 11655 32895
rect 11655 32861 11664 32895
rect 11612 32852 11664 32861
rect 18880 32852 18932 32904
rect 19800 32852 19852 32904
rect 1584 32759 1636 32768
rect 1584 32725 1593 32759
rect 1593 32725 1627 32759
rect 1627 32725 1636 32759
rect 1584 32716 1636 32725
rect 2136 32759 2188 32768
rect 2136 32725 2145 32759
rect 2145 32725 2179 32759
rect 2179 32725 2188 32759
rect 2136 32716 2188 32725
rect 2596 32716 2648 32768
rect 4252 32759 4304 32768
rect 4252 32725 4261 32759
rect 4261 32725 4295 32759
rect 4295 32725 4304 32759
rect 4252 32716 4304 32725
rect 7380 32716 7432 32768
rect 11980 32784 12032 32836
rect 15752 32784 15804 32836
rect 17960 32784 18012 32836
rect 22284 32895 22336 32904
rect 22284 32861 22293 32895
rect 22293 32861 22327 32895
rect 22327 32861 22336 32895
rect 22284 32852 22336 32861
rect 29920 32852 29972 32904
rect 10784 32716 10836 32768
rect 12900 32716 12952 32768
rect 18420 32759 18472 32768
rect 18420 32725 18429 32759
rect 18429 32725 18463 32759
rect 18463 32725 18472 32759
rect 18420 32716 18472 32725
rect 19892 32716 19944 32768
rect 22100 32759 22152 32768
rect 22100 32725 22109 32759
rect 22109 32725 22143 32759
rect 22143 32725 22152 32759
rect 22100 32716 22152 32725
rect 10880 32614 10932 32666
rect 10944 32614 10996 32666
rect 11008 32614 11060 32666
rect 11072 32614 11124 32666
rect 11136 32614 11188 32666
rect 20811 32614 20863 32666
rect 20875 32614 20927 32666
rect 20939 32614 20991 32666
rect 21003 32614 21055 32666
rect 21067 32614 21119 32666
rect 3976 32512 4028 32564
rect 6920 32555 6972 32564
rect 6920 32521 6929 32555
rect 6929 32521 6963 32555
rect 6963 32521 6972 32555
rect 6920 32512 6972 32521
rect 8760 32555 8812 32564
rect 8760 32521 8769 32555
rect 8769 32521 8803 32555
rect 8803 32521 8812 32555
rect 8760 32512 8812 32521
rect 9772 32512 9824 32564
rect 10784 32512 10836 32564
rect 12992 32512 13044 32564
rect 13268 32512 13320 32564
rect 14648 32512 14700 32564
rect 15752 32555 15804 32564
rect 15752 32521 15761 32555
rect 15761 32521 15795 32555
rect 15795 32521 15804 32555
rect 15752 32512 15804 32521
rect 17960 32555 18012 32564
rect 17960 32521 17969 32555
rect 17969 32521 18003 32555
rect 18003 32521 18012 32555
rect 17960 32512 18012 32521
rect 7932 32444 7984 32496
rect 10692 32487 10744 32496
rect 10692 32453 10710 32487
rect 10710 32453 10744 32487
rect 10692 32444 10744 32453
rect 2136 32376 2188 32428
rect 3700 32376 3752 32428
rect 4528 32376 4580 32428
rect 6736 32419 6788 32428
rect 6736 32385 6745 32419
rect 6745 32385 6779 32419
rect 6779 32385 6788 32419
rect 6736 32376 6788 32385
rect 7380 32419 7432 32428
rect 7380 32385 7389 32419
rect 7389 32385 7423 32419
rect 7423 32385 7432 32419
rect 7380 32376 7432 32385
rect 15476 32487 15528 32496
rect 15476 32453 15485 32487
rect 15485 32453 15519 32487
rect 15519 32453 15528 32487
rect 15476 32444 15528 32453
rect 12256 32376 12308 32428
rect 14648 32376 14700 32428
rect 2780 32308 2832 32360
rect 11612 32351 11664 32360
rect 11612 32317 11621 32351
rect 11621 32317 11655 32351
rect 11655 32317 11664 32351
rect 11612 32308 11664 32317
rect 15384 32419 15436 32428
rect 15384 32385 15393 32419
rect 15393 32385 15427 32419
rect 15427 32385 15436 32419
rect 15384 32376 15436 32385
rect 15752 32376 15804 32428
rect 16580 32376 16632 32428
rect 17224 32419 17276 32428
rect 17224 32385 17233 32419
rect 17233 32385 17267 32419
rect 17267 32385 17276 32419
rect 17224 32376 17276 32385
rect 18052 32444 18104 32496
rect 18420 32512 18472 32564
rect 20536 32555 20588 32564
rect 20536 32521 20561 32555
rect 20561 32521 20588 32555
rect 20536 32512 20588 32521
rect 17132 32308 17184 32360
rect 17868 32308 17920 32360
rect 18052 32308 18104 32360
rect 18788 32444 18840 32496
rect 20352 32487 20404 32496
rect 18880 32376 18932 32428
rect 20352 32453 20361 32487
rect 20361 32453 20395 32487
rect 20395 32453 20404 32487
rect 20352 32444 20404 32453
rect 19800 32419 19852 32428
rect 19800 32385 19809 32419
rect 19809 32385 19843 32419
rect 19843 32385 19852 32419
rect 19800 32376 19852 32385
rect 19984 32376 20036 32428
rect 20628 32376 20680 32428
rect 2228 32215 2280 32224
rect 2228 32181 2237 32215
rect 2237 32181 2271 32215
rect 2271 32181 2280 32215
rect 2228 32172 2280 32181
rect 3056 32172 3108 32224
rect 5724 32172 5776 32224
rect 10048 32172 10100 32224
rect 12716 32172 12768 32224
rect 14188 32240 14240 32292
rect 17408 32240 17460 32292
rect 29828 32308 29880 32360
rect 13820 32172 13872 32224
rect 15108 32172 15160 32224
rect 17868 32172 17920 32224
rect 20260 32240 20312 32292
rect 19064 32215 19116 32224
rect 19064 32181 19073 32215
rect 19073 32181 19107 32215
rect 19107 32181 19116 32215
rect 19064 32172 19116 32181
rect 19616 32215 19668 32224
rect 19616 32181 19625 32215
rect 19625 32181 19659 32215
rect 19659 32181 19668 32215
rect 19616 32172 19668 32181
rect 20628 32172 20680 32224
rect 21640 32172 21692 32224
rect 5915 32070 5967 32122
rect 5979 32070 6031 32122
rect 6043 32070 6095 32122
rect 6107 32070 6159 32122
rect 6171 32070 6223 32122
rect 15846 32070 15898 32122
rect 15910 32070 15962 32122
rect 15974 32070 16026 32122
rect 16038 32070 16090 32122
rect 16102 32070 16154 32122
rect 25776 32070 25828 32122
rect 25840 32070 25892 32122
rect 25904 32070 25956 32122
rect 25968 32070 26020 32122
rect 26032 32070 26084 32122
rect 2780 32011 2832 32020
rect 2780 31977 2789 32011
rect 2789 31977 2823 32011
rect 2823 31977 2832 32011
rect 2780 31968 2832 31977
rect 3700 31968 3752 32020
rect 4252 31968 4304 32020
rect 3056 31832 3108 31884
rect 4160 31875 4212 31884
rect 4160 31841 4169 31875
rect 4169 31841 4203 31875
rect 4203 31841 4212 31875
rect 4160 31832 4212 31841
rect 2596 31807 2648 31816
rect 2596 31773 2605 31807
rect 2605 31773 2639 31807
rect 2639 31773 2648 31807
rect 2596 31764 2648 31773
rect 3976 31807 4028 31816
rect 3976 31773 3985 31807
rect 3985 31773 4019 31807
rect 4019 31773 4028 31807
rect 3976 31764 4028 31773
rect 4252 31807 4304 31816
rect 4252 31773 4261 31807
rect 4261 31773 4295 31807
rect 4295 31773 4304 31807
rect 4252 31764 4304 31773
rect 4528 31807 4580 31816
rect 4528 31773 4537 31807
rect 4537 31773 4571 31807
rect 4571 31773 4580 31807
rect 4528 31764 4580 31773
rect 4620 31764 4672 31816
rect 6460 31807 6512 31816
rect 6460 31773 6469 31807
rect 6469 31773 6503 31807
rect 6503 31773 6512 31807
rect 6460 31764 6512 31773
rect 6828 31764 6880 31816
rect 9864 31968 9916 32020
rect 9680 31832 9732 31884
rect 10232 31832 10284 31884
rect 11244 31875 11296 31884
rect 11244 31841 11253 31875
rect 11253 31841 11287 31875
rect 11287 31841 11296 31875
rect 11244 31832 11296 31841
rect 13728 31832 13780 31884
rect 13820 31832 13872 31884
rect 9772 31764 9824 31816
rect 10048 31764 10100 31816
rect 10508 31764 10560 31816
rect 11520 31807 11572 31816
rect 11520 31773 11529 31807
rect 11529 31773 11563 31807
rect 11563 31773 11572 31807
rect 11520 31764 11572 31773
rect 12072 31764 12124 31816
rect 14464 31968 14516 32020
rect 15752 31968 15804 32020
rect 17132 31968 17184 32020
rect 19156 31968 19208 32020
rect 19800 32011 19852 32020
rect 15108 31900 15160 31952
rect 18696 31900 18748 31952
rect 14096 31875 14148 31884
rect 14096 31841 14105 31875
rect 14105 31841 14139 31875
rect 14139 31841 14148 31875
rect 14096 31832 14148 31841
rect 17500 31832 17552 31884
rect 4988 31696 5040 31748
rect 9496 31696 9548 31748
rect 15384 31764 15436 31816
rect 17408 31807 17460 31816
rect 17408 31773 17417 31807
rect 17417 31773 17451 31807
rect 17451 31773 17460 31807
rect 17408 31764 17460 31773
rect 18512 31807 18564 31816
rect 18512 31773 18521 31807
rect 18521 31773 18555 31807
rect 18555 31773 18564 31807
rect 18512 31764 18564 31773
rect 19432 31764 19484 31816
rect 1492 31671 1544 31680
rect 1492 31637 1501 31671
rect 1501 31637 1535 31671
rect 1535 31637 1544 31671
rect 1492 31628 1544 31637
rect 6368 31671 6420 31680
rect 6368 31637 6377 31671
rect 6377 31637 6411 31671
rect 6411 31637 6420 31671
rect 6368 31628 6420 31637
rect 7748 31671 7800 31680
rect 7748 31637 7757 31671
rect 7757 31637 7791 31671
rect 7791 31637 7800 31671
rect 7748 31628 7800 31637
rect 8852 31628 8904 31680
rect 13820 31696 13872 31748
rect 17592 31739 17644 31748
rect 13912 31628 13964 31680
rect 15476 31671 15528 31680
rect 15476 31637 15485 31671
rect 15485 31637 15519 31671
rect 15519 31637 15528 31671
rect 15476 31628 15528 31637
rect 17592 31705 17601 31739
rect 17601 31705 17635 31739
rect 17635 31705 17644 31739
rect 17592 31696 17644 31705
rect 18972 31696 19024 31748
rect 19800 31977 19809 32011
rect 19809 31977 19843 32011
rect 19843 31977 19852 32011
rect 19800 31968 19852 31977
rect 20352 31968 20404 32020
rect 19984 31900 20036 31952
rect 20260 31900 20312 31952
rect 22008 31875 22060 31884
rect 22008 31841 22017 31875
rect 22017 31841 22051 31875
rect 22051 31841 22060 31875
rect 22008 31832 22060 31841
rect 20352 31764 20404 31816
rect 21180 31764 21232 31816
rect 21456 31628 21508 31680
rect 10880 31526 10932 31578
rect 10944 31526 10996 31578
rect 11008 31526 11060 31578
rect 11072 31526 11124 31578
rect 11136 31526 11188 31578
rect 20811 31526 20863 31578
rect 20875 31526 20927 31578
rect 20939 31526 20991 31578
rect 21003 31526 21055 31578
rect 21067 31526 21119 31578
rect 1400 31467 1452 31476
rect 1400 31433 1409 31467
rect 1409 31433 1443 31467
rect 1443 31433 1452 31467
rect 1400 31424 1452 31433
rect 2228 31424 2280 31476
rect 3240 31424 3292 31476
rect 3884 31424 3936 31476
rect 5080 31424 5132 31476
rect 9680 31424 9732 31476
rect 11612 31424 11664 31476
rect 12256 31467 12308 31476
rect 12256 31433 12265 31467
rect 12265 31433 12299 31467
rect 12299 31433 12308 31467
rect 12256 31424 12308 31433
rect 3240 31331 3292 31340
rect 2136 31220 2188 31272
rect 3240 31297 3249 31331
rect 3249 31297 3283 31331
rect 3283 31297 3292 31331
rect 3240 31288 3292 31297
rect 4160 31356 4212 31408
rect 4988 31356 5040 31408
rect 5264 31356 5316 31408
rect 8576 31356 8628 31408
rect 4528 31288 4580 31340
rect 5356 31288 5408 31340
rect 6276 31288 6328 31340
rect 7748 31331 7800 31340
rect 7748 31297 7757 31331
rect 7757 31297 7791 31331
rect 7791 31297 7800 31331
rect 7748 31288 7800 31297
rect 9404 31288 9456 31340
rect 10324 31288 10376 31340
rect 10876 31331 10928 31340
rect 10876 31297 10885 31331
rect 10885 31297 10919 31331
rect 10919 31297 10928 31331
rect 10876 31288 10928 31297
rect 11520 31331 11572 31340
rect 11520 31297 11529 31331
rect 11529 31297 11563 31331
rect 11563 31297 11572 31331
rect 11520 31288 11572 31297
rect 12808 31356 12860 31408
rect 13820 31424 13872 31476
rect 12716 31288 12768 31340
rect 12992 31331 13044 31340
rect 12992 31297 13001 31331
rect 13001 31297 13035 31331
rect 13035 31297 13044 31331
rect 12992 31288 13044 31297
rect 13084 31331 13136 31340
rect 13084 31297 13094 31331
rect 13094 31297 13128 31331
rect 13128 31297 13136 31331
rect 13084 31288 13136 31297
rect 4344 31220 4396 31272
rect 6368 31220 6420 31272
rect 9312 31220 9364 31272
rect 11796 31263 11848 31272
rect 4620 31152 4672 31204
rect 10048 31152 10100 31204
rect 2320 31084 2372 31136
rect 3700 31127 3752 31136
rect 3700 31093 3709 31127
rect 3709 31093 3743 31127
rect 3743 31093 3752 31127
rect 3700 31084 3752 31093
rect 5816 31084 5868 31136
rect 7012 31084 7064 31136
rect 8116 31084 8168 31136
rect 8576 31127 8628 31136
rect 8576 31093 8585 31127
rect 8585 31093 8619 31127
rect 8619 31093 8628 31127
rect 8576 31084 8628 31093
rect 9864 31084 9916 31136
rect 10692 31084 10744 31136
rect 11796 31229 11805 31263
rect 11805 31229 11839 31263
rect 11839 31229 11848 31263
rect 11796 31220 11848 31229
rect 11704 31152 11756 31204
rect 14004 31288 14056 31340
rect 14556 31424 14608 31476
rect 15384 31467 15436 31476
rect 15384 31433 15393 31467
rect 15393 31433 15427 31467
rect 15427 31433 15436 31467
rect 15384 31424 15436 31433
rect 17868 31467 17920 31476
rect 17868 31433 17877 31467
rect 17877 31433 17911 31467
rect 17911 31433 17920 31467
rect 17868 31424 17920 31433
rect 19064 31424 19116 31476
rect 15568 31356 15620 31408
rect 18512 31356 18564 31408
rect 19524 31424 19576 31476
rect 14464 31331 14516 31340
rect 14464 31297 14473 31331
rect 14473 31297 14507 31331
rect 14507 31297 14516 31331
rect 14464 31288 14516 31297
rect 13728 31220 13780 31272
rect 15200 31288 15252 31340
rect 16304 31288 16356 31340
rect 16672 31331 16724 31340
rect 16672 31297 16681 31331
rect 16681 31297 16715 31331
rect 16715 31297 16724 31331
rect 16672 31288 16724 31297
rect 18696 31331 18748 31340
rect 18696 31297 18705 31331
rect 18705 31297 18739 31331
rect 18739 31297 18748 31331
rect 18696 31288 18748 31297
rect 18880 31331 18932 31340
rect 18880 31297 18889 31331
rect 18889 31297 18923 31331
rect 18923 31297 18932 31331
rect 18880 31288 18932 31297
rect 19156 31288 19208 31340
rect 20352 31288 20404 31340
rect 21456 31356 21508 31408
rect 22100 31356 22152 31408
rect 20720 31331 20772 31340
rect 20720 31297 20729 31331
rect 20729 31297 20763 31331
rect 20763 31297 20772 31331
rect 20720 31288 20772 31297
rect 15476 31152 15528 31204
rect 13820 31084 13872 31136
rect 14464 31084 14516 31136
rect 14740 31127 14792 31136
rect 14740 31093 14749 31127
rect 14749 31093 14783 31127
rect 14783 31093 14792 31127
rect 14740 31084 14792 31093
rect 17224 31084 17276 31136
rect 18420 31084 18472 31136
rect 19616 31220 19668 31272
rect 20812 31220 20864 31272
rect 20996 31263 21048 31272
rect 20996 31229 21005 31263
rect 21005 31229 21039 31263
rect 21039 31229 21048 31263
rect 22008 31288 22060 31340
rect 29828 31331 29880 31340
rect 29828 31297 29837 31331
rect 29837 31297 29871 31331
rect 29871 31297 29880 31331
rect 29828 31288 29880 31297
rect 20996 31220 21048 31229
rect 21732 31220 21784 31272
rect 19156 31152 19208 31204
rect 21180 31152 21232 31204
rect 21456 31152 21508 31204
rect 22284 31220 22336 31272
rect 30104 31263 30156 31272
rect 30104 31229 30113 31263
rect 30113 31229 30147 31263
rect 30147 31229 30156 31263
rect 30104 31220 30156 31229
rect 19616 31084 19668 31136
rect 19984 31127 20036 31136
rect 19984 31093 19993 31127
rect 19993 31093 20027 31127
rect 20027 31093 20036 31127
rect 19984 31084 20036 31093
rect 5915 30982 5967 31034
rect 5979 30982 6031 31034
rect 6043 30982 6095 31034
rect 6107 30982 6159 31034
rect 6171 30982 6223 31034
rect 15846 30982 15898 31034
rect 15910 30982 15962 31034
rect 15974 30982 16026 31034
rect 16038 30982 16090 31034
rect 16102 30982 16154 31034
rect 25776 30982 25828 31034
rect 25840 30982 25892 31034
rect 25904 30982 25956 31034
rect 25968 30982 26020 31034
rect 26032 30982 26084 31034
rect 2136 30812 2188 30864
rect 2320 30880 2372 30932
rect 3056 30923 3108 30932
rect 3056 30889 3065 30923
rect 3065 30889 3099 30923
rect 3099 30889 3108 30923
rect 3056 30880 3108 30889
rect 6276 30880 6328 30932
rect 9864 30923 9916 30932
rect 9864 30889 9873 30923
rect 9873 30889 9907 30923
rect 9907 30889 9916 30923
rect 9864 30880 9916 30889
rect 10876 30880 10928 30932
rect 18512 30923 18564 30932
rect 6460 30812 6512 30864
rect 7104 30855 7156 30864
rect 7104 30821 7113 30855
rect 7113 30821 7147 30855
rect 7147 30821 7156 30855
rect 7104 30812 7156 30821
rect 2964 30676 3016 30728
rect 6368 30787 6420 30796
rect 6368 30753 6377 30787
rect 6377 30753 6411 30787
rect 6411 30753 6420 30787
rect 6368 30744 6420 30753
rect 4896 30719 4948 30728
rect 4896 30685 4905 30719
rect 4905 30685 4939 30719
rect 4939 30685 4948 30719
rect 4896 30676 4948 30685
rect 5264 30719 5316 30728
rect 5264 30685 5273 30719
rect 5273 30685 5307 30719
rect 5307 30685 5316 30719
rect 5264 30676 5316 30685
rect 5356 30676 5408 30728
rect 5816 30608 5868 30660
rect 3976 30583 4028 30592
rect 3976 30549 3985 30583
rect 3985 30549 4019 30583
rect 4019 30549 4028 30583
rect 3976 30540 4028 30549
rect 4712 30583 4764 30592
rect 4712 30549 4721 30583
rect 4721 30549 4755 30583
rect 4755 30549 4764 30583
rect 4712 30540 4764 30549
rect 7012 30608 7064 30660
rect 7380 30676 7432 30728
rect 7472 30719 7524 30728
rect 7472 30685 7481 30719
rect 7481 30685 7515 30719
rect 7515 30685 7524 30719
rect 8852 30812 8904 30864
rect 11244 30812 11296 30864
rect 11980 30855 12032 30864
rect 11980 30821 11989 30855
rect 11989 30821 12023 30855
rect 12023 30821 12032 30855
rect 11980 30812 12032 30821
rect 12440 30812 12492 30864
rect 7472 30676 7524 30685
rect 11888 30744 11940 30796
rect 12072 30744 12124 30796
rect 14280 30812 14332 30864
rect 8300 30676 8352 30728
rect 9956 30676 10008 30728
rect 10140 30676 10192 30728
rect 10692 30719 10744 30728
rect 10692 30685 10701 30719
rect 10701 30685 10735 30719
rect 10735 30685 10744 30719
rect 10692 30676 10744 30685
rect 11428 30719 11480 30728
rect 11428 30685 11437 30719
rect 11437 30685 11471 30719
rect 11471 30685 11480 30719
rect 11428 30676 11480 30685
rect 11704 30676 11756 30728
rect 12900 30676 12952 30728
rect 13084 30676 13136 30728
rect 13268 30719 13320 30728
rect 13268 30685 13277 30719
rect 13277 30685 13311 30719
rect 13311 30685 13320 30719
rect 13268 30676 13320 30685
rect 6460 30540 6512 30592
rect 7472 30540 7524 30592
rect 8944 30583 8996 30592
rect 8944 30549 8953 30583
rect 8953 30549 8987 30583
rect 8987 30549 8996 30583
rect 8944 30540 8996 30549
rect 9404 30540 9456 30592
rect 11520 30608 11572 30660
rect 12256 30608 12308 30660
rect 13728 30676 13780 30728
rect 14464 30719 14516 30728
rect 14464 30685 14473 30719
rect 14473 30685 14507 30719
rect 14507 30685 14516 30719
rect 14464 30676 14516 30685
rect 14556 30719 14608 30728
rect 14556 30685 14601 30719
rect 14601 30685 14608 30719
rect 14556 30676 14608 30685
rect 15108 30676 15160 30728
rect 18512 30889 18521 30923
rect 18521 30889 18555 30923
rect 18555 30889 18564 30923
rect 18512 30880 18564 30889
rect 19800 30880 19852 30932
rect 20996 30880 21048 30932
rect 17592 30812 17644 30864
rect 18420 30787 18472 30796
rect 16212 30651 16264 30660
rect 16212 30617 16221 30651
rect 16221 30617 16255 30651
rect 16255 30617 16264 30651
rect 16212 30608 16264 30617
rect 17132 30719 17184 30728
rect 17132 30685 17141 30719
rect 17141 30685 17175 30719
rect 17175 30685 17184 30719
rect 17132 30676 17184 30685
rect 17040 30608 17092 30660
rect 18420 30753 18429 30787
rect 18429 30753 18463 30787
rect 18463 30753 18472 30787
rect 18420 30744 18472 30753
rect 20812 30812 20864 30864
rect 21548 30812 21600 30864
rect 18788 30744 18840 30796
rect 20720 30744 20772 30796
rect 17500 30719 17552 30728
rect 17500 30685 17509 30719
rect 17509 30685 17543 30719
rect 17543 30685 17552 30719
rect 17500 30676 17552 30685
rect 19064 30676 19116 30728
rect 21272 30719 21324 30728
rect 21272 30685 21281 30719
rect 21281 30685 21315 30719
rect 21315 30685 21324 30719
rect 21272 30676 21324 30685
rect 21640 30719 21692 30728
rect 21640 30685 21649 30719
rect 21649 30685 21683 30719
rect 21683 30685 21692 30719
rect 21640 30676 21692 30685
rect 21824 30719 21876 30728
rect 21824 30685 21833 30719
rect 21833 30685 21867 30719
rect 21867 30685 21876 30719
rect 22008 30719 22060 30728
rect 21824 30676 21876 30685
rect 22008 30685 22017 30719
rect 22017 30685 22051 30719
rect 22051 30685 22060 30719
rect 22008 30676 22060 30685
rect 22376 30676 22428 30728
rect 19156 30608 19208 30660
rect 18052 30540 18104 30592
rect 19892 30608 19944 30660
rect 22652 30651 22704 30660
rect 22652 30617 22661 30651
rect 22661 30617 22695 30651
rect 22695 30617 22704 30651
rect 22652 30608 22704 30617
rect 20536 30540 20588 30592
rect 10880 30438 10932 30490
rect 10944 30438 10996 30490
rect 11008 30438 11060 30490
rect 11072 30438 11124 30490
rect 11136 30438 11188 30490
rect 20811 30438 20863 30490
rect 20875 30438 20927 30490
rect 20939 30438 20991 30490
rect 21003 30438 21055 30490
rect 21067 30438 21119 30490
rect 4620 30379 4672 30388
rect 3700 30268 3752 30320
rect 4620 30345 4629 30379
rect 4629 30345 4663 30379
rect 4663 30345 4672 30379
rect 4620 30336 4672 30345
rect 7380 30336 7432 30388
rect 10784 30336 10836 30388
rect 12072 30336 12124 30388
rect 12808 30336 12860 30388
rect 14556 30336 14608 30388
rect 7104 30268 7156 30320
rect 16212 30336 16264 30388
rect 16672 30379 16724 30388
rect 16672 30345 16681 30379
rect 16681 30345 16715 30379
rect 16715 30345 16724 30379
rect 16672 30336 16724 30345
rect 17500 30336 17552 30388
rect 18328 30311 18380 30320
rect 2136 30200 2188 30252
rect 7196 30200 7248 30252
rect 8760 30200 8812 30252
rect 9680 30200 9732 30252
rect 9864 30243 9916 30252
rect 9864 30209 9898 30243
rect 9898 30209 9916 30243
rect 9864 30200 9916 30209
rect 12072 30200 12124 30252
rect 12716 30200 12768 30252
rect 13728 30200 13780 30252
rect 14096 30200 14148 30252
rect 18328 30277 18337 30311
rect 18337 30277 18371 30311
rect 18371 30277 18380 30311
rect 18328 30268 18380 30277
rect 14740 30200 14792 30252
rect 17316 30200 17368 30252
rect 17408 30200 17460 30252
rect 18696 30200 18748 30252
rect 18972 30200 19024 30252
rect 21272 30336 21324 30388
rect 20720 30268 20772 30320
rect 19984 30243 20036 30252
rect 19984 30209 19993 30243
rect 19993 30209 20027 30243
rect 20027 30209 20036 30243
rect 19984 30200 20036 30209
rect 20536 30200 20588 30252
rect 22376 30200 22428 30252
rect 22652 30243 22704 30252
rect 22652 30209 22653 30243
rect 22653 30209 22687 30243
rect 22687 30209 22704 30243
rect 22652 30200 22704 30209
rect 3240 30175 3292 30184
rect 3240 30141 3249 30175
rect 3249 30141 3283 30175
rect 3283 30141 3292 30175
rect 3240 30132 3292 30141
rect 6368 30175 6420 30184
rect 6368 30141 6377 30175
rect 6377 30141 6411 30175
rect 6411 30141 6420 30175
rect 6368 30132 6420 30141
rect 10692 30064 10744 30116
rect 13176 30064 13228 30116
rect 15568 30107 15620 30116
rect 15568 30073 15577 30107
rect 15577 30073 15611 30107
rect 15611 30073 15620 30107
rect 18328 30132 18380 30184
rect 21824 30132 21876 30184
rect 15568 30064 15620 30073
rect 17776 30064 17828 30116
rect 18880 30064 18932 30116
rect 2320 30039 2372 30048
rect 2320 30005 2329 30039
rect 2329 30005 2363 30039
rect 2363 30005 2372 30039
rect 2320 29996 2372 30005
rect 2504 30039 2556 30048
rect 2504 30005 2513 30039
rect 2513 30005 2547 30039
rect 2547 30005 2556 30039
rect 2504 29996 2556 30005
rect 5816 30039 5868 30048
rect 5816 30005 5825 30039
rect 5825 30005 5859 30039
rect 5859 30005 5868 30039
rect 5816 29996 5868 30005
rect 8208 30039 8260 30048
rect 8208 30005 8217 30039
rect 8217 30005 8251 30039
rect 8251 30005 8260 30039
rect 8208 29996 8260 30005
rect 8576 30039 8628 30048
rect 8576 30005 8585 30039
rect 8585 30005 8619 30039
rect 8619 30005 8628 30039
rect 8576 29996 8628 30005
rect 11612 29996 11664 30048
rect 13084 29996 13136 30048
rect 22008 29996 22060 30048
rect 22192 29996 22244 30048
rect 5915 29894 5967 29946
rect 5979 29894 6031 29946
rect 6043 29894 6095 29946
rect 6107 29894 6159 29946
rect 6171 29894 6223 29946
rect 15846 29894 15898 29946
rect 15910 29894 15962 29946
rect 15974 29894 16026 29946
rect 16038 29894 16090 29946
rect 16102 29894 16154 29946
rect 25776 29894 25828 29946
rect 25840 29894 25892 29946
rect 25904 29894 25956 29946
rect 25968 29894 26020 29946
rect 26032 29894 26084 29946
rect 2320 29792 2372 29844
rect 2136 29724 2188 29776
rect 2964 29792 3016 29844
rect 6368 29792 6420 29844
rect 6644 29792 6696 29844
rect 8852 29792 8904 29844
rect 10784 29792 10836 29844
rect 11336 29792 11388 29844
rect 17132 29792 17184 29844
rect 18420 29792 18472 29844
rect 2872 29724 2924 29776
rect 15108 29724 15160 29776
rect 2504 29656 2556 29708
rect 11428 29656 11480 29708
rect 11612 29656 11664 29708
rect 14096 29699 14148 29708
rect 14096 29665 14105 29699
rect 14105 29665 14139 29699
rect 14139 29665 14148 29699
rect 14096 29656 14148 29665
rect 3976 29588 4028 29640
rect 4160 29631 4212 29640
rect 4160 29597 4169 29631
rect 4169 29597 4203 29631
rect 4203 29597 4212 29631
rect 4160 29588 4212 29597
rect 4712 29588 4764 29640
rect 5264 29588 5316 29640
rect 8944 29588 8996 29640
rect 9772 29588 9824 29640
rect 9956 29588 10008 29640
rect 12532 29588 12584 29640
rect 12808 29588 12860 29640
rect 17316 29588 17368 29640
rect 4896 29520 4948 29572
rect 2136 29452 2188 29504
rect 3608 29452 3660 29504
rect 6552 29520 6604 29572
rect 12072 29563 12124 29572
rect 12072 29529 12081 29563
rect 12081 29529 12115 29563
rect 12115 29529 12124 29563
rect 12072 29520 12124 29529
rect 13176 29520 13228 29572
rect 18328 29724 18380 29776
rect 20536 29724 20588 29776
rect 20628 29724 20680 29776
rect 21548 29792 21600 29844
rect 19892 29656 19944 29708
rect 19340 29588 19392 29640
rect 19984 29631 20036 29640
rect 19984 29597 19993 29631
rect 19993 29597 20027 29631
rect 20027 29597 20036 29631
rect 19984 29588 20036 29597
rect 20720 29588 20772 29640
rect 7656 29452 7708 29504
rect 9128 29452 9180 29504
rect 11704 29452 11756 29504
rect 11980 29495 12032 29504
rect 11980 29461 11989 29495
rect 11989 29461 12023 29495
rect 12023 29461 12032 29495
rect 11980 29452 12032 29461
rect 15476 29495 15528 29504
rect 15476 29461 15485 29495
rect 15485 29461 15519 29495
rect 15519 29461 15528 29495
rect 15476 29452 15528 29461
rect 16948 29452 17000 29504
rect 18328 29520 18380 29572
rect 20260 29520 20312 29572
rect 20536 29520 20588 29572
rect 17408 29452 17460 29504
rect 17960 29452 18012 29504
rect 18236 29452 18288 29504
rect 19892 29452 19944 29504
rect 20168 29495 20220 29504
rect 20168 29461 20177 29495
rect 20177 29461 20211 29495
rect 20211 29461 20220 29495
rect 21824 29631 21876 29640
rect 21824 29597 21833 29631
rect 21833 29597 21867 29631
rect 21867 29597 21876 29631
rect 21824 29588 21876 29597
rect 29736 29588 29788 29640
rect 22100 29520 22152 29572
rect 20168 29452 20220 29461
rect 22468 29495 22520 29504
rect 22468 29461 22477 29495
rect 22477 29461 22511 29495
rect 22511 29461 22520 29495
rect 22468 29452 22520 29461
rect 10880 29350 10932 29402
rect 10944 29350 10996 29402
rect 11008 29350 11060 29402
rect 11072 29350 11124 29402
rect 11136 29350 11188 29402
rect 20811 29350 20863 29402
rect 20875 29350 20927 29402
rect 20939 29350 20991 29402
rect 21003 29350 21055 29402
rect 21067 29350 21119 29402
rect 2780 29248 2832 29300
rect 3240 29248 3292 29300
rect 5264 29291 5316 29300
rect 5264 29257 5273 29291
rect 5273 29257 5307 29291
rect 5307 29257 5316 29291
rect 5264 29248 5316 29257
rect 8576 29248 8628 29300
rect 9128 29291 9180 29300
rect 9128 29257 9137 29291
rect 9137 29257 9171 29291
rect 9171 29257 9180 29291
rect 9128 29248 9180 29257
rect 12072 29248 12124 29300
rect 13176 29291 13228 29300
rect 13176 29257 13185 29291
rect 13185 29257 13219 29291
rect 13219 29257 13228 29291
rect 13176 29248 13228 29257
rect 14648 29291 14700 29300
rect 14648 29257 14657 29291
rect 14657 29257 14691 29291
rect 14691 29257 14700 29291
rect 14648 29248 14700 29257
rect 12716 29180 12768 29232
rect 15476 29180 15528 29232
rect 2136 29155 2188 29164
rect 2136 29121 2145 29155
rect 2145 29121 2179 29155
rect 2179 29121 2188 29155
rect 2136 29112 2188 29121
rect 3608 29155 3660 29164
rect 3608 29121 3617 29155
rect 3617 29121 3651 29155
rect 3651 29121 3660 29155
rect 3608 29112 3660 29121
rect 4068 29112 4120 29164
rect 7012 29155 7064 29164
rect 7012 29121 7021 29155
rect 7021 29121 7055 29155
rect 7055 29121 7064 29155
rect 7012 29112 7064 29121
rect 8208 29112 8260 29164
rect 4712 29044 4764 29096
rect 5540 29044 5592 29096
rect 7196 29087 7248 29096
rect 7196 29053 7205 29087
rect 7205 29053 7239 29087
rect 7239 29053 7248 29087
rect 9220 29087 9272 29096
rect 7196 29044 7248 29053
rect 9220 29053 9229 29087
rect 9229 29053 9263 29087
rect 9263 29053 9272 29087
rect 9220 29044 9272 29053
rect 10048 29112 10100 29164
rect 12532 29112 12584 29164
rect 13452 29155 13504 29164
rect 13452 29121 13461 29155
rect 13461 29121 13495 29155
rect 13495 29121 13504 29155
rect 13452 29112 13504 29121
rect 14740 29155 14792 29164
rect 1492 29019 1544 29028
rect 1492 28985 1501 29019
rect 1501 28985 1535 29019
rect 1535 28985 1544 29019
rect 1492 28976 1544 28985
rect 7840 29019 7892 29028
rect 7840 28985 7849 29019
rect 7849 28985 7883 29019
rect 7883 28985 7892 29019
rect 7840 28976 7892 28985
rect 8392 28976 8444 29028
rect 12532 28976 12584 29028
rect 12808 29044 12860 29096
rect 14740 29121 14749 29155
rect 14749 29121 14783 29155
rect 14783 29121 14792 29155
rect 14740 29112 14792 29121
rect 16948 29180 17000 29232
rect 16672 29155 16724 29164
rect 16672 29121 16681 29155
rect 16681 29121 16715 29155
rect 16715 29121 16724 29155
rect 16672 29112 16724 29121
rect 16856 29155 16908 29164
rect 16856 29121 16865 29155
rect 16865 29121 16899 29155
rect 16899 29121 16908 29155
rect 16856 29112 16908 29121
rect 17132 29248 17184 29300
rect 17408 29180 17460 29232
rect 21824 29248 21876 29300
rect 17224 29155 17276 29164
rect 17224 29121 17233 29155
rect 17233 29121 17267 29155
rect 17267 29121 17276 29155
rect 17224 29112 17276 29121
rect 14004 29044 14056 29096
rect 15108 29044 15160 29096
rect 17776 29112 17828 29164
rect 18052 29155 18104 29164
rect 18052 29121 18061 29155
rect 18061 29121 18095 29155
rect 18095 29121 18104 29155
rect 18052 29112 18104 29121
rect 21548 29180 21600 29232
rect 18328 29155 18380 29164
rect 18328 29121 18337 29155
rect 18337 29121 18371 29155
rect 18371 29121 18380 29155
rect 18328 29112 18380 29121
rect 20168 29112 20220 29164
rect 22468 29112 22520 29164
rect 22560 29112 22612 29164
rect 30196 29112 30248 29164
rect 20536 29087 20588 29096
rect 20536 29053 20545 29087
rect 20545 29053 20579 29087
rect 20579 29053 20588 29087
rect 20536 29044 20588 29053
rect 20628 29087 20680 29096
rect 20628 29053 20637 29087
rect 20637 29053 20671 29087
rect 20671 29053 20680 29087
rect 20628 29044 20680 29053
rect 21456 29044 21508 29096
rect 21732 29044 21784 29096
rect 13176 28976 13228 29028
rect 17868 29019 17920 29028
rect 17868 28985 17877 29019
rect 17877 28985 17911 29019
rect 17911 28985 17920 29019
rect 17868 28976 17920 28985
rect 29828 28976 29880 29028
rect 30012 29019 30064 29028
rect 30012 28985 30021 29019
rect 30021 28985 30055 29019
rect 30055 28985 30064 29019
rect 30012 28976 30064 28985
rect 3792 28908 3844 28960
rect 6644 28951 6696 28960
rect 6644 28917 6653 28951
rect 6653 28917 6687 28951
rect 6687 28917 6696 28951
rect 6644 28908 6696 28917
rect 5915 28806 5967 28858
rect 5979 28806 6031 28858
rect 6043 28806 6095 28858
rect 6107 28806 6159 28858
rect 6171 28806 6223 28858
rect 15846 28806 15898 28858
rect 15910 28806 15962 28858
rect 15974 28806 16026 28858
rect 16038 28806 16090 28858
rect 16102 28806 16154 28858
rect 25776 28806 25828 28858
rect 25840 28806 25892 28858
rect 25904 28806 25956 28858
rect 25968 28806 26020 28858
rect 26032 28806 26084 28858
rect 4160 28704 4212 28756
rect 5540 28704 5592 28756
rect 7012 28704 7064 28756
rect 11336 28747 11388 28756
rect 11336 28713 11345 28747
rect 11345 28713 11379 28747
rect 11379 28713 11388 28747
rect 11336 28704 11388 28713
rect 12624 28704 12676 28756
rect 2596 28543 2648 28552
rect 2596 28509 2605 28543
rect 2605 28509 2639 28543
rect 2639 28509 2648 28543
rect 2596 28500 2648 28509
rect 3792 28543 3844 28552
rect 3792 28509 3801 28543
rect 3801 28509 3835 28543
rect 3835 28509 3844 28543
rect 3792 28500 3844 28509
rect 4988 28543 5040 28552
rect 4988 28509 4997 28543
rect 4997 28509 5031 28543
rect 5031 28509 5040 28543
rect 4988 28500 5040 28509
rect 7564 28636 7616 28688
rect 12440 28636 12492 28688
rect 12716 28636 12768 28688
rect 7196 28568 7248 28620
rect 7472 28568 7524 28620
rect 9680 28568 9732 28620
rect 14648 28704 14700 28756
rect 16856 28704 16908 28756
rect 22008 28704 22060 28756
rect 15108 28636 15160 28688
rect 16212 28636 16264 28688
rect 5816 28500 5868 28552
rect 8392 28500 8444 28552
rect 9312 28500 9364 28552
rect 9496 28500 9548 28552
rect 12808 28543 12860 28552
rect 12808 28509 12818 28543
rect 12818 28509 12852 28543
rect 12852 28509 12860 28543
rect 14464 28568 14516 28620
rect 16948 28611 17000 28620
rect 16948 28577 16957 28611
rect 16957 28577 16991 28611
rect 16991 28577 17000 28611
rect 16948 28568 17000 28577
rect 12808 28500 12860 28509
rect 2136 28432 2188 28484
rect 1492 28407 1544 28416
rect 1492 28373 1501 28407
rect 1501 28373 1535 28407
rect 1535 28373 1544 28407
rect 1492 28364 1544 28373
rect 6828 28407 6880 28416
rect 6828 28373 6837 28407
rect 6837 28373 6871 28407
rect 6871 28373 6880 28407
rect 10324 28432 10376 28484
rect 10416 28432 10468 28484
rect 13084 28475 13136 28484
rect 13084 28441 13093 28475
rect 13093 28441 13127 28475
rect 13127 28441 13136 28475
rect 13084 28432 13136 28441
rect 6828 28364 6880 28373
rect 8024 28407 8076 28416
rect 8024 28373 8033 28407
rect 8033 28373 8067 28407
rect 8067 28373 8076 28407
rect 9036 28407 9088 28416
rect 8024 28364 8076 28373
rect 9036 28373 9045 28407
rect 9045 28373 9079 28407
rect 9079 28373 9088 28407
rect 9036 28364 9088 28373
rect 11244 28364 11296 28416
rect 14004 28432 14056 28484
rect 14740 28500 14792 28552
rect 17684 28568 17736 28620
rect 18052 28611 18104 28620
rect 18052 28577 18061 28611
rect 18061 28577 18095 28611
rect 18095 28577 18104 28611
rect 18052 28568 18104 28577
rect 18144 28568 18196 28620
rect 18328 28568 18380 28620
rect 18420 28500 18472 28552
rect 18880 28500 18932 28552
rect 15200 28475 15252 28484
rect 15200 28441 15209 28475
rect 15209 28441 15243 28475
rect 15243 28441 15252 28475
rect 15200 28432 15252 28441
rect 22100 28500 22152 28552
rect 20536 28432 20588 28484
rect 13360 28407 13412 28416
rect 13360 28373 13369 28407
rect 13369 28373 13403 28407
rect 13403 28373 13412 28407
rect 13360 28364 13412 28373
rect 16856 28407 16908 28416
rect 16856 28373 16865 28407
rect 16865 28373 16899 28407
rect 16899 28373 16908 28407
rect 16856 28364 16908 28373
rect 18052 28364 18104 28416
rect 18512 28364 18564 28416
rect 19708 28364 19760 28416
rect 20444 28364 20496 28416
rect 20628 28407 20680 28416
rect 20628 28373 20637 28407
rect 20637 28373 20671 28407
rect 20671 28373 20680 28407
rect 20628 28364 20680 28373
rect 29092 28364 29144 28416
rect 10880 28262 10932 28314
rect 10944 28262 10996 28314
rect 11008 28262 11060 28314
rect 11072 28262 11124 28314
rect 11136 28262 11188 28314
rect 20811 28262 20863 28314
rect 20875 28262 20927 28314
rect 20939 28262 20991 28314
rect 21003 28262 21055 28314
rect 21067 28262 21119 28314
rect 4712 28203 4764 28212
rect 4712 28169 4721 28203
rect 4721 28169 4755 28203
rect 4755 28169 4764 28203
rect 4712 28160 4764 28169
rect 4988 28160 5040 28212
rect 6828 28203 6880 28212
rect 3884 28135 3936 28144
rect 2136 28067 2188 28076
rect 2136 28033 2145 28067
rect 2145 28033 2179 28067
rect 2179 28033 2188 28067
rect 2136 28024 2188 28033
rect 3884 28101 3893 28135
rect 3893 28101 3927 28135
rect 3927 28101 3936 28135
rect 3884 28092 3936 28101
rect 5356 28092 5408 28144
rect 5724 28092 5776 28144
rect 6828 28169 6837 28203
rect 6837 28169 6871 28203
rect 6871 28169 6880 28203
rect 6828 28160 6880 28169
rect 8024 28160 8076 28212
rect 7196 28092 7248 28144
rect 7288 28092 7340 28144
rect 8760 28160 8812 28212
rect 9220 28203 9272 28212
rect 9220 28169 9229 28203
rect 9229 28169 9263 28203
rect 9263 28169 9272 28203
rect 9220 28160 9272 28169
rect 10324 28203 10376 28212
rect 10324 28169 10333 28203
rect 10333 28169 10367 28203
rect 10367 28169 10376 28203
rect 10324 28160 10376 28169
rect 14464 28203 14516 28212
rect 14464 28169 14473 28203
rect 14473 28169 14507 28203
rect 14507 28169 14516 28203
rect 14464 28160 14516 28169
rect 16672 28160 16724 28212
rect 16856 28160 16908 28212
rect 20536 28203 20588 28212
rect 20536 28169 20545 28203
rect 20545 28169 20579 28203
rect 20579 28169 20588 28203
rect 20536 28160 20588 28169
rect 2596 27956 2648 28008
rect 6644 28024 6696 28076
rect 7012 28067 7064 28076
rect 7012 28033 7021 28067
rect 7021 28033 7055 28067
rect 7055 28033 7064 28067
rect 7012 28024 7064 28033
rect 7932 28024 7984 28076
rect 8116 28024 8168 28076
rect 8208 27956 8260 28008
rect 8484 28067 8536 28076
rect 8484 28033 8493 28067
rect 8493 28033 8527 28067
rect 8527 28033 8536 28067
rect 12808 28092 12860 28144
rect 8484 28024 8536 28033
rect 9036 28067 9088 28076
rect 9036 28033 9045 28067
rect 9045 28033 9079 28067
rect 9079 28033 9088 28067
rect 9036 28024 9088 28033
rect 9128 28024 9180 28076
rect 5632 27931 5684 27940
rect 5632 27897 5641 27931
rect 5641 27897 5675 27931
rect 5675 27897 5684 27931
rect 5632 27888 5684 27897
rect 5816 27888 5868 27940
rect 1492 27863 1544 27872
rect 1492 27829 1501 27863
rect 1501 27829 1535 27863
rect 1535 27829 1544 27863
rect 1492 27820 1544 27829
rect 2872 27863 2924 27872
rect 2872 27829 2881 27863
rect 2881 27829 2915 27863
rect 2915 27829 2924 27863
rect 2872 27820 2924 27829
rect 3700 27820 3752 27872
rect 7380 27820 7432 27872
rect 8116 27888 8168 27940
rect 9312 27956 9364 28008
rect 10048 28067 10100 28076
rect 10048 28033 10057 28067
rect 10057 28033 10091 28067
rect 10091 28033 10100 28067
rect 10048 28024 10100 28033
rect 10232 28024 10284 28076
rect 11336 28024 11388 28076
rect 11612 28024 11664 28076
rect 14096 28092 14148 28144
rect 17592 28092 17644 28144
rect 21916 28160 21968 28212
rect 29736 28160 29788 28212
rect 21272 28092 21324 28144
rect 22008 28135 22060 28144
rect 22008 28101 22017 28135
rect 22017 28101 22051 28135
rect 22051 28101 22060 28135
rect 22008 28092 22060 28101
rect 13360 28067 13412 28076
rect 13360 28033 13394 28067
rect 13394 28033 13412 28067
rect 13360 28024 13412 28033
rect 14648 28024 14700 28076
rect 15752 28067 15804 28076
rect 15752 28033 15761 28067
rect 15761 28033 15795 28067
rect 15795 28033 15804 28067
rect 15752 28024 15804 28033
rect 16212 28024 16264 28076
rect 17408 28067 17460 28076
rect 17408 28033 17417 28067
rect 17417 28033 17451 28067
rect 17451 28033 17460 28067
rect 17408 28024 17460 28033
rect 18328 28024 18380 28076
rect 18696 28067 18748 28076
rect 18696 28033 18705 28067
rect 18705 28033 18739 28067
rect 18739 28033 18748 28067
rect 18972 28067 19024 28076
rect 18696 28024 18748 28033
rect 18972 28033 18981 28067
rect 18981 28033 19015 28067
rect 19015 28033 19024 28067
rect 18972 28024 19024 28033
rect 19340 28024 19392 28076
rect 20720 28067 20772 28076
rect 16396 27956 16448 28008
rect 17684 27956 17736 28008
rect 20720 28033 20729 28067
rect 20729 28033 20763 28067
rect 20763 28033 20772 28067
rect 20720 28024 20772 28033
rect 20812 28067 20864 28076
rect 20812 28033 20821 28067
rect 20821 28033 20855 28067
rect 20855 28033 20864 28067
rect 20812 28024 20864 28033
rect 22100 28024 22152 28076
rect 22376 28024 22428 28076
rect 29828 28067 29880 28076
rect 29828 28033 29837 28067
rect 29837 28033 29871 28067
rect 29871 28033 29880 28067
rect 29828 28024 29880 28033
rect 21548 27956 21600 28008
rect 9496 27888 9548 27940
rect 10968 27888 11020 27940
rect 12164 27931 12216 27940
rect 12164 27897 12173 27931
rect 12173 27897 12207 27931
rect 12207 27897 12216 27931
rect 12164 27888 12216 27897
rect 9128 27820 9180 27872
rect 15292 27820 15344 27872
rect 18420 27863 18472 27872
rect 18420 27829 18429 27863
rect 18429 27829 18463 27863
rect 18463 27829 18472 27863
rect 18420 27820 18472 27829
rect 19432 27820 19484 27872
rect 5915 27718 5967 27770
rect 5979 27718 6031 27770
rect 6043 27718 6095 27770
rect 6107 27718 6159 27770
rect 6171 27718 6223 27770
rect 15846 27718 15898 27770
rect 15910 27718 15962 27770
rect 15974 27718 16026 27770
rect 16038 27718 16090 27770
rect 16102 27718 16154 27770
rect 25776 27718 25828 27770
rect 25840 27718 25892 27770
rect 25904 27718 25956 27770
rect 25968 27718 26020 27770
rect 26032 27718 26084 27770
rect 5816 27659 5868 27668
rect 5816 27625 5825 27659
rect 5825 27625 5859 27659
rect 5859 27625 5868 27659
rect 5816 27616 5868 27625
rect 7012 27616 7064 27668
rect 7380 27616 7432 27668
rect 6552 27591 6604 27600
rect 6552 27557 6561 27591
rect 6561 27557 6595 27591
rect 6595 27557 6604 27591
rect 6552 27548 6604 27557
rect 2596 27455 2648 27464
rect 2596 27421 2605 27455
rect 2605 27421 2639 27455
rect 2639 27421 2648 27455
rect 2596 27412 2648 27421
rect 4344 27412 4396 27464
rect 4896 27344 4948 27396
rect 6736 27387 6788 27396
rect 6736 27353 6745 27387
rect 6745 27353 6779 27387
rect 6779 27353 6788 27387
rect 6736 27344 6788 27353
rect 7104 27412 7156 27464
rect 13636 27616 13688 27668
rect 16212 27616 16264 27668
rect 18972 27616 19024 27668
rect 20812 27616 20864 27668
rect 8392 27548 8444 27600
rect 9496 27548 9548 27600
rect 9864 27548 9916 27600
rect 11244 27548 11296 27600
rect 14280 27548 14332 27600
rect 18696 27548 18748 27600
rect 15660 27480 15712 27532
rect 16396 27480 16448 27532
rect 8668 27412 8720 27464
rect 9036 27412 9088 27464
rect 9312 27455 9364 27464
rect 9312 27421 9319 27455
rect 9319 27421 9364 27455
rect 9312 27412 9364 27421
rect 9680 27412 9732 27464
rect 10232 27412 10284 27464
rect 10324 27412 10376 27464
rect 10968 27455 11020 27464
rect 10968 27421 10977 27455
rect 10977 27421 11011 27455
rect 11011 27421 11020 27455
rect 11428 27455 11480 27464
rect 10968 27412 11020 27421
rect 11428 27421 11437 27455
rect 11437 27421 11471 27455
rect 11471 27421 11480 27455
rect 11428 27412 11480 27421
rect 14372 27455 14424 27464
rect 14372 27421 14381 27455
rect 14381 27421 14415 27455
rect 14415 27421 14424 27455
rect 14372 27412 14424 27421
rect 14556 27412 14608 27464
rect 15292 27455 15344 27464
rect 15292 27421 15301 27455
rect 15301 27421 15335 27455
rect 15335 27421 15344 27455
rect 15292 27412 15344 27421
rect 17408 27480 17460 27532
rect 17684 27480 17736 27532
rect 18972 27480 19024 27532
rect 16856 27412 16908 27464
rect 17500 27412 17552 27464
rect 18144 27455 18196 27464
rect 18144 27421 18153 27455
rect 18153 27421 18187 27455
rect 18187 27421 18196 27455
rect 18144 27412 18196 27421
rect 18512 27455 18564 27464
rect 8576 27344 8628 27396
rect 1676 27276 1728 27328
rect 6276 27276 6328 27328
rect 8392 27276 8444 27328
rect 8852 27276 8904 27328
rect 11520 27344 11572 27396
rect 18512 27421 18521 27455
rect 18521 27421 18555 27455
rect 18555 27421 18564 27455
rect 18512 27412 18564 27421
rect 19064 27412 19116 27464
rect 20720 27548 20772 27600
rect 21180 27548 21232 27600
rect 20812 27523 20864 27532
rect 20812 27489 20821 27523
rect 20821 27489 20855 27523
rect 20855 27489 20864 27523
rect 20812 27480 20864 27489
rect 18788 27344 18840 27396
rect 19156 27344 19208 27396
rect 20536 27344 20588 27396
rect 21272 27412 21324 27464
rect 21548 27455 21600 27464
rect 21548 27421 21557 27455
rect 21557 27421 21591 27455
rect 21591 27421 21600 27455
rect 21548 27412 21600 27421
rect 29368 27412 29420 27464
rect 12716 27276 12768 27328
rect 15568 27319 15620 27328
rect 15568 27285 15577 27319
rect 15577 27285 15611 27319
rect 15611 27285 15620 27319
rect 15568 27276 15620 27285
rect 16672 27276 16724 27328
rect 17408 27319 17460 27328
rect 17408 27285 17417 27319
rect 17417 27285 17451 27319
rect 17451 27285 17460 27319
rect 17408 27276 17460 27285
rect 18512 27276 18564 27328
rect 18604 27276 18656 27328
rect 19064 27276 19116 27328
rect 30012 27319 30064 27328
rect 30012 27285 30021 27319
rect 30021 27285 30055 27319
rect 30055 27285 30064 27319
rect 30012 27276 30064 27285
rect 10880 27174 10932 27226
rect 10944 27174 10996 27226
rect 11008 27174 11060 27226
rect 11072 27174 11124 27226
rect 11136 27174 11188 27226
rect 20811 27174 20863 27226
rect 20875 27174 20927 27226
rect 20939 27174 20991 27226
rect 21003 27174 21055 27226
rect 21067 27174 21119 27226
rect 8208 27072 8260 27124
rect 8392 27072 8444 27124
rect 10324 27072 10376 27124
rect 10692 27072 10744 27124
rect 10784 27072 10836 27124
rect 16672 27115 16724 27124
rect 16672 27081 16681 27115
rect 16681 27081 16715 27115
rect 16715 27081 16724 27115
rect 16672 27072 16724 27081
rect 20536 27115 20588 27124
rect 20536 27081 20545 27115
rect 20545 27081 20579 27115
rect 20579 27081 20588 27115
rect 20536 27072 20588 27081
rect 1676 26979 1728 26988
rect 1676 26945 1685 26979
rect 1685 26945 1719 26979
rect 1719 26945 1728 26979
rect 1676 26936 1728 26945
rect 4344 27004 4396 27056
rect 6736 27004 6788 27056
rect 10416 27004 10468 27056
rect 15568 27004 15620 27056
rect 3608 26979 3660 26988
rect 3608 26945 3642 26979
rect 3642 26945 3660 26979
rect 3608 26936 3660 26945
rect 4988 26936 5040 26988
rect 5816 26936 5868 26988
rect 5448 26911 5500 26920
rect 1492 26843 1544 26852
rect 1492 26809 1501 26843
rect 1501 26809 1535 26843
rect 1535 26809 1544 26843
rect 1492 26800 1544 26809
rect 5448 26877 5457 26911
rect 5457 26877 5491 26911
rect 5491 26877 5500 26911
rect 7564 26936 7616 26988
rect 7932 26936 7984 26988
rect 5448 26868 5500 26877
rect 7380 26868 7432 26920
rect 8116 26868 8168 26920
rect 5724 26800 5776 26852
rect 6276 26800 6328 26852
rect 7932 26800 7984 26852
rect 8024 26800 8076 26852
rect 8944 26936 8996 26988
rect 9772 26979 9824 26988
rect 9772 26945 9806 26979
rect 9806 26945 9824 26979
rect 9772 26936 9824 26945
rect 10324 26936 10376 26988
rect 12624 26936 12676 26988
rect 11428 26868 11480 26920
rect 4712 26775 4764 26784
rect 4712 26741 4721 26775
rect 4721 26741 4755 26775
rect 4755 26741 4764 26775
rect 4712 26732 4764 26741
rect 6828 26732 6880 26784
rect 9680 26732 9732 26784
rect 12440 26732 12492 26784
rect 14372 26868 14424 26920
rect 15016 26979 15068 26988
rect 15016 26945 15025 26979
rect 15025 26945 15059 26979
rect 15059 26945 15068 26979
rect 15016 26936 15068 26945
rect 15108 26979 15160 26988
rect 15108 26945 15117 26979
rect 15117 26945 15151 26979
rect 15151 26945 15160 26979
rect 15108 26936 15160 26945
rect 17132 26936 17184 26988
rect 17316 26936 17368 26988
rect 18972 27004 19024 27056
rect 20076 27004 20128 27056
rect 18236 26979 18288 26988
rect 18236 26945 18245 26979
rect 18245 26945 18279 26979
rect 18279 26945 18288 26979
rect 18420 26979 18472 26988
rect 18236 26936 18288 26945
rect 18420 26945 18429 26979
rect 18429 26945 18463 26979
rect 18463 26945 18472 26979
rect 18420 26936 18472 26945
rect 18604 26979 18656 26988
rect 18604 26945 18613 26979
rect 18613 26945 18647 26979
rect 18647 26945 18656 26979
rect 18604 26936 18656 26945
rect 18788 26936 18840 26988
rect 19340 26936 19392 26988
rect 22284 27004 22336 27056
rect 15660 26868 15712 26920
rect 19156 26868 19208 26920
rect 22100 26868 22152 26920
rect 14280 26800 14332 26852
rect 18052 26800 18104 26852
rect 18236 26800 18288 26852
rect 19064 26800 19116 26852
rect 17684 26732 17736 26784
rect 19432 26732 19484 26784
rect 21640 26732 21692 26784
rect 5915 26630 5967 26682
rect 5979 26630 6031 26682
rect 6043 26630 6095 26682
rect 6107 26630 6159 26682
rect 6171 26630 6223 26682
rect 15846 26630 15898 26682
rect 15910 26630 15962 26682
rect 15974 26630 16026 26682
rect 16038 26630 16090 26682
rect 16102 26630 16154 26682
rect 25776 26630 25828 26682
rect 25840 26630 25892 26682
rect 25904 26630 25956 26682
rect 25968 26630 26020 26682
rect 26032 26630 26084 26682
rect 4896 26571 4948 26580
rect 4896 26537 4905 26571
rect 4905 26537 4939 26571
rect 4939 26537 4948 26571
rect 4896 26528 4948 26537
rect 4620 26460 4672 26512
rect 6920 26528 6972 26580
rect 5448 26460 5500 26512
rect 6276 26460 6328 26512
rect 7564 26528 7616 26580
rect 7932 26528 7984 26580
rect 8392 26460 8444 26512
rect 9588 26460 9640 26512
rect 9772 26528 9824 26580
rect 10416 26571 10468 26580
rect 10416 26537 10425 26571
rect 10425 26537 10459 26571
rect 10459 26537 10468 26571
rect 10416 26528 10468 26537
rect 10048 26460 10100 26512
rect 2596 26324 2648 26376
rect 4252 26367 4304 26376
rect 4252 26333 4261 26367
rect 4261 26333 4295 26367
rect 4295 26333 4304 26367
rect 4252 26324 4304 26333
rect 4620 26367 4672 26376
rect 2964 26256 3016 26308
rect 4620 26333 4629 26367
rect 4629 26333 4663 26367
rect 4663 26333 4672 26367
rect 4620 26324 4672 26333
rect 4804 26324 4856 26376
rect 5264 26324 5316 26376
rect 5816 26256 5868 26308
rect 6828 26324 6880 26376
rect 7564 26435 7616 26444
rect 7564 26401 7573 26435
rect 7573 26401 7607 26435
rect 7607 26401 7616 26435
rect 7564 26392 7616 26401
rect 8668 26392 8720 26444
rect 9036 26392 9088 26444
rect 7840 26324 7892 26376
rect 7932 26324 7984 26376
rect 8944 26324 8996 26376
rect 9312 26367 9364 26376
rect 9312 26333 9322 26367
rect 9322 26333 9356 26367
rect 9356 26333 9364 26367
rect 10784 26392 10836 26444
rect 9312 26324 9364 26333
rect 10232 26324 10284 26376
rect 12900 26528 12952 26580
rect 14280 26571 14332 26580
rect 14280 26537 14289 26571
rect 14289 26537 14323 26571
rect 14323 26537 14332 26571
rect 14280 26528 14332 26537
rect 14648 26571 14700 26580
rect 14648 26537 14657 26571
rect 14657 26537 14691 26571
rect 14691 26537 14700 26571
rect 14648 26528 14700 26537
rect 15016 26528 15068 26580
rect 17500 26571 17552 26580
rect 11244 26460 11296 26512
rect 11336 26324 11388 26376
rect 12072 26460 12124 26512
rect 12164 26460 12216 26512
rect 12624 26503 12676 26512
rect 12624 26469 12633 26503
rect 12633 26469 12667 26503
rect 12667 26469 12676 26503
rect 12624 26460 12676 26469
rect 12716 26460 12768 26512
rect 12440 26367 12492 26376
rect 9588 26299 9640 26308
rect 1492 26231 1544 26240
rect 1492 26197 1501 26231
rect 1501 26197 1535 26231
rect 1535 26197 1544 26231
rect 1492 26188 1544 26197
rect 2780 26231 2832 26240
rect 2780 26197 2789 26231
rect 2789 26197 2823 26231
rect 2823 26197 2832 26231
rect 2780 26188 2832 26197
rect 4252 26188 4304 26240
rect 7288 26188 7340 26240
rect 7932 26188 7984 26240
rect 9588 26265 9597 26299
rect 9597 26265 9631 26299
rect 9631 26265 9640 26299
rect 9588 26256 9640 26265
rect 12440 26333 12449 26367
rect 12449 26333 12483 26367
rect 12483 26333 12492 26367
rect 12440 26324 12492 26333
rect 12808 26324 12860 26376
rect 14556 26392 14608 26444
rect 17500 26537 17509 26571
rect 17509 26537 17543 26571
rect 17543 26537 17552 26571
rect 17500 26528 17552 26537
rect 18144 26528 18196 26580
rect 20720 26528 20772 26580
rect 19340 26460 19392 26512
rect 15568 26392 15620 26444
rect 12532 26256 12584 26308
rect 12992 26256 13044 26308
rect 14372 26256 14424 26308
rect 17040 26256 17092 26308
rect 17316 26392 17368 26444
rect 18052 26392 18104 26444
rect 18788 26392 18840 26444
rect 17500 26324 17552 26376
rect 22100 26460 22152 26512
rect 21640 26435 21692 26444
rect 21640 26401 21649 26435
rect 21649 26401 21683 26435
rect 21683 26401 21692 26435
rect 21640 26392 21692 26401
rect 22376 26392 22428 26444
rect 17316 26299 17368 26308
rect 16948 26188 17000 26240
rect 17316 26265 17325 26299
rect 17325 26265 17359 26299
rect 17359 26265 17368 26299
rect 17316 26256 17368 26265
rect 18696 26256 18748 26308
rect 22100 26324 22152 26376
rect 23112 26367 23164 26376
rect 23112 26333 23121 26367
rect 23121 26333 23155 26367
rect 23155 26333 23164 26367
rect 23112 26324 23164 26333
rect 21272 26256 21324 26308
rect 22008 26256 22060 26308
rect 18236 26188 18288 26240
rect 10880 26086 10932 26138
rect 10944 26086 10996 26138
rect 11008 26086 11060 26138
rect 11072 26086 11124 26138
rect 11136 26086 11188 26138
rect 20811 26086 20863 26138
rect 20875 26086 20927 26138
rect 20939 26086 20991 26138
rect 21003 26086 21055 26138
rect 21067 26086 21119 26138
rect 2964 25984 3016 26036
rect 3608 25984 3660 26036
rect 2688 25891 2740 25900
rect 2688 25857 2697 25891
rect 2697 25857 2731 25891
rect 2731 25857 2740 25891
rect 2688 25848 2740 25857
rect 4436 25984 4488 26036
rect 4804 25984 4856 26036
rect 4712 25916 4764 25968
rect 2780 25780 2832 25832
rect 4068 25891 4120 25900
rect 4068 25857 4077 25891
rect 4077 25857 4111 25891
rect 4111 25857 4120 25891
rect 4068 25848 4120 25857
rect 4252 25891 4304 25900
rect 4252 25857 4297 25891
rect 4297 25857 4304 25891
rect 4252 25848 4304 25857
rect 4528 25848 4580 25900
rect 4896 25891 4948 25900
rect 4896 25857 4905 25891
rect 4905 25857 4939 25891
rect 4939 25857 4948 25891
rect 5816 25984 5868 26036
rect 7104 25984 7156 26036
rect 7472 25984 7524 26036
rect 8024 25984 8076 26036
rect 6552 25916 6604 25968
rect 9220 25984 9272 26036
rect 9588 25984 9640 26036
rect 11520 26027 11572 26036
rect 11520 25993 11529 26027
rect 11529 25993 11563 26027
rect 11563 25993 11572 26027
rect 11520 25984 11572 25993
rect 15108 25984 15160 26036
rect 4896 25848 4948 25857
rect 5080 25848 5132 25900
rect 7748 25848 7800 25900
rect 7012 25823 7064 25832
rect 7012 25789 7021 25823
rect 7021 25789 7055 25823
rect 7055 25789 7064 25823
rect 7012 25780 7064 25789
rect 7564 25780 7616 25832
rect 7840 25780 7892 25832
rect 6828 25712 6880 25764
rect 8024 25891 8076 25900
rect 8024 25857 8033 25891
rect 8033 25857 8067 25891
rect 8067 25857 8076 25891
rect 8024 25848 8076 25857
rect 8208 25780 8260 25832
rect 9404 25780 9456 25832
rect 9956 25848 10008 25900
rect 10784 25848 10836 25900
rect 12716 25916 12768 25968
rect 12164 25848 12216 25900
rect 12348 25848 12400 25900
rect 1492 25687 1544 25696
rect 1492 25653 1501 25687
rect 1501 25653 1535 25687
rect 1535 25653 1544 25687
rect 1492 25644 1544 25653
rect 5816 25644 5868 25696
rect 7932 25644 7984 25696
rect 12532 25780 12584 25832
rect 13820 25916 13872 25968
rect 15752 25959 15804 25968
rect 15752 25925 15761 25959
rect 15761 25925 15795 25959
rect 15795 25925 15804 25959
rect 15752 25916 15804 25925
rect 17040 25984 17092 26036
rect 18328 26027 18380 26036
rect 18328 25993 18337 26027
rect 18337 25993 18371 26027
rect 18371 25993 18380 26027
rect 18328 25984 18380 25993
rect 18788 25916 18840 25968
rect 13360 25848 13412 25900
rect 14372 25848 14424 25900
rect 15200 25780 15252 25832
rect 16488 25848 16540 25900
rect 19340 25984 19392 26036
rect 19524 25984 19576 26036
rect 19340 25848 19392 25900
rect 20628 25848 20680 25900
rect 22284 25984 22336 26036
rect 23204 25984 23256 26036
rect 20904 25916 20956 25968
rect 21180 25916 21232 25968
rect 21088 25891 21140 25900
rect 21088 25857 21097 25891
rect 21097 25857 21131 25891
rect 21131 25857 21140 25891
rect 21088 25848 21140 25857
rect 21456 25848 21508 25900
rect 18052 25780 18104 25832
rect 18696 25780 18748 25832
rect 18880 25823 18932 25832
rect 18880 25789 18889 25823
rect 18889 25789 18923 25823
rect 18923 25789 18932 25823
rect 19892 25823 19944 25832
rect 18880 25780 18932 25789
rect 19892 25789 19901 25823
rect 19901 25789 19935 25823
rect 19935 25789 19944 25823
rect 19892 25780 19944 25789
rect 20352 25780 20404 25832
rect 21180 25780 21232 25832
rect 21824 25823 21876 25832
rect 21824 25789 21833 25823
rect 21833 25789 21867 25823
rect 21867 25789 21876 25823
rect 21824 25780 21876 25789
rect 9956 25644 10008 25696
rect 12624 25644 12676 25696
rect 17500 25712 17552 25764
rect 15752 25644 15804 25696
rect 19432 25644 19484 25696
rect 20996 25644 21048 25696
rect 21272 25687 21324 25696
rect 21272 25653 21281 25687
rect 21281 25653 21315 25687
rect 21315 25653 21324 25687
rect 21272 25644 21324 25653
rect 22468 25644 22520 25696
rect 23112 25644 23164 25696
rect 5915 25542 5967 25594
rect 5979 25542 6031 25594
rect 6043 25542 6095 25594
rect 6107 25542 6159 25594
rect 6171 25542 6223 25594
rect 15846 25542 15898 25594
rect 15910 25542 15962 25594
rect 15974 25542 16026 25594
rect 16038 25542 16090 25594
rect 16102 25542 16154 25594
rect 25776 25542 25828 25594
rect 25840 25542 25892 25594
rect 25904 25542 25956 25594
rect 25968 25542 26020 25594
rect 26032 25542 26084 25594
rect 4068 25440 4120 25492
rect 6368 25440 6420 25492
rect 6920 25440 6972 25492
rect 7288 25440 7340 25492
rect 7840 25440 7892 25492
rect 9404 25440 9456 25492
rect 11796 25440 11848 25492
rect 12072 25440 12124 25492
rect 12348 25440 12400 25492
rect 13360 25440 13412 25492
rect 16396 25440 16448 25492
rect 16672 25440 16724 25492
rect 16764 25440 16816 25492
rect 17040 25440 17092 25492
rect 17316 25440 17368 25492
rect 19616 25483 19668 25492
rect 19616 25449 19625 25483
rect 19625 25449 19659 25483
rect 19659 25449 19668 25483
rect 19616 25440 19668 25449
rect 21456 25440 21508 25492
rect 23204 25483 23256 25492
rect 23204 25449 23213 25483
rect 23213 25449 23247 25483
rect 23247 25449 23256 25483
rect 23204 25440 23256 25449
rect 5724 25372 5776 25424
rect 7564 25415 7616 25424
rect 7564 25381 7573 25415
rect 7573 25381 7607 25415
rect 7607 25381 7616 25415
rect 7564 25372 7616 25381
rect 10324 25372 10376 25424
rect 10784 25415 10836 25424
rect 10784 25381 10793 25415
rect 10793 25381 10827 25415
rect 10827 25381 10836 25415
rect 10784 25372 10836 25381
rect 15200 25372 15252 25424
rect 15660 25372 15712 25424
rect 7932 25304 7984 25356
rect 10508 25304 10560 25356
rect 11888 25304 11940 25356
rect 12348 25347 12400 25356
rect 12348 25313 12357 25347
rect 12357 25313 12391 25347
rect 12391 25313 12400 25347
rect 12348 25304 12400 25313
rect 12532 25304 12584 25356
rect 13544 25304 13596 25356
rect 4344 25236 4396 25288
rect 5816 25236 5868 25288
rect 6920 25236 6972 25288
rect 9128 25279 9180 25288
rect 9128 25245 9137 25279
rect 9137 25245 9171 25279
rect 9171 25245 9180 25279
rect 9128 25236 9180 25245
rect 4804 25168 4856 25220
rect 6460 25211 6512 25220
rect 6460 25177 6494 25211
rect 6494 25177 6512 25211
rect 6460 25168 6512 25177
rect 6644 25168 6696 25220
rect 8024 25168 8076 25220
rect 9680 25236 9732 25288
rect 8208 25143 8260 25152
rect 8208 25109 8217 25143
rect 8217 25109 8251 25143
rect 8251 25109 8260 25143
rect 8208 25100 8260 25109
rect 8576 25100 8628 25152
rect 11612 25236 11664 25288
rect 12072 25279 12124 25288
rect 12072 25245 12081 25279
rect 12081 25245 12115 25279
rect 12115 25245 12124 25279
rect 12072 25236 12124 25245
rect 12624 25279 12676 25288
rect 11336 25168 11388 25220
rect 12624 25245 12633 25279
rect 12633 25245 12667 25279
rect 12667 25245 12676 25279
rect 12624 25236 12676 25245
rect 13268 25279 13320 25288
rect 13268 25245 13277 25279
rect 13277 25245 13311 25279
rect 13311 25245 13320 25279
rect 13268 25236 13320 25245
rect 13360 25279 13412 25288
rect 13360 25245 13369 25279
rect 13369 25245 13403 25279
rect 13403 25245 13412 25279
rect 13360 25236 13412 25245
rect 15292 25279 15344 25288
rect 15292 25245 15301 25279
rect 15301 25245 15335 25279
rect 15335 25245 15344 25279
rect 16672 25347 16724 25356
rect 16672 25313 16681 25347
rect 16681 25313 16715 25347
rect 16715 25313 16724 25347
rect 16672 25304 16724 25313
rect 18052 25304 18104 25356
rect 20076 25304 20128 25356
rect 20996 25347 21048 25356
rect 20996 25313 21005 25347
rect 21005 25313 21039 25347
rect 21039 25313 21048 25347
rect 20996 25304 21048 25313
rect 21824 25347 21876 25356
rect 21824 25313 21833 25347
rect 21833 25313 21867 25347
rect 21867 25313 21876 25347
rect 21824 25304 21876 25313
rect 19524 25279 19576 25288
rect 15292 25236 15344 25245
rect 12992 25168 13044 25220
rect 11520 25100 11572 25152
rect 15384 25143 15436 25152
rect 15384 25109 15393 25143
rect 15393 25109 15427 25143
rect 15427 25109 15436 25143
rect 15384 25100 15436 25109
rect 16488 25100 16540 25152
rect 18052 25168 18104 25220
rect 19524 25245 19533 25279
rect 19533 25245 19567 25279
rect 19567 25245 19576 25279
rect 19524 25236 19576 25245
rect 20536 25236 20588 25288
rect 20628 25279 20680 25288
rect 20628 25245 20637 25279
rect 20637 25245 20671 25279
rect 20671 25245 20680 25279
rect 20628 25236 20680 25245
rect 17040 25100 17092 25152
rect 17224 25100 17276 25152
rect 18144 25143 18196 25152
rect 18144 25109 18153 25143
rect 18153 25109 18187 25143
rect 18187 25109 18196 25143
rect 18144 25100 18196 25109
rect 20352 25100 20404 25152
rect 20904 25279 20956 25288
rect 20904 25245 20913 25279
rect 20913 25245 20947 25279
rect 20947 25245 20956 25279
rect 20904 25236 20956 25245
rect 21088 25236 21140 25288
rect 21272 25236 21324 25288
rect 29184 25236 29236 25288
rect 21548 25168 21600 25220
rect 22468 25100 22520 25152
rect 30012 25143 30064 25152
rect 30012 25109 30021 25143
rect 30021 25109 30055 25143
rect 30055 25109 30064 25143
rect 30012 25100 30064 25109
rect 10880 24998 10932 25050
rect 10944 24998 10996 25050
rect 11008 24998 11060 25050
rect 11072 24998 11124 25050
rect 11136 24998 11188 25050
rect 20811 24998 20863 25050
rect 20875 24998 20927 25050
rect 20939 24998 20991 25050
rect 21003 24998 21055 25050
rect 21067 24998 21119 25050
rect 4804 24939 4856 24948
rect 4804 24905 4813 24939
rect 4813 24905 4847 24939
rect 4847 24905 4856 24939
rect 4804 24896 4856 24905
rect 7656 24939 7708 24948
rect 7656 24905 7665 24939
rect 7665 24905 7699 24939
rect 7699 24905 7708 24939
rect 7656 24896 7708 24905
rect 9588 24896 9640 24948
rect 10692 24896 10744 24948
rect 11704 24896 11756 24948
rect 12164 24896 12216 24948
rect 2688 24803 2740 24812
rect 2688 24769 2697 24803
rect 2697 24769 2731 24803
rect 2731 24769 2740 24803
rect 2688 24760 2740 24769
rect 1492 24667 1544 24676
rect 1492 24633 1501 24667
rect 1501 24633 1535 24667
rect 1535 24633 1544 24667
rect 1492 24624 1544 24633
rect 4160 24760 4212 24812
rect 4528 24760 4580 24812
rect 4896 24760 4948 24812
rect 6736 24803 6788 24812
rect 6736 24769 6745 24803
rect 6745 24769 6779 24803
rect 6779 24769 6788 24803
rect 6736 24760 6788 24769
rect 7380 24760 7432 24812
rect 7656 24760 7708 24812
rect 8576 24803 8628 24812
rect 8576 24769 8585 24803
rect 8585 24769 8619 24803
rect 8619 24769 8628 24803
rect 8576 24760 8628 24769
rect 4344 24735 4396 24744
rect 4344 24701 4353 24735
rect 4353 24701 4387 24735
rect 4387 24701 4396 24735
rect 4344 24692 4396 24701
rect 4436 24735 4488 24744
rect 4436 24701 4445 24735
rect 4445 24701 4479 24735
rect 4479 24701 4488 24735
rect 4436 24692 4488 24701
rect 6828 24692 6880 24744
rect 7748 24735 7800 24744
rect 4068 24624 4120 24676
rect 7748 24701 7757 24735
rect 7757 24701 7791 24735
rect 7791 24701 7800 24735
rect 7748 24692 7800 24701
rect 7840 24735 7892 24744
rect 7840 24701 7849 24735
rect 7849 24701 7883 24735
rect 7883 24701 7892 24735
rect 7840 24692 7892 24701
rect 10232 24803 10284 24812
rect 10232 24769 10241 24803
rect 10241 24769 10275 24803
rect 10275 24769 10284 24803
rect 10232 24760 10284 24769
rect 7104 24556 7156 24608
rect 8116 24556 8168 24608
rect 10324 24692 10376 24744
rect 10692 24760 10744 24812
rect 10692 24624 10744 24676
rect 11244 24760 11296 24812
rect 11428 24760 11480 24812
rect 13268 24896 13320 24948
rect 13636 24896 13688 24948
rect 17132 24896 17184 24948
rect 17868 24939 17920 24948
rect 17868 24905 17877 24939
rect 17877 24905 17911 24939
rect 17911 24905 17920 24939
rect 17868 24896 17920 24905
rect 19892 24939 19944 24948
rect 19892 24905 19901 24939
rect 19901 24905 19935 24939
rect 19935 24905 19944 24939
rect 19892 24896 19944 24905
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 15568 24760 15620 24812
rect 17500 24828 17552 24880
rect 18880 24828 18932 24880
rect 21180 24896 21232 24948
rect 20536 24828 20588 24880
rect 15292 24692 15344 24744
rect 15016 24624 15068 24676
rect 15108 24556 15160 24608
rect 15476 24692 15528 24744
rect 18052 24760 18104 24812
rect 19340 24760 19392 24812
rect 16948 24692 17000 24744
rect 17868 24692 17920 24744
rect 19156 24692 19208 24744
rect 19984 24760 20036 24812
rect 20168 24760 20220 24812
rect 21732 24828 21784 24880
rect 19616 24624 19668 24676
rect 20536 24692 20588 24744
rect 15476 24556 15528 24608
rect 18880 24556 18932 24608
rect 18972 24599 19024 24608
rect 18972 24565 18981 24599
rect 18981 24565 19015 24599
rect 19015 24565 19024 24599
rect 20444 24599 20496 24608
rect 18972 24556 19024 24565
rect 20444 24565 20453 24599
rect 20453 24565 20487 24599
rect 20487 24565 20496 24599
rect 20444 24556 20496 24565
rect 5915 24454 5967 24506
rect 5979 24454 6031 24506
rect 6043 24454 6095 24506
rect 6107 24454 6159 24506
rect 6171 24454 6223 24506
rect 15846 24454 15898 24506
rect 15910 24454 15962 24506
rect 15974 24454 16026 24506
rect 16038 24454 16090 24506
rect 16102 24454 16154 24506
rect 25776 24454 25828 24506
rect 25840 24454 25892 24506
rect 25904 24454 25956 24506
rect 25968 24454 26020 24506
rect 26032 24454 26084 24506
rect 2688 24191 2740 24200
rect 2688 24157 2697 24191
rect 2697 24157 2731 24191
rect 2731 24157 2740 24191
rect 2688 24148 2740 24157
rect 5080 24352 5132 24404
rect 6460 24352 6512 24404
rect 6644 24352 6696 24404
rect 4344 24284 4396 24336
rect 4528 24284 4580 24336
rect 5908 24284 5960 24336
rect 5172 24216 5224 24268
rect 4344 24191 4396 24200
rect 3516 24080 3568 24132
rect 1492 24055 1544 24064
rect 1492 24021 1501 24055
rect 1501 24021 1535 24055
rect 1535 24021 1544 24055
rect 1492 24012 1544 24021
rect 3792 24055 3844 24064
rect 3792 24021 3801 24055
rect 3801 24021 3835 24055
rect 3835 24021 3844 24055
rect 3792 24012 3844 24021
rect 4344 24157 4353 24191
rect 4353 24157 4387 24191
rect 4387 24157 4396 24191
rect 4344 24148 4396 24157
rect 4528 24191 4580 24200
rect 4528 24157 4537 24191
rect 4537 24157 4571 24191
rect 4571 24157 4580 24191
rect 4528 24148 4580 24157
rect 5264 24148 5316 24200
rect 5540 24148 5592 24200
rect 6552 24216 6604 24268
rect 5908 24191 5960 24200
rect 5908 24157 5917 24191
rect 5917 24157 5951 24191
rect 5951 24157 5960 24191
rect 5908 24148 5960 24157
rect 7564 24284 7616 24336
rect 7748 24352 7800 24404
rect 10692 24352 10744 24404
rect 11980 24352 12032 24404
rect 14740 24352 14792 24404
rect 17868 24395 17920 24404
rect 8116 24216 8168 24268
rect 10784 24216 10836 24268
rect 12348 24259 12400 24268
rect 7380 24191 7432 24200
rect 7380 24157 7389 24191
rect 7389 24157 7423 24191
rect 7423 24157 7432 24191
rect 7380 24148 7432 24157
rect 4252 24080 4304 24132
rect 4436 24080 4488 24132
rect 7748 24191 7800 24200
rect 7748 24157 7757 24191
rect 7757 24157 7791 24191
rect 7791 24157 7800 24191
rect 7748 24148 7800 24157
rect 9128 24191 9180 24200
rect 9128 24157 9137 24191
rect 9137 24157 9171 24191
rect 9171 24157 9180 24191
rect 12072 24191 12124 24200
rect 9128 24148 9180 24157
rect 12072 24157 12081 24191
rect 12081 24157 12115 24191
rect 12115 24157 12124 24191
rect 12072 24148 12124 24157
rect 12348 24225 12357 24259
rect 12357 24225 12391 24259
rect 12391 24225 12400 24259
rect 12348 24216 12400 24225
rect 12532 24216 12584 24268
rect 17868 24361 17877 24395
rect 17877 24361 17911 24395
rect 17911 24361 17920 24395
rect 17868 24352 17920 24361
rect 9864 24080 9916 24132
rect 12164 24080 12216 24132
rect 14280 24148 14332 24200
rect 14648 24148 14700 24200
rect 15384 24284 15436 24336
rect 15568 24284 15620 24336
rect 18972 24352 19024 24404
rect 19616 24352 19668 24404
rect 15476 24216 15528 24268
rect 15108 24123 15160 24132
rect 15108 24089 15117 24123
rect 15117 24089 15151 24123
rect 15151 24089 15160 24123
rect 15108 24080 15160 24089
rect 4160 24012 4212 24064
rect 5264 24012 5316 24064
rect 6000 24012 6052 24064
rect 8576 24012 8628 24064
rect 11336 24012 11388 24064
rect 11612 24012 11664 24064
rect 13176 24012 13228 24064
rect 15016 24012 15068 24064
rect 15568 24148 15620 24200
rect 16396 24216 16448 24268
rect 18328 24216 18380 24268
rect 17408 24148 17460 24200
rect 18604 24284 18656 24336
rect 21916 24216 21968 24268
rect 22468 24259 22520 24268
rect 22468 24225 22477 24259
rect 22477 24225 22511 24259
rect 22511 24225 22520 24259
rect 22468 24216 22520 24225
rect 20352 24191 20404 24200
rect 16396 24080 16448 24132
rect 16948 24080 17000 24132
rect 20352 24157 20361 24191
rect 20361 24157 20395 24191
rect 20395 24157 20404 24191
rect 20352 24148 20404 24157
rect 16120 24012 16172 24064
rect 16488 24012 16540 24064
rect 16580 24012 16632 24064
rect 17132 24012 17184 24064
rect 18328 24012 18380 24064
rect 21640 24080 21692 24132
rect 22284 24080 22336 24132
rect 21456 24012 21508 24064
rect 10880 23910 10932 23962
rect 10944 23910 10996 23962
rect 11008 23910 11060 23962
rect 11072 23910 11124 23962
rect 11136 23910 11188 23962
rect 20811 23910 20863 23962
rect 20875 23910 20927 23962
rect 20939 23910 20991 23962
rect 21003 23910 21055 23962
rect 21067 23910 21119 23962
rect 4160 23851 4212 23860
rect 4160 23817 4169 23851
rect 4169 23817 4203 23851
rect 4203 23817 4212 23851
rect 4160 23808 4212 23817
rect 7288 23808 7340 23860
rect 7380 23808 7432 23860
rect 2872 23740 2924 23792
rect 4068 23740 4120 23792
rect 3792 23672 3844 23724
rect 4988 23740 5040 23792
rect 5908 23740 5960 23792
rect 7564 23740 7616 23792
rect 1400 23647 1452 23656
rect 1400 23613 1409 23647
rect 1409 23613 1443 23647
rect 1443 23613 1452 23647
rect 1400 23604 1452 23613
rect 2320 23604 2372 23656
rect 4252 23604 4304 23656
rect 4896 23604 4948 23656
rect 5080 23647 5132 23656
rect 5080 23613 5089 23647
rect 5089 23613 5123 23647
rect 5123 23613 5132 23647
rect 5540 23672 5592 23724
rect 6460 23672 6512 23724
rect 5080 23604 5132 23613
rect 5724 23604 5776 23656
rect 4344 23536 4396 23588
rect 6644 23715 6696 23724
rect 6644 23681 6653 23715
rect 6653 23681 6687 23715
rect 6687 23681 6696 23715
rect 6644 23672 6696 23681
rect 6920 23715 6972 23724
rect 6920 23681 6929 23715
rect 6929 23681 6963 23715
rect 6963 23681 6972 23715
rect 6920 23672 6972 23681
rect 7288 23672 7340 23724
rect 9680 23808 9732 23860
rect 9864 23851 9916 23860
rect 9864 23817 9873 23851
rect 9873 23817 9907 23851
rect 9907 23817 9916 23851
rect 9864 23808 9916 23817
rect 10232 23808 10284 23860
rect 11612 23808 11664 23860
rect 12256 23808 12308 23860
rect 14280 23851 14332 23860
rect 14280 23817 14289 23851
rect 14289 23817 14323 23851
rect 14323 23817 14332 23851
rect 14280 23808 14332 23817
rect 14740 23808 14792 23860
rect 18328 23808 18380 23860
rect 20076 23851 20128 23860
rect 20076 23817 20085 23851
rect 20085 23817 20119 23851
rect 20119 23817 20128 23851
rect 20076 23808 20128 23817
rect 8576 23740 8628 23792
rect 8024 23672 8076 23724
rect 8208 23715 8260 23724
rect 8208 23681 8217 23715
rect 8217 23681 8251 23715
rect 8251 23681 8260 23715
rect 8208 23672 8260 23681
rect 9220 23672 9272 23724
rect 9496 23715 9548 23724
rect 9496 23681 9505 23715
rect 9505 23681 9539 23715
rect 9539 23681 9548 23715
rect 9496 23672 9548 23681
rect 11336 23740 11388 23792
rect 11428 23740 11480 23792
rect 10508 23715 10560 23724
rect 10508 23681 10517 23715
rect 10517 23681 10551 23715
rect 10551 23681 10560 23715
rect 10508 23672 10560 23681
rect 12992 23740 13044 23792
rect 13176 23783 13228 23792
rect 13176 23749 13210 23783
rect 13210 23749 13228 23783
rect 13176 23740 13228 23749
rect 15108 23740 15160 23792
rect 16304 23740 16356 23792
rect 19340 23740 19392 23792
rect 20352 23740 20404 23792
rect 12348 23672 12400 23724
rect 14280 23672 14332 23724
rect 16488 23672 16540 23724
rect 16672 23715 16724 23724
rect 16672 23681 16681 23715
rect 16681 23681 16715 23715
rect 16715 23681 16724 23715
rect 16672 23672 16724 23681
rect 17132 23715 17184 23724
rect 17132 23681 17141 23715
rect 17141 23681 17175 23715
rect 17175 23681 17184 23715
rect 17132 23672 17184 23681
rect 17776 23672 17828 23724
rect 17868 23672 17920 23724
rect 20444 23715 20496 23724
rect 9404 23647 9456 23656
rect 4620 23511 4672 23520
rect 4620 23477 4629 23511
rect 4629 23477 4663 23511
rect 4663 23477 4672 23511
rect 4620 23468 4672 23477
rect 6644 23536 6696 23588
rect 9404 23613 9413 23647
rect 9413 23613 9447 23647
rect 9447 23613 9456 23647
rect 9404 23604 9456 23613
rect 9588 23604 9640 23656
rect 9772 23604 9824 23656
rect 10048 23604 10100 23656
rect 15476 23647 15528 23656
rect 15476 23613 15485 23647
rect 15485 23613 15519 23647
rect 15519 23613 15528 23647
rect 15476 23604 15528 23613
rect 15568 23604 15620 23656
rect 16120 23604 16172 23656
rect 17224 23647 17276 23656
rect 8668 23536 8720 23588
rect 16396 23536 16448 23588
rect 17224 23613 17233 23647
rect 17233 23613 17267 23647
rect 17267 23613 17276 23647
rect 17224 23604 17276 23613
rect 17408 23647 17460 23656
rect 17408 23613 17417 23647
rect 17417 23613 17451 23647
rect 17451 23613 17460 23647
rect 17408 23604 17460 23613
rect 18604 23647 18656 23656
rect 18604 23613 18613 23647
rect 18613 23613 18647 23647
rect 18647 23613 18656 23647
rect 18604 23604 18656 23613
rect 19156 23604 19208 23656
rect 20444 23681 20453 23715
rect 20453 23681 20487 23715
rect 20487 23681 20496 23715
rect 20444 23672 20496 23681
rect 22284 23808 22336 23860
rect 21916 23783 21968 23792
rect 21916 23749 21925 23783
rect 21925 23749 21959 23783
rect 21959 23749 21968 23783
rect 21916 23740 21968 23749
rect 22836 23672 22888 23724
rect 20536 23604 20588 23656
rect 20720 23604 20772 23656
rect 22652 23647 22704 23656
rect 22652 23613 22661 23647
rect 22661 23613 22695 23647
rect 22695 23613 22704 23647
rect 22652 23604 22704 23613
rect 22928 23647 22980 23656
rect 22928 23613 22937 23647
rect 22937 23613 22971 23647
rect 22971 23613 22980 23647
rect 22928 23604 22980 23613
rect 20628 23536 20680 23588
rect 6920 23468 6972 23520
rect 7932 23468 7984 23520
rect 8944 23468 8996 23520
rect 9772 23468 9824 23520
rect 16212 23468 16264 23520
rect 16304 23468 16356 23520
rect 18144 23511 18196 23520
rect 18144 23477 18153 23511
rect 18153 23477 18187 23511
rect 18187 23477 18196 23511
rect 18144 23468 18196 23477
rect 19524 23468 19576 23520
rect 5915 23366 5967 23418
rect 5979 23366 6031 23418
rect 6043 23366 6095 23418
rect 6107 23366 6159 23418
rect 6171 23366 6223 23418
rect 15846 23366 15898 23418
rect 15910 23366 15962 23418
rect 15974 23366 16026 23418
rect 16038 23366 16090 23418
rect 16102 23366 16154 23418
rect 25776 23366 25828 23418
rect 25840 23366 25892 23418
rect 25904 23366 25956 23418
rect 25968 23366 26020 23418
rect 26032 23366 26084 23418
rect 4988 23264 5040 23316
rect 5448 23307 5500 23316
rect 5448 23273 5457 23307
rect 5457 23273 5491 23307
rect 5491 23273 5500 23307
rect 5448 23264 5500 23273
rect 5724 23264 5776 23316
rect 7288 23307 7340 23316
rect 7288 23273 7297 23307
rect 7297 23273 7331 23307
rect 7331 23273 7340 23307
rect 7288 23264 7340 23273
rect 7656 23264 7708 23316
rect 4068 23171 4120 23180
rect 4068 23137 4077 23171
rect 4077 23137 4111 23171
rect 4111 23137 4120 23171
rect 4068 23128 4120 23137
rect 5816 23128 5868 23180
rect 7288 23128 7340 23180
rect 7840 23128 7892 23180
rect 2044 23103 2096 23112
rect 2044 23069 2053 23103
rect 2053 23069 2087 23103
rect 2087 23069 2096 23103
rect 2044 23060 2096 23069
rect 4620 23060 4672 23112
rect 6920 23060 6972 23112
rect 9220 23103 9272 23112
rect 2780 22992 2832 23044
rect 1676 22924 1728 22976
rect 4252 22924 4304 22976
rect 7840 22967 7892 22976
rect 7840 22933 7849 22967
rect 7849 22933 7883 22967
rect 7883 22933 7892 22967
rect 7840 22924 7892 22933
rect 9220 23069 9229 23103
rect 9229 23069 9263 23103
rect 9263 23069 9272 23103
rect 9220 23060 9272 23069
rect 9496 23196 9548 23248
rect 11520 23264 11572 23316
rect 13084 23264 13136 23316
rect 15016 23264 15068 23316
rect 15568 23264 15620 23316
rect 16672 23264 16724 23316
rect 19524 23307 19576 23316
rect 19524 23273 19533 23307
rect 19533 23273 19567 23307
rect 19567 23273 19576 23307
rect 19524 23264 19576 23273
rect 22652 23264 22704 23316
rect 10416 23060 10468 23112
rect 11704 23128 11756 23180
rect 12164 23128 12216 23180
rect 12532 23128 12584 23180
rect 12072 23103 12124 23112
rect 9588 22992 9640 23044
rect 12072 23069 12081 23103
rect 12081 23069 12115 23103
rect 12115 23069 12124 23103
rect 12072 23060 12124 23069
rect 12256 23103 12308 23112
rect 12256 23069 12265 23103
rect 12265 23069 12299 23103
rect 12299 23069 12308 23103
rect 12256 23060 12308 23069
rect 14280 23128 14332 23180
rect 16672 23128 16724 23180
rect 17040 23128 17092 23180
rect 13728 23060 13780 23112
rect 15752 23060 15804 23112
rect 16212 23103 16264 23112
rect 16212 23069 16221 23103
rect 16221 23069 16255 23103
rect 16255 23069 16264 23103
rect 16212 23060 16264 23069
rect 16580 23103 16632 23112
rect 8024 22924 8076 22976
rect 12992 22992 13044 23044
rect 14556 23035 14608 23044
rect 14556 23001 14565 23035
rect 14565 23001 14599 23035
rect 14599 23001 14608 23035
rect 14556 22992 14608 23001
rect 14740 23035 14792 23044
rect 14740 23001 14749 23035
rect 14749 23001 14783 23035
rect 14783 23001 14792 23035
rect 14740 22992 14792 23001
rect 16580 23069 16589 23103
rect 16589 23069 16623 23103
rect 16623 23069 16632 23103
rect 16580 23060 16632 23069
rect 18972 23060 19024 23112
rect 19156 23060 19208 23112
rect 19708 23060 19760 23112
rect 20076 23103 20128 23112
rect 20076 23069 20085 23103
rect 20085 23069 20119 23103
rect 20119 23069 20128 23103
rect 20076 23060 20128 23069
rect 20260 23103 20312 23112
rect 20260 23069 20269 23103
rect 20269 23069 20303 23103
rect 20303 23069 20312 23103
rect 20260 23060 20312 23069
rect 20720 23128 20772 23180
rect 21272 23128 21324 23180
rect 21456 23171 21508 23180
rect 21456 23137 21465 23171
rect 21465 23137 21499 23171
rect 21499 23137 21508 23171
rect 21456 23128 21508 23137
rect 21180 23060 21232 23112
rect 22192 23196 22244 23248
rect 22376 23128 22428 23180
rect 22928 23128 22980 23180
rect 22192 23060 22244 23112
rect 29460 23060 29512 23112
rect 20536 22992 20588 23044
rect 10048 22924 10100 22976
rect 11796 22924 11848 22976
rect 12808 22967 12860 22976
rect 12808 22933 12817 22967
rect 12817 22933 12851 22967
rect 12851 22933 12860 22967
rect 12808 22924 12860 22933
rect 19156 22924 19208 22976
rect 20720 22967 20772 22976
rect 20720 22933 20729 22967
rect 20729 22933 20763 22967
rect 20763 22933 20772 22967
rect 20720 22924 20772 22933
rect 22284 22992 22336 23044
rect 22928 23035 22980 23044
rect 22928 23001 22937 23035
rect 22937 23001 22971 23035
rect 22971 23001 22980 23035
rect 22928 22992 22980 23001
rect 23388 22967 23440 22976
rect 23388 22933 23397 22967
rect 23397 22933 23431 22967
rect 23431 22933 23440 22967
rect 23388 22924 23440 22933
rect 30012 22967 30064 22976
rect 30012 22933 30021 22967
rect 30021 22933 30055 22967
rect 30055 22933 30064 22967
rect 30012 22924 30064 22933
rect 10880 22822 10932 22874
rect 10944 22822 10996 22874
rect 11008 22822 11060 22874
rect 11072 22822 11124 22874
rect 11136 22822 11188 22874
rect 20811 22822 20863 22874
rect 20875 22822 20927 22874
rect 20939 22822 20991 22874
rect 21003 22822 21055 22874
rect 21067 22822 21119 22874
rect 7012 22720 7064 22772
rect 9128 22720 9180 22772
rect 9404 22720 9456 22772
rect 12256 22720 12308 22772
rect 13728 22720 13780 22772
rect 14280 22763 14332 22772
rect 14280 22729 14289 22763
rect 14289 22729 14323 22763
rect 14323 22729 14332 22763
rect 14280 22720 14332 22729
rect 15752 22720 15804 22772
rect 16304 22720 16356 22772
rect 16396 22720 16448 22772
rect 17408 22763 17460 22772
rect 17408 22729 17417 22763
rect 17417 22729 17451 22763
rect 17451 22729 17460 22763
rect 17408 22720 17460 22729
rect 18604 22720 18656 22772
rect 19800 22763 19852 22772
rect 19800 22729 19809 22763
rect 19809 22729 19843 22763
rect 19843 22729 19852 22763
rect 19800 22720 19852 22729
rect 20076 22720 20128 22772
rect 21180 22720 21232 22772
rect 22008 22720 22060 22772
rect 22192 22763 22244 22772
rect 22192 22729 22201 22763
rect 22201 22729 22235 22763
rect 22235 22729 22244 22763
rect 22192 22720 22244 22729
rect 1860 22584 1912 22636
rect 2964 22584 3016 22636
rect 5080 22584 5132 22636
rect 3148 22516 3200 22568
rect 5264 22559 5316 22568
rect 5264 22525 5273 22559
rect 5273 22525 5307 22559
rect 5307 22525 5316 22559
rect 5264 22516 5316 22525
rect 5724 22516 5776 22568
rect 9220 22652 9272 22704
rect 12808 22652 12860 22704
rect 19340 22652 19392 22704
rect 19616 22652 19668 22704
rect 20536 22652 20588 22704
rect 22468 22652 22520 22704
rect 22928 22720 22980 22772
rect 22836 22695 22888 22704
rect 22836 22661 22845 22695
rect 22845 22661 22879 22695
rect 22879 22661 22888 22695
rect 22836 22652 22888 22661
rect 23020 22695 23072 22704
rect 23020 22661 23029 22695
rect 23029 22661 23063 22695
rect 23063 22661 23072 22695
rect 23020 22652 23072 22661
rect 23388 22652 23440 22704
rect 6460 22584 6512 22636
rect 7840 22627 7892 22636
rect 7840 22593 7849 22627
rect 7849 22593 7883 22627
rect 7883 22593 7892 22627
rect 7840 22584 7892 22593
rect 8208 22627 8260 22636
rect 8208 22593 8217 22627
rect 8217 22593 8251 22627
rect 8251 22593 8260 22627
rect 8208 22584 8260 22593
rect 9128 22584 9180 22636
rect 9496 22584 9548 22636
rect 12348 22584 12400 22636
rect 12532 22584 12584 22636
rect 15660 22627 15712 22636
rect 15660 22593 15669 22627
rect 15669 22593 15703 22627
rect 15703 22593 15712 22627
rect 15660 22584 15712 22593
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 17040 22584 17092 22593
rect 18328 22627 18380 22636
rect 18328 22593 18337 22627
rect 18337 22593 18371 22627
rect 18371 22593 18380 22627
rect 18328 22584 18380 22593
rect 19156 22627 19208 22636
rect 19156 22593 19165 22627
rect 19165 22593 19199 22627
rect 19199 22593 19208 22627
rect 19156 22584 19208 22593
rect 19984 22584 20036 22636
rect 20720 22627 20772 22636
rect 20720 22593 20729 22627
rect 20729 22593 20763 22627
rect 20763 22593 20772 22627
rect 20720 22584 20772 22593
rect 21272 22584 21324 22636
rect 7932 22516 7984 22568
rect 8300 22516 8352 22568
rect 10324 22516 10376 22568
rect 17408 22516 17460 22568
rect 18420 22516 18472 22568
rect 8944 22448 8996 22500
rect 19708 22448 19760 22500
rect 21548 22448 21600 22500
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 1768 22380 1820 22432
rect 3976 22380 4028 22432
rect 19064 22380 19116 22432
rect 5915 22278 5967 22330
rect 5979 22278 6031 22330
rect 6043 22278 6095 22330
rect 6107 22278 6159 22330
rect 6171 22278 6223 22330
rect 15846 22278 15898 22330
rect 15910 22278 15962 22330
rect 15974 22278 16026 22330
rect 16038 22278 16090 22330
rect 16102 22278 16154 22330
rect 25776 22278 25828 22330
rect 25840 22278 25892 22330
rect 25904 22278 25956 22330
rect 25968 22278 26020 22330
rect 26032 22278 26084 22330
rect 7380 22176 7432 22228
rect 8392 22176 8444 22228
rect 11520 22176 11572 22228
rect 12992 22219 13044 22228
rect 12992 22185 13001 22219
rect 13001 22185 13035 22219
rect 13035 22185 13044 22219
rect 12992 22176 13044 22185
rect 18328 22176 18380 22228
rect 20720 22176 20772 22228
rect 22100 22176 22152 22228
rect 22836 22176 22888 22228
rect 7564 22108 7616 22160
rect 8116 22108 8168 22160
rect 8668 22108 8720 22160
rect 15476 22108 15528 22160
rect 15844 22108 15896 22160
rect 4988 22040 5040 22092
rect 8208 22040 8260 22092
rect 8300 22040 8352 22092
rect 9680 22040 9732 22092
rect 15568 22040 15620 22092
rect 2872 21972 2924 22024
rect 2136 21947 2188 21956
rect 2136 21913 2170 21947
rect 2170 21913 2188 21947
rect 5448 21972 5500 22024
rect 7104 21972 7156 22024
rect 7564 21972 7616 22024
rect 2136 21904 2188 21913
rect 5264 21904 5316 21956
rect 3056 21836 3108 21888
rect 6736 21836 6788 21888
rect 7840 21836 7892 21888
rect 8300 21904 8352 21956
rect 9404 21972 9456 22024
rect 10048 22015 10100 22024
rect 10048 21981 10082 22015
rect 10082 21981 10100 22015
rect 10048 21972 10100 21981
rect 11520 21972 11572 22024
rect 12348 21972 12400 22024
rect 15476 22015 15528 22024
rect 15476 21981 15490 22015
rect 15490 21981 15524 22015
rect 15524 21981 15528 22015
rect 17868 22108 17920 22160
rect 16580 22083 16632 22092
rect 16580 22049 16589 22083
rect 16589 22049 16623 22083
rect 16623 22049 16632 22083
rect 16580 22040 16632 22049
rect 17224 22040 17276 22092
rect 19156 22108 19208 22160
rect 18052 22040 18104 22092
rect 18604 22083 18656 22092
rect 18604 22049 18613 22083
rect 18613 22049 18647 22083
rect 18647 22049 18656 22083
rect 18604 22040 18656 22049
rect 19248 22040 19300 22092
rect 19892 22083 19944 22092
rect 19892 22049 19901 22083
rect 19901 22049 19935 22083
rect 19935 22049 19944 22083
rect 19892 22040 19944 22049
rect 20812 22040 20864 22092
rect 22008 22040 22060 22092
rect 16488 22015 16540 22024
rect 15476 21972 15528 21981
rect 16488 21981 16497 22015
rect 16497 21981 16531 22015
rect 16531 21981 16540 22015
rect 16488 21972 16540 21981
rect 8576 21836 8628 21888
rect 9956 21904 10008 21956
rect 11888 21947 11940 21956
rect 11888 21913 11922 21947
rect 11922 21913 11940 21947
rect 11888 21904 11940 21913
rect 15292 21947 15344 21956
rect 14372 21836 14424 21888
rect 15292 21913 15301 21947
rect 15301 21913 15335 21947
rect 15335 21913 15344 21947
rect 15292 21904 15344 21913
rect 15384 21947 15436 21956
rect 15384 21913 15393 21947
rect 15393 21913 15427 21947
rect 15427 21913 15436 21947
rect 16856 21972 16908 22024
rect 17868 21972 17920 22024
rect 15384 21904 15436 21913
rect 17132 21904 17184 21956
rect 19432 21972 19484 22024
rect 19984 21972 20036 22024
rect 20720 22015 20772 22024
rect 20720 21981 20729 22015
rect 20729 21981 20763 22015
rect 20763 21981 20772 22015
rect 20720 21972 20772 21981
rect 22100 21972 22152 22024
rect 19708 21904 19760 21956
rect 21456 21904 21508 21956
rect 22376 21904 22428 21956
rect 19524 21836 19576 21888
rect 10880 21734 10932 21786
rect 10944 21734 10996 21786
rect 11008 21734 11060 21786
rect 11072 21734 11124 21786
rect 11136 21734 11188 21786
rect 20811 21734 20863 21786
rect 20875 21734 20927 21786
rect 20939 21734 20991 21786
rect 21003 21734 21055 21786
rect 21067 21734 21119 21786
rect 7748 21632 7800 21684
rect 8208 21632 8260 21684
rect 2872 21564 2924 21616
rect 5448 21564 5500 21616
rect 7564 21564 7616 21616
rect 2228 21539 2280 21548
rect 2228 21505 2262 21539
rect 2262 21505 2280 21539
rect 2228 21496 2280 21505
rect 2964 21292 3016 21344
rect 6552 21539 6604 21548
rect 6552 21505 6556 21539
rect 6556 21505 6590 21539
rect 6590 21505 6604 21539
rect 6552 21496 6604 21505
rect 6460 21428 6512 21480
rect 6828 21539 6880 21548
rect 6828 21505 6873 21539
rect 6873 21505 6880 21539
rect 6828 21496 6880 21505
rect 8208 21496 8260 21548
rect 6276 21292 6328 21344
rect 6552 21292 6604 21344
rect 7840 21428 7892 21480
rect 8392 21360 8444 21412
rect 9220 21496 9272 21548
rect 9496 21496 9548 21548
rect 10508 21496 10560 21548
rect 12532 21632 12584 21684
rect 15292 21632 15344 21684
rect 16488 21632 16540 21684
rect 17868 21675 17920 21684
rect 17868 21641 17877 21675
rect 17877 21641 17911 21675
rect 17911 21641 17920 21675
rect 17868 21632 17920 21641
rect 18144 21632 18196 21684
rect 19340 21632 19392 21684
rect 20444 21632 20496 21684
rect 9404 21471 9456 21480
rect 9404 21437 9413 21471
rect 9413 21437 9447 21471
rect 9447 21437 9456 21471
rect 9404 21428 9456 21437
rect 8668 21360 8720 21412
rect 7380 21292 7432 21344
rect 7656 21292 7708 21344
rect 11612 21496 11664 21548
rect 12992 21564 13044 21616
rect 11796 21539 11848 21548
rect 11796 21505 11805 21539
rect 11805 21505 11839 21539
rect 11839 21505 11848 21539
rect 11796 21496 11848 21505
rect 13728 21496 13780 21548
rect 15292 21539 15344 21548
rect 15292 21505 15301 21539
rect 15301 21505 15335 21539
rect 15335 21505 15344 21539
rect 15292 21496 15344 21505
rect 15568 21496 15620 21548
rect 16764 21496 16816 21548
rect 17776 21564 17828 21616
rect 17224 21539 17276 21548
rect 17224 21505 17233 21539
rect 17233 21505 17267 21539
rect 17267 21505 17276 21539
rect 17224 21496 17276 21505
rect 17868 21496 17920 21548
rect 11888 21471 11940 21480
rect 11888 21437 11897 21471
rect 11897 21437 11931 21471
rect 11931 21437 11940 21471
rect 11888 21428 11940 21437
rect 15844 21428 15896 21480
rect 16488 21428 16540 21480
rect 19064 21539 19116 21548
rect 19064 21505 19073 21539
rect 19073 21505 19107 21539
rect 19107 21505 19116 21539
rect 19064 21496 19116 21505
rect 18420 21471 18472 21480
rect 18420 21437 18429 21471
rect 18429 21437 18463 21471
rect 18463 21437 18472 21471
rect 18420 21428 18472 21437
rect 18604 21428 18656 21480
rect 19340 21539 19392 21548
rect 19340 21505 19349 21539
rect 19349 21505 19383 21539
rect 19383 21505 19392 21539
rect 19340 21496 19392 21505
rect 19524 21496 19576 21548
rect 20260 21539 20312 21548
rect 20260 21505 20269 21539
rect 20269 21505 20303 21539
rect 20303 21505 20312 21539
rect 20260 21496 20312 21505
rect 21456 21496 21508 21548
rect 29920 21496 29972 21548
rect 19892 21428 19944 21480
rect 15108 21360 15160 21412
rect 15568 21360 15620 21412
rect 19156 21360 19208 21412
rect 16948 21292 17000 21344
rect 17868 21292 17920 21344
rect 19248 21292 19300 21344
rect 19524 21335 19576 21344
rect 19524 21301 19533 21335
rect 19533 21301 19567 21335
rect 19567 21301 19576 21335
rect 19524 21292 19576 21301
rect 20536 21292 20588 21344
rect 30012 21335 30064 21344
rect 30012 21301 30021 21335
rect 30021 21301 30055 21335
rect 30055 21301 30064 21335
rect 30012 21292 30064 21301
rect 5915 21190 5967 21242
rect 5979 21190 6031 21242
rect 6043 21190 6095 21242
rect 6107 21190 6159 21242
rect 6171 21190 6223 21242
rect 15846 21190 15898 21242
rect 15910 21190 15962 21242
rect 15974 21190 16026 21242
rect 16038 21190 16090 21242
rect 16102 21190 16154 21242
rect 25776 21190 25828 21242
rect 25840 21190 25892 21242
rect 25904 21190 25956 21242
rect 25968 21190 26020 21242
rect 26032 21190 26084 21242
rect 2228 21088 2280 21140
rect 5448 21131 5500 21140
rect 5448 21097 5457 21131
rect 5457 21097 5491 21131
rect 5491 21097 5500 21131
rect 5448 21088 5500 21097
rect 6644 21088 6696 21140
rect 6828 21088 6880 21140
rect 8208 21131 8260 21140
rect 8208 21097 8217 21131
rect 8217 21097 8251 21131
rect 8251 21097 8260 21131
rect 8208 21088 8260 21097
rect 8484 21088 8536 21140
rect 9220 21088 9272 21140
rect 10324 21088 10376 21140
rect 16764 21131 16816 21140
rect 16764 21097 16773 21131
rect 16773 21097 16807 21131
rect 16807 21097 16816 21131
rect 16764 21088 16816 21097
rect 17132 21088 17184 21140
rect 17868 21088 17920 21140
rect 7932 21020 7984 21072
rect 1952 20995 2004 21004
rect 1952 20961 1961 20995
rect 1961 20961 1995 20995
rect 1995 20961 2004 20995
rect 1952 20952 2004 20961
rect 4436 20952 4488 21004
rect 7380 20952 7432 21004
rect 8484 20952 8536 21004
rect 9588 20952 9640 21004
rect 17592 21020 17644 21072
rect 17408 20952 17460 21004
rect 18420 21020 18472 21072
rect 19340 21088 19392 21140
rect 19708 21131 19760 21140
rect 19708 21097 19717 21131
rect 19717 21097 19751 21131
rect 19751 21097 19760 21131
rect 19708 21088 19760 21097
rect 20720 21020 20772 21072
rect 1768 20927 1820 20936
rect 1400 20748 1452 20800
rect 1768 20893 1777 20927
rect 1777 20893 1811 20927
rect 1811 20893 1820 20927
rect 1768 20884 1820 20893
rect 1860 20927 1912 20936
rect 1860 20893 1869 20927
rect 1869 20893 1903 20927
rect 1903 20893 1912 20927
rect 1860 20884 1912 20893
rect 2964 20884 3016 20936
rect 3056 20927 3108 20936
rect 3056 20893 3065 20927
rect 3065 20893 3099 20927
rect 3099 20893 3108 20927
rect 3056 20884 3108 20893
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 5172 20884 5224 20936
rect 6552 20927 6604 20936
rect 6552 20893 6570 20927
rect 6570 20893 6604 20927
rect 6552 20884 6604 20893
rect 6736 20884 6788 20936
rect 6920 20884 6972 20936
rect 7932 20927 7984 20936
rect 7932 20893 7941 20927
rect 7941 20893 7975 20927
rect 7975 20893 7984 20927
rect 7932 20884 7984 20893
rect 9312 20884 9364 20936
rect 13360 20927 13412 20936
rect 13360 20893 13369 20927
rect 13369 20893 13403 20927
rect 13403 20893 13412 20927
rect 13360 20884 13412 20893
rect 3332 20816 3384 20868
rect 4160 20816 4212 20868
rect 7104 20816 7156 20868
rect 9680 20816 9732 20868
rect 10416 20816 10468 20868
rect 10600 20859 10652 20868
rect 10600 20825 10609 20859
rect 10609 20825 10643 20859
rect 10643 20825 10652 20859
rect 10600 20816 10652 20825
rect 4528 20791 4580 20800
rect 4528 20757 4537 20791
rect 4537 20757 4571 20791
rect 4571 20757 4580 20791
rect 4528 20748 4580 20757
rect 6276 20748 6328 20800
rect 6736 20748 6788 20800
rect 8668 20748 8720 20800
rect 14832 20791 14884 20800
rect 14832 20757 14841 20791
rect 14841 20757 14875 20791
rect 14875 20757 14884 20791
rect 14832 20748 14884 20757
rect 15292 20791 15344 20800
rect 15292 20757 15301 20791
rect 15301 20757 15335 20791
rect 15335 20757 15344 20791
rect 16212 20816 16264 20868
rect 16488 20816 16540 20868
rect 17408 20816 17460 20868
rect 18328 20952 18380 21004
rect 19340 20952 19392 21004
rect 19984 20952 20036 21004
rect 20444 20952 20496 21004
rect 18144 20884 18196 20936
rect 18972 20884 19024 20936
rect 19800 20927 19852 20936
rect 19800 20893 19809 20927
rect 19809 20893 19843 20927
rect 19843 20893 19852 20927
rect 19800 20884 19852 20893
rect 21364 20884 21416 20936
rect 22008 20884 22060 20936
rect 22376 20884 22428 20936
rect 20168 20816 20220 20868
rect 15292 20748 15344 20757
rect 16580 20748 16632 20800
rect 16764 20748 16816 20800
rect 16948 20748 17000 20800
rect 18512 20791 18564 20800
rect 18512 20757 18521 20791
rect 18521 20757 18555 20791
rect 18555 20757 18564 20791
rect 18512 20748 18564 20757
rect 19984 20748 20036 20800
rect 20720 20748 20772 20800
rect 10880 20646 10932 20698
rect 10944 20646 10996 20698
rect 11008 20646 11060 20698
rect 11072 20646 11124 20698
rect 11136 20646 11188 20698
rect 20811 20646 20863 20698
rect 20875 20646 20927 20698
rect 20939 20646 20991 20698
rect 21003 20646 21055 20698
rect 21067 20646 21119 20698
rect 2136 20544 2188 20596
rect 5172 20587 5224 20596
rect 5172 20553 5181 20587
rect 5181 20553 5215 20587
rect 5215 20553 5224 20587
rect 5172 20544 5224 20553
rect 8024 20587 8076 20596
rect 8024 20553 8033 20587
rect 8033 20553 8067 20587
rect 8067 20553 8076 20587
rect 8024 20544 8076 20553
rect 8392 20544 8444 20596
rect 9312 20587 9364 20596
rect 9312 20553 9321 20587
rect 9321 20553 9355 20587
rect 9355 20553 9364 20587
rect 9312 20544 9364 20553
rect 15292 20544 15344 20596
rect 17224 20544 17276 20596
rect 18512 20544 18564 20596
rect 19248 20587 19300 20596
rect 19248 20553 19257 20587
rect 19257 20553 19291 20587
rect 19291 20553 19300 20587
rect 20260 20587 20312 20596
rect 19248 20544 19300 20553
rect 20260 20553 20269 20587
rect 20269 20553 20303 20587
rect 20303 20553 20312 20587
rect 20260 20544 20312 20553
rect 20628 20544 20680 20596
rect 22284 20587 22336 20596
rect 22284 20553 22293 20587
rect 22293 20553 22327 20587
rect 22327 20553 22336 20587
rect 22284 20544 22336 20553
rect 1400 20408 1452 20460
rect 1676 20451 1728 20460
rect 1676 20417 1685 20451
rect 1685 20417 1719 20451
rect 1719 20417 1728 20451
rect 1676 20408 1728 20417
rect 1860 20476 1912 20528
rect 3056 20476 3108 20528
rect 4528 20476 4580 20528
rect 2964 20408 3016 20460
rect 7012 20476 7064 20528
rect 6920 20451 6972 20460
rect 6920 20417 6954 20451
rect 6954 20417 6972 20451
rect 6920 20408 6972 20417
rect 8300 20408 8352 20460
rect 1952 20340 2004 20392
rect 3792 20383 3844 20392
rect 3792 20349 3801 20383
rect 3801 20349 3835 20383
rect 3835 20349 3844 20383
rect 3792 20340 3844 20349
rect 6644 20383 6696 20392
rect 6644 20349 6653 20383
rect 6653 20349 6687 20383
rect 6687 20349 6696 20383
rect 6644 20340 6696 20349
rect 8944 20408 8996 20460
rect 10232 20476 10284 20528
rect 10600 20476 10652 20528
rect 10692 20476 10744 20528
rect 12164 20476 12216 20528
rect 10324 20340 10376 20392
rect 7656 20272 7708 20324
rect 7932 20272 7984 20324
rect 19064 20476 19116 20528
rect 19892 20476 19944 20528
rect 22008 20476 22060 20528
rect 22376 20476 22428 20528
rect 12440 20451 12492 20460
rect 12440 20417 12449 20451
rect 12449 20417 12483 20451
rect 12483 20417 12492 20451
rect 12440 20408 12492 20417
rect 13084 20408 13136 20460
rect 13452 20451 13504 20460
rect 13452 20417 13461 20451
rect 13461 20417 13495 20451
rect 13495 20417 13504 20451
rect 13452 20408 13504 20417
rect 16212 20408 16264 20460
rect 16764 20408 16816 20460
rect 14924 20340 14976 20392
rect 17408 20383 17460 20392
rect 17408 20349 17417 20383
rect 17417 20349 17451 20383
rect 17451 20349 17460 20383
rect 17408 20340 17460 20349
rect 17776 20408 17828 20460
rect 20720 20408 20772 20460
rect 19064 20383 19116 20392
rect 19064 20349 19073 20383
rect 19073 20349 19107 20383
rect 19107 20349 19116 20383
rect 19064 20340 19116 20349
rect 20444 20340 20496 20392
rect 21916 20340 21968 20392
rect 14096 20272 14148 20324
rect 14556 20272 14608 20324
rect 1860 20204 1912 20256
rect 6552 20204 6604 20256
rect 8944 20204 8996 20256
rect 9956 20204 10008 20256
rect 11612 20247 11664 20256
rect 11612 20213 11621 20247
rect 11621 20213 11655 20247
rect 11655 20213 11664 20247
rect 11612 20204 11664 20213
rect 13268 20204 13320 20256
rect 14464 20204 14516 20256
rect 16948 20204 17000 20256
rect 19432 20204 19484 20256
rect 5915 20102 5967 20154
rect 5979 20102 6031 20154
rect 6043 20102 6095 20154
rect 6107 20102 6159 20154
rect 6171 20102 6223 20154
rect 15846 20102 15898 20154
rect 15910 20102 15962 20154
rect 15974 20102 16026 20154
rect 16038 20102 16090 20154
rect 16102 20102 16154 20154
rect 25776 20102 25828 20154
rect 25840 20102 25892 20154
rect 25904 20102 25956 20154
rect 25968 20102 26020 20154
rect 26032 20102 26084 20154
rect 6920 20000 6972 20052
rect 7196 20000 7248 20052
rect 3240 19975 3292 19984
rect 3240 19941 3249 19975
rect 3249 19941 3283 19975
rect 3283 19941 3292 19975
rect 3240 19932 3292 19941
rect 4436 19907 4488 19916
rect 4436 19873 4445 19907
rect 4445 19873 4479 19907
rect 4479 19873 4488 19907
rect 4436 19864 4488 19873
rect 2872 19796 2924 19848
rect 4252 19839 4304 19848
rect 2228 19728 2280 19780
rect 4252 19805 4261 19839
rect 4261 19805 4295 19839
rect 4295 19805 4304 19839
rect 4252 19796 4304 19805
rect 4344 19839 4396 19848
rect 4344 19805 4353 19839
rect 4353 19805 4387 19839
rect 4387 19805 4396 19839
rect 4344 19796 4396 19805
rect 5172 19796 5224 19848
rect 4712 19728 4764 19780
rect 5816 19864 5868 19916
rect 7012 19932 7064 19984
rect 9128 20000 9180 20052
rect 9772 20000 9824 20052
rect 8208 19932 8260 19984
rect 9680 19932 9732 19984
rect 6368 19839 6420 19848
rect 6368 19805 6377 19839
rect 6377 19805 6411 19839
rect 6411 19805 6420 19839
rect 6368 19796 6420 19805
rect 6828 19864 6880 19916
rect 7196 19864 7248 19916
rect 10324 19864 10376 19916
rect 7932 19796 7984 19848
rect 8024 19839 8076 19848
rect 8024 19805 8033 19839
rect 8033 19805 8067 19839
rect 8067 19805 8076 19839
rect 8024 19796 8076 19805
rect 8392 19796 8444 19848
rect 8760 19796 8812 19848
rect 9312 19796 9364 19848
rect 9680 19839 9732 19848
rect 9680 19805 9689 19839
rect 9689 19805 9723 19839
rect 9723 19805 9732 19839
rect 9680 19796 9732 19805
rect 12532 20000 12584 20052
rect 13360 20000 13412 20052
rect 11428 19932 11480 19984
rect 14464 19975 14516 19984
rect 14464 19941 14473 19975
rect 14473 19941 14507 19975
rect 14507 19941 14516 19975
rect 16212 20000 16264 20052
rect 17224 20000 17276 20052
rect 17868 20000 17920 20052
rect 20168 20000 20220 20052
rect 14464 19932 14516 19941
rect 11520 19907 11572 19916
rect 11520 19873 11529 19907
rect 11529 19873 11563 19907
rect 11563 19873 11572 19907
rect 11520 19864 11572 19873
rect 1676 19660 1728 19712
rect 3424 19660 3476 19712
rect 4804 19703 4856 19712
rect 4804 19669 4813 19703
rect 4813 19669 4847 19703
rect 4847 19669 4856 19703
rect 4804 19660 4856 19669
rect 6276 19660 6328 19712
rect 8944 19728 8996 19780
rect 13544 19839 13596 19848
rect 9864 19728 9916 19780
rect 10048 19728 10100 19780
rect 10600 19728 10652 19780
rect 12256 19728 12308 19780
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 14096 19839 14148 19848
rect 14096 19805 14105 19839
rect 14105 19805 14139 19839
rect 14139 19805 14148 19839
rect 14096 19796 14148 19805
rect 14740 19864 14792 19916
rect 15752 19907 15804 19916
rect 15752 19873 15761 19907
rect 15761 19873 15795 19907
rect 15795 19873 15804 19907
rect 15752 19864 15804 19873
rect 16028 19907 16080 19916
rect 16028 19873 16037 19907
rect 16037 19873 16071 19907
rect 16071 19873 16080 19907
rect 16028 19864 16080 19873
rect 16672 19864 16724 19916
rect 17592 19864 17644 19916
rect 19064 19864 19116 19916
rect 21640 19932 21692 19984
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 13452 19771 13504 19780
rect 13452 19737 13461 19771
rect 13461 19737 13495 19771
rect 13495 19737 13504 19771
rect 13452 19728 13504 19737
rect 15844 19839 15896 19848
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 15844 19796 15896 19805
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 16948 19796 17000 19848
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 19800 19796 19852 19848
rect 20260 19839 20312 19848
rect 20260 19805 20269 19839
rect 20269 19805 20303 19839
rect 20303 19805 20312 19839
rect 20260 19796 20312 19805
rect 20628 19796 20680 19848
rect 21916 19839 21968 19848
rect 21916 19805 21925 19839
rect 21925 19805 21959 19839
rect 21959 19805 21968 19839
rect 21916 19796 21968 19805
rect 22468 19796 22520 19848
rect 23020 19796 23072 19848
rect 7196 19660 7248 19712
rect 8024 19660 8076 19712
rect 11336 19660 11388 19712
rect 14740 19703 14792 19712
rect 14740 19669 14749 19703
rect 14749 19669 14783 19703
rect 14783 19669 14792 19703
rect 14740 19660 14792 19669
rect 15292 19660 15344 19712
rect 18604 19728 18656 19780
rect 17132 19660 17184 19712
rect 17592 19660 17644 19712
rect 20260 19660 20312 19712
rect 10880 19558 10932 19610
rect 10944 19558 10996 19610
rect 11008 19558 11060 19610
rect 11072 19558 11124 19610
rect 11136 19558 11188 19610
rect 20811 19558 20863 19610
rect 20875 19558 20927 19610
rect 20939 19558 20991 19610
rect 21003 19558 21055 19610
rect 21067 19558 21119 19610
rect 1308 19456 1360 19508
rect 1676 19184 1728 19236
rect 2504 19363 2556 19372
rect 2504 19329 2538 19363
rect 2538 19329 2556 19363
rect 4804 19388 4856 19440
rect 8392 19388 8444 19440
rect 9312 19431 9364 19440
rect 9312 19397 9321 19431
rect 9321 19397 9355 19431
rect 9355 19397 9364 19431
rect 9312 19388 9364 19397
rect 10048 19431 10100 19440
rect 10048 19397 10057 19431
rect 10057 19397 10091 19431
rect 10091 19397 10100 19431
rect 10048 19388 10100 19397
rect 10232 19431 10284 19440
rect 10232 19397 10241 19431
rect 10241 19397 10275 19431
rect 10275 19397 10284 19431
rect 10232 19388 10284 19397
rect 2504 19320 2556 19329
rect 2872 19320 2924 19372
rect 3792 19320 3844 19372
rect 5172 19320 5224 19372
rect 6460 19363 6512 19372
rect 6460 19329 6469 19363
rect 6469 19329 6503 19363
rect 6503 19329 6512 19363
rect 8760 19363 8812 19372
rect 6460 19320 6512 19329
rect 8760 19329 8769 19363
rect 8769 19329 8803 19363
rect 8803 19329 8812 19363
rect 8760 19320 8812 19329
rect 9772 19320 9824 19372
rect 11428 19388 11480 19440
rect 12900 19456 12952 19508
rect 13176 19499 13228 19508
rect 13176 19465 13185 19499
rect 13185 19465 13219 19499
rect 13219 19465 13228 19499
rect 13176 19456 13228 19465
rect 13544 19456 13596 19508
rect 13268 19388 13320 19440
rect 15936 19456 15988 19508
rect 16304 19456 16356 19508
rect 16764 19456 16816 19508
rect 17592 19499 17644 19508
rect 14740 19388 14792 19440
rect 10692 19320 10744 19372
rect 10784 19320 10836 19372
rect 11336 19320 11388 19372
rect 15660 19320 15712 19372
rect 15752 19320 15804 19372
rect 2596 19116 2648 19168
rect 2872 19116 2924 19168
rect 3608 19159 3660 19168
rect 3608 19125 3617 19159
rect 3617 19125 3651 19159
rect 3651 19125 3660 19159
rect 3608 19116 3660 19125
rect 14188 19116 14240 19168
rect 17224 19320 17276 19372
rect 17592 19465 17601 19499
rect 17601 19465 17635 19499
rect 17635 19465 17644 19499
rect 17592 19456 17644 19465
rect 18788 19499 18840 19508
rect 18788 19465 18797 19499
rect 18797 19465 18831 19499
rect 18831 19465 18840 19499
rect 18788 19456 18840 19465
rect 21916 19456 21968 19508
rect 18236 19388 18288 19440
rect 19340 19388 19392 19440
rect 17592 19320 17644 19372
rect 17960 19363 18012 19372
rect 17960 19329 17969 19363
rect 17969 19329 18003 19363
rect 18003 19329 18012 19363
rect 17960 19320 18012 19329
rect 19984 19363 20036 19372
rect 19984 19329 19993 19363
rect 19993 19329 20027 19363
rect 20027 19329 20036 19363
rect 19984 19320 20036 19329
rect 20260 19363 20312 19372
rect 20260 19329 20269 19363
rect 20269 19329 20303 19363
rect 20303 19329 20312 19363
rect 20260 19320 20312 19329
rect 20444 19388 20496 19440
rect 20628 19388 20680 19440
rect 20536 19363 20588 19372
rect 18144 19252 18196 19304
rect 19248 19252 19300 19304
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 22008 19388 22060 19440
rect 22468 19363 22520 19372
rect 22468 19329 22477 19363
rect 22477 19329 22511 19363
rect 22511 19329 22520 19363
rect 22468 19320 22520 19329
rect 30104 19388 30156 19440
rect 29828 19363 29880 19372
rect 29828 19329 29837 19363
rect 29837 19329 29871 19363
rect 29871 19329 29880 19363
rect 29828 19320 29880 19329
rect 16764 19159 16816 19168
rect 16764 19125 16773 19159
rect 16773 19125 16807 19159
rect 16807 19125 16816 19159
rect 16764 19116 16816 19125
rect 19524 19116 19576 19168
rect 19984 19116 20036 19168
rect 20352 19116 20404 19168
rect 20444 19116 20496 19168
rect 30012 19159 30064 19168
rect 30012 19125 30021 19159
rect 30021 19125 30055 19159
rect 30055 19125 30064 19159
rect 30012 19116 30064 19125
rect 5915 19014 5967 19066
rect 5979 19014 6031 19066
rect 6043 19014 6095 19066
rect 6107 19014 6159 19066
rect 6171 19014 6223 19066
rect 15846 19014 15898 19066
rect 15910 19014 15962 19066
rect 15974 19014 16026 19066
rect 16038 19014 16090 19066
rect 16102 19014 16154 19066
rect 25776 19014 25828 19066
rect 25840 19014 25892 19066
rect 25904 19014 25956 19066
rect 25968 19014 26020 19066
rect 26032 19014 26084 19066
rect 2228 18955 2280 18964
rect 2228 18921 2237 18955
rect 2237 18921 2271 18955
rect 2271 18921 2280 18955
rect 2228 18912 2280 18921
rect 3792 18912 3844 18964
rect 12256 18955 12308 18964
rect 1676 18844 1728 18896
rect 3332 18844 3384 18896
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 1952 18776 2004 18828
rect 3608 18776 3660 18828
rect 1584 18708 1636 18760
rect 3240 18708 3292 18760
rect 3792 18751 3844 18760
rect 3792 18717 3801 18751
rect 3801 18717 3835 18751
rect 3835 18717 3844 18751
rect 3792 18708 3844 18717
rect 6368 18776 6420 18828
rect 6184 18751 6236 18760
rect 6184 18717 6193 18751
rect 6193 18717 6227 18751
rect 6227 18717 6236 18751
rect 6184 18708 6236 18717
rect 3332 18640 3384 18692
rect 4068 18640 4120 18692
rect 9036 18776 9088 18828
rect 7656 18751 7708 18760
rect 7656 18717 7665 18751
rect 7665 18717 7699 18751
rect 7699 18717 7708 18751
rect 7656 18708 7708 18717
rect 8024 18751 8076 18760
rect 8024 18717 8033 18751
rect 8033 18717 8067 18751
rect 8067 18717 8076 18751
rect 8024 18708 8076 18717
rect 6736 18640 6788 18692
rect 8392 18708 8444 18760
rect 9312 18751 9364 18760
rect 8852 18640 8904 18692
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 12256 18921 12265 18955
rect 12265 18921 12299 18955
rect 12299 18921 12308 18955
rect 12256 18912 12308 18921
rect 12440 18912 12492 18964
rect 16764 18912 16816 18964
rect 17960 18912 18012 18964
rect 19340 18955 19392 18964
rect 19340 18921 19349 18955
rect 19349 18921 19383 18955
rect 19383 18921 19392 18955
rect 19340 18912 19392 18921
rect 19984 18912 20036 18964
rect 20536 18912 20588 18964
rect 29920 18955 29972 18964
rect 29920 18921 29929 18955
rect 29929 18921 29963 18955
rect 29963 18921 29972 18955
rect 29920 18912 29972 18921
rect 11060 18887 11112 18896
rect 11060 18853 11069 18887
rect 11069 18853 11103 18887
rect 11103 18853 11112 18887
rect 11060 18844 11112 18853
rect 11980 18844 12032 18896
rect 14924 18844 14976 18896
rect 11428 18776 11480 18828
rect 11888 18819 11940 18828
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 3056 18615 3108 18624
rect 3056 18581 3065 18615
rect 3065 18581 3099 18615
rect 3099 18581 3108 18615
rect 3056 18572 3108 18581
rect 5540 18615 5592 18624
rect 5540 18581 5549 18615
rect 5549 18581 5583 18615
rect 5583 18581 5592 18615
rect 5540 18572 5592 18581
rect 7472 18615 7524 18624
rect 7472 18581 7481 18615
rect 7481 18581 7515 18615
rect 7515 18581 7524 18615
rect 7472 18572 7524 18581
rect 9956 18572 10008 18624
rect 10784 18640 10836 18692
rect 11612 18708 11664 18760
rect 11888 18785 11897 18819
rect 11897 18785 11931 18819
rect 11931 18785 11940 18819
rect 11888 18776 11940 18785
rect 12164 18776 12216 18828
rect 12532 18708 12584 18760
rect 12716 18751 12768 18760
rect 12716 18717 12725 18751
rect 12725 18717 12759 18751
rect 12759 18717 12768 18751
rect 12716 18708 12768 18717
rect 14188 18751 14240 18760
rect 14188 18717 14197 18751
rect 14197 18717 14231 18751
rect 14231 18717 14240 18751
rect 14188 18708 14240 18717
rect 17040 18776 17092 18828
rect 17316 18819 17368 18828
rect 17316 18785 17325 18819
rect 17325 18785 17359 18819
rect 17359 18785 17368 18819
rect 17316 18776 17368 18785
rect 18052 18844 18104 18896
rect 18144 18776 18196 18828
rect 19064 18776 19116 18828
rect 20444 18819 20496 18828
rect 16948 18708 17000 18760
rect 18788 18708 18840 18760
rect 18144 18640 18196 18692
rect 20444 18785 20453 18819
rect 20453 18785 20487 18819
rect 20487 18785 20496 18819
rect 20444 18776 20496 18785
rect 20352 18751 20404 18760
rect 20352 18717 20361 18751
rect 20361 18717 20395 18751
rect 20395 18717 20404 18751
rect 20352 18708 20404 18717
rect 21916 18776 21968 18828
rect 22008 18751 22060 18760
rect 22008 18717 22017 18751
rect 22017 18717 22051 18751
rect 22051 18717 22060 18751
rect 22008 18708 22060 18717
rect 22468 18708 22520 18760
rect 29644 18708 29696 18760
rect 30104 18751 30156 18760
rect 30104 18717 30113 18751
rect 30113 18717 30147 18751
rect 30147 18717 30156 18751
rect 30104 18708 30156 18717
rect 13636 18572 13688 18624
rect 15384 18572 15436 18624
rect 19800 18572 19852 18624
rect 10880 18470 10932 18522
rect 10944 18470 10996 18522
rect 11008 18470 11060 18522
rect 11072 18470 11124 18522
rect 11136 18470 11188 18522
rect 20811 18470 20863 18522
rect 20875 18470 20927 18522
rect 20939 18470 20991 18522
rect 21003 18470 21055 18522
rect 21067 18470 21119 18522
rect 2504 18368 2556 18420
rect 4436 18368 4488 18420
rect 5724 18411 5776 18420
rect 5724 18377 5733 18411
rect 5733 18377 5767 18411
rect 5767 18377 5776 18411
rect 5724 18368 5776 18377
rect 7656 18368 7708 18420
rect 8760 18368 8812 18420
rect 9496 18368 9548 18420
rect 12072 18411 12124 18420
rect 12072 18377 12081 18411
rect 12081 18377 12115 18411
rect 12115 18377 12124 18411
rect 12072 18368 12124 18377
rect 15384 18411 15436 18420
rect 15384 18377 15393 18411
rect 15393 18377 15427 18411
rect 15427 18377 15436 18411
rect 15384 18368 15436 18377
rect 18972 18411 19024 18420
rect 18972 18377 18981 18411
rect 18981 18377 19015 18411
rect 19015 18377 19024 18411
rect 18972 18368 19024 18377
rect 19340 18411 19392 18420
rect 19340 18377 19349 18411
rect 19349 18377 19383 18411
rect 19383 18377 19392 18411
rect 19340 18368 19392 18377
rect 19708 18368 19760 18420
rect 20628 18368 20680 18420
rect 20720 18368 20772 18420
rect 29828 18368 29880 18420
rect 1676 18275 1728 18284
rect 1676 18241 1685 18275
rect 1685 18241 1719 18275
rect 1719 18241 1728 18275
rect 1676 18232 1728 18241
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 2872 18232 2924 18284
rect 2964 18232 3016 18284
rect 5816 18300 5868 18352
rect 6184 18300 6236 18352
rect 7472 18300 7524 18352
rect 7564 18300 7616 18352
rect 8024 18300 8076 18352
rect 9680 18300 9732 18352
rect 4068 18232 4120 18284
rect 4160 18232 4212 18284
rect 1768 18164 1820 18216
rect 3148 18164 3200 18216
rect 2596 18096 2648 18148
rect 3884 18164 3936 18216
rect 6644 18232 6696 18284
rect 9956 18275 10008 18284
rect 10784 18300 10836 18352
rect 12716 18300 12768 18352
rect 15292 18343 15344 18352
rect 15292 18309 15301 18343
rect 15301 18309 15335 18343
rect 15335 18309 15344 18343
rect 15292 18300 15344 18309
rect 19524 18300 19576 18352
rect 9956 18241 9974 18275
rect 9974 18241 10008 18275
rect 9956 18232 10008 18241
rect 10600 18096 10652 18148
rect 12624 18232 12676 18284
rect 14004 18232 14056 18284
rect 17684 18232 17736 18284
rect 19156 18232 19208 18284
rect 19708 18232 19760 18284
rect 21824 18232 21876 18284
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 29276 18232 29328 18284
rect 30104 18275 30156 18284
rect 30104 18241 30113 18275
rect 30113 18241 30147 18275
rect 30147 18241 30156 18275
rect 30104 18232 30156 18241
rect 16672 18164 16724 18216
rect 16764 18164 16816 18216
rect 17408 18164 17460 18216
rect 19248 18164 19300 18216
rect 16212 18096 16264 18148
rect 17592 18096 17644 18148
rect 2872 18071 2924 18080
rect 2872 18037 2881 18071
rect 2881 18037 2915 18071
rect 2915 18037 2924 18071
rect 2872 18028 2924 18037
rect 5724 18028 5776 18080
rect 6644 18028 6696 18080
rect 7288 18028 7340 18080
rect 7840 18028 7892 18080
rect 14648 18028 14700 18080
rect 5915 17926 5967 17978
rect 5979 17926 6031 17978
rect 6043 17926 6095 17978
rect 6107 17926 6159 17978
rect 6171 17926 6223 17978
rect 15846 17926 15898 17978
rect 15910 17926 15962 17978
rect 15974 17926 16026 17978
rect 16038 17926 16090 17978
rect 16102 17926 16154 17978
rect 25776 17926 25828 17978
rect 25840 17926 25892 17978
rect 25904 17926 25956 17978
rect 25968 17926 26020 17978
rect 26032 17926 26084 17978
rect 5816 17824 5868 17876
rect 7932 17867 7984 17876
rect 7932 17833 7941 17867
rect 7941 17833 7975 17867
rect 7975 17833 7984 17867
rect 7932 17824 7984 17833
rect 11244 17824 11296 17876
rect 4620 17756 4672 17808
rect 3792 17731 3844 17740
rect 3792 17697 3801 17731
rect 3801 17697 3835 17731
rect 3835 17697 3844 17731
rect 3792 17688 3844 17697
rect 3976 17688 4028 17740
rect 15752 17824 15804 17876
rect 17040 17824 17092 17876
rect 19248 17824 19300 17876
rect 22008 17824 22060 17876
rect 14464 17799 14516 17808
rect 14464 17765 14473 17799
rect 14473 17765 14507 17799
rect 14507 17765 14516 17799
rect 14464 17756 14516 17765
rect 1676 17620 1728 17672
rect 2872 17620 2924 17672
rect 4068 17663 4120 17672
rect 4068 17629 4077 17663
rect 4077 17629 4111 17663
rect 4111 17629 4120 17663
rect 4068 17620 4120 17629
rect 3884 17552 3936 17604
rect 7656 17620 7708 17672
rect 9680 17620 9732 17672
rect 7472 17552 7524 17604
rect 9128 17552 9180 17604
rect 13268 17663 13320 17672
rect 13268 17629 13277 17663
rect 13277 17629 13311 17663
rect 13311 17629 13320 17663
rect 14096 17663 14148 17672
rect 13268 17620 13320 17629
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 14372 17731 14424 17740
rect 14372 17697 14381 17731
rect 14381 17697 14415 17731
rect 14415 17697 14424 17731
rect 14372 17688 14424 17697
rect 18052 17756 18104 17808
rect 18236 17756 18288 17808
rect 15476 17688 15528 17740
rect 2964 17527 3016 17536
rect 2964 17493 2973 17527
rect 2973 17493 3007 17527
rect 3007 17493 3016 17527
rect 2964 17484 3016 17493
rect 5080 17527 5132 17536
rect 5080 17493 5089 17527
rect 5089 17493 5123 17527
rect 5123 17493 5132 17527
rect 5080 17484 5132 17493
rect 8760 17484 8812 17536
rect 9220 17484 9272 17536
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 13544 17552 13596 17604
rect 16764 17688 16816 17740
rect 19340 17688 19392 17740
rect 16304 17620 16356 17672
rect 17868 17663 17920 17672
rect 17868 17629 17877 17663
rect 17877 17629 17911 17663
rect 17911 17629 17920 17663
rect 17868 17620 17920 17629
rect 18144 17663 18196 17672
rect 18144 17629 18153 17663
rect 18153 17629 18187 17663
rect 18187 17629 18196 17663
rect 18144 17620 18196 17629
rect 19524 17756 19576 17808
rect 17040 17552 17092 17604
rect 16672 17484 16724 17536
rect 20168 17688 20220 17740
rect 19984 17620 20036 17672
rect 20628 17620 20680 17672
rect 21272 17620 21324 17672
rect 21272 17484 21324 17536
rect 10880 17382 10932 17434
rect 10944 17382 10996 17434
rect 11008 17382 11060 17434
rect 11072 17382 11124 17434
rect 11136 17382 11188 17434
rect 20811 17382 20863 17434
rect 20875 17382 20927 17434
rect 20939 17382 20991 17434
rect 21003 17382 21055 17434
rect 21067 17382 21119 17434
rect 7472 17323 7524 17332
rect 7472 17289 7481 17323
rect 7481 17289 7515 17323
rect 7515 17289 7524 17323
rect 7472 17280 7524 17289
rect 9128 17323 9180 17332
rect 9128 17289 9137 17323
rect 9137 17289 9171 17323
rect 9171 17289 9180 17323
rect 9128 17280 9180 17289
rect 9404 17280 9456 17332
rect 9588 17323 9640 17332
rect 9588 17289 9597 17323
rect 9597 17289 9631 17323
rect 9631 17289 9640 17323
rect 9588 17280 9640 17289
rect 13268 17280 13320 17332
rect 13728 17280 13780 17332
rect 14556 17280 14608 17332
rect 15200 17280 15252 17332
rect 16948 17323 17000 17332
rect 16948 17289 16957 17323
rect 16957 17289 16991 17323
rect 16991 17289 17000 17323
rect 16948 17280 17000 17289
rect 19248 17280 19300 17332
rect 20168 17280 20220 17332
rect 21824 17280 21876 17332
rect 1400 17187 1452 17196
rect 1400 17153 1409 17187
rect 1409 17153 1443 17187
rect 1443 17153 1452 17187
rect 1400 17144 1452 17153
rect 2596 17187 2648 17196
rect 2596 17153 2605 17187
rect 2605 17153 2639 17187
rect 2639 17153 2648 17187
rect 2596 17144 2648 17153
rect 4528 17144 4580 17196
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 6736 17144 6788 17153
rect 7196 17144 7248 17196
rect 7932 17144 7984 17196
rect 8392 17187 8444 17196
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 8760 17212 8812 17264
rect 8852 17144 8904 17196
rect 11244 17212 11296 17264
rect 12532 17212 12584 17264
rect 13912 17212 13964 17264
rect 10876 17144 10928 17196
rect 14004 17187 14056 17196
rect 14004 17153 14013 17187
rect 14013 17153 14047 17187
rect 14047 17153 14056 17187
rect 14004 17144 14056 17153
rect 15292 17212 15344 17264
rect 17224 17212 17276 17264
rect 17868 17212 17920 17264
rect 19340 17212 19392 17264
rect 17040 17144 17092 17196
rect 17776 17144 17828 17196
rect 3240 17076 3292 17128
rect 3700 17076 3752 17128
rect 3884 17119 3936 17128
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 8760 17119 8812 17128
rect 8760 17085 8769 17119
rect 8769 17085 8803 17119
rect 8803 17085 8812 17119
rect 8760 17076 8812 17085
rect 9036 17076 9088 17128
rect 11704 17119 11756 17128
rect 11704 17085 11713 17119
rect 11713 17085 11747 17119
rect 11747 17085 11756 17119
rect 11704 17076 11756 17085
rect 14188 17076 14240 17128
rect 17224 17119 17276 17128
rect 17224 17085 17233 17119
rect 17233 17085 17267 17119
rect 17267 17085 17276 17119
rect 18604 17144 18656 17196
rect 17224 17076 17276 17085
rect 18512 17076 18564 17128
rect 19340 17076 19392 17128
rect 19156 17008 19208 17060
rect 19800 17008 19852 17060
rect 21272 17144 21324 17196
rect 21824 17187 21876 17196
rect 21824 17153 21833 17187
rect 21833 17153 21867 17187
rect 21867 17153 21876 17187
rect 21824 17144 21876 17153
rect 29920 17144 29972 17196
rect 20352 17076 20404 17128
rect 20628 17119 20680 17128
rect 20628 17085 20637 17119
rect 20637 17085 20671 17119
rect 20671 17085 20680 17119
rect 20628 17076 20680 17085
rect 2320 16940 2372 16992
rect 4988 16940 5040 16992
rect 12808 16940 12860 16992
rect 13728 16940 13780 16992
rect 15108 16940 15160 16992
rect 20444 16940 20496 16992
rect 30012 16983 30064 16992
rect 30012 16949 30021 16983
rect 30021 16949 30055 16983
rect 30055 16949 30064 16983
rect 30012 16940 30064 16949
rect 5915 16838 5967 16890
rect 5979 16838 6031 16890
rect 6043 16838 6095 16890
rect 6107 16838 6159 16890
rect 6171 16838 6223 16890
rect 15846 16838 15898 16890
rect 15910 16838 15962 16890
rect 15974 16838 16026 16890
rect 16038 16838 16090 16890
rect 16102 16838 16154 16890
rect 25776 16838 25828 16890
rect 25840 16838 25892 16890
rect 25904 16838 25956 16890
rect 25968 16838 26020 16890
rect 26032 16838 26084 16890
rect 2964 16736 3016 16788
rect 3700 16600 3752 16652
rect 1216 16532 1268 16584
rect 2872 16532 2924 16584
rect 3240 16575 3292 16584
rect 3240 16541 3249 16575
rect 3249 16541 3283 16575
rect 3283 16541 3292 16575
rect 3240 16532 3292 16541
rect 3424 16532 3476 16584
rect 3976 16532 4028 16584
rect 10876 16736 10928 16788
rect 14464 16736 14516 16788
rect 17224 16779 17276 16788
rect 17224 16745 17233 16779
rect 17233 16745 17267 16779
rect 17267 16745 17276 16779
rect 17224 16736 17276 16745
rect 20352 16736 20404 16788
rect 21824 16736 21876 16788
rect 8852 16668 8904 16720
rect 8760 16600 8812 16652
rect 9312 16600 9364 16652
rect 13360 16668 13412 16720
rect 13452 16668 13504 16720
rect 15108 16711 15160 16720
rect 15108 16677 15117 16711
rect 15117 16677 15151 16711
rect 15151 16677 15160 16711
rect 15108 16668 15160 16677
rect 19984 16668 20036 16720
rect 4252 16464 4304 16516
rect 9404 16464 9456 16516
rect 10140 16532 10192 16584
rect 10416 16575 10468 16584
rect 10416 16541 10425 16575
rect 10425 16541 10459 16575
rect 10459 16541 10468 16575
rect 10416 16532 10468 16541
rect 11980 16575 12032 16584
rect 2688 16396 2740 16448
rect 5724 16439 5776 16448
rect 5724 16405 5733 16439
rect 5733 16405 5767 16439
rect 5767 16405 5776 16439
rect 5724 16396 5776 16405
rect 6276 16439 6328 16448
rect 6276 16405 6285 16439
rect 6285 16405 6319 16439
rect 6319 16405 6328 16439
rect 6276 16396 6328 16405
rect 7748 16396 7800 16448
rect 9588 16396 9640 16448
rect 11980 16541 11989 16575
rect 11989 16541 12023 16575
rect 12023 16541 12032 16575
rect 11980 16532 12032 16541
rect 12808 16532 12860 16584
rect 16948 16600 17000 16652
rect 13912 16532 13964 16584
rect 14556 16575 14608 16584
rect 13084 16464 13136 16516
rect 14556 16541 14565 16575
rect 14565 16541 14599 16575
rect 14599 16541 14608 16575
rect 14556 16532 14608 16541
rect 15292 16575 15344 16584
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15292 16532 15344 16541
rect 16764 16532 16816 16584
rect 17040 16575 17092 16584
rect 17040 16541 17049 16575
rect 17049 16541 17083 16575
rect 17083 16541 17092 16575
rect 17040 16532 17092 16541
rect 18144 16532 18196 16584
rect 19616 16600 19668 16652
rect 19524 16532 19576 16584
rect 20444 16532 20496 16584
rect 11244 16396 11296 16448
rect 13360 16396 13412 16448
rect 16304 16396 16356 16448
rect 16856 16396 16908 16448
rect 19248 16464 19300 16516
rect 18604 16396 18656 16448
rect 10880 16294 10932 16346
rect 10944 16294 10996 16346
rect 11008 16294 11060 16346
rect 11072 16294 11124 16346
rect 11136 16294 11188 16346
rect 20811 16294 20863 16346
rect 20875 16294 20927 16346
rect 20939 16294 20991 16346
rect 21003 16294 21055 16346
rect 21067 16294 21119 16346
rect 1768 16056 1820 16108
rect 3792 16192 3844 16244
rect 4068 16192 4120 16244
rect 4252 16235 4304 16244
rect 4252 16201 4261 16235
rect 4261 16201 4295 16235
rect 4295 16201 4304 16235
rect 4252 16192 4304 16201
rect 5172 16192 5224 16244
rect 7196 16235 7248 16244
rect 5080 16124 5132 16176
rect 4988 16099 5040 16108
rect 1676 16031 1728 16040
rect 1676 15997 1685 16031
rect 1685 15997 1719 16031
rect 1719 15997 1728 16031
rect 1676 15988 1728 15997
rect 2872 15988 2924 16040
rect 3884 16031 3936 16040
rect 3884 15997 3893 16031
rect 3893 15997 3927 16031
rect 3927 15997 3936 16031
rect 4988 16065 4997 16099
rect 4997 16065 5031 16099
rect 5031 16065 5040 16099
rect 4988 16056 5040 16065
rect 7196 16201 7205 16235
rect 7205 16201 7239 16235
rect 7239 16201 7248 16235
rect 7196 16192 7248 16201
rect 9588 16192 9640 16244
rect 11428 16192 11480 16244
rect 14004 16192 14056 16244
rect 18144 16192 18196 16244
rect 19064 16192 19116 16244
rect 7472 16124 7524 16176
rect 11244 16124 11296 16176
rect 3884 15988 3936 15997
rect 5724 15988 5776 16040
rect 1952 15852 2004 15904
rect 8116 16056 8168 16108
rect 9680 16056 9732 16108
rect 9864 16099 9916 16108
rect 9864 16065 9898 16099
rect 9898 16065 9916 16099
rect 12808 16099 12860 16108
rect 9864 16056 9916 16065
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 14096 16056 14148 16108
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 19524 16124 19576 16176
rect 14464 16056 14516 16065
rect 17224 16099 17276 16108
rect 17224 16065 17258 16099
rect 17258 16065 17276 16099
rect 17224 16056 17276 16065
rect 18236 16056 18288 16108
rect 19064 16099 19116 16108
rect 19064 16065 19073 16099
rect 19073 16065 19107 16099
rect 19107 16065 19116 16099
rect 19064 16056 19116 16065
rect 19248 16099 19300 16108
rect 19248 16065 19257 16099
rect 19257 16065 19291 16099
rect 19291 16065 19300 16099
rect 19248 16056 19300 16065
rect 19432 16099 19484 16108
rect 19432 16065 19441 16099
rect 19441 16065 19475 16099
rect 19475 16065 19484 16099
rect 19432 16056 19484 16065
rect 29368 16192 29420 16244
rect 20352 16124 20404 16176
rect 21272 16124 21324 16176
rect 20812 16056 20864 16108
rect 21180 16099 21232 16108
rect 21180 16065 21189 16099
rect 21189 16065 21223 16099
rect 21223 16065 21232 16099
rect 21180 16056 21232 16065
rect 21640 16056 21692 16108
rect 29000 16056 29052 16108
rect 30104 16099 30156 16108
rect 30104 16065 30113 16099
rect 30113 16065 30147 16099
rect 30147 16065 30156 16099
rect 30104 16056 30156 16065
rect 8852 15988 8904 16040
rect 13360 15988 13412 16040
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 19340 15988 19392 16040
rect 5080 15895 5132 15904
rect 5080 15861 5089 15895
rect 5089 15861 5123 15895
rect 5123 15861 5132 15895
rect 5080 15852 5132 15861
rect 6920 15920 6972 15972
rect 7012 15852 7064 15904
rect 7196 15852 7248 15904
rect 10508 15852 10560 15904
rect 13268 15852 13320 15904
rect 13452 15852 13504 15904
rect 15108 15852 15160 15904
rect 16212 15852 16264 15904
rect 16764 15852 16816 15904
rect 17316 15852 17368 15904
rect 19708 15852 19760 15904
rect 20720 15852 20772 15904
rect 5915 15750 5967 15802
rect 5979 15750 6031 15802
rect 6043 15750 6095 15802
rect 6107 15750 6159 15802
rect 6171 15750 6223 15802
rect 15846 15750 15898 15802
rect 15910 15750 15962 15802
rect 15974 15750 16026 15802
rect 16038 15750 16090 15802
rect 16102 15750 16154 15802
rect 25776 15750 25828 15802
rect 25840 15750 25892 15802
rect 25904 15750 25956 15802
rect 25968 15750 26020 15802
rect 26032 15750 26084 15802
rect 1768 15691 1820 15700
rect 1768 15657 1777 15691
rect 1777 15657 1811 15691
rect 1811 15657 1820 15691
rect 1768 15648 1820 15657
rect 4528 15691 4580 15700
rect 4528 15657 4537 15691
rect 4537 15657 4571 15691
rect 4571 15657 4580 15691
rect 4528 15648 4580 15657
rect 3148 15580 3200 15632
rect 1952 15487 2004 15496
rect 1952 15453 1961 15487
rect 1961 15453 1995 15487
rect 1995 15453 2004 15487
rect 1952 15444 2004 15453
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2780 15512 2832 15564
rect 3884 15512 3936 15564
rect 2320 15444 2372 15453
rect 3148 15487 3200 15496
rect 3148 15453 3157 15487
rect 3157 15453 3191 15487
rect 3191 15453 3200 15487
rect 3148 15444 3200 15453
rect 3792 15487 3844 15496
rect 3792 15453 3801 15487
rect 3801 15453 3835 15487
rect 3835 15453 3844 15487
rect 3792 15444 3844 15453
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 2872 15376 2924 15428
rect 4988 15444 5040 15496
rect 5080 15487 5132 15496
rect 5080 15453 5089 15487
rect 5089 15453 5123 15487
rect 5123 15453 5132 15487
rect 5080 15444 5132 15453
rect 5448 15444 5500 15496
rect 6460 15648 6512 15700
rect 6644 15648 6696 15700
rect 7656 15580 7708 15632
rect 9864 15648 9916 15700
rect 14740 15648 14792 15700
rect 16304 15648 16356 15700
rect 10140 15580 10192 15632
rect 6644 15512 6696 15564
rect 6184 15444 6236 15496
rect 8760 15512 8812 15564
rect 9404 15555 9456 15564
rect 7656 15487 7708 15496
rect 7656 15453 7666 15487
rect 7666 15453 7700 15487
rect 7700 15453 7708 15487
rect 7656 15444 7708 15453
rect 9404 15521 9413 15555
rect 9413 15521 9447 15555
rect 9447 15521 9456 15555
rect 9404 15512 9456 15521
rect 14096 15512 14148 15564
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 15200 15512 15252 15564
rect 9128 15444 9180 15496
rect 9588 15487 9640 15496
rect 6736 15376 6788 15428
rect 7380 15376 7432 15428
rect 7932 15419 7984 15428
rect 7932 15385 7941 15419
rect 7941 15385 7975 15419
rect 7975 15385 7984 15419
rect 9588 15453 9597 15487
rect 9597 15453 9631 15487
rect 9631 15453 9640 15487
rect 9588 15444 9640 15453
rect 9680 15444 9732 15496
rect 10048 15444 10100 15496
rect 13360 15444 13412 15496
rect 14740 15487 14792 15496
rect 14740 15453 14749 15487
rect 14749 15453 14783 15487
rect 14783 15453 14792 15487
rect 14740 15444 14792 15453
rect 7932 15376 7984 15385
rect 10324 15376 10376 15428
rect 11244 15376 11296 15428
rect 16580 15444 16632 15496
rect 16856 15580 16908 15632
rect 17224 15648 17276 15700
rect 20812 15691 20864 15700
rect 20812 15657 20821 15691
rect 20821 15657 20855 15691
rect 20855 15657 20864 15691
rect 20812 15648 20864 15657
rect 29460 15648 29512 15700
rect 19340 15512 19392 15564
rect 2964 15351 3016 15360
rect 2964 15317 2973 15351
rect 2973 15317 3007 15351
rect 3007 15317 3016 15351
rect 2964 15308 3016 15317
rect 5816 15308 5868 15360
rect 6460 15351 6512 15360
rect 6460 15317 6469 15351
rect 6469 15317 6503 15351
rect 6503 15317 6512 15351
rect 6460 15308 6512 15317
rect 7656 15308 7708 15360
rect 8116 15308 8168 15360
rect 8760 15308 8812 15360
rect 9312 15308 9364 15360
rect 9680 15308 9732 15360
rect 9864 15308 9916 15360
rect 10600 15308 10652 15360
rect 12532 15308 12584 15360
rect 14832 15308 14884 15360
rect 15108 15308 15160 15360
rect 16396 15376 16448 15428
rect 17040 15487 17092 15496
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 17224 15487 17276 15496
rect 17224 15453 17233 15487
rect 17233 15453 17267 15487
rect 17267 15453 17276 15487
rect 17224 15444 17276 15453
rect 17408 15444 17460 15496
rect 18604 15487 18656 15496
rect 18236 15376 18288 15428
rect 18604 15453 18613 15487
rect 18613 15453 18647 15487
rect 18647 15453 18656 15487
rect 18604 15444 18656 15453
rect 19524 15444 19576 15496
rect 19708 15487 19760 15496
rect 19708 15453 19742 15487
rect 19742 15453 19760 15487
rect 19708 15444 19760 15453
rect 21456 15444 21508 15496
rect 29920 15487 29972 15496
rect 29920 15453 29929 15487
rect 29929 15453 29963 15487
rect 29963 15453 29972 15487
rect 29920 15444 29972 15453
rect 30104 15487 30156 15496
rect 30104 15453 30113 15487
rect 30113 15453 30147 15487
rect 30147 15453 30156 15487
rect 30104 15444 30156 15453
rect 16948 15308 17000 15360
rect 19248 15308 19300 15360
rect 21824 15308 21876 15360
rect 10880 15206 10932 15258
rect 10944 15206 10996 15258
rect 11008 15206 11060 15258
rect 11072 15206 11124 15258
rect 11136 15206 11188 15258
rect 20811 15206 20863 15258
rect 20875 15206 20927 15258
rect 20939 15206 20991 15258
rect 21003 15206 21055 15258
rect 21067 15206 21119 15258
rect 1492 15104 1544 15156
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 3056 15036 3108 15088
rect 7380 15104 7432 15156
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 2504 14968 2556 15020
rect 2780 15011 2832 15020
rect 2780 14977 2789 15011
rect 2789 14977 2823 15011
rect 2823 14977 2832 15011
rect 2964 15011 3016 15020
rect 2780 14968 2832 14977
rect 2964 14977 2973 15011
rect 2973 14977 3007 15011
rect 3007 14977 3016 15011
rect 2964 14968 3016 14977
rect 8760 15079 8812 15088
rect 8760 15045 8778 15079
rect 8778 15045 8812 15079
rect 8760 15036 8812 15045
rect 9588 15036 9640 15088
rect 10048 15036 10100 15088
rect 10324 15036 10376 15088
rect 14832 15104 14884 15156
rect 16948 15104 17000 15156
rect 29920 15104 29972 15156
rect 1492 14764 1544 14816
rect 2872 14900 2924 14952
rect 2780 14764 2832 14816
rect 5724 14968 5776 15020
rect 6552 15011 6604 15020
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 6552 14968 6604 14977
rect 6644 15011 6696 15020
rect 6644 14977 6653 15011
rect 6653 14977 6687 15011
rect 6687 14977 6696 15011
rect 6920 15011 6972 15020
rect 6644 14968 6696 14977
rect 6920 14977 6929 15011
rect 6929 14977 6963 15011
rect 6963 14977 6972 15011
rect 6920 14968 6972 14977
rect 7104 14968 7156 15020
rect 3792 14900 3844 14952
rect 6736 14943 6788 14952
rect 6736 14909 6745 14943
rect 6745 14909 6779 14943
rect 6779 14909 6788 14943
rect 9312 14968 9364 15020
rect 13820 15036 13872 15088
rect 12348 14968 12400 15020
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 13268 15011 13320 15020
rect 12532 14968 12584 14977
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 13544 14968 13596 15020
rect 14464 15011 14516 15020
rect 14464 14977 14473 15011
rect 14473 14977 14507 15011
rect 14507 14977 14516 15011
rect 14464 14968 14516 14977
rect 14556 14968 14608 15020
rect 17040 15036 17092 15088
rect 18880 15036 18932 15088
rect 19432 15036 19484 15088
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 17224 14968 17276 15020
rect 6736 14900 6788 14909
rect 12808 14900 12860 14952
rect 16304 14900 16356 14952
rect 17868 14968 17920 15020
rect 18512 15011 18564 15020
rect 17960 14900 18012 14952
rect 18512 14977 18521 15011
rect 18521 14977 18555 15011
rect 18555 14977 18564 15011
rect 18512 14968 18564 14977
rect 18604 15011 18656 15020
rect 18604 14977 18618 15011
rect 18618 14977 18652 15011
rect 18652 14977 18656 15011
rect 18604 14968 18656 14977
rect 19616 14968 19668 15020
rect 19800 14968 19852 15020
rect 20536 14968 20588 15020
rect 21824 15011 21876 15020
rect 20628 14900 20680 14952
rect 21824 14977 21833 15011
rect 21833 14977 21867 15011
rect 21867 14977 21876 15011
rect 21824 14968 21876 14977
rect 5908 14832 5960 14884
rect 6552 14832 6604 14884
rect 5080 14764 5132 14816
rect 6460 14764 6512 14816
rect 8024 14764 8076 14816
rect 10600 14764 10652 14816
rect 13268 14807 13320 14816
rect 13268 14773 13277 14807
rect 13277 14773 13311 14807
rect 13311 14773 13320 14807
rect 13268 14764 13320 14773
rect 29920 14968 29972 15020
rect 30104 14900 30156 14952
rect 29184 14875 29236 14884
rect 29184 14841 29193 14875
rect 29193 14841 29227 14875
rect 29227 14841 29236 14875
rect 29184 14832 29236 14841
rect 30012 14875 30064 14884
rect 30012 14841 30021 14875
rect 30021 14841 30055 14875
rect 30055 14841 30064 14875
rect 30012 14832 30064 14841
rect 16212 14764 16264 14816
rect 16948 14764 17000 14816
rect 17316 14764 17368 14816
rect 18604 14764 18656 14816
rect 19340 14764 19392 14816
rect 5915 14662 5967 14714
rect 5979 14662 6031 14714
rect 6043 14662 6095 14714
rect 6107 14662 6159 14714
rect 6171 14662 6223 14714
rect 15846 14662 15898 14714
rect 15910 14662 15962 14714
rect 15974 14662 16026 14714
rect 16038 14662 16090 14714
rect 16102 14662 16154 14714
rect 25776 14662 25828 14714
rect 25840 14662 25892 14714
rect 25904 14662 25956 14714
rect 25968 14662 26020 14714
rect 26032 14662 26084 14714
rect 2136 14560 2188 14612
rect 5172 14603 5224 14612
rect 2872 14492 2924 14544
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 2688 14399 2740 14408
rect 2688 14365 2697 14399
rect 2697 14365 2731 14399
rect 2731 14365 2740 14399
rect 2688 14356 2740 14365
rect 2964 14356 3016 14408
rect 5172 14569 5181 14603
rect 5181 14569 5215 14603
rect 5215 14569 5224 14603
rect 5172 14560 5224 14569
rect 5908 14467 5960 14476
rect 5908 14433 5917 14467
rect 5917 14433 5951 14467
rect 5951 14433 5960 14467
rect 5908 14424 5960 14433
rect 3792 14399 3844 14408
rect 3792 14365 3801 14399
rect 3801 14365 3835 14399
rect 3835 14365 3844 14399
rect 3792 14356 3844 14365
rect 5540 14356 5592 14408
rect 5816 14399 5868 14408
rect 5816 14365 5825 14399
rect 5825 14365 5859 14399
rect 5859 14365 5868 14399
rect 5816 14356 5868 14365
rect 6828 14560 6880 14612
rect 7196 14560 7248 14612
rect 7380 14560 7432 14612
rect 8116 14603 8168 14612
rect 8116 14569 8125 14603
rect 8125 14569 8159 14603
rect 8159 14569 8168 14603
rect 8116 14560 8168 14569
rect 9588 14603 9640 14612
rect 9588 14569 9597 14603
rect 9597 14569 9631 14603
rect 9631 14569 9640 14603
rect 9588 14560 9640 14569
rect 8024 14492 8076 14544
rect 6920 14424 6972 14476
rect 7104 14467 7156 14476
rect 7104 14433 7113 14467
rect 7113 14433 7147 14467
rect 7147 14433 7156 14467
rect 7104 14424 7156 14433
rect 8116 14424 8168 14476
rect 6736 14356 6788 14408
rect 7012 14399 7064 14408
rect 7012 14365 7021 14399
rect 7021 14365 7055 14399
rect 7055 14365 7064 14399
rect 7012 14356 7064 14365
rect 7196 14399 7248 14408
rect 7196 14365 7205 14399
rect 7205 14365 7239 14399
rect 7239 14365 7248 14399
rect 7196 14356 7248 14365
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 8944 14399 8996 14408
rect 8944 14365 8953 14399
rect 8953 14365 8987 14399
rect 8987 14365 8996 14399
rect 8944 14356 8996 14365
rect 9588 14424 9640 14476
rect 12072 14492 12124 14544
rect 13360 14492 13412 14544
rect 14556 14560 14608 14612
rect 16672 14560 16724 14612
rect 18604 14560 18656 14612
rect 20720 14560 20772 14612
rect 29920 14603 29972 14612
rect 29920 14569 29929 14603
rect 29929 14569 29963 14603
rect 29963 14569 29972 14603
rect 29920 14560 29972 14569
rect 29000 14492 29052 14544
rect 8300 14288 8352 14340
rect 7564 14263 7616 14272
rect 7564 14229 7573 14263
rect 7573 14229 7607 14263
rect 7607 14229 7616 14263
rect 7564 14220 7616 14229
rect 8484 14288 8536 14340
rect 9404 14399 9456 14408
rect 9404 14365 9418 14399
rect 9418 14365 9452 14399
rect 9452 14365 9456 14399
rect 9404 14356 9456 14365
rect 9496 14288 9548 14340
rect 10600 14424 10652 14476
rect 11704 14424 11756 14476
rect 12164 14467 12216 14476
rect 12164 14433 12173 14467
rect 12173 14433 12207 14467
rect 12207 14433 12216 14467
rect 12164 14424 12216 14433
rect 14924 14467 14976 14476
rect 14924 14433 14933 14467
rect 14933 14433 14967 14467
rect 14967 14433 14976 14467
rect 14924 14424 14976 14433
rect 10048 14356 10100 14408
rect 10876 14356 10928 14408
rect 11520 14399 11572 14408
rect 11520 14365 11529 14399
rect 11529 14365 11563 14399
rect 11563 14365 11572 14399
rect 11520 14356 11572 14365
rect 13268 14356 13320 14408
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 14832 14399 14884 14408
rect 14832 14365 14841 14399
rect 14841 14365 14875 14399
rect 14875 14365 14884 14399
rect 14832 14356 14884 14365
rect 16120 14424 16172 14476
rect 16304 14467 16356 14476
rect 16304 14433 16313 14467
rect 16313 14433 16347 14467
rect 16347 14433 16356 14467
rect 16304 14424 16356 14433
rect 15200 14399 15252 14408
rect 15200 14365 15209 14399
rect 15209 14365 15243 14399
rect 15243 14365 15252 14399
rect 15200 14356 15252 14365
rect 16396 14356 16448 14408
rect 16764 14424 16816 14476
rect 17224 14424 17276 14476
rect 17408 14467 17460 14476
rect 17408 14433 17417 14467
rect 17417 14433 17451 14467
rect 17451 14433 17460 14467
rect 17408 14424 17460 14433
rect 29644 14424 29696 14476
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 17592 14399 17644 14408
rect 17592 14365 17601 14399
rect 17601 14365 17635 14399
rect 17635 14365 17644 14399
rect 17592 14356 17644 14365
rect 17960 14356 18012 14408
rect 18328 14399 18380 14408
rect 18328 14365 18337 14399
rect 18337 14365 18371 14399
rect 18371 14365 18380 14399
rect 18328 14356 18380 14365
rect 19800 14399 19852 14408
rect 19800 14365 19809 14399
rect 19809 14365 19843 14399
rect 19843 14365 19852 14399
rect 19800 14356 19852 14365
rect 20076 14399 20128 14408
rect 20076 14365 20085 14399
rect 20085 14365 20119 14399
rect 20119 14365 20128 14399
rect 20076 14356 20128 14365
rect 20628 14356 20680 14408
rect 21180 14356 21232 14408
rect 10140 14331 10192 14340
rect 10140 14297 10149 14331
rect 10149 14297 10183 14331
rect 10183 14297 10192 14331
rect 10140 14288 10192 14297
rect 10324 14331 10376 14340
rect 10324 14297 10333 14331
rect 10333 14297 10367 14331
rect 10367 14297 10376 14331
rect 10324 14288 10376 14297
rect 13084 14288 13136 14340
rect 30104 14399 30156 14408
rect 30104 14365 30113 14399
rect 30113 14365 30147 14399
rect 30147 14365 30156 14399
rect 30104 14356 30156 14365
rect 9680 14220 9732 14272
rect 10600 14220 10652 14272
rect 12440 14220 12492 14272
rect 16212 14220 16264 14272
rect 18328 14220 18380 14272
rect 20720 14220 20772 14272
rect 10880 14118 10932 14170
rect 10944 14118 10996 14170
rect 11008 14118 11060 14170
rect 11072 14118 11124 14170
rect 11136 14118 11188 14170
rect 20811 14118 20863 14170
rect 20875 14118 20927 14170
rect 20939 14118 20991 14170
rect 21003 14118 21055 14170
rect 21067 14118 21119 14170
rect 1676 14016 1728 14068
rect 1768 14016 1820 14068
rect 3792 13948 3844 14000
rect 1492 13880 1544 13932
rect 3056 13880 3108 13932
rect 5908 14016 5960 14068
rect 11428 14016 11480 14068
rect 11520 14016 11572 14068
rect 6460 13948 6512 14000
rect 7564 13948 7616 14000
rect 17592 14016 17644 14068
rect 18420 14016 18472 14068
rect 29828 14016 29880 14068
rect 12808 13991 12860 14000
rect 12808 13957 12817 13991
rect 12817 13957 12851 13991
rect 12851 13957 12860 13991
rect 12808 13948 12860 13957
rect 13820 13948 13872 14000
rect 14556 13948 14608 14000
rect 15476 13948 15528 14000
rect 4988 13923 5040 13932
rect 4988 13889 4997 13923
rect 4997 13889 5031 13923
rect 5031 13889 5040 13923
rect 4988 13880 5040 13889
rect 3424 13812 3476 13864
rect 6644 13923 6696 13932
rect 6644 13889 6653 13923
rect 6653 13889 6687 13923
rect 6687 13889 6696 13923
rect 6644 13880 6696 13889
rect 6828 13880 6880 13932
rect 8760 13880 8812 13932
rect 9680 13880 9732 13932
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 10508 13880 10560 13932
rect 6460 13812 6512 13864
rect 7012 13812 7064 13864
rect 7564 13812 7616 13864
rect 7840 13812 7892 13864
rect 3976 13676 4028 13728
rect 7380 13676 7432 13728
rect 8392 13812 8444 13864
rect 8852 13812 8904 13864
rect 9588 13812 9640 13864
rect 9956 13812 10008 13864
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 13084 13880 13136 13932
rect 13728 13880 13780 13932
rect 15108 13923 15160 13932
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 16856 13923 16908 13932
rect 15108 13880 15160 13889
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 17040 13880 17092 13932
rect 18328 13880 18380 13932
rect 18512 13880 18564 13932
rect 21180 13948 21232 14000
rect 19800 13880 19852 13932
rect 20352 13880 20404 13932
rect 13360 13812 13412 13864
rect 16580 13812 16632 13864
rect 17868 13812 17920 13864
rect 20720 13880 20772 13932
rect 29920 13923 29972 13932
rect 29920 13889 29929 13923
rect 29929 13889 29963 13923
rect 29963 13889 29972 13923
rect 29920 13880 29972 13889
rect 30104 13923 30156 13932
rect 30104 13889 30113 13923
rect 30113 13889 30147 13923
rect 30147 13889 30156 13923
rect 30104 13880 30156 13889
rect 29276 13812 29328 13864
rect 8024 13744 8076 13796
rect 8208 13744 8260 13796
rect 15752 13744 15804 13796
rect 11244 13676 11296 13728
rect 12808 13676 12860 13728
rect 16672 13719 16724 13728
rect 16672 13685 16681 13719
rect 16681 13685 16715 13719
rect 16715 13685 16724 13719
rect 16672 13676 16724 13685
rect 18420 13744 18472 13796
rect 18604 13744 18656 13796
rect 17224 13676 17276 13728
rect 17776 13676 17828 13728
rect 18512 13719 18564 13728
rect 18512 13685 18521 13719
rect 18521 13685 18555 13719
rect 18555 13685 18564 13719
rect 18512 13676 18564 13685
rect 5915 13574 5967 13626
rect 5979 13574 6031 13626
rect 6043 13574 6095 13626
rect 6107 13574 6159 13626
rect 6171 13574 6223 13626
rect 15846 13574 15898 13626
rect 15910 13574 15962 13626
rect 15974 13574 16026 13626
rect 16038 13574 16090 13626
rect 16102 13574 16154 13626
rect 25776 13574 25828 13626
rect 25840 13574 25892 13626
rect 25904 13574 25956 13626
rect 25968 13574 26020 13626
rect 26032 13574 26084 13626
rect 5356 13472 5408 13524
rect 9312 13472 9364 13524
rect 9588 13472 9640 13524
rect 10048 13472 10100 13524
rect 12072 13472 12124 13524
rect 16304 13472 16356 13524
rect 17500 13472 17552 13524
rect 18512 13472 18564 13524
rect 19708 13515 19760 13524
rect 19708 13481 19717 13515
rect 19717 13481 19751 13515
rect 19751 13481 19760 13515
rect 19708 13472 19760 13481
rect 20260 13472 20312 13524
rect 14464 13447 14516 13456
rect 14464 13413 14473 13447
rect 14473 13413 14507 13447
rect 14507 13413 14516 13447
rect 14464 13404 14516 13413
rect 15752 13447 15804 13456
rect 15752 13413 15761 13447
rect 15761 13413 15795 13447
rect 15795 13413 15804 13447
rect 15752 13404 15804 13413
rect 3240 13336 3292 13388
rect 3976 13336 4028 13388
rect 6644 13336 6696 13388
rect 7380 13336 7432 13388
rect 9864 13336 9916 13388
rect 13820 13336 13872 13388
rect 19616 13404 19668 13456
rect 16028 13336 16080 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 3516 13268 3568 13320
rect 4252 13268 4304 13320
rect 5908 13311 5960 13320
rect 5172 13243 5224 13252
rect 5172 13209 5181 13243
rect 5181 13209 5215 13243
rect 5215 13209 5224 13243
rect 5172 13200 5224 13209
rect 5908 13277 5917 13311
rect 5917 13277 5951 13311
rect 5951 13277 5960 13311
rect 5908 13268 5960 13277
rect 6092 13311 6144 13320
rect 6092 13277 6101 13311
rect 6101 13277 6135 13311
rect 6135 13277 6144 13311
rect 6276 13311 6328 13320
rect 6092 13268 6144 13277
rect 6276 13277 6285 13311
rect 6285 13277 6319 13311
rect 6319 13277 6328 13311
rect 6276 13268 6328 13277
rect 8208 13268 8260 13320
rect 8484 13268 8536 13320
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 10600 13311 10652 13320
rect 10600 13277 10634 13311
rect 10634 13277 10652 13311
rect 10600 13268 10652 13277
rect 11336 13268 11388 13320
rect 15016 13268 15068 13320
rect 16672 13268 16724 13320
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 17500 13311 17552 13320
rect 6368 13200 6420 13252
rect 7196 13200 7248 13252
rect 9496 13243 9548 13252
rect 9496 13209 9505 13243
rect 9505 13209 9539 13243
rect 9539 13209 9548 13243
rect 9496 13200 9548 13209
rect 9588 13200 9640 13252
rect 12808 13243 12860 13252
rect 2688 13132 2740 13184
rect 3792 13132 3844 13184
rect 7012 13132 7064 13184
rect 8392 13132 8444 13184
rect 9864 13132 9916 13184
rect 10048 13132 10100 13184
rect 12808 13209 12817 13243
rect 12817 13209 12851 13243
rect 12851 13209 12860 13243
rect 12808 13200 12860 13209
rect 14280 13243 14332 13252
rect 14280 13209 14289 13243
rect 14289 13209 14323 13243
rect 14323 13209 14332 13243
rect 14280 13200 14332 13209
rect 14648 13200 14700 13252
rect 15108 13243 15160 13252
rect 15108 13209 15117 13243
rect 15117 13209 15151 13243
rect 15151 13209 15160 13243
rect 15108 13200 15160 13209
rect 12624 13132 12676 13184
rect 15476 13132 15528 13184
rect 16580 13200 16632 13252
rect 17040 13200 17092 13252
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 19432 13268 19484 13320
rect 19892 13268 19944 13320
rect 20352 13311 20404 13320
rect 20352 13277 20361 13311
rect 20361 13277 20395 13311
rect 20395 13277 20404 13311
rect 20352 13268 20404 13277
rect 16856 13132 16908 13184
rect 17316 13132 17368 13184
rect 18972 13200 19024 13252
rect 20720 13311 20772 13320
rect 20720 13277 20729 13311
rect 20729 13277 20763 13311
rect 20763 13277 20772 13311
rect 20720 13268 20772 13277
rect 30104 13268 30156 13320
rect 29920 13200 29972 13252
rect 18604 13175 18656 13184
rect 18604 13141 18613 13175
rect 18613 13141 18647 13175
rect 18647 13141 18656 13175
rect 18604 13132 18656 13141
rect 30012 13175 30064 13184
rect 30012 13141 30021 13175
rect 30021 13141 30055 13175
rect 30055 13141 30064 13175
rect 30012 13132 30064 13141
rect 10880 13030 10932 13082
rect 10944 13030 10996 13082
rect 11008 13030 11060 13082
rect 11072 13030 11124 13082
rect 11136 13030 11188 13082
rect 20811 13030 20863 13082
rect 20875 13030 20927 13082
rect 20939 13030 20991 13082
rect 21003 13030 21055 13082
rect 21067 13030 21119 13082
rect 5172 12928 5224 12980
rect 10140 12928 10192 12980
rect 8300 12860 8352 12912
rect 16028 12928 16080 12980
rect 2780 12835 2832 12844
rect 2780 12801 2789 12835
rect 2789 12801 2823 12835
rect 2823 12801 2832 12835
rect 2780 12792 2832 12801
rect 3148 12792 3200 12844
rect 3700 12792 3752 12844
rect 5816 12792 5868 12844
rect 1400 12656 1452 12708
rect 2780 12588 2832 12640
rect 5632 12724 5684 12776
rect 6644 12835 6696 12844
rect 6644 12801 6653 12835
rect 6653 12801 6687 12835
rect 6687 12801 6696 12835
rect 6920 12835 6972 12844
rect 6644 12792 6696 12801
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 10508 12860 10560 12912
rect 12164 12860 12216 12912
rect 15568 12860 15620 12912
rect 6092 12656 6144 12708
rect 8024 12724 8076 12776
rect 8760 12767 8812 12776
rect 7564 12656 7616 12708
rect 8760 12733 8769 12767
rect 8769 12733 8803 12767
rect 8803 12733 8812 12767
rect 8760 12724 8812 12733
rect 9404 12724 9456 12776
rect 9588 12792 9640 12844
rect 9864 12792 9916 12844
rect 11796 12792 11848 12844
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 12992 12792 13044 12844
rect 14280 12792 14332 12844
rect 15016 12835 15068 12844
rect 15016 12801 15025 12835
rect 15025 12801 15059 12835
rect 15059 12801 15068 12835
rect 15016 12792 15068 12801
rect 11980 12724 12032 12776
rect 11336 12656 11388 12708
rect 11888 12656 11940 12708
rect 16212 12792 16264 12844
rect 18236 12860 18288 12912
rect 17316 12835 17368 12844
rect 16488 12724 16540 12776
rect 16672 12767 16724 12776
rect 16672 12733 16681 12767
rect 16681 12733 16715 12767
rect 16715 12733 16724 12767
rect 16672 12724 16724 12733
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 18420 12928 18472 12980
rect 18696 12928 18748 12980
rect 19340 12860 19392 12912
rect 19984 12860 20036 12912
rect 19616 12792 19668 12844
rect 30196 12928 30248 12980
rect 21640 12792 21692 12844
rect 29920 12835 29972 12844
rect 29920 12801 29929 12835
rect 29929 12801 29963 12835
rect 29963 12801 29972 12835
rect 29920 12792 29972 12801
rect 30104 12835 30156 12844
rect 30104 12801 30113 12835
rect 30113 12801 30147 12835
rect 30147 12801 30156 12835
rect 30104 12792 30156 12801
rect 17040 12656 17092 12708
rect 3792 12588 3844 12640
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 9772 12588 9824 12640
rect 10784 12588 10836 12640
rect 12624 12631 12676 12640
rect 12624 12597 12633 12631
rect 12633 12597 12667 12631
rect 12667 12597 12676 12631
rect 12624 12588 12676 12597
rect 15476 12588 15528 12640
rect 16488 12588 16540 12640
rect 18052 12588 18104 12640
rect 5915 12486 5967 12538
rect 5979 12486 6031 12538
rect 6043 12486 6095 12538
rect 6107 12486 6159 12538
rect 6171 12486 6223 12538
rect 15846 12486 15898 12538
rect 15910 12486 15962 12538
rect 15974 12486 16026 12538
rect 16038 12486 16090 12538
rect 16102 12486 16154 12538
rect 25776 12486 25828 12538
rect 25840 12486 25892 12538
rect 25904 12486 25956 12538
rect 25968 12486 26020 12538
rect 26032 12486 26084 12538
rect 6276 12384 6328 12436
rect 7104 12384 7156 12436
rect 3056 12316 3108 12368
rect 3792 12291 3844 12300
rect 3792 12257 3801 12291
rect 3801 12257 3835 12291
rect 3835 12257 3844 12291
rect 3792 12248 3844 12257
rect 1216 12180 1268 12232
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 2872 12112 2924 12164
rect 2964 12044 3016 12096
rect 5356 12180 5408 12232
rect 7196 12248 7248 12300
rect 7564 12248 7616 12300
rect 8208 12248 8260 12300
rect 8944 12248 8996 12300
rect 14280 12384 14332 12436
rect 12164 12316 12216 12368
rect 16672 12384 16724 12436
rect 16948 12384 17000 12436
rect 18328 12316 18380 12368
rect 15660 12248 15712 12300
rect 19340 12248 19392 12300
rect 4896 12112 4948 12164
rect 5632 12044 5684 12096
rect 7748 12180 7800 12232
rect 10232 12180 10284 12232
rect 12256 12180 12308 12232
rect 12992 12180 13044 12232
rect 16304 12180 16356 12232
rect 16396 12180 16448 12232
rect 18604 12180 18656 12232
rect 19064 12180 19116 12232
rect 19708 12180 19760 12232
rect 20352 12180 20404 12232
rect 8392 12044 8444 12096
rect 9036 12044 9088 12096
rect 9588 12112 9640 12164
rect 11244 12155 11296 12164
rect 11244 12121 11278 12155
rect 11278 12121 11296 12155
rect 11244 12112 11296 12121
rect 14188 12112 14240 12164
rect 29920 12248 29972 12300
rect 20628 12180 20680 12232
rect 20812 12223 20864 12232
rect 20812 12189 20821 12223
rect 20821 12189 20855 12223
rect 20855 12189 20864 12223
rect 21456 12223 21508 12232
rect 20812 12180 20864 12189
rect 21456 12189 21465 12223
rect 21465 12189 21499 12223
rect 21499 12189 21508 12223
rect 21456 12180 21508 12189
rect 21640 12155 21692 12164
rect 11336 12044 11388 12096
rect 12348 12087 12400 12096
rect 12348 12053 12357 12087
rect 12357 12053 12391 12087
rect 12391 12053 12400 12087
rect 12348 12044 12400 12053
rect 12900 12044 12952 12096
rect 21640 12121 21649 12155
rect 21649 12121 21683 12155
rect 21683 12121 21692 12155
rect 21640 12112 21692 12121
rect 15660 12044 15712 12096
rect 18052 12087 18104 12096
rect 18052 12053 18061 12087
rect 18061 12053 18095 12087
rect 18095 12053 18104 12087
rect 18052 12044 18104 12053
rect 19892 12044 19944 12096
rect 22192 12044 22244 12096
rect 10880 11942 10932 11994
rect 10944 11942 10996 11994
rect 11008 11942 11060 11994
rect 11072 11942 11124 11994
rect 11136 11942 11188 11994
rect 20811 11942 20863 11994
rect 20875 11942 20927 11994
rect 20939 11942 20991 11994
rect 21003 11942 21055 11994
rect 21067 11942 21119 11994
rect 3700 11840 3752 11892
rect 4804 11883 4856 11892
rect 4804 11849 4813 11883
rect 4813 11849 4847 11883
rect 4847 11849 4856 11883
rect 4804 11840 4856 11849
rect 6920 11840 6972 11892
rect 8852 11883 8904 11892
rect 8852 11849 8861 11883
rect 8861 11849 8895 11883
rect 8895 11849 8904 11883
rect 8852 11840 8904 11849
rect 2504 11772 2556 11824
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 3792 11772 3844 11824
rect 4620 11772 4672 11824
rect 11244 11840 11296 11892
rect 11336 11840 11388 11892
rect 12900 11840 12952 11892
rect 12992 11840 13044 11892
rect 17408 11840 17460 11892
rect 18052 11840 18104 11892
rect 20628 11883 20680 11892
rect 20628 11849 20637 11883
rect 20637 11849 20671 11883
rect 20671 11849 20680 11883
rect 20628 11840 20680 11849
rect 2780 11747 2832 11756
rect 2780 11713 2789 11747
rect 2789 11713 2823 11747
rect 2823 11713 2832 11747
rect 2780 11704 2832 11713
rect 3056 11704 3108 11756
rect 4988 11704 5040 11756
rect 5356 11704 5408 11756
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 9956 11772 10008 11824
rect 2872 11679 2924 11688
rect 2872 11645 2881 11679
rect 2881 11645 2915 11679
rect 2915 11645 2924 11679
rect 2872 11636 2924 11645
rect 4068 11636 4120 11688
rect 2228 11568 2280 11620
rect 7564 11679 7616 11688
rect 7564 11645 7573 11679
rect 7573 11645 7607 11679
rect 7607 11645 7616 11679
rect 7564 11636 7616 11645
rect 8484 11704 8536 11756
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 8852 11704 8904 11756
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 10416 11747 10468 11756
rect 10416 11713 10425 11747
rect 10425 11713 10459 11747
rect 10459 11713 10468 11747
rect 10416 11704 10468 11713
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 12348 11772 12400 11824
rect 12624 11772 12676 11824
rect 14464 11772 14516 11824
rect 19064 11815 19116 11824
rect 19064 11781 19073 11815
rect 19073 11781 19107 11815
rect 19107 11781 19116 11815
rect 19064 11772 19116 11781
rect 19984 11772 20036 11824
rect 10508 11704 10560 11713
rect 12256 11747 12308 11756
rect 12256 11713 12265 11747
rect 12265 11713 12299 11747
rect 12299 11713 12308 11747
rect 12256 11704 12308 11713
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 14372 11747 14424 11756
rect 14372 11713 14406 11747
rect 14406 11713 14424 11747
rect 14372 11704 14424 11713
rect 15292 11704 15344 11756
rect 11888 11636 11940 11688
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 2964 11500 3016 11552
rect 3976 11500 4028 11552
rect 7288 11500 7340 11552
rect 9037 11500 9089 11552
rect 9312 11500 9364 11552
rect 9864 11568 9916 11620
rect 11244 11568 11296 11620
rect 16948 11704 17000 11756
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 19892 11747 19944 11756
rect 19892 11713 19901 11747
rect 19901 11713 19935 11747
rect 19935 11713 19944 11747
rect 19892 11704 19944 11713
rect 20352 11704 20404 11756
rect 20444 11747 20496 11756
rect 20444 11713 20453 11747
rect 20453 11713 20487 11747
rect 20487 11713 20496 11747
rect 22192 11747 22244 11756
rect 20444 11704 20496 11713
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 18420 11679 18472 11688
rect 12440 11500 12492 11552
rect 14832 11500 14884 11552
rect 18420 11645 18429 11679
rect 18429 11645 18463 11679
rect 18463 11645 18472 11679
rect 18420 11636 18472 11645
rect 20168 11679 20220 11688
rect 20168 11645 20177 11679
rect 20177 11645 20211 11679
rect 20211 11645 20220 11679
rect 20168 11636 20220 11645
rect 20260 11679 20312 11688
rect 20260 11645 20269 11679
rect 20269 11645 20303 11679
rect 20303 11645 20312 11679
rect 20260 11636 20312 11645
rect 29828 11636 29880 11688
rect 16856 11568 16908 11620
rect 17316 11500 17368 11552
rect 20628 11500 20680 11552
rect 5915 11398 5967 11450
rect 5979 11398 6031 11450
rect 6043 11398 6095 11450
rect 6107 11398 6159 11450
rect 6171 11398 6223 11450
rect 15846 11398 15898 11450
rect 15910 11398 15962 11450
rect 15974 11398 16026 11450
rect 16038 11398 16090 11450
rect 16102 11398 16154 11450
rect 25776 11398 25828 11450
rect 25840 11398 25892 11450
rect 25904 11398 25956 11450
rect 25968 11398 26020 11450
rect 26032 11398 26084 11450
rect 8484 11296 8536 11348
rect 17868 11339 17920 11348
rect 2964 11228 3016 11280
rect 2780 11092 2832 11144
rect 2136 11024 2188 11076
rect 1768 10956 1820 11008
rect 2044 10956 2096 11008
rect 3792 11135 3844 11144
rect 3792 11101 3801 11135
rect 3801 11101 3835 11135
rect 3835 11101 3844 11135
rect 3792 11092 3844 11101
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 4068 11135 4120 11144
rect 4068 11101 4077 11135
rect 4077 11101 4111 11135
rect 4111 11101 4120 11135
rect 4344 11135 4396 11144
rect 4068 11092 4120 11101
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 8024 11228 8076 11280
rect 5448 11203 5500 11212
rect 5448 11169 5457 11203
rect 5457 11169 5491 11203
rect 5491 11169 5500 11203
rect 5448 11160 5500 11169
rect 7012 11203 7064 11212
rect 7012 11169 7021 11203
rect 7021 11169 7055 11203
rect 7055 11169 7064 11203
rect 7012 11160 7064 11169
rect 9588 11160 9640 11212
rect 11796 11160 11848 11212
rect 12992 11228 13044 11280
rect 7288 11135 7340 11144
rect 7288 11101 7322 11135
rect 7322 11101 7340 11135
rect 7288 11092 7340 11101
rect 8852 11092 8904 11144
rect 9312 11092 9364 11144
rect 9772 11092 9824 11144
rect 10232 11092 10284 11144
rect 5172 11024 5224 11076
rect 5356 11024 5408 11076
rect 6276 11024 6328 11076
rect 7196 11024 7248 11076
rect 12164 11092 12216 11144
rect 13728 11160 13780 11212
rect 14096 11203 14148 11212
rect 14096 11169 14105 11203
rect 14105 11169 14139 11203
rect 14139 11169 14148 11203
rect 14096 11160 14148 11169
rect 12900 11092 12952 11144
rect 13268 11092 13320 11144
rect 16948 11228 17000 11280
rect 17868 11305 17877 11339
rect 17877 11305 17911 11339
rect 17911 11305 17920 11339
rect 17868 11296 17920 11305
rect 18420 11339 18472 11348
rect 18420 11305 18429 11339
rect 18429 11305 18463 11339
rect 18463 11305 18472 11339
rect 18420 11296 18472 11305
rect 20076 11296 20128 11348
rect 20352 11296 20404 11348
rect 15660 11160 15712 11212
rect 16304 11203 16356 11212
rect 15752 11092 15804 11144
rect 16304 11169 16313 11203
rect 16313 11169 16347 11203
rect 16347 11169 16356 11203
rect 16304 11160 16356 11169
rect 17040 11160 17092 11212
rect 18328 11160 18380 11212
rect 16488 11135 16540 11144
rect 10692 11024 10744 11076
rect 14556 11024 14608 11076
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 16764 11092 16816 11144
rect 17132 11135 17184 11144
rect 17132 11101 17141 11135
rect 17141 11101 17175 11135
rect 17175 11101 17184 11135
rect 17132 11092 17184 11101
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 16948 11024 17000 11076
rect 18052 11092 18104 11144
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 20168 11160 20220 11212
rect 19524 11092 19576 11144
rect 20260 11135 20312 11144
rect 20260 11101 20269 11135
rect 20269 11101 20303 11135
rect 20303 11101 20312 11135
rect 20260 11092 20312 11101
rect 20628 11135 20680 11144
rect 20628 11101 20637 11135
rect 20637 11101 20671 11135
rect 20671 11101 20680 11135
rect 20628 11092 20680 11101
rect 21364 11092 21416 11144
rect 29828 11135 29880 11144
rect 29828 11101 29837 11135
rect 29837 11101 29871 11135
rect 29871 11101 29880 11135
rect 29828 11092 29880 11101
rect 20720 11024 20772 11076
rect 4528 10999 4580 11008
rect 4528 10965 4537 10999
rect 4537 10965 4571 10999
rect 4571 10965 4580 10999
rect 4528 10956 4580 10965
rect 11520 10999 11572 11008
rect 11520 10965 11529 10999
rect 11529 10965 11563 10999
rect 11563 10965 11572 10999
rect 11520 10956 11572 10965
rect 11612 10956 11664 11008
rect 13820 10956 13872 11008
rect 15016 10956 15068 11008
rect 30012 10999 30064 11008
rect 30012 10965 30021 10999
rect 30021 10965 30055 10999
rect 30055 10965 30064 10999
rect 30012 10956 30064 10965
rect 10880 10854 10932 10906
rect 10944 10854 10996 10906
rect 11008 10854 11060 10906
rect 11072 10854 11124 10906
rect 11136 10854 11188 10906
rect 20811 10854 20863 10906
rect 20875 10854 20927 10906
rect 20939 10854 20991 10906
rect 21003 10854 21055 10906
rect 21067 10854 21119 10906
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 2964 10752 3016 10804
rect 2136 10727 2188 10736
rect 2136 10693 2145 10727
rect 2145 10693 2179 10727
rect 2179 10693 2188 10727
rect 2136 10684 2188 10693
rect 4528 10684 4580 10736
rect 5172 10684 5224 10736
rect 6552 10752 6604 10804
rect 6920 10752 6972 10804
rect 10692 10795 10744 10804
rect 10692 10761 10701 10795
rect 10701 10761 10735 10795
rect 10735 10761 10744 10795
rect 10692 10752 10744 10761
rect 10784 10752 10836 10804
rect 12716 10752 12768 10804
rect 14372 10752 14424 10804
rect 16580 10752 16632 10804
rect 18052 10795 18104 10804
rect 18052 10761 18061 10795
rect 18061 10761 18095 10795
rect 18095 10761 18104 10795
rect 18052 10752 18104 10761
rect 20536 10795 20588 10804
rect 20536 10761 20545 10795
rect 20545 10761 20579 10795
rect 20579 10761 20588 10795
rect 20536 10752 20588 10761
rect 20720 10752 20772 10804
rect 1492 10548 1544 10600
rect 1768 10591 1820 10600
rect 1768 10557 1777 10591
rect 1777 10557 1811 10591
rect 1811 10557 1820 10591
rect 1768 10548 1820 10557
rect 2780 10659 2832 10668
rect 2780 10625 2789 10659
rect 2789 10625 2823 10659
rect 2823 10625 2832 10659
rect 2780 10616 2832 10625
rect 3884 10616 3936 10668
rect 5448 10616 5500 10668
rect 2688 10548 2740 10600
rect 4896 10548 4948 10600
rect 4344 10480 4396 10532
rect 11612 10684 11664 10736
rect 12348 10684 12400 10736
rect 6276 10616 6328 10668
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 8116 10616 8168 10668
rect 9864 10616 9916 10668
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 10140 10659 10192 10668
rect 9956 10616 10008 10625
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 10140 10616 10192 10625
rect 11428 10616 11480 10668
rect 11704 10659 11756 10668
rect 5724 10480 5776 10532
rect 8300 10480 8352 10532
rect 10508 10480 10560 10532
rect 3516 10412 3568 10464
rect 6552 10412 6604 10464
rect 7564 10412 7616 10464
rect 10968 10480 11020 10532
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 11980 10616 12032 10668
rect 12624 10616 12676 10668
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 13452 10616 13504 10668
rect 14832 10616 14884 10668
rect 15016 10659 15068 10668
rect 15016 10625 15025 10659
rect 15025 10625 15059 10659
rect 15059 10625 15068 10659
rect 15016 10616 15068 10625
rect 15660 10659 15712 10668
rect 15660 10625 15669 10659
rect 15669 10625 15703 10659
rect 15703 10625 15712 10659
rect 15660 10616 15712 10625
rect 18972 10684 19024 10736
rect 11888 10591 11940 10600
rect 11888 10557 11897 10591
rect 11897 10557 11931 10591
rect 11931 10557 11940 10591
rect 11888 10548 11940 10557
rect 13268 10591 13320 10600
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 13268 10548 13320 10557
rect 13728 10548 13780 10600
rect 15752 10591 15804 10600
rect 15752 10557 15761 10591
rect 15761 10557 15795 10591
rect 15795 10557 15804 10591
rect 15752 10548 15804 10557
rect 12256 10455 12308 10464
rect 12256 10421 12265 10455
rect 12265 10421 12299 10455
rect 12299 10421 12308 10455
rect 12256 10412 12308 10421
rect 16580 10616 16632 10668
rect 16856 10659 16908 10668
rect 16856 10625 16865 10659
rect 16865 10625 16899 10659
rect 16899 10625 16908 10659
rect 16856 10616 16908 10625
rect 16948 10659 17000 10668
rect 16948 10625 16957 10659
rect 16957 10625 16991 10659
rect 16991 10625 17000 10659
rect 17224 10659 17276 10668
rect 16948 10616 17000 10625
rect 17224 10625 17233 10659
rect 17233 10625 17267 10659
rect 17267 10625 17276 10659
rect 17224 10616 17276 10625
rect 17960 10659 18012 10668
rect 17960 10625 17969 10659
rect 17969 10625 18003 10659
rect 18003 10625 18012 10659
rect 17960 10616 18012 10625
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 19984 10659 20036 10668
rect 17040 10591 17092 10600
rect 17040 10557 17049 10591
rect 17049 10557 17083 10591
rect 17083 10557 17092 10591
rect 17040 10548 17092 10557
rect 19984 10625 19993 10659
rect 19993 10625 20027 10659
rect 20027 10625 20036 10659
rect 19984 10616 20036 10625
rect 20352 10659 20404 10668
rect 20352 10625 20361 10659
rect 20361 10625 20395 10659
rect 20395 10625 20404 10659
rect 20352 10616 20404 10625
rect 21456 10616 21508 10668
rect 20076 10591 20128 10600
rect 20076 10557 20085 10591
rect 20085 10557 20119 10591
rect 20119 10557 20128 10591
rect 20076 10548 20128 10557
rect 20260 10548 20312 10600
rect 18604 10412 18656 10464
rect 19064 10455 19116 10464
rect 19064 10421 19073 10455
rect 19073 10421 19107 10455
rect 19107 10421 19116 10455
rect 19064 10412 19116 10421
rect 5915 10310 5967 10362
rect 5979 10310 6031 10362
rect 6043 10310 6095 10362
rect 6107 10310 6159 10362
rect 6171 10310 6223 10362
rect 15846 10310 15898 10362
rect 15910 10310 15962 10362
rect 15974 10310 16026 10362
rect 16038 10310 16090 10362
rect 16102 10310 16154 10362
rect 25776 10310 25828 10362
rect 25840 10310 25892 10362
rect 25904 10310 25956 10362
rect 25968 10310 26020 10362
rect 26032 10310 26084 10362
rect 8576 10208 8628 10260
rect 10232 10208 10284 10260
rect 11520 10208 11572 10260
rect 15752 10208 15804 10260
rect 17684 10208 17736 10260
rect 19984 10208 20036 10260
rect 1492 10140 1544 10192
rect 2596 10140 2648 10192
rect 6276 10140 6328 10192
rect 8760 10140 8812 10192
rect 9956 10140 10008 10192
rect 10968 10140 11020 10192
rect 12624 10183 12676 10192
rect 12624 10149 12633 10183
rect 12633 10149 12667 10183
rect 12667 10149 12676 10183
rect 28724 10208 28776 10260
rect 12624 10140 12676 10149
rect 2044 10004 2096 10056
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 5080 10004 5132 10056
rect 6644 10072 6696 10124
rect 13728 10072 13780 10124
rect 6000 10004 6052 10056
rect 3516 9936 3568 9988
rect 4988 9936 5040 9988
rect 5356 9936 5408 9988
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 7196 10004 7248 10056
rect 10784 10004 10836 10056
rect 12440 10004 12492 10056
rect 12992 10004 13044 10056
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 14556 10004 14608 10056
rect 16396 10072 16448 10124
rect 16580 10115 16632 10124
rect 16580 10081 16589 10115
rect 16589 10081 16623 10115
rect 16623 10081 16632 10115
rect 16580 10072 16632 10081
rect 17132 10072 17184 10124
rect 15752 10004 15804 10056
rect 16672 10047 16724 10056
rect 16672 10013 16717 10047
rect 16717 10013 16724 10047
rect 16672 10004 16724 10013
rect 6552 9936 6604 9988
rect 7012 9936 7064 9988
rect 1952 9868 2004 9920
rect 2412 9911 2464 9920
rect 2412 9877 2421 9911
rect 2421 9877 2455 9911
rect 2455 9877 2464 9911
rect 2412 9868 2464 9877
rect 5264 9911 5316 9920
rect 5264 9877 5273 9911
rect 5273 9877 5307 9911
rect 5307 9877 5316 9911
rect 5264 9868 5316 9877
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 6276 9868 6328 9920
rect 9496 9936 9548 9988
rect 10232 9979 10284 9988
rect 10232 9945 10241 9979
rect 10241 9945 10275 9979
rect 10275 9945 10284 9979
rect 10232 9936 10284 9945
rect 12256 9936 12308 9988
rect 9956 9868 10008 9920
rect 10692 9868 10744 9920
rect 14188 9936 14240 9988
rect 15568 9979 15620 9988
rect 15568 9945 15577 9979
rect 15577 9945 15611 9979
rect 15611 9945 15620 9979
rect 15568 9936 15620 9945
rect 15660 9936 15712 9988
rect 17408 9979 17460 9988
rect 12624 9868 12676 9920
rect 14648 9868 14700 9920
rect 14832 9911 14884 9920
rect 14832 9877 14841 9911
rect 14841 9877 14875 9911
rect 14875 9877 14884 9911
rect 14832 9868 14884 9877
rect 17408 9945 17417 9979
rect 17417 9945 17451 9979
rect 17451 9945 17460 9979
rect 17408 9936 17460 9945
rect 17684 10047 17736 10056
rect 17684 10013 17693 10047
rect 17693 10013 17727 10047
rect 17727 10013 17736 10047
rect 17684 10004 17736 10013
rect 18144 10004 18196 10056
rect 18696 10072 18748 10124
rect 18880 10004 18932 10056
rect 19248 10004 19300 10056
rect 19892 10004 19944 10056
rect 21272 10047 21324 10056
rect 21272 10013 21281 10047
rect 21281 10013 21315 10047
rect 21315 10013 21324 10047
rect 21272 10004 21324 10013
rect 20720 9936 20772 9988
rect 21180 9936 21232 9988
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 10880 9766 10932 9818
rect 10944 9766 10996 9818
rect 11008 9766 11060 9818
rect 11072 9766 11124 9818
rect 11136 9766 11188 9818
rect 20811 9766 20863 9818
rect 20875 9766 20927 9818
rect 20939 9766 20991 9818
rect 21003 9766 21055 9818
rect 21067 9766 21119 9818
rect 3516 9707 3568 9716
rect 3516 9673 3525 9707
rect 3525 9673 3559 9707
rect 3559 9673 3568 9707
rect 3516 9664 3568 9673
rect 13176 9664 13228 9716
rect 13268 9664 13320 9716
rect 2412 9639 2464 9648
rect 2412 9605 2446 9639
rect 2446 9605 2464 9639
rect 2412 9596 2464 9605
rect 3056 9596 3108 9648
rect 7104 9596 7156 9648
rect 8300 9596 8352 9648
rect 9864 9596 9916 9648
rect 10692 9639 10744 9648
rect 10692 9605 10701 9639
rect 10701 9605 10735 9639
rect 10735 9605 10744 9639
rect 10692 9596 10744 9605
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 4068 9571 4120 9580
rect 4068 9537 4077 9571
rect 4077 9537 4111 9571
rect 4111 9537 4120 9571
rect 4068 9528 4120 9537
rect 4528 9528 4580 9580
rect 5540 9528 5592 9580
rect 1676 9460 1728 9512
rect 4436 9503 4488 9512
rect 4436 9469 4445 9503
rect 4445 9469 4479 9503
rect 4479 9469 4488 9503
rect 4436 9460 4488 9469
rect 5356 9460 5408 9512
rect 6552 9528 6604 9580
rect 7012 9571 7064 9580
rect 7012 9537 7021 9571
rect 7021 9537 7055 9571
rect 7055 9537 7064 9571
rect 7012 9528 7064 9537
rect 8116 9528 8168 9580
rect 8208 9503 8260 9512
rect 4712 9392 4764 9444
rect 1492 9324 1544 9376
rect 4804 9367 4856 9376
rect 4804 9333 4813 9367
rect 4813 9333 4847 9367
rect 4847 9333 4856 9367
rect 4804 9324 4856 9333
rect 5080 9392 5132 9444
rect 6736 9392 6788 9444
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 8484 9503 8536 9512
rect 8484 9469 8493 9503
rect 8493 9469 8527 9503
rect 8527 9469 8536 9503
rect 8484 9460 8536 9469
rect 10232 9528 10284 9580
rect 13728 9596 13780 9648
rect 17224 9664 17276 9716
rect 17408 9664 17460 9716
rect 19064 9664 19116 9716
rect 19248 9707 19300 9716
rect 19248 9673 19257 9707
rect 19257 9673 19291 9707
rect 19291 9673 19300 9707
rect 19248 9664 19300 9673
rect 20352 9664 20404 9716
rect 13636 9528 13688 9580
rect 12992 9460 13044 9512
rect 13084 9392 13136 9444
rect 15108 9571 15160 9580
rect 15108 9537 15117 9571
rect 15117 9537 15151 9571
rect 15151 9537 15160 9571
rect 15292 9571 15344 9580
rect 15108 9528 15160 9537
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 16488 9596 16540 9648
rect 18144 9639 18196 9648
rect 18144 9605 18178 9639
rect 18178 9605 18196 9639
rect 18144 9596 18196 9605
rect 15660 9528 15712 9580
rect 17224 9571 17276 9580
rect 17224 9537 17233 9571
rect 17233 9537 17267 9571
rect 17267 9537 17276 9571
rect 17224 9528 17276 9537
rect 15752 9460 15804 9512
rect 17868 9503 17920 9512
rect 17868 9469 17877 9503
rect 17877 9469 17911 9503
rect 17911 9469 17920 9503
rect 17868 9460 17920 9469
rect 7380 9324 7432 9376
rect 7564 9367 7616 9376
rect 7564 9333 7573 9367
rect 7573 9333 7607 9367
rect 7607 9333 7616 9367
rect 7564 9324 7616 9333
rect 9588 9367 9640 9376
rect 9588 9333 9597 9367
rect 9597 9333 9631 9367
rect 9631 9333 9640 9367
rect 9588 9324 9640 9333
rect 9956 9324 10008 9376
rect 13268 9324 13320 9376
rect 16304 9324 16356 9376
rect 19432 9324 19484 9376
rect 20260 9324 20312 9376
rect 21272 9324 21324 9376
rect 21548 9324 21600 9376
rect 5915 9222 5967 9274
rect 5979 9222 6031 9274
rect 6043 9222 6095 9274
rect 6107 9222 6159 9274
rect 6171 9222 6223 9274
rect 15846 9222 15898 9274
rect 15910 9222 15962 9274
rect 15974 9222 16026 9274
rect 16038 9222 16090 9274
rect 16102 9222 16154 9274
rect 25776 9222 25828 9274
rect 25840 9222 25892 9274
rect 25904 9222 25956 9274
rect 25968 9222 26020 9274
rect 26032 9222 26084 9274
rect 3608 9120 3660 9172
rect 3240 8984 3292 9036
rect 3792 9027 3844 9036
rect 3792 8993 3801 9027
rect 3801 8993 3835 9027
rect 3835 8993 3844 9027
rect 3792 8984 3844 8993
rect 5080 9027 5132 9036
rect 5080 8993 5089 9027
rect 5089 8993 5123 9027
rect 5123 8993 5132 9027
rect 5080 8984 5132 8993
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 5724 8916 5776 8968
rect 6644 9120 6696 9172
rect 6828 9120 6880 9172
rect 8484 9120 8536 9172
rect 10140 9120 10192 9172
rect 13544 9120 13596 9172
rect 17868 9120 17920 9172
rect 20444 9120 20496 9172
rect 21180 9120 21232 9172
rect 11336 9052 11388 9104
rect 16396 9052 16448 9104
rect 9772 8984 9824 9036
rect 11888 8984 11940 9036
rect 18236 9052 18288 9104
rect 20260 8984 20312 9036
rect 21272 8984 21324 9036
rect 21548 9027 21600 9036
rect 21548 8993 21557 9027
rect 21557 8993 21591 9027
rect 21591 8993 21600 9027
rect 21548 8984 21600 8993
rect 8300 8959 8352 8968
rect 6276 8848 6328 8900
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 3608 8780 3660 8832
rect 7104 8780 7156 8832
rect 7288 8848 7340 8900
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 8300 8916 8352 8925
rect 8392 8916 8444 8968
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 9588 8916 9640 8968
rect 11428 8916 11480 8968
rect 11980 8916 12032 8968
rect 13268 8959 13320 8968
rect 13268 8925 13286 8959
rect 13286 8925 13320 8959
rect 13544 8959 13596 8968
rect 13268 8916 13320 8925
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 14096 8848 14148 8900
rect 14832 8848 14884 8900
rect 15568 8916 15620 8968
rect 17776 8959 17828 8968
rect 17776 8925 17785 8959
rect 17785 8925 17819 8959
rect 17819 8925 17828 8959
rect 17776 8916 17828 8925
rect 8116 8780 8168 8832
rect 10232 8780 10284 8832
rect 11520 8823 11572 8832
rect 11520 8789 11529 8823
rect 11529 8789 11563 8823
rect 11563 8789 11572 8823
rect 11520 8780 11572 8789
rect 12164 8823 12216 8832
rect 12164 8789 12173 8823
rect 12173 8789 12207 8823
rect 12207 8789 12216 8823
rect 12164 8780 12216 8789
rect 12900 8780 12952 8832
rect 15292 8780 15344 8832
rect 16488 8780 16540 8832
rect 18144 8916 18196 8968
rect 18328 8959 18380 8968
rect 18328 8925 18337 8959
rect 18337 8925 18371 8959
rect 18371 8925 18380 8959
rect 18328 8916 18380 8925
rect 20352 8959 20404 8968
rect 18788 8848 18840 8900
rect 18880 8848 18932 8900
rect 20352 8925 20361 8959
rect 20361 8925 20395 8959
rect 20395 8925 20404 8959
rect 20352 8916 20404 8925
rect 20536 8959 20588 8968
rect 20536 8925 20545 8959
rect 20545 8925 20579 8959
rect 20579 8925 20588 8959
rect 20536 8916 20588 8925
rect 20720 8959 20772 8968
rect 20720 8925 20729 8959
rect 20729 8925 20763 8959
rect 20763 8925 20772 8959
rect 20720 8916 20772 8925
rect 20904 8959 20956 8968
rect 20904 8925 20913 8959
rect 20913 8925 20947 8959
rect 20947 8925 20956 8959
rect 29828 8959 29880 8968
rect 20904 8916 20956 8925
rect 29828 8925 29837 8959
rect 29837 8925 29871 8959
rect 29871 8925 29880 8959
rect 29828 8916 29880 8925
rect 19800 8848 19852 8900
rect 21640 8848 21692 8900
rect 21824 8891 21876 8900
rect 21824 8857 21858 8891
rect 21858 8857 21876 8891
rect 21824 8848 21876 8857
rect 18420 8780 18472 8832
rect 18696 8780 18748 8832
rect 19064 8780 19116 8832
rect 22008 8780 22060 8832
rect 30012 8823 30064 8832
rect 30012 8789 30021 8823
rect 30021 8789 30055 8823
rect 30055 8789 30064 8823
rect 30012 8780 30064 8789
rect 10880 8678 10932 8730
rect 10944 8678 10996 8730
rect 11008 8678 11060 8730
rect 11072 8678 11124 8730
rect 11136 8678 11188 8730
rect 20811 8678 20863 8730
rect 20875 8678 20927 8730
rect 20939 8678 20991 8730
rect 21003 8678 21055 8730
rect 21067 8678 21119 8730
rect 3056 8619 3108 8628
rect 3056 8585 3065 8619
rect 3065 8585 3099 8619
rect 3099 8585 3108 8619
rect 3056 8576 3108 8585
rect 3608 8619 3660 8628
rect 3608 8585 3617 8619
rect 3617 8585 3651 8619
rect 3651 8585 3660 8619
rect 3608 8576 3660 8585
rect 3792 8576 3844 8628
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 2228 8440 2280 8492
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 4160 8440 4212 8492
rect 5080 8508 5132 8560
rect 5540 8576 5592 8628
rect 8300 8576 8352 8628
rect 11704 8576 11756 8628
rect 12164 8576 12216 8628
rect 12900 8576 12952 8628
rect 6552 8508 6604 8560
rect 7564 8508 7616 8560
rect 11336 8508 11388 8560
rect 4804 8440 4856 8492
rect 6828 8440 6880 8492
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 10692 8440 10744 8492
rect 12900 8440 12952 8492
rect 13636 8508 13688 8560
rect 13544 8440 13596 8492
rect 5632 8372 5684 8424
rect 6552 8372 6604 8424
rect 8392 8372 8444 8424
rect 9312 8372 9364 8424
rect 9680 8304 9732 8356
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 2412 8236 2464 8288
rect 9404 8236 9456 8288
rect 10140 8279 10192 8288
rect 10140 8245 10149 8279
rect 10149 8245 10183 8279
rect 10183 8245 10192 8279
rect 10140 8236 10192 8245
rect 11888 8304 11940 8356
rect 14004 8372 14056 8424
rect 14648 8483 14700 8492
rect 14648 8449 14682 8483
rect 14682 8449 14700 8483
rect 14648 8440 14700 8449
rect 18420 8576 18472 8628
rect 19800 8619 19852 8628
rect 19800 8585 19809 8619
rect 19809 8585 19843 8619
rect 19843 8585 19852 8619
rect 19800 8576 19852 8585
rect 20352 8576 20404 8628
rect 21824 8619 21876 8628
rect 17316 8440 17368 8492
rect 17776 8440 17828 8492
rect 17868 8440 17920 8492
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 21364 8508 21416 8560
rect 21824 8585 21833 8619
rect 21833 8585 21867 8619
rect 21867 8585 21876 8619
rect 21824 8576 21876 8585
rect 29828 8576 29880 8628
rect 21180 8440 21232 8492
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 22192 8483 22244 8492
rect 22192 8449 22201 8483
rect 22201 8449 22235 8483
rect 22235 8449 22244 8483
rect 22376 8483 22428 8492
rect 22192 8440 22244 8449
rect 22376 8449 22385 8483
rect 22385 8449 22419 8483
rect 22419 8449 22428 8483
rect 22376 8440 22428 8449
rect 29920 8483 29972 8492
rect 29920 8449 29929 8483
rect 29929 8449 29963 8483
rect 29963 8449 29972 8483
rect 29920 8440 29972 8449
rect 30104 8483 30156 8492
rect 30104 8449 30113 8483
rect 30113 8449 30147 8483
rect 30147 8449 30156 8483
rect 30104 8440 30156 8449
rect 15752 8347 15804 8356
rect 15752 8313 15761 8347
rect 15761 8313 15795 8347
rect 15795 8313 15804 8347
rect 15752 8304 15804 8313
rect 19432 8372 19484 8424
rect 20444 8372 20496 8424
rect 20720 8304 20772 8356
rect 21272 8304 21324 8356
rect 15292 8236 15344 8288
rect 20536 8279 20588 8288
rect 20536 8245 20545 8279
rect 20545 8245 20579 8279
rect 20579 8245 20588 8279
rect 20536 8236 20588 8245
rect 22192 8236 22244 8288
rect 5915 8134 5967 8186
rect 5979 8134 6031 8186
rect 6043 8134 6095 8186
rect 6107 8134 6159 8186
rect 6171 8134 6223 8186
rect 15846 8134 15898 8186
rect 15910 8134 15962 8186
rect 15974 8134 16026 8186
rect 16038 8134 16090 8186
rect 16102 8134 16154 8186
rect 25776 8134 25828 8186
rect 25840 8134 25892 8186
rect 25904 8134 25956 8186
rect 25968 8134 26020 8186
rect 26032 8134 26084 8186
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 4988 8032 5040 8084
rect 6736 8032 6788 8084
rect 7288 8075 7340 8084
rect 2044 7964 2096 8016
rect 5448 7964 5500 8016
rect 5816 7964 5868 8016
rect 7288 8041 7297 8075
rect 7297 8041 7331 8075
rect 7331 8041 7340 8075
rect 7288 8032 7340 8041
rect 10048 8075 10100 8084
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 4436 7896 4488 7948
rect 9220 7964 9272 8016
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 11980 8032 12032 8084
rect 12072 8032 12124 8084
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 10140 7964 10192 8016
rect 11520 7896 11572 7948
rect 11888 7896 11940 7948
rect 1584 7828 1636 7880
rect 1952 7828 2004 7880
rect 3056 7828 3108 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 2596 7760 2648 7812
rect 5080 7760 5132 7812
rect 5356 7760 5408 7812
rect 6276 7828 6328 7880
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 7104 7871 7156 7880
rect 6828 7828 6880 7837
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 7932 7828 7984 7880
rect 10232 7871 10284 7880
rect 7840 7803 7892 7812
rect 7840 7769 7849 7803
rect 7849 7769 7883 7803
rect 7883 7769 7892 7803
rect 7840 7760 7892 7769
rect 8484 7760 8536 7812
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 14556 7896 14608 7948
rect 10324 7828 10376 7837
rect 14096 7871 14148 7880
rect 10692 7760 10744 7812
rect 11704 7760 11756 7812
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 14372 7828 14424 7880
rect 14832 7873 14884 7880
rect 14004 7760 14056 7812
rect 14832 7839 14841 7873
rect 14841 7839 14875 7873
rect 14875 7839 14884 7873
rect 14832 7828 14884 7839
rect 15200 7871 15252 7880
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 18880 8032 18932 8084
rect 21364 8032 21416 8084
rect 19432 7964 19484 8016
rect 19708 7828 19760 7880
rect 20536 7828 20588 7880
rect 15476 7760 15528 7812
rect 16488 7760 16540 7812
rect 18052 7760 18104 7812
rect 1584 7692 1636 7744
rect 4804 7692 4856 7744
rect 6644 7692 6696 7744
rect 6736 7692 6788 7744
rect 7196 7692 7248 7744
rect 9036 7692 9088 7744
rect 9496 7692 9548 7744
rect 10600 7692 10652 7744
rect 11796 7735 11848 7744
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 11888 7735 11940 7744
rect 11888 7701 11897 7735
rect 11897 7701 11931 7735
rect 11931 7701 11940 7735
rect 11888 7692 11940 7701
rect 10880 7590 10932 7642
rect 10944 7590 10996 7642
rect 11008 7590 11060 7642
rect 11072 7590 11124 7642
rect 11136 7590 11188 7642
rect 20811 7590 20863 7642
rect 20875 7590 20927 7642
rect 20939 7590 20991 7642
rect 21003 7590 21055 7642
rect 21067 7590 21119 7642
rect 2044 7488 2096 7540
rect 4344 7488 4396 7540
rect 1768 7420 1820 7472
rect 3792 7420 3844 7472
rect 7840 7488 7892 7540
rect 10140 7531 10192 7540
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 10324 7488 10376 7540
rect 5816 7463 5868 7472
rect 5816 7429 5825 7463
rect 5825 7429 5859 7463
rect 5859 7429 5868 7463
rect 5816 7420 5868 7429
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 5172 7352 5224 7404
rect 7380 7420 7432 7472
rect 9680 7420 9732 7472
rect 9956 7420 10008 7472
rect 14648 7488 14700 7540
rect 15200 7488 15252 7540
rect 17960 7531 18012 7540
rect 6644 7352 6696 7404
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 7472 7352 7524 7404
rect 8392 7352 8444 7404
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 9036 7395 9088 7404
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9036 7352 9088 7361
rect 11428 7420 11480 7472
rect 15016 7420 15068 7472
rect 11704 7395 11756 7404
rect 4436 7284 4488 7336
rect 6828 7284 6880 7336
rect 3516 7216 3568 7268
rect 7656 7216 7708 7268
rect 8484 7216 8536 7268
rect 9312 7284 9364 7336
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 12900 7352 12952 7404
rect 14004 7395 14056 7404
rect 10600 7284 10652 7336
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 9772 7216 9824 7268
rect 9956 7216 10008 7268
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 14464 7352 14516 7404
rect 13544 7284 13596 7336
rect 14832 7352 14884 7404
rect 15200 7395 15252 7404
rect 15200 7361 15209 7395
rect 15209 7361 15243 7395
rect 15243 7361 15252 7395
rect 15200 7352 15252 7361
rect 15384 7395 15436 7404
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 15292 7284 15344 7336
rect 17960 7497 17969 7531
rect 17969 7497 18003 7531
rect 18003 7497 18012 7531
rect 17960 7488 18012 7497
rect 18604 7488 18656 7540
rect 17316 7463 17368 7472
rect 17316 7429 17325 7463
rect 17325 7429 17359 7463
rect 17359 7429 17368 7463
rect 17316 7420 17368 7429
rect 18052 7420 18104 7472
rect 16948 7352 17000 7404
rect 18236 7352 18288 7404
rect 20352 7352 20404 7404
rect 15108 7216 15160 7268
rect 19708 7284 19760 7336
rect 17500 7259 17552 7268
rect 17500 7225 17509 7259
rect 17509 7225 17543 7259
rect 17543 7225 17552 7259
rect 17500 7216 17552 7225
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 20904 7352 20956 7361
rect 21640 7352 21692 7404
rect 29552 7352 29604 7404
rect 20812 7327 20864 7336
rect 20812 7293 20821 7327
rect 20821 7293 20855 7327
rect 20855 7293 20864 7327
rect 20812 7284 20864 7293
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 9220 7191 9272 7200
rect 9220 7157 9229 7191
rect 9229 7157 9263 7191
rect 9263 7157 9272 7191
rect 9220 7148 9272 7157
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 12992 7191 13044 7200
rect 12992 7157 13001 7191
rect 13001 7157 13035 7191
rect 13035 7157 13044 7191
rect 12992 7148 13044 7157
rect 13636 7148 13688 7200
rect 15752 7148 15804 7200
rect 16856 7148 16908 7200
rect 17592 7148 17644 7200
rect 20812 7148 20864 7200
rect 21272 7148 21324 7200
rect 22100 7148 22152 7200
rect 30012 7191 30064 7200
rect 30012 7157 30021 7191
rect 30021 7157 30055 7191
rect 30055 7157 30064 7191
rect 30012 7148 30064 7157
rect 5915 7046 5967 7098
rect 5979 7046 6031 7098
rect 6043 7046 6095 7098
rect 6107 7046 6159 7098
rect 6171 7046 6223 7098
rect 15846 7046 15898 7098
rect 15910 7046 15962 7098
rect 15974 7046 16026 7098
rect 16038 7046 16090 7098
rect 16102 7046 16154 7098
rect 25776 7046 25828 7098
rect 25840 7046 25892 7098
rect 25904 7046 25956 7098
rect 25968 7046 26020 7098
rect 26032 7046 26084 7098
rect 6368 6944 6420 6996
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 1492 6740 1544 6792
rect 1860 6740 1912 6792
rect 2780 6740 2832 6792
rect 5264 6876 5316 6928
rect 5448 6808 5500 6860
rect 6736 6808 6788 6860
rect 4068 6740 4120 6792
rect 2872 6672 2924 6724
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 5172 6715 5224 6724
rect 5172 6681 5181 6715
rect 5181 6681 5215 6715
rect 5215 6681 5224 6715
rect 5172 6672 5224 6681
rect 1584 6604 1636 6656
rect 1952 6604 2004 6656
rect 2136 6647 2188 6656
rect 2136 6613 2145 6647
rect 2145 6613 2179 6647
rect 2179 6613 2188 6647
rect 2136 6604 2188 6613
rect 3700 6604 3752 6656
rect 3884 6604 3936 6656
rect 4344 6604 4396 6656
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 5356 6740 5408 6792
rect 5632 6740 5684 6792
rect 5816 6740 5868 6792
rect 5448 6672 5500 6724
rect 5908 6672 5960 6724
rect 6920 6740 6972 6792
rect 7472 6944 7524 6996
rect 7656 6944 7708 6996
rect 11888 6944 11940 6996
rect 18420 6944 18472 6996
rect 12808 6919 12860 6928
rect 12808 6885 12817 6919
rect 12817 6885 12851 6919
rect 12851 6885 12860 6919
rect 12808 6876 12860 6885
rect 14004 6876 14056 6928
rect 18788 6876 18840 6928
rect 9680 6808 9732 6860
rect 7748 6740 7800 6792
rect 8300 6740 8352 6792
rect 9956 6740 10008 6792
rect 6276 6604 6328 6656
rect 6368 6604 6420 6656
rect 6644 6604 6696 6656
rect 11428 6740 11480 6792
rect 11796 6740 11848 6792
rect 12716 6740 12768 6792
rect 12992 6740 13044 6792
rect 13728 6808 13780 6860
rect 15016 6851 15068 6860
rect 15016 6817 15025 6851
rect 15025 6817 15059 6851
rect 15059 6817 15068 6851
rect 15016 6808 15068 6817
rect 15200 6808 15252 6860
rect 15568 6808 15620 6860
rect 16856 6851 16908 6860
rect 13636 6740 13688 6792
rect 15292 6783 15344 6792
rect 12532 6672 12584 6724
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 16856 6817 16865 6851
rect 16865 6817 16899 6851
rect 16899 6817 16908 6851
rect 16856 6808 16908 6817
rect 16948 6808 17000 6860
rect 19524 6851 19576 6860
rect 16672 6783 16724 6792
rect 14832 6672 14884 6724
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 17040 6783 17092 6792
rect 17040 6749 17049 6783
rect 17049 6749 17083 6783
rect 17083 6749 17092 6783
rect 17040 6740 17092 6749
rect 17224 6740 17276 6792
rect 19524 6817 19533 6851
rect 19533 6817 19567 6851
rect 19567 6817 19576 6851
rect 19524 6808 19576 6817
rect 21272 6740 21324 6792
rect 21640 6740 21692 6792
rect 17776 6672 17828 6724
rect 18052 6672 18104 6724
rect 20720 6672 20772 6724
rect 14556 6604 14608 6656
rect 17224 6647 17276 6656
rect 17224 6613 17233 6647
rect 17233 6613 17267 6647
rect 17267 6613 17276 6647
rect 17224 6604 17276 6613
rect 21456 6647 21508 6656
rect 21456 6613 21465 6647
rect 21465 6613 21499 6647
rect 21499 6613 21508 6647
rect 21456 6604 21508 6613
rect 10880 6502 10932 6554
rect 10944 6502 10996 6554
rect 11008 6502 11060 6554
rect 11072 6502 11124 6554
rect 11136 6502 11188 6554
rect 20811 6502 20863 6554
rect 20875 6502 20927 6554
rect 20939 6502 20991 6554
rect 21003 6502 21055 6554
rect 21067 6502 21119 6554
rect 1676 6400 1728 6452
rect 2872 6443 2924 6452
rect 2872 6409 2881 6443
rect 2881 6409 2915 6443
rect 2915 6409 2924 6443
rect 2872 6400 2924 6409
rect 7012 6400 7064 6452
rect 9036 6400 9088 6452
rect 2136 6332 2188 6384
rect 3700 6332 3752 6384
rect 2044 6264 2096 6316
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 3792 6264 3844 6316
rect 5264 6307 5316 6316
rect 1860 6060 1912 6112
rect 4068 6196 4120 6248
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 6092 6264 6144 6316
rect 6276 6264 6328 6316
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 8300 6332 8352 6384
rect 30104 6400 30156 6452
rect 5356 6196 5408 6248
rect 4344 6128 4396 6180
rect 5080 6128 5132 6180
rect 5724 6128 5776 6180
rect 5908 6128 5960 6180
rect 9220 6264 9272 6316
rect 10600 6332 10652 6384
rect 10784 6375 10836 6384
rect 10784 6341 10793 6375
rect 10793 6341 10827 6375
rect 10827 6341 10836 6375
rect 10784 6332 10836 6341
rect 10968 6332 11020 6384
rect 12624 6332 12676 6384
rect 12808 6332 12860 6384
rect 13544 6332 13596 6384
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 16488 6332 16540 6384
rect 10968 6196 11020 6248
rect 11980 6196 12032 6248
rect 12348 6239 12400 6248
rect 12348 6205 12357 6239
rect 12357 6205 12391 6239
rect 12391 6205 12400 6239
rect 12348 6196 12400 6205
rect 12624 6196 12676 6248
rect 14924 6264 14976 6316
rect 17224 6264 17276 6316
rect 19708 6332 19760 6384
rect 12440 6128 12492 6180
rect 13084 6128 13136 6180
rect 15660 6171 15712 6180
rect 15660 6137 15669 6171
rect 15669 6137 15703 6171
rect 15703 6137 15712 6171
rect 15660 6128 15712 6137
rect 17040 6128 17092 6180
rect 4068 6103 4120 6112
rect 4068 6069 4077 6103
rect 4077 6069 4111 6103
rect 4111 6069 4120 6103
rect 4068 6060 4120 6069
rect 4436 6060 4488 6112
rect 13636 6103 13688 6112
rect 13636 6069 13645 6103
rect 13645 6069 13679 6103
rect 13679 6069 13688 6103
rect 13636 6060 13688 6069
rect 15292 6060 15344 6112
rect 19432 6264 19484 6316
rect 20260 6264 20312 6316
rect 20628 6264 20680 6316
rect 18420 6196 18472 6248
rect 5915 5958 5967 6010
rect 5979 5958 6031 6010
rect 6043 5958 6095 6010
rect 6107 5958 6159 6010
rect 6171 5958 6223 6010
rect 15846 5958 15898 6010
rect 15910 5958 15962 6010
rect 15974 5958 16026 6010
rect 16038 5958 16090 6010
rect 16102 5958 16154 6010
rect 25776 5958 25828 6010
rect 25840 5958 25892 6010
rect 25904 5958 25956 6010
rect 25968 5958 26020 6010
rect 26032 5958 26084 6010
rect 3792 5856 3844 5908
rect 5816 5788 5868 5840
rect 1676 5720 1728 5772
rect 4160 5763 4212 5772
rect 4160 5729 4169 5763
rect 4169 5729 4203 5763
rect 4203 5729 4212 5763
rect 4160 5720 4212 5729
rect 4436 5695 4488 5704
rect 4436 5661 4470 5695
rect 4470 5661 4488 5695
rect 4436 5652 4488 5661
rect 5356 5652 5408 5704
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 9312 5856 9364 5908
rect 10416 5856 10468 5908
rect 13452 5899 13504 5908
rect 13452 5865 13461 5899
rect 13461 5865 13495 5899
rect 13495 5865 13504 5899
rect 13452 5856 13504 5865
rect 16948 5899 17000 5908
rect 6460 5831 6512 5840
rect 6460 5797 6469 5831
rect 6469 5797 6503 5831
rect 6503 5797 6512 5831
rect 6460 5788 6512 5797
rect 8484 5788 8536 5840
rect 16948 5865 16957 5899
rect 16957 5865 16991 5899
rect 16991 5865 17000 5899
rect 16948 5856 17000 5865
rect 18052 5856 18104 5908
rect 18236 5899 18288 5908
rect 18236 5865 18245 5899
rect 18245 5865 18279 5899
rect 18279 5865 18288 5899
rect 18236 5856 18288 5865
rect 20720 5899 20772 5908
rect 20720 5865 20729 5899
rect 20729 5865 20763 5899
rect 20763 5865 20772 5899
rect 20720 5856 20772 5865
rect 6920 5720 6972 5772
rect 17776 5788 17828 5840
rect 19984 5788 20036 5840
rect 12440 5720 12492 5772
rect 4068 5584 4120 5636
rect 11244 5652 11296 5704
rect 11796 5652 11848 5704
rect 12900 5720 12952 5772
rect 13636 5720 13688 5772
rect 17592 5720 17644 5772
rect 17960 5720 18012 5772
rect 20260 5763 20312 5772
rect 20260 5729 20269 5763
rect 20269 5729 20303 5763
rect 20303 5729 20312 5763
rect 20260 5720 20312 5729
rect 20444 5720 20496 5772
rect 13544 5652 13596 5704
rect 13728 5652 13780 5704
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 16396 5652 16448 5704
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 6920 5584 6972 5636
rect 11520 5584 11572 5636
rect 13360 5584 13412 5636
rect 15752 5584 15804 5636
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 19432 5695 19484 5704
rect 19432 5661 19441 5695
rect 19441 5661 19475 5695
rect 19475 5661 19484 5695
rect 19432 5652 19484 5661
rect 19800 5652 19852 5704
rect 17960 5584 18012 5636
rect 21456 5652 21508 5704
rect 20444 5584 20496 5636
rect 2504 5516 2556 5568
rect 9128 5516 9180 5568
rect 11244 5559 11296 5568
rect 11244 5525 11253 5559
rect 11253 5525 11287 5559
rect 11287 5525 11296 5559
rect 11244 5516 11296 5525
rect 13084 5559 13136 5568
rect 13084 5525 13093 5559
rect 13093 5525 13127 5559
rect 13127 5525 13136 5559
rect 13084 5516 13136 5525
rect 10880 5414 10932 5466
rect 10944 5414 10996 5466
rect 11008 5414 11060 5466
rect 11072 5414 11124 5466
rect 11136 5414 11188 5466
rect 20811 5414 20863 5466
rect 20875 5414 20927 5466
rect 20939 5414 20991 5466
rect 21003 5414 21055 5466
rect 21067 5414 21119 5466
rect 4160 5244 4212 5296
rect 5264 5312 5316 5364
rect 6368 5312 6420 5364
rect 3884 5219 3936 5228
rect 3884 5185 3918 5219
rect 3918 5185 3936 5219
rect 3884 5176 3936 5185
rect 6828 5244 6880 5296
rect 6460 5176 6512 5228
rect 7012 5312 7064 5364
rect 11520 5355 11572 5364
rect 11520 5321 11529 5355
rect 11529 5321 11563 5355
rect 11563 5321 11572 5355
rect 11520 5312 11572 5321
rect 13084 5312 13136 5364
rect 14924 5355 14976 5364
rect 14924 5321 14933 5355
rect 14933 5321 14967 5355
rect 14967 5321 14976 5355
rect 14924 5312 14976 5321
rect 19892 5355 19944 5364
rect 19892 5321 19901 5355
rect 19901 5321 19935 5355
rect 19935 5321 19944 5355
rect 19892 5312 19944 5321
rect 8392 5219 8444 5228
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 6000 5108 6052 5160
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 8576 5219 8628 5228
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 9680 5244 9732 5296
rect 10600 5244 10652 5296
rect 14004 5244 14056 5296
rect 10048 5176 10100 5228
rect 9956 5108 10008 5160
rect 11244 5176 11296 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 12900 5176 12952 5228
rect 13912 5219 13964 5228
rect 11520 5108 11572 5160
rect 12808 5151 12860 5160
rect 12808 5117 12817 5151
rect 12817 5117 12851 5151
rect 12851 5117 12860 5151
rect 12808 5108 12860 5117
rect 5540 5040 5592 5092
rect 12532 5040 12584 5092
rect 13912 5185 13921 5219
rect 13921 5185 13955 5219
rect 13955 5185 13964 5219
rect 13912 5176 13964 5185
rect 15752 5244 15804 5296
rect 15016 5108 15068 5160
rect 15568 5176 15620 5228
rect 16304 5176 16356 5228
rect 18144 5176 18196 5228
rect 20628 5176 20680 5228
rect 21272 5219 21324 5228
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 29736 5176 29788 5228
rect 16580 5108 16632 5160
rect 18236 5108 18288 5160
rect 18972 5108 19024 5160
rect 17592 5040 17644 5092
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 13636 4972 13688 5024
rect 15108 4972 15160 5024
rect 18052 4972 18104 5024
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 30012 5015 30064 5024
rect 30012 4981 30021 5015
rect 30021 4981 30055 5015
rect 30055 4981 30064 5015
rect 30012 4972 30064 4981
rect 5915 4870 5967 4922
rect 5979 4870 6031 4922
rect 6043 4870 6095 4922
rect 6107 4870 6159 4922
rect 6171 4870 6223 4922
rect 15846 4870 15898 4922
rect 15910 4870 15962 4922
rect 15974 4870 16026 4922
rect 16038 4870 16090 4922
rect 16102 4870 16154 4922
rect 25776 4870 25828 4922
rect 25840 4870 25892 4922
rect 25904 4870 25956 4922
rect 25968 4870 26020 4922
rect 26032 4870 26084 4922
rect 5172 4768 5224 4820
rect 6460 4768 6512 4820
rect 6920 4768 6972 4820
rect 5908 4700 5960 4752
rect 9864 4768 9916 4820
rect 10692 4768 10744 4820
rect 14188 4768 14240 4820
rect 15384 4768 15436 4820
rect 18696 4768 18748 4820
rect 19340 4811 19392 4820
rect 19340 4777 19349 4811
rect 19349 4777 19383 4811
rect 19383 4777 19392 4811
rect 19340 4768 19392 4777
rect 1216 4632 1268 4684
rect 4620 4632 4672 4684
rect 5448 4632 5500 4684
rect 6644 4632 6696 4684
rect 8300 4632 8352 4684
rect 9680 4632 9732 4684
rect 5632 4564 5684 4616
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6368 4564 6420 4616
rect 6552 4564 6604 4616
rect 8392 4564 8444 4616
rect 6736 4496 6788 4548
rect 7104 4496 7156 4548
rect 9036 4564 9088 4616
rect 9312 4496 9364 4548
rect 9772 4564 9824 4616
rect 10508 4564 10560 4616
rect 18052 4700 18104 4752
rect 20260 4768 20312 4820
rect 20628 4811 20680 4820
rect 20628 4777 20637 4811
rect 20637 4777 20671 4811
rect 20671 4777 20680 4811
rect 20628 4768 20680 4777
rect 13084 4632 13136 4684
rect 14096 4632 14148 4684
rect 14556 4675 14608 4684
rect 14556 4641 14565 4675
rect 14565 4641 14599 4675
rect 14599 4641 14608 4675
rect 14556 4632 14608 4641
rect 5540 4428 5592 4480
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 9864 4496 9916 4548
rect 11612 4539 11664 4548
rect 9956 4428 10008 4480
rect 10416 4428 10468 4480
rect 11612 4505 11621 4539
rect 11621 4505 11655 4539
rect 11655 4505 11664 4539
rect 11612 4496 11664 4505
rect 11888 4496 11940 4548
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 13636 4564 13688 4616
rect 15936 4632 15988 4684
rect 17776 4632 17828 4684
rect 19892 4700 19944 4752
rect 16396 4564 16448 4616
rect 16764 4564 16816 4616
rect 12440 4496 12492 4548
rect 15016 4496 15068 4548
rect 16028 4496 16080 4548
rect 17500 4564 17552 4616
rect 12072 4428 12124 4480
rect 12532 4471 12584 4480
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 15568 4428 15620 4480
rect 15752 4471 15804 4480
rect 15752 4437 15761 4471
rect 15761 4437 15795 4471
rect 15795 4437 15804 4471
rect 16488 4471 16540 4480
rect 15752 4428 15804 4437
rect 16488 4437 16497 4471
rect 16497 4437 16531 4471
rect 16531 4437 16540 4471
rect 16488 4428 16540 4437
rect 18052 4564 18104 4616
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 19340 4564 19392 4616
rect 19800 4564 19852 4616
rect 20076 4607 20128 4616
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 19984 4496 20036 4548
rect 20260 4607 20312 4616
rect 20260 4573 20269 4607
rect 20269 4573 20303 4607
rect 20303 4573 20312 4607
rect 20260 4564 20312 4573
rect 20536 4496 20588 4548
rect 19432 4428 19484 4480
rect 29644 4428 29696 4480
rect 10880 4326 10932 4378
rect 10944 4326 10996 4378
rect 11008 4326 11060 4378
rect 11072 4326 11124 4378
rect 11136 4326 11188 4378
rect 20811 4326 20863 4378
rect 20875 4326 20927 4378
rect 20939 4326 20991 4378
rect 21003 4326 21055 4378
rect 21067 4326 21119 4378
rect 1860 4199 1912 4208
rect 1860 4165 1869 4199
rect 1869 4165 1903 4199
rect 1903 4165 1912 4199
rect 1860 4156 1912 4165
rect 5908 4224 5960 4276
rect 6736 4224 6788 4276
rect 7104 4267 7156 4276
rect 7104 4233 7113 4267
rect 7113 4233 7147 4267
rect 7147 4233 7156 4267
rect 7104 4224 7156 4233
rect 10048 4224 10100 4276
rect 15568 4267 15620 4276
rect 15568 4233 15577 4267
rect 15577 4233 15611 4267
rect 15611 4233 15620 4267
rect 15568 4224 15620 4233
rect 16580 4224 16632 4276
rect 18512 4224 18564 4276
rect 2780 4131 2832 4140
rect 2780 4097 2789 4131
rect 2789 4097 2823 4131
rect 2823 4097 2832 4131
rect 2780 4088 2832 4097
rect 3148 4088 3200 4140
rect 2596 4020 2648 4072
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5356 4131 5408 4140
rect 5172 4088 5224 4097
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 6368 4131 6420 4140
rect 5080 4020 5132 4072
rect 3056 3995 3108 4004
rect 3056 3961 3065 3995
rect 3065 3961 3099 3995
rect 3099 3961 3108 3995
rect 3056 3952 3108 3961
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 9128 4156 9180 4208
rect 13360 4156 13412 4208
rect 17040 4199 17092 4208
rect 6736 4131 6788 4140
rect 6736 4097 6745 4131
rect 6745 4097 6779 4131
rect 6779 4097 6788 4131
rect 6920 4131 6972 4140
rect 6736 4088 6788 4097
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 5816 4020 5868 4072
rect 7564 4020 7616 4072
rect 9864 4088 9916 4140
rect 9312 4020 9364 4072
rect 4804 3884 4856 3936
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 6736 3884 6788 3936
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 10784 4088 10836 4140
rect 12072 4088 12124 4140
rect 12532 4088 12584 4140
rect 13728 4088 13780 4140
rect 17040 4165 17049 4199
rect 17049 4165 17083 4199
rect 17083 4165 17092 4199
rect 17040 4156 17092 4165
rect 19340 4156 19392 4208
rect 15384 4088 15436 4140
rect 15752 4131 15804 4140
rect 15752 4097 15761 4131
rect 15761 4097 15795 4131
rect 15795 4097 15804 4131
rect 15752 4088 15804 4097
rect 15936 4131 15988 4140
rect 15936 4097 15945 4131
rect 15945 4097 15979 4131
rect 15979 4097 15988 4131
rect 15936 4088 15988 4097
rect 16028 4131 16080 4140
rect 16028 4097 16037 4131
rect 16037 4097 16071 4131
rect 16071 4097 16080 4131
rect 16028 4088 16080 4097
rect 17316 4088 17368 4140
rect 19432 4131 19484 4140
rect 19432 4097 19450 4131
rect 19450 4097 19484 4131
rect 19708 4131 19760 4140
rect 19432 4088 19484 4097
rect 19708 4097 19717 4131
rect 19717 4097 19751 4131
rect 19751 4097 19760 4131
rect 19708 4088 19760 4097
rect 19800 4088 19852 4140
rect 20352 4131 20404 4140
rect 20352 4097 20361 4131
rect 20361 4097 20395 4131
rect 20395 4097 20404 4131
rect 20352 4088 20404 4097
rect 21364 4088 21416 4140
rect 30104 4131 30156 4140
rect 10600 4020 10652 4072
rect 11888 4063 11940 4072
rect 11888 4029 11897 4063
rect 11897 4029 11931 4063
rect 11931 4029 11940 4063
rect 11888 4020 11940 4029
rect 12164 4020 12216 4072
rect 12624 4020 12676 4072
rect 12808 4020 12860 4072
rect 15292 4020 15344 4072
rect 16396 4020 16448 4072
rect 17224 4063 17276 4072
rect 17224 4029 17233 4063
rect 17233 4029 17267 4063
rect 17267 4029 17276 4063
rect 17224 4020 17276 4029
rect 19984 4020 20036 4072
rect 20536 4063 20588 4072
rect 20536 4029 20545 4063
rect 20545 4029 20579 4063
rect 20579 4029 20588 4063
rect 30104 4097 30113 4131
rect 30113 4097 30147 4131
rect 30147 4097 30156 4131
rect 30104 4088 30156 4097
rect 20536 4020 20588 4029
rect 31576 4020 31628 4072
rect 11796 3952 11848 4004
rect 12532 3952 12584 4004
rect 13912 3952 13964 4004
rect 14188 3952 14240 4004
rect 16304 3952 16356 4004
rect 20076 3952 20128 4004
rect 20628 3952 20680 4004
rect 21456 3952 21508 4004
rect 10876 3927 10928 3936
rect 10876 3893 10885 3927
rect 10885 3893 10919 3927
rect 10919 3893 10928 3927
rect 10876 3884 10928 3893
rect 12440 3884 12492 3936
rect 20904 3927 20956 3936
rect 20904 3893 20913 3927
rect 20913 3893 20947 3927
rect 20947 3893 20956 3927
rect 20904 3884 20956 3893
rect 21180 3884 21232 3936
rect 21548 3884 21600 3936
rect 29552 3884 29604 3936
rect 30012 3884 30064 3936
rect 5915 3782 5967 3834
rect 5979 3782 6031 3834
rect 6043 3782 6095 3834
rect 6107 3782 6159 3834
rect 6171 3782 6223 3834
rect 15846 3782 15898 3834
rect 15910 3782 15962 3834
rect 15974 3782 16026 3834
rect 16038 3782 16090 3834
rect 16102 3782 16154 3834
rect 25776 3782 25828 3834
rect 25840 3782 25892 3834
rect 25904 3782 25956 3834
rect 25968 3782 26020 3834
rect 26032 3782 26084 3834
rect 2320 3680 2372 3732
rect 2412 3723 2464 3732
rect 2412 3689 2421 3723
rect 2421 3689 2455 3723
rect 2455 3689 2464 3723
rect 2412 3680 2464 3689
rect 4252 3680 4304 3732
rect 5632 3680 5684 3732
rect 10140 3680 10192 3732
rect 10784 3723 10836 3732
rect 6552 3612 6604 3664
rect 6828 3612 6880 3664
rect 8944 3612 8996 3664
rect 4160 3544 4212 3596
rect 8300 3544 8352 3596
rect 9220 3544 9272 3596
rect 10784 3689 10793 3723
rect 10793 3689 10827 3723
rect 10827 3689 10836 3723
rect 10784 3680 10836 3689
rect 12440 3680 12492 3732
rect 13636 3680 13688 3732
rect 15476 3680 15528 3732
rect 16672 3680 16724 3732
rect 17960 3723 18012 3732
rect 17960 3689 17969 3723
rect 17969 3689 18003 3723
rect 18003 3689 18012 3723
rect 17960 3680 18012 3689
rect 19340 3680 19392 3732
rect 20444 3680 20496 3732
rect 10784 3544 10836 3596
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 2504 3519 2556 3528
rect 2504 3485 2513 3519
rect 2513 3485 2547 3519
rect 2547 3485 2556 3519
rect 2504 3476 2556 3485
rect 5540 3519 5592 3528
rect 5540 3485 5574 3519
rect 5574 3485 5592 3519
rect 5540 3476 5592 3485
rect 10876 3476 10928 3528
rect 13176 3544 13228 3596
rect 13728 3544 13780 3596
rect 16212 3612 16264 3664
rect 21548 3680 21600 3732
rect 22928 3612 22980 3664
rect 17224 3544 17276 3596
rect 18512 3587 18564 3596
rect 18512 3553 18521 3587
rect 18521 3553 18555 3587
rect 18555 3553 18564 3587
rect 18512 3544 18564 3553
rect 21180 3544 21232 3596
rect 21456 3587 21508 3596
rect 21456 3553 21465 3587
rect 21465 3553 21499 3587
rect 21499 3553 21508 3587
rect 21456 3544 21508 3553
rect 2872 3408 2924 3460
rect 4252 3408 4304 3460
rect 9588 3408 9640 3460
rect 11888 3476 11940 3528
rect 12440 3476 12492 3528
rect 12992 3476 13044 3528
rect 16488 3476 16540 3528
rect 20904 3476 20956 3528
rect 21088 3476 21140 3528
rect 11520 3408 11572 3460
rect 13268 3408 13320 3460
rect 16764 3408 16816 3460
rect 17960 3408 18012 3460
rect 19248 3408 19300 3460
rect 19432 3408 19484 3460
rect 22468 3476 22520 3528
rect 27896 3476 27948 3528
rect 28540 3476 28592 3528
rect 29276 3476 29328 3528
rect 21824 3408 21876 3460
rect 8116 3340 8168 3392
rect 12164 3340 12216 3392
rect 17132 3383 17184 3392
rect 17132 3349 17141 3383
rect 17141 3349 17175 3383
rect 17175 3349 17184 3383
rect 17132 3340 17184 3349
rect 17224 3383 17276 3392
rect 17224 3349 17233 3383
rect 17233 3349 17267 3383
rect 17267 3349 17276 3383
rect 18328 3383 18380 3392
rect 17224 3340 17276 3349
rect 18328 3349 18337 3383
rect 18337 3349 18371 3383
rect 18371 3349 18380 3383
rect 18328 3340 18380 3349
rect 20720 3340 20772 3392
rect 21272 3340 21324 3392
rect 27804 3340 27856 3392
rect 27988 3340 28040 3392
rect 29920 3340 29972 3392
rect 10880 3238 10932 3290
rect 10944 3238 10996 3290
rect 11008 3238 11060 3290
rect 11072 3238 11124 3290
rect 11136 3238 11188 3290
rect 20811 3238 20863 3290
rect 20875 3238 20927 3290
rect 20939 3238 20991 3290
rect 21003 3238 21055 3290
rect 21067 3238 21119 3290
rect 2964 3068 3016 3120
rect 3148 3111 3200 3120
rect 3148 3077 3157 3111
rect 3157 3077 3191 3111
rect 3191 3077 3200 3111
rect 3148 3068 3200 3077
rect 4988 3068 5040 3120
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 3424 3000 3476 3052
rect 4160 3000 4212 3052
rect 5172 3000 5224 3052
rect 6460 3000 6512 3052
rect 7196 3000 7248 3052
rect 9588 3136 9640 3188
rect 9772 3136 9824 3188
rect 11612 3136 11664 3188
rect 14280 3136 14332 3188
rect 16764 3136 16816 3188
rect 9680 3068 9732 3120
rect 10784 3068 10836 3120
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 18052 3136 18104 3188
rect 18236 3136 18288 3188
rect 18328 3136 18380 3188
rect 17960 3068 18012 3120
rect 21272 3136 21324 3188
rect 22100 3136 22152 3188
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 14096 3043 14148 3052
rect 13084 3000 13136 3009
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 14096 3000 14148 3009
rect 14556 3000 14608 3052
rect 15108 3043 15160 3052
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 16396 3000 16448 3052
rect 17224 3000 17276 3052
rect 18144 3000 18196 3052
rect 20352 3068 20404 3120
rect 21824 3068 21876 3120
rect 19248 3043 19300 3052
rect 11796 2932 11848 2984
rect 6736 2907 6788 2916
rect 6736 2873 6745 2907
rect 6745 2873 6779 2907
rect 6779 2873 6788 2907
rect 6736 2864 6788 2873
rect 9036 2864 9088 2916
rect 13636 2932 13688 2984
rect 14004 2975 14056 2984
rect 14004 2941 14013 2975
rect 14013 2941 14047 2975
rect 14047 2941 14056 2975
rect 14004 2932 14056 2941
rect 15200 2932 15252 2984
rect 19248 3009 19257 3043
rect 19257 3009 19291 3043
rect 19291 3009 19300 3043
rect 19248 3000 19300 3009
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 21180 3000 21232 3052
rect 18512 2932 18564 2984
rect 18972 2975 19024 2984
rect 18972 2941 18981 2975
rect 18981 2941 19015 2975
rect 19015 2941 19024 2975
rect 18972 2932 19024 2941
rect 21916 3000 21968 3052
rect 22376 3068 22428 3120
rect 25044 3068 25096 3120
rect 27988 3068 28040 3120
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22100 3000 22152 3009
rect 22560 3000 22612 3052
rect 7104 2796 7156 2848
rect 8116 2839 8168 2848
rect 8116 2805 8125 2839
rect 8125 2805 8159 2839
rect 8159 2805 8168 2839
rect 8116 2796 8168 2805
rect 8760 2796 8812 2848
rect 21732 2932 21784 2984
rect 23204 3000 23256 3052
rect 27160 3000 27212 3052
rect 29552 3043 29604 3052
rect 29552 3009 29561 3043
rect 29561 3009 29595 3043
rect 29595 3009 29604 3043
rect 29552 3000 29604 3009
rect 29920 3043 29972 3052
rect 29920 3009 29929 3043
rect 29929 3009 29963 3043
rect 29963 3009 29972 3043
rect 29920 3000 29972 3009
rect 30012 3043 30064 3052
rect 30012 3009 30021 3043
rect 30021 3009 30055 3043
rect 30055 3009 30064 3043
rect 30012 3000 30064 3009
rect 27620 2975 27672 2984
rect 27620 2941 27629 2975
rect 27629 2941 27663 2975
rect 27663 2941 27672 2975
rect 27620 2932 27672 2941
rect 12992 2796 13044 2848
rect 22008 2864 22060 2916
rect 24400 2864 24452 2916
rect 15200 2839 15252 2848
rect 15200 2805 15209 2839
rect 15209 2805 15243 2839
rect 15243 2805 15252 2839
rect 15200 2796 15252 2805
rect 17316 2839 17368 2848
rect 17316 2805 17325 2839
rect 17325 2805 17359 2839
rect 17359 2805 17368 2839
rect 17316 2796 17368 2805
rect 17684 2796 17736 2848
rect 18144 2796 18196 2848
rect 18696 2796 18748 2848
rect 20444 2839 20496 2848
rect 20444 2805 20453 2839
rect 20453 2805 20487 2839
rect 20487 2805 20496 2839
rect 20444 2796 20496 2805
rect 21088 2796 21140 2848
rect 21180 2796 21232 2848
rect 22284 2839 22336 2848
rect 22284 2805 22293 2839
rect 22293 2805 22327 2839
rect 22327 2805 22336 2839
rect 22284 2796 22336 2805
rect 22928 2839 22980 2848
rect 22928 2805 22937 2839
rect 22937 2805 22971 2839
rect 22971 2805 22980 2839
rect 22928 2796 22980 2805
rect 27804 2839 27856 2848
rect 27804 2805 27813 2839
rect 27813 2805 27847 2839
rect 27847 2805 27856 2839
rect 27804 2796 27856 2805
rect 28632 2839 28684 2848
rect 28632 2805 28641 2839
rect 28641 2805 28675 2839
rect 28675 2805 28684 2839
rect 28632 2796 28684 2805
rect 29644 2839 29696 2848
rect 29644 2805 29653 2839
rect 29653 2805 29687 2839
rect 29687 2805 29696 2839
rect 29644 2796 29696 2805
rect 30840 2796 30892 2848
rect 5915 2694 5967 2746
rect 5979 2694 6031 2746
rect 6043 2694 6095 2746
rect 6107 2694 6159 2746
rect 6171 2694 6223 2746
rect 15846 2694 15898 2746
rect 15910 2694 15962 2746
rect 15974 2694 16026 2746
rect 16038 2694 16090 2746
rect 16102 2694 16154 2746
rect 25776 2694 25828 2746
rect 25840 2694 25892 2746
rect 25904 2694 25956 2746
rect 25968 2694 26020 2746
rect 26032 2694 26084 2746
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 6828 2592 6880 2644
rect 8760 2592 8812 2644
rect 11704 2592 11756 2644
rect 14096 2635 14148 2644
rect 14096 2601 14105 2635
rect 14105 2601 14139 2635
rect 14139 2601 14148 2635
rect 14096 2592 14148 2601
rect 15016 2635 15068 2644
rect 15016 2601 15025 2635
rect 15025 2601 15059 2635
rect 15059 2601 15068 2635
rect 15016 2592 15068 2601
rect 15384 2592 15436 2644
rect 17132 2592 17184 2644
rect 17684 2592 17736 2644
rect 20720 2592 20772 2644
rect 21088 2635 21140 2644
rect 21088 2601 21097 2635
rect 21097 2601 21131 2635
rect 21131 2601 21140 2635
rect 21088 2592 21140 2601
rect 21916 2635 21968 2644
rect 21916 2601 21925 2635
rect 21925 2601 21959 2635
rect 21959 2601 21968 2635
rect 21916 2592 21968 2601
rect 22560 2592 22612 2644
rect 27160 2635 27212 2644
rect 27160 2601 27169 2635
rect 27169 2601 27203 2635
rect 27203 2601 27212 2635
rect 27160 2592 27212 2601
rect 27620 2635 27672 2644
rect 27620 2601 27629 2635
rect 27629 2601 27663 2635
rect 27663 2601 27672 2635
rect 27620 2592 27672 2601
rect 30012 2635 30064 2644
rect 30012 2601 30021 2635
rect 30021 2601 30055 2635
rect 30055 2601 30064 2635
rect 30012 2592 30064 2601
rect 8576 2524 8628 2576
rect 2504 2456 2556 2508
rect 11428 2524 11480 2576
rect 15292 2524 15344 2576
rect 17224 2524 17276 2576
rect 9956 2456 10008 2508
rect 11980 2456 12032 2508
rect 16212 2456 16264 2508
rect 17040 2456 17092 2508
rect 1860 2388 1912 2440
rect 388 2320 440 2372
rect 4896 2388 4948 2440
rect 2780 2320 2832 2372
rect 5724 2388 5776 2440
rect 7932 2388 7984 2440
rect 8668 2388 8720 2440
rect 8760 2388 8812 2440
rect 9496 2388 9548 2440
rect 10232 2388 10284 2440
rect 13728 2388 13780 2440
rect 14004 2388 14056 2440
rect 15108 2388 15160 2440
rect 15292 2388 15344 2440
rect 15568 2388 15620 2440
rect 17684 2388 17736 2440
rect 20260 2524 20312 2576
rect 24400 2567 24452 2576
rect 17868 2456 17920 2508
rect 17960 2431 18012 2440
rect 17960 2397 17969 2431
rect 17969 2397 18003 2431
rect 18003 2397 18012 2431
rect 17960 2388 18012 2397
rect 18696 2431 18748 2440
rect 9404 2320 9456 2372
rect 14372 2320 14424 2372
rect 18696 2397 18705 2431
rect 18705 2397 18739 2431
rect 18739 2397 18748 2431
rect 18696 2388 18748 2397
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 21824 2456 21876 2508
rect 23296 2456 23348 2508
rect 18972 2320 19024 2372
rect 22284 2388 22336 2440
rect 22652 2388 22704 2440
rect 22836 2431 22888 2440
rect 22836 2397 22845 2431
rect 22845 2397 22879 2431
rect 22879 2397 22888 2431
rect 22836 2388 22888 2397
rect 24400 2533 24409 2567
rect 24409 2533 24443 2567
rect 24443 2533 24452 2567
rect 24400 2524 24452 2533
rect 25044 2567 25096 2576
rect 25044 2533 25053 2567
rect 25053 2533 25087 2567
rect 25087 2533 25096 2567
rect 25044 2524 25096 2533
rect 23940 2388 23992 2440
rect 24768 2388 24820 2440
rect 25504 2388 25556 2440
rect 26240 2388 26292 2440
rect 27068 2388 27120 2440
rect 28724 2431 28776 2440
rect 28724 2397 28733 2431
rect 28733 2397 28767 2431
rect 28767 2397 28776 2431
rect 28724 2388 28776 2397
rect 29092 2388 29144 2440
rect 12072 2252 12124 2304
rect 16856 2252 16908 2304
rect 18328 2252 18380 2304
rect 20168 2252 20220 2304
rect 28632 2320 28684 2372
rect 22560 2252 22612 2304
rect 22652 2295 22704 2304
rect 22652 2261 22661 2295
rect 22661 2261 22695 2295
rect 22695 2261 22704 2295
rect 23296 2295 23348 2304
rect 22652 2252 22704 2261
rect 23296 2261 23305 2295
rect 23305 2261 23339 2295
rect 23339 2261 23348 2295
rect 23296 2252 23348 2261
rect 28908 2295 28960 2304
rect 28908 2261 28917 2295
rect 28917 2261 28951 2295
rect 28951 2261 28960 2295
rect 28908 2252 28960 2261
rect 10880 2150 10932 2202
rect 10944 2150 10996 2202
rect 11008 2150 11060 2202
rect 11072 2150 11124 2202
rect 11136 2150 11188 2202
rect 20811 2150 20863 2202
rect 20875 2150 20927 2202
rect 20939 2150 20991 2202
rect 21003 2150 21055 2202
rect 21067 2150 21119 2202
rect 16856 2048 16908 2100
rect 18328 2048 18380 2100
rect 18604 2048 18656 2100
rect 22836 2048 22888 2100
rect 13084 1912 13136 1964
rect 20168 1912 20220 1964
rect 9404 1368 9456 1420
rect 11060 1368 11112 1420
rect 17132 1368 17184 1420
rect 18696 1368 18748 1420
<< metal2 >>
rect 2778 47560 2834 47569
rect 2778 47495 2834 47504
rect 1676 45484 1728 45490
rect 1676 45426 1728 45432
rect 1492 44736 1544 44742
rect 1492 44678 1544 44684
rect 1504 44577 1532 44678
rect 1490 44568 1546 44577
rect 1490 44503 1546 44512
rect 1492 44192 1544 44198
rect 1492 44134 1544 44140
rect 1504 43897 1532 44134
rect 1490 43888 1546 43897
rect 1490 43823 1546 43832
rect 1492 43648 1544 43654
rect 1492 43590 1544 43596
rect 1400 43104 1452 43110
rect 1504 43081 1532 43590
rect 1400 43046 1452 43052
rect 1490 43072 1546 43081
rect 1412 42401 1440 43046
rect 1490 43007 1546 43016
rect 1492 42560 1544 42566
rect 1492 42502 1544 42508
rect 1398 42392 1454 42401
rect 1398 42327 1454 42336
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1308 41472 1360 41478
rect 1308 41414 1360 41420
rect 1320 40225 1348 41414
rect 1412 40905 1440 41958
rect 1504 41721 1532 42502
rect 1490 41712 1546 41721
rect 1490 41647 1546 41656
rect 1398 40896 1454 40905
rect 1398 40831 1454 40840
rect 1492 40384 1544 40390
rect 1492 40326 1544 40332
rect 1306 40216 1362 40225
rect 1306 40151 1362 40160
rect 1400 39840 1452 39846
rect 1400 39782 1452 39788
rect 1412 38729 1440 39782
rect 1504 39409 1532 40326
rect 1490 39400 1546 39409
rect 1490 39335 1546 39344
rect 1398 38720 1454 38729
rect 1398 38655 1454 38664
rect 1492 37664 1544 37670
rect 1492 37606 1544 37612
rect 1504 36553 1532 37606
rect 1490 36544 1546 36553
rect 1490 36479 1546 36488
rect 1492 36032 1544 36038
rect 1492 35974 1544 35980
rect 1504 35057 1532 35974
rect 1490 35048 1546 35057
rect 1490 34983 1546 34992
rect 1492 33312 1544 33318
rect 1492 33254 1544 33260
rect 1400 32904 1452 32910
rect 1400 32846 1452 32852
rect 1412 31482 1440 32846
rect 1504 32745 1532 33254
rect 1584 32768 1636 32774
rect 1490 32736 1546 32745
rect 1584 32710 1636 32716
rect 1490 32671 1546 32680
rect 1596 32065 1624 32710
rect 1582 32056 1638 32065
rect 1582 31991 1638 32000
rect 1492 31680 1544 31686
rect 1492 31622 1544 31628
rect 1400 31476 1452 31482
rect 1400 31418 1452 31424
rect 1504 31385 1532 31622
rect 1490 31376 1546 31385
rect 1490 31311 1546 31320
rect 1490 29064 1546 29073
rect 1490 28999 1492 29008
rect 1544 28999 1546 29008
rect 1492 28970 1544 28976
rect 1688 28608 1716 45426
rect 2226 45384 2282 45393
rect 2226 45319 2228 45328
rect 2280 45319 2282 45328
rect 2228 45290 2280 45296
rect 2792 45286 2820 47495
rect 30010 47016 30066 47025
rect 30010 46951 30066 46960
rect 2870 46880 2926 46889
rect 2870 46815 2926 46824
rect 2780 45280 2832 45286
rect 2780 45222 2832 45228
rect 2884 45082 2912 46815
rect 2962 46064 3018 46073
rect 2962 45999 3018 46008
rect 2976 45354 3004 45999
rect 10880 45724 11188 45744
rect 10880 45722 10886 45724
rect 10942 45722 10966 45724
rect 11022 45722 11046 45724
rect 11102 45722 11126 45724
rect 11182 45722 11188 45724
rect 10942 45670 10944 45722
rect 11124 45670 11126 45722
rect 10880 45668 10886 45670
rect 10942 45668 10966 45670
rect 11022 45668 11046 45670
rect 11102 45668 11126 45670
rect 11182 45668 11188 45670
rect 10880 45648 11188 45668
rect 20811 45724 21119 45744
rect 20811 45722 20817 45724
rect 20873 45722 20897 45724
rect 20953 45722 20977 45724
rect 21033 45722 21057 45724
rect 21113 45722 21119 45724
rect 20873 45670 20875 45722
rect 21055 45670 21057 45722
rect 20811 45668 20817 45670
rect 20873 45668 20897 45670
rect 20953 45668 20977 45670
rect 21033 45668 21057 45670
rect 21113 45668 21119 45670
rect 20811 45648 21119 45668
rect 4528 45484 4580 45490
rect 4528 45426 4580 45432
rect 4896 45484 4948 45490
rect 4896 45426 4948 45432
rect 5448 45484 5500 45490
rect 5448 45426 5500 45432
rect 6460 45484 6512 45490
rect 6460 45426 6512 45432
rect 7288 45484 7340 45490
rect 7288 45426 7340 45432
rect 2964 45348 3016 45354
rect 2964 45290 3016 45296
rect 3792 45280 3844 45286
rect 3792 45222 3844 45228
rect 4436 45280 4488 45286
rect 4436 45222 4488 45228
rect 2872 45076 2924 45082
rect 2872 45018 2924 45024
rect 2412 44872 2464 44878
rect 2410 44840 2412 44849
rect 3148 44872 3200 44878
rect 2464 44840 2466 44849
rect 3148 44814 3200 44820
rect 2410 44775 2466 44784
rect 2872 44736 2924 44742
rect 2872 44678 2924 44684
rect 2320 44396 2372 44402
rect 2320 44338 2372 44344
rect 1768 44192 1820 44198
rect 1768 44134 1820 44140
rect 1780 40526 1808 44134
rect 1860 43308 1912 43314
rect 1860 43250 1912 43256
rect 1768 40520 1820 40526
rect 1768 40462 1820 40468
rect 1872 39114 1900 43250
rect 2136 43104 2188 43110
rect 2136 43046 2188 43052
rect 2148 41138 2176 43046
rect 2228 42696 2280 42702
rect 2228 42638 2280 42644
rect 2240 42090 2268 42638
rect 2228 42084 2280 42090
rect 2228 42026 2280 42032
rect 2240 41614 2268 42026
rect 2228 41608 2280 41614
rect 2228 41550 2280 41556
rect 2136 41132 2188 41138
rect 2136 41074 2188 41080
rect 2148 39574 2176 41074
rect 2240 40662 2268 41550
rect 2228 40656 2280 40662
rect 2228 40598 2280 40604
rect 2332 39624 2360 44338
rect 2884 43858 2912 44678
rect 2964 44396 3016 44402
rect 2964 44338 3016 44344
rect 2872 43852 2924 43858
rect 2872 43794 2924 43800
rect 2596 43784 2648 43790
rect 2596 43726 2648 43732
rect 2504 43648 2556 43654
rect 2504 43590 2556 43596
rect 2516 42906 2544 43590
rect 2504 42900 2556 42906
rect 2504 42842 2556 42848
rect 2516 42022 2544 42842
rect 2504 42016 2556 42022
rect 2504 41958 2556 41964
rect 2516 41818 2544 41958
rect 2504 41812 2556 41818
rect 2424 41772 2504 41800
rect 2424 40934 2452 41772
rect 2504 41754 2556 41760
rect 2412 40928 2464 40934
rect 2412 40870 2464 40876
rect 2424 40730 2452 40870
rect 2412 40724 2464 40730
rect 2412 40666 2464 40672
rect 2412 39636 2464 39642
rect 2332 39596 2412 39624
rect 2412 39578 2464 39584
rect 2136 39568 2188 39574
rect 2136 39510 2188 39516
rect 1780 39086 1900 39114
rect 1780 36786 1808 39086
rect 2148 38962 2176 39510
rect 2412 39500 2464 39506
rect 2412 39442 2464 39448
rect 1860 38956 1912 38962
rect 1860 38898 1912 38904
rect 2136 38956 2188 38962
rect 2136 38898 2188 38904
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1780 36310 1808 36722
rect 1768 36304 1820 36310
rect 1768 36246 1820 36252
rect 1872 34746 1900 38898
rect 2148 38486 2176 38898
rect 2424 38758 2452 39442
rect 2504 39024 2556 39030
rect 2504 38966 2556 38972
rect 2412 38752 2464 38758
rect 2412 38694 2464 38700
rect 2424 38554 2452 38694
rect 2412 38548 2464 38554
rect 2412 38490 2464 38496
rect 2136 38480 2188 38486
rect 2136 38422 2188 38428
rect 1952 37256 2004 37262
rect 1952 37198 2004 37204
rect 1964 36922 1992 37198
rect 1952 36916 2004 36922
rect 1952 36858 2004 36864
rect 1964 35698 1992 36858
rect 2148 36786 2176 38422
rect 2424 37466 2452 38490
rect 2516 38418 2544 38966
rect 2608 38554 2636 43726
rect 2780 43308 2832 43314
rect 2780 43250 2832 43256
rect 2688 42152 2740 42158
rect 2688 42094 2740 42100
rect 2700 41614 2728 42094
rect 2688 41608 2740 41614
rect 2688 41550 2740 41556
rect 2792 38962 2820 43250
rect 2976 43194 3004 44338
rect 3056 44192 3108 44198
rect 3056 44134 3108 44140
rect 2884 43166 3004 43194
rect 2884 40730 2912 43166
rect 2964 43104 3016 43110
rect 2964 43046 3016 43052
rect 2872 40724 2924 40730
rect 2872 40666 2924 40672
rect 2780 38956 2832 38962
rect 2780 38898 2832 38904
rect 2780 38820 2832 38826
rect 2780 38762 2832 38768
rect 2596 38548 2648 38554
rect 2596 38490 2648 38496
rect 2504 38412 2556 38418
rect 2504 38354 2556 38360
rect 2516 38010 2544 38354
rect 2504 38004 2556 38010
rect 2504 37946 2556 37952
rect 2412 37460 2464 37466
rect 2412 37402 2464 37408
rect 2136 36780 2188 36786
rect 2136 36722 2188 36728
rect 2424 36582 2452 37402
rect 2412 36576 2464 36582
rect 2412 36518 2464 36524
rect 2320 36304 2372 36310
rect 2320 36246 2372 36252
rect 2228 36032 2280 36038
rect 2228 35974 2280 35980
rect 2240 35737 2268 35974
rect 2226 35728 2282 35737
rect 1952 35692 2004 35698
rect 2226 35663 2282 35672
rect 1952 35634 2004 35640
rect 1964 35222 1992 35634
rect 2228 35488 2280 35494
rect 2228 35430 2280 35436
rect 2240 35290 2268 35430
rect 2228 35284 2280 35290
rect 2228 35226 2280 35232
rect 1952 35216 2004 35222
rect 1952 35158 2004 35164
rect 1860 34740 1912 34746
rect 1860 34682 1912 34688
rect 1964 34610 1992 35158
rect 1952 34604 2004 34610
rect 1952 34546 2004 34552
rect 1964 34134 1992 34546
rect 2240 34406 2268 35226
rect 2228 34400 2280 34406
rect 2228 34342 2280 34348
rect 2240 34202 2268 34342
rect 2228 34196 2280 34202
rect 2228 34138 2280 34144
rect 1952 34128 2004 34134
rect 1952 34070 2004 34076
rect 2136 32768 2188 32774
rect 2136 32710 2188 32716
rect 2148 32434 2176 32710
rect 2136 32428 2188 32434
rect 2136 32370 2188 32376
rect 2148 31278 2176 32370
rect 2240 32230 2268 34138
rect 2332 32910 2360 36246
rect 2792 35086 2820 38762
rect 2872 38752 2924 38758
rect 2872 38694 2924 38700
rect 2884 36242 2912 38694
rect 2976 38350 3004 43046
rect 3068 42362 3096 44134
rect 3160 42566 3188 44814
rect 3804 44470 3832 45222
rect 4252 45076 4304 45082
rect 4252 45018 4304 45024
rect 4068 44872 4120 44878
rect 4068 44814 4120 44820
rect 3792 44464 3844 44470
rect 3792 44406 3844 44412
rect 4080 43994 4108 44814
rect 4264 44742 4292 45018
rect 4448 44946 4476 45222
rect 4436 44940 4488 44946
rect 4436 44882 4488 44888
rect 4252 44736 4304 44742
rect 4252 44678 4304 44684
rect 4264 44198 4292 44678
rect 4434 44568 4490 44577
rect 4434 44503 4436 44512
rect 4488 44503 4490 44512
rect 4436 44474 4488 44480
rect 4252 44192 4304 44198
rect 4252 44134 4304 44140
rect 4068 43988 4120 43994
rect 4068 43930 4120 43936
rect 3332 43920 3384 43926
rect 3332 43862 3384 43868
rect 3148 42560 3200 42566
rect 3148 42502 3200 42508
rect 3056 42356 3108 42362
rect 3056 42298 3108 42304
rect 3240 42220 3292 42226
rect 3240 42162 3292 42168
rect 3056 40044 3108 40050
rect 3056 39986 3108 39992
rect 3068 39642 3096 39986
rect 3056 39636 3108 39642
rect 3056 39578 3108 39584
rect 3252 39438 3280 42162
rect 3240 39432 3292 39438
rect 3240 39374 3292 39380
rect 3056 38956 3108 38962
rect 3056 38898 3108 38904
rect 2964 38344 3016 38350
rect 2964 38286 3016 38292
rect 2964 37120 3016 37126
rect 2964 37062 3016 37068
rect 2976 36582 3004 37062
rect 3068 36922 3096 38898
rect 3148 38208 3200 38214
rect 3148 38150 3200 38156
rect 3160 37913 3188 38150
rect 3146 37904 3202 37913
rect 3146 37839 3202 37848
rect 3252 37262 3280 39374
rect 3240 37256 3292 37262
rect 3146 37224 3202 37233
rect 3240 37198 3292 37204
rect 3344 37194 3372 43862
rect 3976 43784 4028 43790
rect 3976 43726 4028 43732
rect 3792 43648 3844 43654
rect 3792 43590 3844 43596
rect 3608 43308 3660 43314
rect 3608 43250 3660 43256
rect 3424 43104 3476 43110
rect 3424 43046 3476 43052
rect 3516 43104 3568 43110
rect 3516 43046 3568 43052
rect 3436 40186 3464 43046
rect 3528 41682 3556 43046
rect 3516 41676 3568 41682
rect 3516 41618 3568 41624
rect 3516 41064 3568 41070
rect 3516 41006 3568 41012
rect 3528 40633 3556 41006
rect 3514 40624 3570 40633
rect 3514 40559 3570 40568
rect 3424 40180 3476 40186
rect 3424 40122 3476 40128
rect 3620 39098 3648 43250
rect 3804 42770 3832 43590
rect 3884 43308 3936 43314
rect 3884 43250 3936 43256
rect 3792 42764 3844 42770
rect 3792 42706 3844 42712
rect 3700 42696 3752 42702
rect 3700 42638 3752 42644
rect 3712 42362 3740 42638
rect 3792 42560 3844 42566
rect 3792 42502 3844 42508
rect 3700 42356 3752 42362
rect 3700 42298 3752 42304
rect 3804 41682 3832 42502
rect 3792 41676 3844 41682
rect 3792 41618 3844 41624
rect 3792 41472 3844 41478
rect 3792 41414 3844 41420
rect 3804 41138 3832 41414
rect 3896 41274 3924 43250
rect 3988 41818 4016 43726
rect 4344 43308 4396 43314
rect 4344 43250 4396 43256
rect 4356 42022 4384 43250
rect 4540 42566 4568 45426
rect 4908 44538 4936 45426
rect 5356 44872 5408 44878
rect 5356 44814 5408 44820
rect 4896 44532 4948 44538
rect 4896 44474 4948 44480
rect 5368 44266 5396 44814
rect 5356 44260 5408 44266
rect 5356 44202 5408 44208
rect 5264 44192 5316 44198
rect 5264 44134 5316 44140
rect 5276 43994 5304 44134
rect 4988 43988 5040 43994
rect 4988 43930 5040 43936
rect 5264 43988 5316 43994
rect 5264 43930 5316 43936
rect 4528 42560 4580 42566
rect 4528 42502 4580 42508
rect 4712 42560 4764 42566
rect 4712 42502 4764 42508
rect 4344 42016 4396 42022
rect 4344 41958 4396 41964
rect 4724 41818 4752 42502
rect 4896 42016 4948 42022
rect 4896 41958 4948 41964
rect 3976 41812 4028 41818
rect 3976 41754 4028 41760
rect 4712 41812 4764 41818
rect 4712 41754 4764 41760
rect 4068 41540 4120 41546
rect 4068 41482 4120 41488
rect 4080 41274 4108 41482
rect 3884 41268 3936 41274
rect 3884 41210 3936 41216
rect 4068 41268 4120 41274
rect 4068 41210 4120 41216
rect 3700 41132 3752 41138
rect 3700 41074 3752 41080
rect 3792 41132 3844 41138
rect 3792 41074 3844 41080
rect 4344 41132 4396 41138
rect 4344 41074 4396 41080
rect 3712 40662 3740 41074
rect 4160 41064 4212 41070
rect 4160 41006 4212 41012
rect 3700 40656 3752 40662
rect 3700 40598 3752 40604
rect 3608 39092 3660 39098
rect 3608 39034 3660 39040
rect 3712 38978 3740 40598
rect 3976 40180 4028 40186
rect 3976 40122 4028 40128
rect 3792 40044 3844 40050
rect 3792 39986 3844 39992
rect 3804 39642 3832 39986
rect 3792 39636 3844 39642
rect 3792 39578 3844 39584
rect 3988 39438 4016 40122
rect 4172 39506 4200 41006
rect 4356 40730 4384 41074
rect 4528 40996 4580 41002
rect 4528 40938 4580 40944
rect 4436 40928 4488 40934
rect 4436 40870 4488 40876
rect 4344 40724 4396 40730
rect 4344 40666 4396 40672
rect 4250 40624 4306 40633
rect 4250 40559 4306 40568
rect 4160 39500 4212 39506
rect 4160 39442 4212 39448
rect 4264 39438 4292 40559
rect 4448 40526 4476 40870
rect 4436 40520 4488 40526
rect 4436 40462 4488 40468
rect 4344 39908 4396 39914
rect 4344 39850 4396 39856
rect 4356 39438 4384 39850
rect 4540 39438 4568 40938
rect 4802 40624 4858 40633
rect 4802 40559 4804 40568
rect 4856 40559 4858 40568
rect 4804 40530 4856 40536
rect 4712 40520 4764 40526
rect 4712 40462 4764 40468
rect 4724 39506 4752 40462
rect 4908 40118 4936 41958
rect 5000 41414 5028 43930
rect 5276 42906 5304 43930
rect 5368 43790 5396 44202
rect 5460 43994 5488 45426
rect 5915 45180 6223 45200
rect 5915 45178 5921 45180
rect 5977 45178 6001 45180
rect 6057 45178 6081 45180
rect 6137 45178 6161 45180
rect 6217 45178 6223 45180
rect 5977 45126 5979 45178
rect 6159 45126 6161 45178
rect 5915 45124 5921 45126
rect 5977 45124 6001 45126
rect 6057 45124 6081 45126
rect 6137 45124 6161 45126
rect 6217 45124 6223 45126
rect 5915 45104 6223 45124
rect 5724 44872 5776 44878
rect 5724 44814 5776 44820
rect 5540 44736 5592 44742
rect 5540 44678 5592 44684
rect 5448 43988 5500 43994
rect 5448 43930 5500 43936
rect 5356 43784 5408 43790
rect 5356 43726 5408 43732
rect 5264 42900 5316 42906
rect 5264 42842 5316 42848
rect 5080 42696 5132 42702
rect 5080 42638 5132 42644
rect 5092 42158 5120 42638
rect 5080 42152 5132 42158
rect 5080 42094 5132 42100
rect 5092 41682 5120 42094
rect 5080 41676 5132 41682
rect 5080 41618 5132 41624
rect 5000 41386 5120 41414
rect 4896 40112 4948 40118
rect 4896 40054 4948 40060
rect 4712 39500 4764 39506
rect 4712 39442 4764 39448
rect 3976 39432 4028 39438
rect 3976 39374 4028 39380
rect 4252 39432 4304 39438
rect 4252 39374 4304 39380
rect 4344 39432 4396 39438
rect 4344 39374 4396 39380
rect 4528 39432 4580 39438
rect 4528 39374 4580 39380
rect 3516 38956 3568 38962
rect 3516 38898 3568 38904
rect 3620 38950 3740 38978
rect 3976 38956 4028 38962
rect 3146 37159 3202 37168
rect 3332 37188 3384 37194
rect 3160 37126 3188 37159
rect 3332 37130 3384 37136
rect 3148 37120 3200 37126
rect 3148 37062 3200 37068
rect 3424 37120 3476 37126
rect 3424 37062 3476 37068
rect 3056 36916 3108 36922
rect 3056 36858 3108 36864
rect 3436 36786 3464 37062
rect 3424 36780 3476 36786
rect 3424 36722 3476 36728
rect 2964 36576 3016 36582
rect 2964 36518 3016 36524
rect 2872 36236 2924 36242
rect 2872 36178 2924 36184
rect 2964 36168 3016 36174
rect 2964 36110 3016 36116
rect 2872 36032 2924 36038
rect 2872 35974 2924 35980
rect 2780 35080 2832 35086
rect 2780 35022 2832 35028
rect 2884 33590 2912 35974
rect 2976 33946 3004 36110
rect 3148 36032 3200 36038
rect 3148 35974 3200 35980
rect 3056 34944 3108 34950
rect 3056 34886 3108 34892
rect 3068 34241 3096 34886
rect 3054 34232 3110 34241
rect 3054 34167 3110 34176
rect 3160 33998 3188 35974
rect 3240 35760 3292 35766
rect 3240 35702 3292 35708
rect 3148 33992 3200 33998
rect 2976 33918 3096 33946
rect 3148 33934 3200 33940
rect 2964 33856 3016 33862
rect 2964 33798 3016 33804
rect 2872 33584 2924 33590
rect 2976 33561 3004 33798
rect 2872 33526 2924 33532
rect 2962 33552 3018 33561
rect 2962 33487 3018 33496
rect 2320 32904 2372 32910
rect 2320 32846 2372 32852
rect 2596 32768 2648 32774
rect 2596 32710 2648 32716
rect 2228 32224 2280 32230
rect 2228 32166 2280 32172
rect 2240 31482 2268 32166
rect 2608 31822 2636 32710
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2792 32026 2820 32302
rect 3068 32230 3096 33918
rect 3252 33522 3280 35702
rect 3528 35290 3556 38898
rect 3516 35284 3568 35290
rect 3516 35226 3568 35232
rect 3620 35170 3648 38950
rect 3976 38898 4028 38904
rect 3792 38208 3844 38214
rect 3792 38150 3844 38156
rect 3804 37942 3832 38150
rect 3792 37936 3844 37942
rect 3792 37878 3844 37884
rect 3700 37800 3752 37806
rect 3700 37742 3752 37748
rect 3712 36922 3740 37742
rect 3792 37256 3844 37262
rect 3792 37198 3844 37204
rect 3804 36922 3832 37198
rect 3700 36916 3752 36922
rect 3700 36858 3752 36864
rect 3792 36916 3844 36922
rect 3792 36858 3844 36864
rect 3804 36174 3832 36858
rect 3988 36378 4016 38898
rect 4160 38752 4212 38758
rect 4160 38694 4212 38700
rect 4172 37874 4200 38694
rect 4264 38554 4292 39374
rect 4252 38548 4304 38554
rect 4252 38490 4304 38496
rect 4264 38350 4292 38490
rect 4252 38344 4304 38350
rect 4252 38286 4304 38292
rect 4160 37868 4212 37874
rect 4160 37810 4212 37816
rect 3976 36372 4028 36378
rect 3976 36314 4028 36320
rect 3792 36168 3844 36174
rect 3792 36110 3844 36116
rect 3976 36168 4028 36174
rect 3976 36110 4028 36116
rect 3792 35488 3844 35494
rect 3792 35430 3844 35436
rect 3436 35142 3648 35170
rect 3804 35154 3832 35430
rect 3792 35148 3844 35154
rect 3436 34610 3464 35142
rect 3792 35090 3844 35096
rect 3792 34944 3844 34950
rect 3792 34886 3844 34892
rect 3804 34610 3832 34886
rect 3424 34604 3476 34610
rect 3424 34546 3476 34552
rect 3516 34604 3568 34610
rect 3516 34546 3568 34552
rect 3792 34604 3844 34610
rect 3792 34546 3844 34552
rect 3240 33516 3292 33522
rect 3240 33458 3292 33464
rect 3252 32910 3280 33458
rect 3528 33386 3556 34546
rect 3608 34536 3660 34542
rect 3608 34478 3660 34484
rect 3620 33454 3648 34478
rect 3988 34202 4016 36110
rect 4068 35012 4120 35018
rect 4068 34954 4120 34960
rect 4080 34746 4108 34954
rect 4068 34740 4120 34746
rect 4068 34682 4120 34688
rect 3976 34196 4028 34202
rect 3976 34138 4028 34144
rect 3792 33992 3844 33998
rect 3792 33934 3844 33940
rect 3804 33658 3832 33934
rect 3884 33924 3936 33930
rect 3884 33866 3936 33872
rect 4160 33924 4212 33930
rect 4160 33866 4212 33872
rect 3792 33652 3844 33658
rect 3792 33594 3844 33600
rect 3896 33522 3924 33866
rect 3884 33516 3936 33522
rect 3884 33458 3936 33464
rect 4172 33454 4200 33866
rect 4356 33522 4384 39374
rect 4540 38654 4568 39374
rect 4540 38626 4660 38654
rect 4632 38350 4660 38626
rect 4724 38418 4752 39442
rect 5092 39438 5120 41386
rect 5172 40928 5224 40934
rect 5172 40870 5224 40876
rect 5184 40526 5212 40870
rect 5368 40526 5396 43726
rect 5552 43382 5580 44678
rect 5736 43450 5764 44814
rect 5816 44736 5868 44742
rect 5816 44678 5868 44684
rect 5828 43858 5856 44678
rect 5915 44092 6223 44112
rect 5915 44090 5921 44092
rect 5977 44090 6001 44092
rect 6057 44090 6081 44092
rect 6137 44090 6161 44092
rect 6217 44090 6223 44092
rect 5977 44038 5979 44090
rect 6159 44038 6161 44090
rect 5915 44036 5921 44038
rect 5977 44036 6001 44038
rect 6057 44036 6081 44038
rect 6137 44036 6161 44038
rect 6217 44036 6223 44038
rect 5915 44016 6223 44036
rect 5816 43852 5868 43858
rect 5816 43794 5868 43800
rect 5724 43444 5776 43450
rect 5724 43386 5776 43392
rect 5540 43376 5592 43382
rect 5540 43318 5592 43324
rect 5724 43308 5776 43314
rect 5724 43250 5776 43256
rect 5736 42702 5764 43250
rect 6472 43178 6500 45426
rect 6736 45280 6788 45286
rect 6736 45222 6788 45228
rect 6644 44872 6696 44878
rect 6644 44814 6696 44820
rect 6656 44538 6684 44814
rect 6644 44532 6696 44538
rect 6644 44474 6696 44480
rect 6748 44402 6776 45222
rect 7300 45082 7328 45426
rect 29000 45280 29052 45286
rect 29000 45222 29052 45228
rect 15846 45180 16154 45200
rect 15846 45178 15852 45180
rect 15908 45178 15932 45180
rect 15988 45178 16012 45180
rect 16068 45178 16092 45180
rect 16148 45178 16154 45180
rect 15908 45126 15910 45178
rect 16090 45126 16092 45178
rect 15846 45124 15852 45126
rect 15908 45124 15932 45126
rect 15988 45124 16012 45126
rect 16068 45124 16092 45126
rect 16148 45124 16154 45126
rect 15846 45104 16154 45124
rect 25776 45180 26084 45200
rect 25776 45178 25782 45180
rect 25838 45178 25862 45180
rect 25918 45178 25942 45180
rect 25998 45178 26022 45180
rect 26078 45178 26084 45180
rect 25838 45126 25840 45178
rect 26020 45126 26022 45178
rect 25776 45124 25782 45126
rect 25838 45124 25862 45126
rect 25918 45124 25942 45126
rect 25998 45124 26022 45126
rect 26078 45124 26084 45126
rect 25776 45104 26084 45124
rect 7288 45076 7340 45082
rect 7288 45018 7340 45024
rect 7380 45008 7432 45014
rect 7380 44950 7432 44956
rect 7196 44872 7248 44878
rect 7196 44814 7248 44820
rect 6828 44736 6880 44742
rect 6828 44678 6880 44684
rect 6840 44470 6868 44678
rect 7208 44470 7236 44814
rect 6828 44464 6880 44470
rect 6828 44406 6880 44412
rect 7196 44464 7248 44470
rect 7196 44406 7248 44412
rect 6736 44396 6788 44402
rect 6736 44338 6788 44344
rect 6644 43716 6696 43722
rect 6644 43658 6696 43664
rect 6460 43172 6512 43178
rect 6460 43114 6512 43120
rect 5915 43004 6223 43024
rect 5915 43002 5921 43004
rect 5977 43002 6001 43004
rect 6057 43002 6081 43004
rect 6137 43002 6161 43004
rect 6217 43002 6223 43004
rect 5977 42950 5979 43002
rect 6159 42950 6161 43002
rect 5915 42948 5921 42950
rect 5977 42948 6001 42950
rect 6057 42948 6081 42950
rect 6137 42948 6161 42950
rect 6217 42948 6223 42950
rect 5915 42928 6223 42948
rect 6656 42906 6684 43658
rect 6828 43648 6880 43654
rect 6828 43590 6880 43596
rect 6644 42900 6696 42906
rect 6644 42842 6696 42848
rect 6840 42702 6868 43590
rect 7012 43240 7064 43246
rect 7012 43182 7064 43188
rect 5724 42696 5776 42702
rect 5724 42638 5776 42644
rect 6828 42696 6880 42702
rect 6828 42638 6880 42644
rect 5736 42226 5764 42638
rect 7024 42634 7052 43182
rect 7208 43178 7236 44406
rect 7392 43314 7420 44950
rect 7472 44872 7524 44878
rect 8208 44872 8260 44878
rect 7472 44814 7524 44820
rect 8022 44840 8078 44849
rect 7380 43308 7432 43314
rect 7380 43250 7432 43256
rect 7196 43172 7248 43178
rect 7196 43114 7248 43120
rect 7208 42838 7236 43114
rect 7196 42832 7248 42838
rect 7196 42774 7248 42780
rect 6736 42628 6788 42634
rect 6736 42570 6788 42576
rect 7012 42628 7064 42634
rect 7012 42570 7064 42576
rect 6552 42560 6604 42566
rect 6552 42502 6604 42508
rect 5724 42220 5776 42226
rect 5724 42162 5776 42168
rect 6460 42220 6512 42226
rect 6460 42162 6512 42168
rect 5632 41608 5684 41614
rect 5632 41550 5684 41556
rect 5644 40594 5672 41550
rect 5632 40588 5684 40594
rect 5632 40530 5684 40536
rect 5172 40520 5224 40526
rect 5172 40462 5224 40468
rect 5356 40520 5408 40526
rect 5356 40462 5408 40468
rect 5632 40044 5684 40050
rect 5632 39986 5684 39992
rect 5644 39642 5672 39986
rect 5632 39636 5684 39642
rect 5632 39578 5684 39584
rect 5736 39438 5764 42162
rect 5915 41916 6223 41936
rect 5915 41914 5921 41916
rect 5977 41914 6001 41916
rect 6057 41914 6081 41916
rect 6137 41914 6161 41916
rect 6217 41914 6223 41916
rect 5977 41862 5979 41914
rect 6159 41862 6161 41914
rect 5915 41860 5921 41862
rect 5977 41860 6001 41862
rect 6057 41860 6081 41862
rect 6137 41860 6161 41862
rect 6217 41860 6223 41862
rect 5915 41840 6223 41860
rect 6276 41540 6328 41546
rect 6276 41482 6328 41488
rect 5816 41064 5868 41070
rect 5816 41006 5868 41012
rect 5828 40186 5856 41006
rect 5915 40828 6223 40848
rect 5915 40826 5921 40828
rect 5977 40826 6001 40828
rect 6057 40826 6081 40828
rect 6137 40826 6161 40828
rect 6217 40826 6223 40828
rect 5977 40774 5979 40826
rect 6159 40774 6161 40826
rect 5915 40772 5921 40774
rect 5977 40772 6001 40774
rect 6057 40772 6081 40774
rect 6137 40772 6161 40774
rect 6217 40772 6223 40774
rect 5915 40752 6223 40772
rect 6288 40610 6316 41482
rect 6288 40582 6408 40610
rect 6276 40520 6328 40526
rect 6276 40462 6328 40468
rect 5816 40180 5868 40186
rect 5816 40122 5868 40128
rect 5816 39840 5868 39846
rect 5816 39782 5868 39788
rect 5080 39432 5132 39438
rect 5080 39374 5132 39380
rect 5724 39432 5776 39438
rect 5724 39374 5776 39380
rect 4712 38412 4764 38418
rect 4712 38354 4764 38360
rect 4620 38344 4672 38350
rect 4620 38286 4672 38292
rect 4528 38208 4580 38214
rect 4528 38150 4580 38156
rect 4436 37868 4488 37874
rect 4436 37810 4488 37816
rect 4448 36854 4476 37810
rect 4436 36848 4488 36854
rect 4436 36790 4488 36796
rect 4540 36718 4568 38150
rect 4632 37330 4660 38286
rect 4620 37324 4672 37330
rect 4620 37266 4672 37272
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 4632 36786 4660 37062
rect 4620 36780 4672 36786
rect 4620 36722 4672 36728
rect 4528 36712 4580 36718
rect 4528 36654 4580 36660
rect 4724 36650 4752 38354
rect 4896 38276 4948 38282
rect 4896 38218 4948 38224
rect 4804 37324 4856 37330
rect 4804 37266 4856 37272
rect 4816 36786 4844 37266
rect 4804 36780 4856 36786
rect 4804 36722 4856 36728
rect 4712 36644 4764 36650
rect 4712 36586 4764 36592
rect 4908 36530 4936 38218
rect 4988 37120 5040 37126
rect 4988 37062 5040 37068
rect 4632 36502 4936 36530
rect 4436 35080 4488 35086
rect 4436 35022 4488 35028
rect 4448 34746 4476 35022
rect 4436 34740 4488 34746
rect 4436 34682 4488 34688
rect 4528 34536 4580 34542
rect 4528 34478 4580 34484
rect 4436 33992 4488 33998
rect 4436 33934 4488 33940
rect 4344 33516 4396 33522
rect 4344 33458 4396 33464
rect 3608 33448 3660 33454
rect 3608 33390 3660 33396
rect 4160 33448 4212 33454
rect 4160 33390 4212 33396
rect 3516 33380 3568 33386
rect 3516 33322 3568 33328
rect 3240 32904 3292 32910
rect 3240 32846 3292 32852
rect 4068 32904 4120 32910
rect 4068 32846 4120 32852
rect 3976 32564 4028 32570
rect 3976 32506 4028 32512
rect 3700 32428 3752 32434
rect 3700 32370 3752 32376
rect 3056 32224 3108 32230
rect 3056 32166 3108 32172
rect 3712 32026 3740 32370
rect 2780 32020 2832 32026
rect 2780 31962 2832 31968
rect 3700 32020 3752 32026
rect 3700 31962 3752 31968
rect 3056 31884 3108 31890
rect 3056 31826 3108 31832
rect 2596 31816 2648 31822
rect 2596 31758 2648 31764
rect 2228 31476 2280 31482
rect 2228 31418 2280 31424
rect 2136 31272 2188 31278
rect 2136 31214 2188 31220
rect 2148 30870 2176 31214
rect 2320 31136 2372 31142
rect 2320 31078 2372 31084
rect 2332 30938 2360 31078
rect 3068 30938 3096 31826
rect 3988 31822 4016 32506
rect 3976 31816 4028 31822
rect 3976 31758 4028 31764
rect 3240 31476 3292 31482
rect 3240 31418 3292 31424
rect 3884 31476 3936 31482
rect 3884 31418 3936 31424
rect 3252 31346 3280 31418
rect 3240 31340 3292 31346
rect 3240 31282 3292 31288
rect 3700 31136 3752 31142
rect 3700 31078 3752 31084
rect 2320 30932 2372 30938
rect 2320 30874 2372 30880
rect 3056 30932 3108 30938
rect 3056 30874 3108 30880
rect 2136 30864 2188 30870
rect 2136 30806 2188 30812
rect 2148 30258 2176 30806
rect 2136 30252 2188 30258
rect 2136 30194 2188 30200
rect 2148 29782 2176 30194
rect 2332 30054 2360 30874
rect 2964 30728 3016 30734
rect 2964 30670 3016 30676
rect 2320 30048 2372 30054
rect 2320 29990 2372 29996
rect 2504 30048 2556 30054
rect 2504 29990 2556 29996
rect 2332 29850 2360 29990
rect 2320 29844 2372 29850
rect 2320 29786 2372 29792
rect 2136 29776 2188 29782
rect 2136 29718 2188 29724
rect 2516 29714 2544 29990
rect 2778 29880 2834 29889
rect 2976 29850 3004 30670
rect 3712 30326 3740 31078
rect 3700 30320 3752 30326
rect 3700 30262 3752 30268
rect 3240 30184 3292 30190
rect 3240 30126 3292 30132
rect 2778 29815 2834 29824
rect 2964 29844 3016 29850
rect 2504 29708 2556 29714
rect 2504 29650 2556 29656
rect 2136 29504 2188 29510
rect 2136 29446 2188 29452
rect 2148 29170 2176 29446
rect 2792 29306 2820 29815
rect 2964 29786 3016 29792
rect 2872 29776 2924 29782
rect 2872 29718 2924 29724
rect 2780 29300 2832 29306
rect 2780 29242 2832 29248
rect 2136 29164 2188 29170
rect 2136 29106 2188 29112
rect 1596 28580 1716 28608
rect 1492 28416 1544 28422
rect 1490 28384 1492 28393
rect 1544 28384 1546 28393
rect 1490 28319 1546 28328
rect 1492 27872 1544 27878
rect 1492 27814 1544 27820
rect 1504 27577 1532 27814
rect 1490 27568 1546 27577
rect 1490 27503 1546 27512
rect 1490 26888 1546 26897
rect 1490 26823 1492 26832
rect 1544 26823 1546 26832
rect 1492 26794 1544 26800
rect 1492 26240 1544 26246
rect 1490 26208 1492 26217
rect 1544 26208 1546 26217
rect 1490 26143 1546 26152
rect 1492 25696 1544 25702
rect 1492 25638 1544 25644
rect 1504 25401 1532 25638
rect 1490 25392 1546 25401
rect 1490 25327 1546 25336
rect 1490 24712 1546 24721
rect 1490 24647 1492 24656
rect 1544 24647 1546 24656
rect 1492 24618 1544 24624
rect 1492 24064 1544 24070
rect 1492 24006 1544 24012
rect 1504 23905 1532 24006
rect 1490 23896 1546 23905
rect 1490 23831 1546 23840
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1412 23225 1440 23598
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 1596 22522 1624 28580
rect 2596 28552 2648 28558
rect 2596 28494 2648 28500
rect 2136 28484 2188 28490
rect 2136 28426 2188 28432
rect 2148 28082 2176 28426
rect 2136 28076 2188 28082
rect 2136 28018 2188 28024
rect 2608 28014 2636 28494
rect 2596 28008 2648 28014
rect 2596 27950 2648 27956
rect 2608 27470 2636 27950
rect 2884 27878 2912 29718
rect 3252 29306 3280 30126
rect 3608 29504 3660 29510
rect 3608 29446 3660 29452
rect 3240 29300 3292 29306
rect 3240 29242 3292 29248
rect 3620 29170 3648 29446
rect 3608 29164 3660 29170
rect 3608 29106 3660 29112
rect 3792 28960 3844 28966
rect 3792 28902 3844 28908
rect 3804 28558 3832 28902
rect 3792 28552 3844 28558
rect 3792 28494 3844 28500
rect 3896 28150 3924 31418
rect 3976 30592 4028 30598
rect 3974 30560 3976 30569
rect 4028 30560 4030 30569
rect 3974 30495 4030 30504
rect 3976 29640 4028 29646
rect 4080 29628 4108 32846
rect 4172 31890 4200 33390
rect 4344 33380 4396 33386
rect 4448 33368 4476 33934
rect 4540 33522 4568 34478
rect 4528 33516 4580 33522
rect 4528 33458 4580 33464
rect 4396 33340 4476 33368
rect 4344 33322 4396 33328
rect 4252 32768 4304 32774
rect 4252 32710 4304 32716
rect 4264 32026 4292 32710
rect 4252 32020 4304 32026
rect 4252 31962 4304 31968
rect 4160 31884 4212 31890
rect 4160 31826 4212 31832
rect 4172 31414 4200 31826
rect 4252 31816 4304 31822
rect 4356 31804 4384 33322
rect 4540 32434 4568 33458
rect 4632 33046 4660 36502
rect 4896 35488 4948 35494
rect 4896 35430 4948 35436
rect 4712 34672 4764 34678
rect 4712 34614 4764 34620
rect 4724 33114 4752 34614
rect 4712 33108 4764 33114
rect 4712 33050 4764 33056
rect 4620 33040 4672 33046
rect 4620 32982 4672 32988
rect 4528 32428 4580 32434
rect 4528 32370 4580 32376
rect 4540 31822 4568 32370
rect 4632 31822 4660 32982
rect 4908 32910 4936 35430
rect 4896 32904 4948 32910
rect 4896 32846 4948 32852
rect 4304 31776 4384 31804
rect 4252 31758 4304 31764
rect 4160 31408 4212 31414
rect 4160 31350 4212 31356
rect 4356 31278 4384 31776
rect 4528 31816 4580 31822
rect 4528 31758 4580 31764
rect 4620 31816 4672 31822
rect 4620 31758 4672 31764
rect 4540 31346 4568 31758
rect 5000 31754 5028 37062
rect 4988 31748 5040 31754
rect 4988 31690 5040 31696
rect 5000 31414 5028 31690
rect 5092 31482 5120 39374
rect 5736 39098 5764 39374
rect 5724 39092 5776 39098
rect 5724 39034 5776 39040
rect 5828 38962 5856 39782
rect 5915 39740 6223 39760
rect 5915 39738 5921 39740
rect 5977 39738 6001 39740
rect 6057 39738 6081 39740
rect 6137 39738 6161 39740
rect 6217 39738 6223 39740
rect 5977 39686 5979 39738
rect 6159 39686 6161 39738
rect 5915 39684 5921 39686
rect 5977 39684 6001 39686
rect 6057 39684 6081 39686
rect 6137 39684 6161 39686
rect 6217 39684 6223 39686
rect 5915 39664 6223 39684
rect 5632 38956 5684 38962
rect 5632 38898 5684 38904
rect 5816 38956 5868 38962
rect 5816 38898 5868 38904
rect 5644 38282 5672 38898
rect 5915 38652 6223 38672
rect 5915 38650 5921 38652
rect 5977 38650 6001 38652
rect 6057 38650 6081 38652
rect 6137 38650 6161 38652
rect 6217 38650 6223 38652
rect 5977 38598 5979 38650
rect 6159 38598 6161 38650
rect 5915 38596 5921 38598
rect 5977 38596 6001 38598
rect 6057 38596 6081 38598
rect 6137 38596 6161 38598
rect 6217 38596 6223 38598
rect 5915 38576 6223 38596
rect 5632 38276 5684 38282
rect 5632 38218 5684 38224
rect 5632 37732 5684 37738
rect 5632 37674 5684 37680
rect 5540 37664 5592 37670
rect 5540 37606 5592 37612
rect 5552 36854 5580 37606
rect 5644 37330 5672 37674
rect 5915 37564 6223 37584
rect 5915 37562 5921 37564
rect 5977 37562 6001 37564
rect 6057 37562 6081 37564
rect 6137 37562 6161 37564
rect 6217 37562 6223 37564
rect 5977 37510 5979 37562
rect 6159 37510 6161 37562
rect 5915 37508 5921 37510
rect 5977 37508 6001 37510
rect 6057 37508 6081 37510
rect 6137 37508 6161 37510
rect 6217 37508 6223 37510
rect 5915 37488 6223 37508
rect 5632 37324 5684 37330
rect 5632 37266 5684 37272
rect 5816 37324 5868 37330
rect 5816 37266 5868 37272
rect 5724 37256 5776 37262
rect 5724 37198 5776 37204
rect 5540 36848 5592 36854
rect 5540 36790 5592 36796
rect 5632 36780 5684 36786
rect 5632 36722 5684 36728
rect 5540 36168 5592 36174
rect 5540 36110 5592 36116
rect 5552 35834 5580 36110
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 5540 35692 5592 35698
rect 5540 35634 5592 35640
rect 5172 33856 5224 33862
rect 5172 33798 5224 33804
rect 5184 33590 5212 33798
rect 5552 33658 5580 35634
rect 5644 35290 5672 36722
rect 5736 36378 5764 37198
rect 5724 36372 5776 36378
rect 5724 36314 5776 36320
rect 5632 35284 5684 35290
rect 5632 35226 5684 35232
rect 5828 35170 5856 37266
rect 5915 36476 6223 36496
rect 5915 36474 5921 36476
rect 5977 36474 6001 36476
rect 6057 36474 6081 36476
rect 6137 36474 6161 36476
rect 6217 36474 6223 36476
rect 5977 36422 5979 36474
rect 6159 36422 6161 36474
rect 5915 36420 5921 36422
rect 5977 36420 6001 36422
rect 6057 36420 6081 36422
rect 6137 36420 6161 36422
rect 6217 36420 6223 36422
rect 5915 36400 6223 36420
rect 6288 35494 6316 40462
rect 6380 37874 6408 40582
rect 6472 40050 6500 42162
rect 6564 41614 6592 42502
rect 6552 41608 6604 41614
rect 6552 41550 6604 41556
rect 6748 41274 6776 42570
rect 7024 42158 7052 42570
rect 7208 42158 7236 42774
rect 7392 42702 7420 43250
rect 7380 42696 7432 42702
rect 7380 42638 7432 42644
rect 7288 42356 7340 42362
rect 7288 42298 7340 42304
rect 7012 42152 7064 42158
rect 7012 42094 7064 42100
rect 7196 42152 7248 42158
rect 7196 42094 7248 42100
rect 6920 42016 6972 42022
rect 6920 41958 6972 41964
rect 6736 41268 6788 41274
rect 6736 41210 6788 41216
rect 6552 40520 6604 40526
rect 6552 40462 6604 40468
rect 6460 40044 6512 40050
rect 6460 39986 6512 39992
rect 6472 39370 6500 39986
rect 6460 39364 6512 39370
rect 6460 39306 6512 39312
rect 6368 37868 6420 37874
rect 6368 37810 6420 37816
rect 6380 37754 6408 37810
rect 6380 37726 6500 37754
rect 6368 37664 6420 37670
rect 6368 37606 6420 37612
rect 6380 37262 6408 37606
rect 6472 37466 6500 37726
rect 6460 37460 6512 37466
rect 6460 37402 6512 37408
rect 6368 37256 6420 37262
rect 6368 37198 6420 37204
rect 6564 36174 6592 40462
rect 6748 40118 6776 41210
rect 6736 40112 6788 40118
rect 6736 40054 6788 40060
rect 6644 39976 6696 39982
rect 6644 39918 6696 39924
rect 6656 39438 6684 39918
rect 6932 39438 6960 41958
rect 7024 41274 7052 42094
rect 7012 41268 7064 41274
rect 7012 41210 7064 41216
rect 7104 41132 7156 41138
rect 7104 41074 7156 41080
rect 7012 40520 7064 40526
rect 7012 40462 7064 40468
rect 7024 39982 7052 40462
rect 7116 40050 7144 41074
rect 7208 40594 7236 42094
rect 7196 40588 7248 40594
rect 7196 40530 7248 40536
rect 7104 40044 7156 40050
rect 7104 39986 7156 39992
rect 7012 39976 7064 39982
rect 7012 39918 7064 39924
rect 7024 39506 7052 39918
rect 7012 39500 7064 39506
rect 7012 39442 7064 39448
rect 6644 39432 6696 39438
rect 6644 39374 6696 39380
rect 6920 39432 6972 39438
rect 6920 39374 6972 39380
rect 6656 39302 6684 39374
rect 6828 39364 6880 39370
rect 6828 39306 6880 39312
rect 6644 39296 6696 39302
rect 6644 39238 6696 39244
rect 6656 37806 6684 39238
rect 6736 38752 6788 38758
rect 6736 38694 6788 38700
rect 6748 38418 6776 38694
rect 6736 38412 6788 38418
rect 6736 38354 6788 38360
rect 6644 37800 6696 37806
rect 6644 37742 6696 37748
rect 6840 37482 6868 39306
rect 6932 39098 6960 39374
rect 6920 39092 6972 39098
rect 6920 39034 6972 39040
rect 7024 37942 7052 39442
rect 7104 39296 7156 39302
rect 7104 39238 7156 39244
rect 7116 38962 7144 39238
rect 7104 38956 7156 38962
rect 7104 38898 7156 38904
rect 7012 37936 7064 37942
rect 7012 37878 7064 37884
rect 7104 37868 7156 37874
rect 7104 37810 7156 37816
rect 7116 37482 7144 37810
rect 6748 37454 7144 37482
rect 6552 36168 6604 36174
rect 6552 36110 6604 36116
rect 6276 35488 6328 35494
rect 6276 35430 6328 35436
rect 5915 35388 6223 35408
rect 5915 35386 5921 35388
rect 5977 35386 6001 35388
rect 6057 35386 6081 35388
rect 6137 35386 6161 35388
rect 6217 35386 6223 35388
rect 5977 35334 5979 35386
rect 6159 35334 6161 35386
rect 5915 35332 5921 35334
rect 5977 35332 6001 35334
rect 6057 35332 6081 35334
rect 6137 35332 6161 35334
rect 6217 35332 6223 35334
rect 5915 35312 6223 35332
rect 5644 35142 5856 35170
rect 5540 33652 5592 33658
rect 5540 33594 5592 33600
rect 5172 33584 5224 33590
rect 5172 33526 5224 33532
rect 5080 31476 5132 31482
rect 5080 31418 5132 31424
rect 4988 31408 5040 31414
rect 4988 31350 5040 31356
rect 5264 31408 5316 31414
rect 5264 31350 5316 31356
rect 4528 31340 4580 31346
rect 4528 31282 4580 31288
rect 4344 31272 4396 31278
rect 4344 31214 4396 31220
rect 4620 31204 4672 31210
rect 4620 31146 4672 31152
rect 4632 30394 4660 31146
rect 5276 30734 5304 31350
rect 5356 31340 5408 31346
rect 5356 31282 5408 31288
rect 5368 30734 5396 31282
rect 4896 30728 4948 30734
rect 4896 30670 4948 30676
rect 5264 30728 5316 30734
rect 5264 30670 5316 30676
rect 5356 30728 5408 30734
rect 5356 30670 5408 30676
rect 4712 30592 4764 30598
rect 4712 30534 4764 30540
rect 4620 30388 4672 30394
rect 4620 30330 4672 30336
rect 4724 29646 4752 30534
rect 4028 29600 4108 29628
rect 3976 29582 4028 29588
rect 4080 29170 4108 29600
rect 4160 29640 4212 29646
rect 4160 29582 4212 29588
rect 4712 29640 4764 29646
rect 4712 29582 4764 29588
rect 4068 29164 4120 29170
rect 4068 29106 4120 29112
rect 4172 28762 4200 29582
rect 4908 29578 4936 30670
rect 5264 29640 5316 29646
rect 5264 29582 5316 29588
rect 4896 29572 4948 29578
rect 4896 29514 4948 29520
rect 5276 29306 5304 29582
rect 5264 29300 5316 29306
rect 5264 29242 5316 29248
rect 4712 29096 4764 29102
rect 4712 29038 4764 29044
rect 5540 29096 5592 29102
rect 5540 29038 5592 29044
rect 4160 28756 4212 28762
rect 4160 28698 4212 28704
rect 4724 28218 4752 29038
rect 5552 28762 5580 29038
rect 5540 28756 5592 28762
rect 5540 28698 5592 28704
rect 4988 28552 5040 28558
rect 4988 28494 5040 28500
rect 5000 28218 5028 28494
rect 4712 28212 4764 28218
rect 4712 28154 4764 28160
rect 4988 28212 5040 28218
rect 4988 28154 5040 28160
rect 3884 28144 3936 28150
rect 3884 28086 3936 28092
rect 5356 28144 5408 28150
rect 5356 28086 5408 28092
rect 2872 27872 2924 27878
rect 2872 27814 2924 27820
rect 3700 27872 3752 27878
rect 3700 27814 3752 27820
rect 2596 27464 2648 27470
rect 2596 27406 2648 27412
rect 1676 27328 1728 27334
rect 1676 27270 1728 27276
rect 1688 26994 1716 27270
rect 1676 26988 1728 26994
rect 1676 26930 1728 26936
rect 2608 26382 2636 27406
rect 3608 26988 3660 26994
rect 3608 26930 3660 26936
rect 2596 26376 2648 26382
rect 2596 26318 2648 26324
rect 2608 26234 2636 26318
rect 2964 26308 3016 26314
rect 2964 26250 3016 26256
rect 2780 26240 2832 26246
rect 2608 26206 2728 26234
rect 2700 25906 2728 26206
rect 2780 26182 2832 26188
rect 2688 25900 2740 25906
rect 2688 25842 2740 25848
rect 2700 24818 2728 25842
rect 2792 25838 2820 26182
rect 2976 26042 3004 26250
rect 3620 26042 3648 26930
rect 2964 26036 3016 26042
rect 2964 25978 3016 25984
rect 3608 26036 3660 26042
rect 3608 25978 3660 25984
rect 2780 25832 2832 25838
rect 2780 25774 2832 25780
rect 2688 24812 2740 24818
rect 2688 24754 2740 24760
rect 2700 24206 2728 24754
rect 2688 24200 2740 24206
rect 2688 24142 2740 24148
rect 3516 24132 3568 24138
rect 3516 24074 3568 24080
rect 2872 23792 2924 23798
rect 2872 23734 2924 23740
rect 2320 23656 2372 23662
rect 2320 23598 2372 23604
rect 2044 23112 2096 23118
rect 2044 23054 2096 23060
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1504 22494 1624 22522
rect 1400 20800 1452 20806
rect 1400 20742 1452 20748
rect 1412 20466 1440 20742
rect 1400 20460 1452 20466
rect 1400 20402 1452 20408
rect 1308 19508 1360 19514
rect 1308 19450 1360 19456
rect 1216 16584 1268 16590
rect 1216 16526 1268 16532
rect 1228 14385 1256 16526
rect 1214 14376 1270 14385
rect 1214 14311 1270 14320
rect 1216 12232 1268 12238
rect 1216 12174 1268 12180
rect 1228 11393 1256 12174
rect 1214 11384 1270 11393
rect 1214 11319 1270 11328
rect 1214 5536 1270 5545
rect 1214 5471 1270 5480
rect 1228 4690 1256 5471
rect 1216 4684 1268 4690
rect 1216 4626 1268 4632
rect 1320 2774 1348 19450
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 1412 15881 1440 17138
rect 1398 15872 1454 15881
rect 1398 15807 1454 15816
rect 1504 15162 1532 22494
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 18766 1624 22374
rect 1688 20466 1716 22918
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 1768 22432 1820 22438
rect 1768 22374 1820 22380
rect 1780 20942 1808 22374
rect 1872 21049 1900 22578
rect 2056 22409 2084 23054
rect 2042 22400 2098 22409
rect 2042 22335 2098 22344
rect 2136 21956 2188 21962
rect 2136 21898 2188 21904
rect 1858 21040 1914 21049
rect 1858 20975 1914 20984
rect 1952 21004 2004 21010
rect 1952 20946 2004 20952
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1872 20534 1900 20878
rect 1860 20528 1912 20534
rect 1860 20470 1912 20476
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 1872 20346 1900 20470
rect 1964 20398 1992 20946
rect 2148 20602 2176 21898
rect 2228 21548 2280 21554
rect 2228 21490 2280 21496
rect 2240 21146 2268 21490
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 2136 20596 2188 20602
rect 2136 20538 2188 20544
rect 1780 20318 1900 20346
rect 1952 20392 2004 20398
rect 1952 20334 2004 20340
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 19242 1716 19654
rect 1676 19236 1728 19242
rect 1676 19178 1728 19184
rect 1676 18896 1728 18902
rect 1676 18838 1728 18844
rect 1584 18760 1636 18766
rect 1584 18702 1636 18708
rect 1688 18290 1716 18838
rect 1780 18834 1808 20318
rect 1860 20256 1912 20262
rect 1860 20198 1912 20204
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1676 18284 1728 18290
rect 1676 18226 1728 18232
rect 1780 18222 1808 18770
rect 1872 18290 1900 20198
rect 1964 18834 1992 20334
rect 2228 19780 2280 19786
rect 2228 19722 2280 19728
rect 2240 18970 2268 19722
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2332 18850 2360 23598
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2792 20233 2820 22986
rect 2884 22030 2912 23734
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 2872 22024 2924 22030
rect 2872 21966 2924 21972
rect 2884 21622 2912 21966
rect 2976 21729 3004 22578
rect 3148 22568 3200 22574
rect 3148 22510 3200 22516
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 2962 21720 3018 21729
rect 2962 21655 3018 21664
rect 2872 21616 2924 21622
rect 2872 21558 2924 21564
rect 2778 20224 2834 20233
rect 2778 20159 2834 20168
rect 2884 19854 2912 21558
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2976 20942 3004 21286
rect 3068 20942 3096 21830
rect 2964 20936 3016 20942
rect 2964 20878 3016 20884
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 3068 20534 3096 20878
rect 3056 20528 3108 20534
rect 3056 20470 3108 20476
rect 2964 20460 3016 20466
rect 2964 20402 3016 20408
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2884 19378 2912 19790
rect 2504 19372 2556 19378
rect 2504 19314 2556 19320
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 2240 18822 2360 18850
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1688 16046 1716 17614
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 13569 1440 14350
rect 1504 13938 1532 14758
rect 1688 14074 1716 15982
rect 1780 15706 1808 16050
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1964 15502 1992 15846
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 1780 14074 1808 14962
rect 2148 14618 2176 14962
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1398 13560 1454 13569
rect 1398 13495 1454 13504
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 12889 1440 13262
rect 1398 12880 1454 12889
rect 1398 12815 1454 12824
rect 1400 12708 1452 12714
rect 1400 12650 1452 12656
rect 1412 12073 1440 12650
rect 1398 12064 1454 12073
rect 1398 11999 1454 12008
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1412 10713 1440 11698
rect 2240 11626 2268 18822
rect 2516 18426 2544 19314
rect 2596 19168 2648 19174
rect 2872 19168 2924 19174
rect 2648 19116 2820 19122
rect 2596 19110 2820 19116
rect 2872 19110 2924 19116
rect 2608 19094 2820 19110
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2596 18148 2648 18154
rect 2596 18090 2648 18096
rect 2608 17202 2636 18090
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 2332 15502 2360 16934
rect 2792 16561 2820 19094
rect 2884 18290 2912 19110
rect 2976 18737 3004 20402
rect 3160 19553 3188 22510
rect 3332 20868 3384 20874
rect 3332 20810 3384 20816
rect 3240 19984 3292 19990
rect 3240 19926 3292 19932
rect 3146 19544 3202 19553
rect 3146 19479 3202 19488
rect 3252 18766 3280 19926
rect 3344 18902 3372 20810
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3332 18896 3384 18902
rect 3332 18838 3384 18844
rect 3240 18760 3292 18766
rect 2962 18728 3018 18737
rect 3240 18702 3292 18708
rect 2962 18663 3018 18672
rect 3332 18692 3384 18698
rect 3332 18634 3384 18640
rect 3056 18624 3108 18630
rect 3108 18584 3188 18612
rect 3056 18566 3108 18572
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2884 17678 2912 18022
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2976 17542 3004 18226
rect 3160 18222 3188 18584
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2976 16794 3004 17478
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2872 16584 2924 16590
rect 2778 16552 2834 16561
rect 2872 16526 2924 16532
rect 2778 16487 2834 16496
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2516 14414 2544 14962
rect 2700 14414 2728 16390
rect 2884 16046 2912 16526
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2792 15026 2820 15506
rect 2884 15434 2912 15982
rect 3160 15638 3188 18158
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 3252 16590 3280 17070
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3252 16289 3280 16526
rect 3344 16436 3372 18634
rect 3436 16590 3464 19654
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 3344 16408 3464 16436
rect 3238 16280 3294 16289
rect 3238 16215 3294 16224
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 2872 15428 2924 15434
rect 2872 15370 2924 15376
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 2884 14958 2912 15370
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2976 15026 3004 15302
rect 3056 15088 3108 15094
rect 3160 15065 3188 15438
rect 3056 15030 3108 15036
rect 3146 15056 3202 15065
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2516 13326 2544 14350
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2516 12238 2544 13262
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2700 12238 2728 13126
rect 2792 12850 2820 14758
rect 2884 14550 2912 14894
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2964 14408 3016 14414
rect 3068 14396 3096 15030
rect 3146 14991 3202 15000
rect 3252 14940 3280 16215
rect 3016 14368 3096 14396
rect 2964 14350 3016 14356
rect 3068 13938 3096 14368
rect 3160 14912 3280 14940
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2792 12730 2820 12786
rect 2792 12702 2912 12730
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2516 11830 2544 12174
rect 2504 11824 2556 11830
rect 2504 11766 2556 11772
rect 2792 11762 2820 12582
rect 2884 12170 2912 12702
rect 3068 12374 3096 13874
rect 3160 12850 3188 14912
rect 3436 13870 3464 16408
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2884 11694 2912 12106
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2228 11620 2280 11626
rect 2228 11562 2280 11568
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1398 10704 1454 10713
rect 1596 10674 1624 11494
rect 2884 11370 2912 11630
rect 2976 11558 3004 12038
rect 3068 11762 3096 12310
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2792 11342 2912 11370
rect 2792 11234 2820 11342
rect 2700 11206 2820 11234
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 1768 11008 1820 11014
rect 1768 10950 1820 10956
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 1398 10639 1454 10648
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1780 10606 1808 10950
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1504 10198 1532 10542
rect 1492 10192 1544 10198
rect 1492 10134 1544 10140
rect 2056 10062 2084 10950
rect 2148 10742 2176 11018
rect 2136 10736 2188 10742
rect 2136 10678 2188 10684
rect 2700 10606 2728 11206
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2792 10674 2820 11086
rect 2976 10810 3004 11222
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 9217 1440 9522
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 8401 1440 8910
rect 1398 8392 1454 8401
rect 1398 8327 1454 8336
rect 1398 7712 1454 7721
rect 1398 7647 1454 7656
rect 1412 7410 1440 7647
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1504 6798 1532 9318
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1596 7886 1624 8774
rect 1688 8498 1716 9454
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1596 6662 1624 7686
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1688 6458 1716 8434
rect 1964 7886 1992 9862
rect 2056 8022 2084 9998
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2424 9654 2452 9862
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2318 9480 2374 9489
rect 2318 9415 2374 9424
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 2240 8090 2268 8434
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2044 8016 2096 8022
rect 2044 7958 2096 7964
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1768 7472 1820 7478
rect 1768 7414 1820 7420
rect 1780 6866 1808 7414
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1860 6792 1912 6798
rect 1964 6780 1992 7822
rect 2056 7546 2084 7958
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2056 6905 2084 7346
rect 2042 6896 2098 6905
rect 2042 6831 2098 6840
rect 1912 6752 1992 6780
rect 1860 6734 1912 6740
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1688 5778 1716 6394
rect 1872 6118 1900 6734
rect 1952 6656 2004 6662
rect 2136 6656 2188 6662
rect 2004 6616 2084 6644
rect 1952 6598 2004 6604
rect 2056 6322 2084 6616
rect 2136 6598 2188 6604
rect 2148 6390 2176 6598
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1412 4729 1440 5102
rect 1398 4720 1454 4729
rect 1398 4655 1454 4664
rect 1860 4208 1912 4214
rect 1860 4150 1912 4156
rect 1398 4040 1454 4049
rect 1398 3975 1454 3984
rect 1412 3534 1440 3975
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1136 2746 1348 2774
rect 388 2372 440 2378
rect 388 2314 440 2320
rect 400 800 428 2314
rect 1136 800 1164 2746
rect 1872 2553 1900 4150
rect 2332 3738 2360 9415
rect 2608 8974 2636 10134
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3068 9897 3096 9998
rect 3054 9888 3110 9897
rect 3054 9823 3110 9832
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2424 3738 2452 8230
rect 2608 7818 2636 8910
rect 3068 8634 3096 9590
rect 3252 9042 3280 13330
rect 3436 9058 3464 13806
rect 3528 13326 3556 24074
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3620 18834 3648 19110
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3712 17252 3740 27814
rect 4344 27464 4396 27470
rect 4344 27406 4396 27412
rect 4356 27062 4384 27406
rect 4896 27396 4948 27402
rect 4896 27338 4948 27344
rect 4344 27056 4396 27062
rect 4344 26998 4396 27004
rect 4252 26376 4304 26382
rect 4250 26344 4252 26353
rect 4304 26344 4306 26353
rect 4250 26279 4306 26288
rect 4252 26240 4304 26246
rect 4252 26182 4304 26188
rect 4264 25906 4292 26182
rect 4068 25900 4120 25906
rect 4068 25842 4120 25848
rect 4252 25900 4304 25906
rect 4252 25842 4304 25848
rect 4080 25498 4108 25842
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 4264 25106 4292 25842
rect 4356 25294 4384 26998
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4620 26512 4672 26518
rect 4620 26454 4672 26460
rect 4632 26382 4660 26454
rect 4620 26376 4672 26382
rect 4526 26344 4582 26353
rect 4620 26318 4672 26324
rect 4526 26279 4582 26288
rect 4436 26036 4488 26042
rect 4436 25978 4488 25984
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4264 25078 4384 25106
rect 4160 24812 4212 24818
rect 4160 24754 4212 24760
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 3792 24064 3844 24070
rect 3792 24006 3844 24012
rect 3804 23730 3832 24006
rect 4080 23798 4108 24618
rect 4172 24177 4200 24754
rect 4356 24750 4384 25078
rect 4448 24750 4476 25978
rect 4540 25906 4568 26279
rect 4724 25974 4752 26726
rect 4908 26586 4936 27338
rect 4988 26988 5040 26994
rect 4988 26930 5040 26936
rect 4896 26580 4948 26586
rect 4896 26522 4948 26528
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 4816 26042 4844 26318
rect 4804 26036 4856 26042
rect 4804 25978 4856 25984
rect 4712 25968 4764 25974
rect 4712 25910 4764 25916
rect 4528 25900 4580 25906
rect 4528 25842 4580 25848
rect 4896 25900 4948 25906
rect 4896 25842 4948 25848
rect 4804 25220 4856 25226
rect 4804 25162 4856 25168
rect 4816 24954 4844 25162
rect 4804 24948 4856 24954
rect 4804 24890 4856 24896
rect 4908 24818 4936 25842
rect 4528 24812 4580 24818
rect 4528 24754 4580 24760
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4344 24744 4396 24750
rect 4344 24686 4396 24692
rect 4436 24744 4488 24750
rect 4436 24686 4488 24692
rect 4356 24342 4384 24686
rect 4344 24336 4396 24342
rect 4344 24278 4396 24284
rect 4344 24200 4396 24206
rect 4158 24168 4214 24177
rect 4344 24142 4396 24148
rect 4158 24103 4214 24112
rect 4252 24132 4304 24138
rect 4252 24074 4304 24080
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 4172 23866 4200 24006
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 4080 23186 4108 23734
rect 4264 23662 4292 24074
rect 4252 23656 4304 23662
rect 4252 23598 4304 23604
rect 4356 23594 4384 24142
rect 4448 24138 4476 24686
rect 4540 24342 4568 24754
rect 4528 24336 4580 24342
rect 4528 24278 4580 24284
rect 4528 24200 4580 24206
rect 4526 24168 4528 24177
rect 4580 24168 4582 24177
rect 4436 24132 4488 24138
rect 4526 24103 4582 24112
rect 4436 24074 4488 24080
rect 5000 23798 5028 26930
rect 5264 26376 5316 26382
rect 5264 26318 5316 26324
rect 5080 25900 5132 25906
rect 5080 25842 5132 25848
rect 5092 24410 5120 25842
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 5172 24268 5224 24274
rect 5092 24228 5172 24256
rect 4988 23792 5040 23798
rect 4988 23734 5040 23740
rect 4896 23656 4948 23662
rect 4896 23598 4948 23604
rect 4344 23588 4396 23594
rect 4344 23530 4396 23536
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4068 23180 4120 23186
rect 4068 23122 4120 23128
rect 4632 23118 4660 23462
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4252 22976 4304 22982
rect 4252 22918 4304 22924
rect 3976 22432 4028 22438
rect 3976 22374 4028 22380
rect 3988 20942 4016 22374
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 4160 20868 4212 20874
rect 4160 20810 4212 20816
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3804 19378 3832 20334
rect 4172 19666 4200 20810
rect 4264 19854 4292 22918
rect 4908 22094 4936 23598
rect 5000 23322 5028 23734
rect 5092 23662 5120 24228
rect 5172 24210 5224 24216
rect 5276 24206 5304 26318
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 5276 24070 5304 24142
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 4988 23316 5040 23322
rect 4988 23258 5040 23264
rect 5092 22642 5120 23598
rect 5080 22636 5132 22642
rect 5080 22578 5132 22584
rect 5264 22568 5316 22574
rect 5264 22510 5316 22516
rect 4988 22094 5040 22098
rect 4908 22092 5040 22094
rect 4908 22066 4988 22092
rect 4988 22034 5040 22040
rect 5276 21962 5304 22510
rect 5264 21956 5316 21962
rect 5264 21898 5316 21904
rect 4436 21004 4488 21010
rect 4436 20946 4488 20952
rect 4448 19922 4476 20946
rect 5172 20936 5224 20942
rect 5172 20878 5224 20884
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4540 20534 4568 20742
rect 5184 20602 5212 20878
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 4528 20528 4580 20534
rect 4528 20470 4580 20476
rect 4436 19916 4488 19922
rect 4436 19858 4488 19864
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4344 19848 4396 19854
rect 4344 19790 4396 19796
rect 4356 19666 4384 19790
rect 4172 19638 4384 19666
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 3804 18766 3832 18906
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3804 17746 3832 18702
rect 4068 18692 4120 18698
rect 4068 18634 4120 18640
rect 4080 18408 4108 18634
rect 4448 18426 4476 19858
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 4436 18420 4488 18426
rect 4080 18380 4200 18408
rect 4172 18290 4200 18380
rect 4436 18362 4488 18368
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3896 18057 3924 18158
rect 3882 18048 3938 18057
rect 3882 17983 3938 17992
rect 3792 17740 3844 17746
rect 3792 17682 3844 17688
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3884 17604 3936 17610
rect 3884 17546 3936 17552
rect 3620 17224 3740 17252
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3528 9994 3556 10406
rect 3516 9988 3568 9994
rect 3516 9930 3568 9936
rect 3528 9722 3556 9930
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3620 9178 3648 17224
rect 3896 17134 3924 17546
rect 3988 17241 4016 17682
rect 4080 17678 4108 18226
rect 4620 17808 4672 17814
rect 4620 17750 4672 17756
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 3974 17232 4030 17241
rect 3974 17167 4030 17176
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3712 16658 3740 17070
rect 3700 16652 3752 16658
rect 3700 16594 3752 16600
rect 3712 14940 3740 16594
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3804 15502 3832 16186
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3896 15570 3924 15982
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3988 15502 4016 16526
rect 4080 16250 4108 17614
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 4264 16250 4292 16458
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4540 15706 4568 17138
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3792 14952 3844 14958
rect 3712 14912 3792 14940
rect 3792 14894 3844 14900
rect 3804 14414 3832 14894
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3804 14006 3832 14350
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 3804 13190 3832 13942
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 13394 4016 13670
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3712 11898 3740 12786
rect 3804 12646 3832 13126
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3804 12306 3832 12582
rect 3792 12300 3844 12306
rect 3844 12260 3924 12288
rect 3792 12242 3844 12248
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3804 11150 3832 11766
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3896 10674 3924 12260
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3988 11150 4016 11494
rect 4080 11150 4108 11630
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3240 9036 3292 9042
rect 3436 9030 3648 9058
rect 3240 8978 3292 8984
rect 3620 8838 3648 9030
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3620 8634 3648 8774
rect 3804 8634 3832 8978
rect 4080 8974 4108 9522
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3068 7886 3096 8570
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3804 7886 3832 8434
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 3804 7478 3832 7822
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2792 6225 2820 6734
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2884 6458 2912 6666
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 3528 6322 3556 7210
rect 4080 6798 4108 7890
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3712 6390 3740 6598
rect 3700 6384 3752 6390
rect 3700 6326 3752 6332
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 2778 6216 2834 6225
rect 2778 6151 2834 6160
rect 3804 5914 3832 6258
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2516 3534 2544 5510
rect 3896 5234 3924 6598
rect 4080 6254 4108 6734
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5642 4108 6054
rect 4172 5778 4200 8434
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 4172 5302 4200 5714
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 1858 2544 1914 2553
rect 2516 2514 2544 3470
rect 1858 2479 1914 2488
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1872 800 1900 2382
rect 2608 800 2636 4014
rect 2792 3233 2820 4082
rect 3054 4040 3110 4049
rect 3054 3975 3056 3984
rect 3108 3975 3110 3984
rect 3056 3946 3108 3952
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2778 3224 2834 3233
rect 2778 3159 2834 3168
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2792 2530 2820 2994
rect 2884 2650 2912 3402
rect 3160 3126 3188 4082
rect 4172 3602 4200 5238
rect 4264 3738 4292 13262
rect 4632 11830 4660 17750
rect 4724 11880 4752 19722
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4816 19446 4844 19654
rect 4804 19440 4856 19446
rect 4804 19382 4856 19388
rect 5184 19378 5212 19790
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5000 16114 5028 16934
rect 5092 16182 5120 17478
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5080 16176 5132 16182
rect 5080 16118 5132 16124
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 5000 15502 5028 16050
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 5092 15609 5120 15846
rect 5078 15600 5134 15609
rect 5078 15535 5134 15544
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 5092 14822 5120 15438
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5184 14618 5212 16186
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 4986 13968 5042 13977
rect 4986 13903 4988 13912
rect 5040 13903 5042 13912
rect 4988 13874 5040 13880
rect 5368 13530 5396 28086
rect 5644 27946 5672 35142
rect 6644 35080 6696 35086
rect 6644 35022 6696 35028
rect 5816 34740 5868 34746
rect 5816 34682 5868 34688
rect 5724 34604 5776 34610
rect 5724 34546 5776 34552
rect 5736 34202 5764 34546
rect 5724 34196 5776 34202
rect 5724 34138 5776 34144
rect 5828 33998 5856 34682
rect 6656 34649 6684 35022
rect 6642 34640 6698 34649
rect 6276 34604 6328 34610
rect 6642 34575 6698 34584
rect 6276 34546 6328 34552
rect 5915 34300 6223 34320
rect 5915 34298 5921 34300
rect 5977 34298 6001 34300
rect 6057 34298 6081 34300
rect 6137 34298 6161 34300
rect 6217 34298 6223 34300
rect 5977 34246 5979 34298
rect 6159 34246 6161 34298
rect 5915 34244 5921 34246
rect 5977 34244 6001 34246
rect 6057 34244 6081 34246
rect 6137 34244 6161 34246
rect 6217 34244 6223 34246
rect 5915 34224 6223 34244
rect 6182 34096 6238 34105
rect 6182 34031 6238 34040
rect 6196 33998 6224 34031
rect 5816 33992 5868 33998
rect 5816 33934 5868 33940
rect 6184 33992 6236 33998
rect 6184 33934 6236 33940
rect 6288 33522 6316 34546
rect 6368 33992 6420 33998
rect 6368 33934 6420 33940
rect 6276 33516 6328 33522
rect 6276 33458 6328 33464
rect 5915 33212 6223 33232
rect 5915 33210 5921 33212
rect 5977 33210 6001 33212
rect 6057 33210 6081 33212
rect 6137 33210 6161 33212
rect 6217 33210 6223 33212
rect 5977 33158 5979 33210
rect 6159 33158 6161 33210
rect 5915 33156 5921 33158
rect 5977 33156 6001 33158
rect 6057 33156 6081 33158
rect 6137 33156 6161 33158
rect 6217 33156 6223 33158
rect 5915 33136 6223 33156
rect 6380 33046 6408 33934
rect 6368 33040 6420 33046
rect 6368 32982 6420 32988
rect 5724 32836 5776 32842
rect 5724 32778 5776 32784
rect 5736 32230 5764 32778
rect 5724 32224 5776 32230
rect 5724 32166 5776 32172
rect 5736 28150 5764 32166
rect 5915 32124 6223 32144
rect 5915 32122 5921 32124
rect 5977 32122 6001 32124
rect 6057 32122 6081 32124
rect 6137 32122 6161 32124
rect 6217 32122 6223 32124
rect 5977 32070 5979 32122
rect 6159 32070 6161 32122
rect 5915 32068 5921 32070
rect 5977 32068 6001 32070
rect 6057 32068 6081 32070
rect 6137 32068 6161 32070
rect 6217 32068 6223 32070
rect 5915 32048 6223 32068
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6368 31680 6420 31686
rect 6368 31622 6420 31628
rect 6276 31340 6328 31346
rect 6276 31282 6328 31288
rect 5816 31136 5868 31142
rect 5816 31078 5868 31084
rect 5828 30666 5856 31078
rect 5915 31036 6223 31056
rect 5915 31034 5921 31036
rect 5977 31034 6001 31036
rect 6057 31034 6081 31036
rect 6137 31034 6161 31036
rect 6217 31034 6223 31036
rect 5977 30982 5979 31034
rect 6159 30982 6161 31034
rect 5915 30980 5921 30982
rect 5977 30980 6001 30982
rect 6057 30980 6081 30982
rect 6137 30980 6161 30982
rect 6217 30980 6223 30982
rect 5915 30960 6223 30980
rect 6288 30938 6316 31282
rect 6380 31278 6408 31622
rect 6368 31272 6420 31278
rect 6368 31214 6420 31220
rect 6276 30932 6328 30938
rect 6276 30874 6328 30880
rect 6380 30802 6408 31214
rect 6472 30870 6500 31758
rect 6460 30864 6512 30870
rect 6460 30806 6512 30812
rect 6368 30796 6420 30802
rect 6368 30738 6420 30744
rect 5816 30660 5868 30666
rect 5816 30602 5868 30608
rect 6472 30598 6500 30806
rect 6460 30592 6512 30598
rect 6460 30534 6512 30540
rect 6368 30184 6420 30190
rect 6368 30126 6420 30132
rect 5816 30048 5868 30054
rect 5816 29990 5868 29996
rect 5828 28558 5856 29990
rect 5915 29948 6223 29968
rect 5915 29946 5921 29948
rect 5977 29946 6001 29948
rect 6057 29946 6081 29948
rect 6137 29946 6161 29948
rect 6217 29946 6223 29948
rect 5977 29894 5979 29946
rect 6159 29894 6161 29946
rect 5915 29892 5921 29894
rect 5977 29892 6001 29894
rect 6057 29892 6081 29894
rect 6137 29892 6161 29894
rect 6217 29892 6223 29894
rect 5915 29872 6223 29892
rect 6380 29850 6408 30126
rect 6656 29850 6684 34575
rect 6748 33998 6776 37454
rect 7300 37126 7328 42298
rect 7484 42106 7512 44814
rect 8208 44814 8260 44820
rect 8022 44775 8078 44784
rect 8036 44742 8064 44775
rect 7656 44736 7708 44742
rect 7656 44678 7708 44684
rect 8024 44736 8076 44742
rect 8024 44678 8076 44684
rect 7668 43994 7696 44678
rect 8220 44577 8248 44814
rect 10880 44636 11188 44656
rect 10880 44634 10886 44636
rect 10942 44634 10966 44636
rect 11022 44634 11046 44636
rect 11102 44634 11126 44636
rect 11182 44634 11188 44636
rect 10942 44582 10944 44634
rect 11124 44582 11126 44634
rect 10880 44580 10886 44582
rect 10942 44580 10966 44582
rect 11022 44580 11046 44582
rect 11102 44580 11126 44582
rect 11182 44580 11188 44582
rect 8206 44568 8262 44577
rect 10880 44560 11188 44580
rect 20811 44636 21119 44656
rect 20811 44634 20817 44636
rect 20873 44634 20897 44636
rect 20953 44634 20977 44636
rect 21033 44634 21057 44636
rect 21113 44634 21119 44636
rect 20873 44582 20875 44634
rect 21055 44582 21057 44634
rect 20811 44580 20817 44582
rect 20873 44580 20897 44582
rect 20953 44580 20977 44582
rect 21033 44580 21057 44582
rect 21113 44580 21119 44582
rect 20811 44560 21119 44580
rect 8206 44503 8262 44512
rect 9864 44396 9916 44402
rect 9864 44338 9916 44344
rect 20076 44396 20128 44402
rect 20076 44338 20128 44344
rect 8852 44328 8904 44334
rect 8852 44270 8904 44276
rect 9496 44328 9548 44334
rect 9496 44270 9548 44276
rect 8576 44192 8628 44198
rect 8576 44134 8628 44140
rect 7656 43988 7708 43994
rect 7656 43930 7708 43936
rect 7668 43246 7696 43930
rect 8116 43716 8168 43722
rect 8116 43658 8168 43664
rect 8024 43648 8076 43654
rect 8024 43590 8076 43596
rect 8036 43382 8064 43590
rect 8128 43450 8156 43658
rect 8116 43444 8168 43450
rect 8116 43386 8168 43392
rect 8588 43382 8616 44134
rect 8864 43994 8892 44270
rect 8852 43988 8904 43994
rect 8852 43930 8904 43936
rect 8024 43376 8076 43382
rect 8024 43318 8076 43324
rect 8576 43376 8628 43382
rect 8576 43318 8628 43324
rect 9128 43308 9180 43314
rect 9128 43250 9180 43256
rect 7656 43240 7708 43246
rect 7656 43182 7708 43188
rect 8024 43240 8076 43246
rect 8024 43182 8076 43188
rect 8576 43240 8628 43246
rect 8576 43182 8628 43188
rect 8036 42838 8064 43182
rect 8588 42906 8616 43182
rect 8576 42900 8628 42906
rect 8576 42842 8628 42848
rect 8024 42832 8076 42838
rect 8024 42774 8076 42780
rect 7656 42628 7708 42634
rect 7656 42570 7708 42576
rect 7484 42078 7604 42106
rect 7472 42016 7524 42022
rect 7472 41958 7524 41964
rect 7484 41546 7512 41958
rect 7472 41540 7524 41546
rect 7472 41482 7524 41488
rect 7576 38214 7604 42078
rect 7668 41478 7696 42570
rect 7748 42220 7800 42226
rect 7748 42162 7800 42168
rect 7760 41818 7788 42162
rect 7748 41812 7800 41818
rect 7748 41754 7800 41760
rect 7656 41472 7708 41478
rect 7656 41414 7708 41420
rect 7668 39914 7696 41414
rect 8036 40662 8064 42774
rect 9140 42702 9168 43250
rect 9128 42696 9180 42702
rect 9128 42638 9180 42644
rect 8392 42016 8444 42022
rect 8392 41958 8444 41964
rect 8404 41682 8432 41958
rect 8392 41676 8444 41682
rect 8392 41618 8444 41624
rect 8944 41472 8996 41478
rect 8944 41414 8996 41420
rect 8956 41138 8984 41414
rect 8944 41132 8996 41138
rect 8944 41074 8996 41080
rect 8484 41064 8536 41070
rect 8484 41006 8536 41012
rect 8024 40656 8076 40662
rect 8024 40598 8076 40604
rect 8300 40520 8352 40526
rect 8300 40462 8352 40468
rect 8312 40118 8340 40462
rect 8300 40112 8352 40118
rect 8300 40054 8352 40060
rect 7656 39908 7708 39914
rect 7656 39850 7708 39856
rect 8116 39432 8168 39438
rect 8116 39374 8168 39380
rect 8024 39024 8076 39030
rect 8024 38966 8076 38972
rect 8036 38350 8064 38966
rect 8024 38344 8076 38350
rect 8024 38286 8076 38292
rect 7564 38208 7616 38214
rect 7564 38150 7616 38156
rect 7748 37868 7800 37874
rect 7748 37810 7800 37816
rect 7760 37194 7788 37810
rect 7932 37800 7984 37806
rect 7932 37742 7984 37748
rect 7944 37194 7972 37742
rect 7748 37188 7800 37194
rect 7748 37130 7800 37136
rect 7932 37188 7984 37194
rect 7932 37130 7984 37136
rect 7288 37120 7340 37126
rect 7288 37062 7340 37068
rect 7472 36780 7524 36786
rect 8036 36768 8064 38286
rect 8128 37126 8156 39374
rect 8208 39296 8260 39302
rect 8208 39238 8260 39244
rect 8220 37874 8248 39238
rect 8312 38554 8340 40054
rect 8496 39370 8524 41006
rect 9140 40526 9168 42638
rect 9128 40520 9180 40526
rect 9128 40462 9180 40468
rect 9036 40452 9088 40458
rect 9036 40394 9088 40400
rect 8944 40384 8996 40390
rect 8944 40326 8996 40332
rect 8956 40118 8984 40326
rect 9048 40118 9076 40394
rect 9508 40118 9536 44270
rect 9772 43716 9824 43722
rect 9772 43658 9824 43664
rect 9784 42838 9812 43658
rect 9772 42832 9824 42838
rect 9772 42774 9824 42780
rect 9588 40520 9640 40526
rect 9588 40462 9640 40468
rect 9600 40186 9628 40462
rect 9588 40180 9640 40186
rect 9588 40122 9640 40128
rect 8944 40112 8996 40118
rect 8944 40054 8996 40060
rect 9036 40112 9088 40118
rect 9036 40054 9088 40060
rect 9496 40112 9548 40118
rect 9496 40054 9548 40060
rect 9680 40044 9732 40050
rect 9680 39986 9732 39992
rect 8760 39976 8812 39982
rect 8760 39918 8812 39924
rect 8576 39840 8628 39846
rect 8576 39782 8628 39788
rect 8588 39506 8616 39782
rect 8576 39500 8628 39506
rect 8576 39442 8628 39448
rect 8484 39364 8536 39370
rect 8484 39306 8536 39312
rect 8772 38962 8800 39918
rect 9496 39840 9548 39846
rect 9496 39782 9548 39788
rect 9036 39636 9088 39642
rect 9036 39578 9088 39584
rect 8576 38956 8628 38962
rect 8760 38956 8812 38962
rect 8576 38898 8628 38904
rect 8680 38916 8760 38944
rect 8300 38548 8352 38554
rect 8300 38490 8352 38496
rect 8208 37868 8260 37874
rect 8208 37810 8260 37816
rect 8312 37262 8340 38490
rect 8588 38350 8616 38898
rect 8576 38344 8628 38350
rect 8576 38286 8628 38292
rect 8300 37256 8352 37262
rect 8300 37198 8352 37204
rect 8116 37120 8168 37126
rect 8116 37062 8168 37068
rect 8300 37120 8352 37126
rect 8300 37062 8352 37068
rect 8116 36780 8168 36786
rect 7472 36722 7524 36728
rect 7852 36740 8116 36768
rect 7196 36576 7248 36582
rect 7196 36518 7248 36524
rect 7208 36378 7236 36518
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 7196 36032 7248 36038
rect 7196 35974 7248 35980
rect 6828 34740 6880 34746
rect 6828 34682 6880 34688
rect 6736 33992 6788 33998
rect 6736 33934 6788 33940
rect 6736 33312 6788 33318
rect 6736 33254 6788 33260
rect 6748 32434 6776 33254
rect 6840 32978 6868 34682
rect 7012 33992 7064 33998
rect 7012 33934 7064 33940
rect 7024 33590 7052 33934
rect 7012 33584 7064 33590
rect 7012 33526 7064 33532
rect 7104 33312 7156 33318
rect 7104 33254 7156 33260
rect 6828 32972 6880 32978
rect 6828 32914 6880 32920
rect 6736 32428 6788 32434
rect 6736 32370 6788 32376
rect 6840 31822 6868 32914
rect 6920 32904 6972 32910
rect 6920 32846 6972 32852
rect 6932 32570 6960 32846
rect 7116 32842 7144 33254
rect 7104 32836 7156 32842
rect 7104 32778 7156 32784
rect 6920 32564 6972 32570
rect 6920 32506 6972 32512
rect 6828 31816 6880 31822
rect 6828 31758 6880 31764
rect 7012 31136 7064 31142
rect 7012 31078 7064 31084
rect 7024 30666 7052 31078
rect 7104 30864 7156 30870
rect 7104 30806 7156 30812
rect 7012 30660 7064 30666
rect 7012 30602 7064 30608
rect 7116 30326 7144 30806
rect 7104 30320 7156 30326
rect 7104 30262 7156 30268
rect 7208 30258 7236 35974
rect 7484 35834 7512 36722
rect 7564 36644 7616 36650
rect 7564 36586 7616 36592
rect 7472 35828 7524 35834
rect 7472 35770 7524 35776
rect 7288 33856 7340 33862
rect 7288 33798 7340 33804
rect 7300 32910 7328 33798
rect 7288 32904 7340 32910
rect 7288 32846 7340 32852
rect 7380 32768 7432 32774
rect 7380 32710 7432 32716
rect 7392 32434 7420 32710
rect 7380 32428 7432 32434
rect 7380 32370 7432 32376
rect 7380 30728 7432 30734
rect 7380 30670 7432 30676
rect 7472 30728 7524 30734
rect 7472 30670 7524 30676
rect 7392 30394 7420 30670
rect 7484 30598 7512 30670
rect 7472 30592 7524 30598
rect 7472 30534 7524 30540
rect 7380 30388 7432 30394
rect 7380 30330 7432 30336
rect 7196 30252 7248 30258
rect 7196 30194 7248 30200
rect 6368 29844 6420 29850
rect 6368 29786 6420 29792
rect 6644 29844 6696 29850
rect 6644 29786 6696 29792
rect 6552 29572 6604 29578
rect 6552 29514 6604 29520
rect 5915 28860 6223 28880
rect 5915 28858 5921 28860
rect 5977 28858 6001 28860
rect 6057 28858 6081 28860
rect 6137 28858 6161 28860
rect 6217 28858 6223 28860
rect 5977 28806 5979 28858
rect 6159 28806 6161 28858
rect 5915 28804 5921 28806
rect 5977 28804 6001 28806
rect 6057 28804 6081 28806
rect 6137 28804 6161 28806
rect 6217 28804 6223 28806
rect 5915 28784 6223 28804
rect 5816 28552 5868 28558
rect 5816 28494 5868 28500
rect 5724 28144 5776 28150
rect 5724 28086 5776 28092
rect 5632 27940 5684 27946
rect 5632 27882 5684 27888
rect 5816 27940 5868 27946
rect 5816 27882 5868 27888
rect 5448 26920 5500 26926
rect 5448 26862 5500 26868
rect 5460 26518 5488 26862
rect 5448 26512 5500 26518
rect 5448 26454 5500 26460
rect 5540 24200 5592 24206
rect 5538 24168 5540 24177
rect 5592 24168 5594 24177
rect 5538 24103 5594 24112
rect 5552 23730 5580 24103
rect 5540 23724 5592 23730
rect 5540 23666 5592 23672
rect 5448 23316 5500 23322
rect 5448 23258 5500 23264
rect 5460 22030 5488 23258
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5448 21616 5500 21622
rect 5448 21558 5500 21564
rect 5460 21146 5488 21558
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 5184 12986 5212 13194
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4804 11892 4856 11898
rect 4724 11852 4804 11880
rect 4804 11834 4856 11840
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4356 10538 4384 11086
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4540 10742 4568 10950
rect 4528 10736 4580 10742
rect 4528 10678 4580 10684
rect 4908 10606 4936 12106
rect 5000 11762 5028 12582
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5368 11762 5396 12174
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5460 11218 5488 15438
rect 5552 14498 5580 18566
rect 5644 17252 5672 27882
rect 5828 27674 5856 27882
rect 5915 27772 6223 27792
rect 5915 27770 5921 27772
rect 5977 27770 6001 27772
rect 6057 27770 6081 27772
rect 6137 27770 6161 27772
rect 6217 27770 6223 27772
rect 5977 27718 5979 27770
rect 6159 27718 6161 27770
rect 5915 27716 5921 27718
rect 5977 27716 6001 27718
rect 6057 27716 6081 27718
rect 6137 27716 6161 27718
rect 6217 27716 6223 27718
rect 5915 27696 6223 27716
rect 5816 27668 5868 27674
rect 5816 27610 5868 27616
rect 5828 26994 5856 27610
rect 6564 27606 6592 29514
rect 7012 29164 7064 29170
rect 7012 29106 7064 29112
rect 6644 28960 6696 28966
rect 6644 28902 6696 28908
rect 6656 28082 6684 28902
rect 7024 28762 7052 29106
rect 7196 29096 7248 29102
rect 7196 29038 7248 29044
rect 7012 28756 7064 28762
rect 7012 28698 7064 28704
rect 7208 28626 7236 29038
rect 7576 28694 7604 36586
rect 7748 36576 7800 36582
rect 7748 36518 7800 36524
rect 7656 35080 7708 35086
rect 7656 35022 7708 35028
rect 7668 34542 7696 35022
rect 7656 34536 7708 34542
rect 7656 34478 7708 34484
rect 7656 34400 7708 34406
rect 7656 34342 7708 34348
rect 7668 33590 7696 34342
rect 7656 33584 7708 33590
rect 7656 33526 7708 33532
rect 7760 31754 7788 36518
rect 7852 34746 7880 36740
rect 8116 36722 8168 36728
rect 8024 36644 8076 36650
rect 8024 36586 8076 36592
rect 7932 36032 7984 36038
rect 7932 35974 7984 35980
rect 7944 35698 7972 35974
rect 7932 35692 7984 35698
rect 7932 35634 7984 35640
rect 8036 35290 8064 36586
rect 8116 36168 8168 36174
rect 8116 36110 8168 36116
rect 8024 35284 8076 35290
rect 8024 35226 8076 35232
rect 7932 35012 7984 35018
rect 7932 34954 7984 34960
rect 7840 34740 7892 34746
rect 7840 34682 7892 34688
rect 7944 34082 7972 34954
rect 8036 34610 8064 35226
rect 8024 34604 8076 34610
rect 8024 34546 8076 34552
rect 8128 34202 8156 36110
rect 8208 35828 8260 35834
rect 8208 35770 8260 35776
rect 8220 35086 8248 35770
rect 8312 35222 8340 37062
rect 8484 36168 8536 36174
rect 8484 36110 8536 36116
rect 8392 35692 8444 35698
rect 8392 35634 8444 35640
rect 8404 35290 8432 35634
rect 8496 35494 8524 36110
rect 8484 35488 8536 35494
rect 8484 35430 8536 35436
rect 8680 35306 8708 38916
rect 8760 38898 8812 38904
rect 9048 38350 9076 39578
rect 9312 39364 9364 39370
rect 9312 39306 9364 39312
rect 9128 39296 9180 39302
rect 9128 39238 9180 39244
rect 9140 38962 9168 39238
rect 9324 39098 9352 39306
rect 9312 39092 9364 39098
rect 9312 39034 9364 39040
rect 9128 38956 9180 38962
rect 9128 38898 9180 38904
rect 9140 38486 9168 38898
rect 9312 38888 9364 38894
rect 9312 38830 9364 38836
rect 9220 38752 9272 38758
rect 9220 38694 9272 38700
rect 9128 38480 9180 38486
rect 9128 38422 9180 38428
rect 9232 38418 9260 38694
rect 9220 38412 9272 38418
rect 9220 38354 9272 38360
rect 9036 38344 9088 38350
rect 9036 38286 9088 38292
rect 8944 37868 8996 37874
rect 8944 37810 8996 37816
rect 8956 37466 8984 37810
rect 8944 37460 8996 37466
rect 8944 37402 8996 37408
rect 8392 35284 8444 35290
rect 8392 35226 8444 35232
rect 8496 35278 8708 35306
rect 8300 35216 8352 35222
rect 8496 35170 8524 35278
rect 8300 35158 8352 35164
rect 8404 35142 8524 35170
rect 8852 35216 8904 35222
rect 8852 35158 8904 35164
rect 8208 35080 8260 35086
rect 8208 35022 8260 35028
rect 8116 34196 8168 34202
rect 8116 34138 8168 34144
rect 8300 34128 8352 34134
rect 8298 34096 8300 34105
rect 8352 34096 8354 34105
rect 7944 34066 8248 34082
rect 7932 34060 8248 34066
rect 7984 34054 8248 34060
rect 7932 34002 7984 34008
rect 8116 33992 8168 33998
rect 8116 33934 8168 33940
rect 8128 33862 8156 33934
rect 8116 33856 8168 33862
rect 8116 33798 8168 33804
rect 7932 33312 7984 33318
rect 7932 33254 7984 33260
rect 7944 32502 7972 33254
rect 7932 32496 7984 32502
rect 7932 32438 7984 32444
rect 7760 31726 7880 31754
rect 7748 31680 7800 31686
rect 7748 31622 7800 31628
rect 7760 31346 7788 31622
rect 7748 31340 7800 31346
rect 7748 31282 7800 31288
rect 7656 29504 7708 29510
rect 7656 29446 7708 29452
rect 7564 28688 7616 28694
rect 7564 28630 7616 28636
rect 7196 28620 7248 28626
rect 7196 28562 7248 28568
rect 7472 28620 7524 28626
rect 7472 28562 7524 28568
rect 6828 28416 6880 28422
rect 6828 28358 6880 28364
rect 6840 28218 6868 28358
rect 6828 28212 6880 28218
rect 6828 28154 6880 28160
rect 7196 28144 7248 28150
rect 7196 28086 7248 28092
rect 7288 28144 7340 28150
rect 7288 28086 7340 28092
rect 6644 28076 6696 28082
rect 6644 28018 6696 28024
rect 7012 28076 7064 28082
rect 7012 28018 7064 28024
rect 7024 27674 7052 28018
rect 7012 27668 7064 27674
rect 7012 27610 7064 27616
rect 6552 27600 6604 27606
rect 6552 27542 6604 27548
rect 6276 27328 6328 27334
rect 6276 27270 6328 27276
rect 5816 26988 5868 26994
rect 5816 26930 5868 26936
rect 5724 26852 5776 26858
rect 5724 26794 5776 26800
rect 5736 26058 5764 26794
rect 5828 26314 5856 26930
rect 6288 26858 6316 27270
rect 6276 26852 6328 26858
rect 6276 26794 6328 26800
rect 5915 26684 6223 26704
rect 5915 26682 5921 26684
rect 5977 26682 6001 26684
rect 6057 26682 6081 26684
rect 6137 26682 6161 26684
rect 6217 26682 6223 26684
rect 5977 26630 5979 26682
rect 6159 26630 6161 26682
rect 5915 26628 5921 26630
rect 5977 26628 6001 26630
rect 6057 26628 6081 26630
rect 6137 26628 6161 26630
rect 6217 26628 6223 26630
rect 5915 26608 6223 26628
rect 6288 26518 6316 26794
rect 6276 26512 6328 26518
rect 6276 26454 6328 26460
rect 5816 26308 5868 26314
rect 5816 26250 5868 26256
rect 5736 26042 5856 26058
rect 5736 26036 5868 26042
rect 5736 26030 5816 26036
rect 5736 25430 5764 26030
rect 5816 25978 5868 25984
rect 6564 25974 6592 27542
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 6736 27396 6788 27402
rect 6736 27338 6788 27344
rect 6748 27062 6776 27338
rect 6736 27056 6788 27062
rect 6736 26998 6788 27004
rect 6552 25968 6604 25974
rect 6552 25910 6604 25916
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 5724 25424 5776 25430
rect 5724 25366 5776 25372
rect 5828 25294 5856 25638
rect 5915 25596 6223 25616
rect 5915 25594 5921 25596
rect 5977 25594 6001 25596
rect 6057 25594 6081 25596
rect 6137 25594 6161 25596
rect 6217 25594 6223 25596
rect 5977 25542 5979 25594
rect 6159 25542 6161 25594
rect 5915 25540 5921 25542
rect 5977 25540 6001 25542
rect 6057 25540 6081 25542
rect 6137 25540 6161 25542
rect 6217 25540 6223 25542
rect 5915 25520 6223 25540
rect 6368 25492 6420 25498
rect 6368 25434 6420 25440
rect 5816 25288 5868 25294
rect 5816 25230 5868 25236
rect 5724 23656 5776 23662
rect 5724 23598 5776 23604
rect 5736 23322 5764 23598
rect 5724 23316 5776 23322
rect 5724 23258 5776 23264
rect 5736 22658 5764 23258
rect 5828 23186 5856 25230
rect 5915 24508 6223 24528
rect 5915 24506 5921 24508
rect 5977 24506 6001 24508
rect 6057 24506 6081 24508
rect 6137 24506 6161 24508
rect 6217 24506 6223 24508
rect 5977 24454 5979 24506
rect 6159 24454 6161 24506
rect 5915 24452 5921 24454
rect 5977 24452 6001 24454
rect 6057 24452 6081 24454
rect 6137 24452 6161 24454
rect 6217 24452 6223 24454
rect 5915 24432 6223 24452
rect 5908 24336 5960 24342
rect 5960 24296 6040 24324
rect 5908 24278 5960 24284
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 5920 23798 5948 24142
rect 6012 24070 6040 24296
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 5908 23792 5960 23798
rect 5908 23734 5960 23740
rect 5915 23420 6223 23440
rect 5915 23418 5921 23420
rect 5977 23418 6001 23420
rect 6057 23418 6081 23420
rect 6137 23418 6161 23420
rect 6217 23418 6223 23420
rect 5977 23366 5979 23418
rect 6159 23366 6161 23418
rect 5915 23364 5921 23366
rect 5977 23364 6001 23366
rect 6057 23364 6081 23366
rect 6137 23364 6161 23366
rect 6217 23364 6223 23366
rect 5915 23344 6223 23364
rect 5816 23180 5868 23186
rect 5816 23122 5868 23128
rect 5736 22630 5856 22658
rect 5724 22568 5776 22574
rect 5724 22510 5776 22516
rect 5736 18426 5764 22510
rect 5828 19922 5856 22630
rect 5915 22332 6223 22352
rect 5915 22330 5921 22332
rect 5977 22330 6001 22332
rect 6057 22330 6081 22332
rect 6137 22330 6161 22332
rect 6217 22330 6223 22332
rect 5977 22278 5979 22330
rect 6159 22278 6161 22330
rect 5915 22276 5921 22278
rect 5977 22276 6001 22278
rect 6057 22276 6081 22278
rect 6137 22276 6161 22278
rect 6217 22276 6223 22278
rect 5915 22256 6223 22276
rect 6380 22094 6408 25434
rect 6460 25220 6512 25226
rect 6460 25162 6512 25168
rect 6644 25220 6696 25226
rect 6644 25162 6696 25168
rect 6472 24410 6500 25162
rect 6656 24410 6684 25162
rect 6748 24818 6776 26998
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6840 26382 6868 26726
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 6828 25764 6880 25770
rect 6828 25706 6880 25712
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6840 24750 6868 25706
rect 6932 25498 6960 26522
rect 7116 26042 7144 27406
rect 7104 26036 7156 26042
rect 7104 25978 7156 25984
rect 7012 25832 7064 25838
rect 7012 25774 7064 25780
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6828 24744 6880 24750
rect 6828 24686 6880 24692
rect 6460 24404 6512 24410
rect 6460 24346 6512 24352
rect 6644 24404 6696 24410
rect 6644 24346 6696 24352
rect 6552 24268 6604 24274
rect 6552 24210 6604 24216
rect 6460 23724 6512 23730
rect 6460 23666 6512 23672
rect 6472 22642 6500 23666
rect 6564 23576 6592 24210
rect 6932 23730 6960 25230
rect 6644 23724 6696 23730
rect 6920 23724 6972 23730
rect 6696 23684 6868 23712
rect 6644 23666 6696 23672
rect 6644 23588 6696 23594
rect 6564 23548 6644 23576
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 6380 22066 6500 22094
rect 6472 21486 6500 22066
rect 6564 21554 6592 23548
rect 6644 23530 6696 23536
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6552 21548 6604 21554
rect 6604 21508 6684 21536
rect 6552 21490 6604 21496
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 6276 21344 6328 21350
rect 6276 21286 6328 21292
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 5915 21244 6223 21264
rect 5915 21242 5921 21244
rect 5977 21242 6001 21244
rect 6057 21242 6081 21244
rect 6137 21242 6161 21244
rect 6217 21242 6223 21244
rect 5977 21190 5979 21242
rect 6159 21190 6161 21242
rect 5915 21188 5921 21190
rect 5977 21188 6001 21190
rect 6057 21188 6081 21190
rect 6137 21188 6161 21190
rect 6217 21188 6223 21190
rect 5915 21168 6223 21188
rect 6288 20806 6316 21286
rect 6564 20942 6592 21286
rect 6656 21146 6684 21508
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 6748 20942 6776 21830
rect 6840 21554 6868 23684
rect 6920 23666 6972 23672
rect 6920 23520 6972 23526
rect 6920 23462 6972 23468
rect 6932 23118 6960 23462
rect 6920 23112 6972 23118
rect 6920 23054 6972 23060
rect 7024 22778 7052 25774
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7012 22772 7064 22778
rect 7012 22714 7064 22720
rect 7116 22030 7144 24550
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 6828 21548 6880 21554
rect 6880 21508 6960 21536
rect 6828 21490 6880 21496
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 6552 20936 6604 20942
rect 6736 20936 6788 20942
rect 6552 20878 6604 20884
rect 6656 20896 6736 20924
rect 6276 20800 6328 20806
rect 6276 20742 6328 20748
rect 6656 20398 6684 20896
rect 6736 20878 6788 20884
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 5915 20156 6223 20176
rect 5915 20154 5921 20156
rect 5977 20154 6001 20156
rect 6057 20154 6081 20156
rect 6137 20154 6161 20156
rect 6217 20154 6223 20156
rect 5977 20102 5979 20154
rect 6159 20102 6161 20154
rect 5915 20100 5921 20102
rect 5977 20100 6001 20102
rect 6057 20100 6081 20102
rect 6137 20100 6161 20102
rect 6217 20100 6223 20102
rect 5915 20080 6223 20100
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6276 19712 6328 19718
rect 6276 19654 6328 19660
rect 5915 19068 6223 19088
rect 5915 19066 5921 19068
rect 5977 19066 6001 19068
rect 6057 19066 6081 19068
rect 6137 19066 6161 19068
rect 6217 19066 6223 19068
rect 5977 19014 5979 19066
rect 6159 19014 6161 19066
rect 5915 19012 5921 19014
rect 5977 19012 6001 19014
rect 6057 19012 6081 19014
rect 6137 19012 6161 19014
rect 6217 19012 6223 19014
rect 5915 18992 6223 19012
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5736 18086 5764 18362
rect 6196 18358 6224 18702
rect 5816 18352 5868 18358
rect 5816 18294 5868 18300
rect 6184 18352 6236 18358
rect 6184 18294 6236 18300
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 5828 17882 5856 18294
rect 5915 17980 6223 18000
rect 5915 17978 5921 17980
rect 5977 17978 6001 17980
rect 6057 17978 6081 17980
rect 6137 17978 6161 17980
rect 6217 17978 6223 17980
rect 5977 17926 5979 17978
rect 6159 17926 6161 17978
rect 5915 17924 5921 17926
rect 5977 17924 6001 17926
rect 6057 17924 6081 17926
rect 6137 17924 6161 17926
rect 6217 17924 6223 17926
rect 5915 17904 6223 17924
rect 5816 17876 5868 17882
rect 5816 17818 5868 17824
rect 5644 17224 5856 17252
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 16046 5764 16390
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5828 15586 5856 17224
rect 5915 16892 6223 16912
rect 5915 16890 5921 16892
rect 5977 16890 6001 16892
rect 6057 16890 6081 16892
rect 6137 16890 6161 16892
rect 6217 16890 6223 16892
rect 5977 16838 5979 16890
rect 6159 16838 6161 16890
rect 5915 16836 5921 16838
rect 5977 16836 6001 16838
rect 6057 16836 6081 16838
rect 6137 16836 6161 16838
rect 6217 16836 6223 16838
rect 5915 16816 6223 16836
rect 6288 16640 6316 19654
rect 6380 18834 6408 19790
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6288 16612 6408 16640
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 5915 15804 6223 15824
rect 5915 15802 5921 15804
rect 5977 15802 6001 15804
rect 6057 15802 6081 15804
rect 6137 15802 6161 15804
rect 6217 15802 6223 15804
rect 5977 15750 5979 15802
rect 6159 15750 6161 15802
rect 5915 15748 5921 15750
rect 5977 15748 6001 15750
rect 6057 15748 6081 15750
rect 6137 15748 6161 15750
rect 6217 15748 6223 15750
rect 5915 15728 6223 15748
rect 6182 15600 6238 15609
rect 5828 15558 5948 15586
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5552 14470 5672 14498
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5172 11076 5224 11082
rect 5356 11076 5408 11082
rect 5172 11018 5224 11024
rect 5276 11036 5356 11064
rect 5184 10742 5212 11018
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4540 9466 4568 9522
rect 4448 7954 4476 9454
rect 4540 9450 4752 9466
rect 4540 9444 4764 9450
rect 4540 9438 4712 9444
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4356 6798 4384 7482
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4344 6656 4396 6662
rect 4448 6610 4476 7278
rect 4396 6604 4476 6610
rect 4344 6598 4476 6604
rect 4356 6582 4476 6598
rect 4356 6186 4384 6582
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4448 5710 4476 6054
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4632 4690 4660 9438
rect 4712 9386 4764 9392
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4816 8498 4844 9318
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 5000 8090 5028 9930
rect 5092 9450 5120 9998
rect 5276 9926 5304 11036
rect 5356 11018 5408 11024
rect 5552 10792 5580 14350
rect 5644 12782 5672 14470
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5644 11762 5672 12038
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5552 10764 5672 10792
rect 5448 10668 5500 10674
rect 5500 10628 5580 10656
rect 5448 10610 5500 10616
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 5092 9042 5120 9386
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5092 8566 5120 8978
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5276 7886 5304 9862
rect 5368 9518 5396 9930
rect 5446 9616 5502 9625
rect 5552 9586 5580 10628
rect 5446 9551 5502 9560
rect 5540 9580 5592 9586
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5368 7818 5396 9454
rect 5460 8022 5488 9551
rect 5540 9522 5592 9528
rect 5552 8634 5580 9522
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5644 8514 5672 10764
rect 5736 10538 5764 14962
rect 5828 14414 5856 15302
rect 5920 14890 5948 15558
rect 6182 15535 6238 15544
rect 6196 15502 6224 15535
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 5908 14884 5960 14890
rect 5908 14826 5960 14832
rect 5915 14716 6223 14736
rect 5915 14714 5921 14716
rect 5977 14714 6001 14716
rect 6057 14714 6081 14716
rect 6137 14714 6161 14716
rect 6217 14714 6223 14716
rect 5977 14662 5979 14714
rect 6159 14662 6161 14714
rect 5915 14660 5921 14662
rect 5977 14660 6001 14662
rect 6057 14660 6081 14662
rect 6137 14660 6161 14662
rect 6217 14660 6223 14662
rect 5915 14640 6223 14660
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5816 14408 5868 14414
rect 5920 14385 5948 14418
rect 5816 14350 5868 14356
rect 5906 14376 5962 14385
rect 5906 14311 5962 14320
rect 5920 14074 5948 14311
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 5915 13628 6223 13648
rect 5915 13626 5921 13628
rect 5977 13626 6001 13628
rect 6057 13626 6081 13628
rect 6137 13626 6161 13628
rect 6217 13626 6223 13628
rect 5977 13574 5979 13626
rect 6159 13574 6161 13626
rect 5915 13572 5921 13574
rect 5977 13572 6001 13574
rect 6057 13572 6081 13574
rect 6137 13572 6161 13574
rect 6217 13572 6223 13574
rect 5915 13552 6223 13572
rect 6288 13410 6316 16390
rect 6380 13988 6408 16612
rect 6472 15706 6500 19314
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6472 14822 6500 15302
rect 6564 15026 6592 20198
rect 6656 18290 6684 20334
rect 6748 18952 6776 20742
rect 6840 19922 6868 21082
rect 6932 20942 6960 21508
rect 6920 20936 6972 20942
rect 6972 20896 7052 20924
rect 6920 20878 6972 20884
rect 7024 20534 7052 20896
rect 7104 20868 7156 20874
rect 7104 20810 7156 20816
rect 7012 20528 7064 20534
rect 7012 20470 7064 20476
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 6932 20058 6960 20402
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 7024 19990 7052 20470
rect 7012 19984 7064 19990
rect 7012 19926 7064 19932
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6748 18924 6868 18952
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6644 18080 6696 18086
rect 6644 18022 6696 18028
rect 6656 15706 6684 18022
rect 6748 17202 6776 18634
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6656 15026 6684 15506
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6460 14000 6512 14006
rect 6380 13960 6460 13988
rect 6460 13942 6512 13948
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 5920 13382 6316 13410
rect 5920 13326 5948 13382
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5736 8974 5764 9862
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5828 8786 5856 12786
rect 6104 12714 6132 13262
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 5915 12540 6223 12560
rect 5915 12538 5921 12540
rect 5977 12538 6001 12540
rect 6057 12538 6081 12540
rect 6137 12538 6161 12540
rect 6217 12538 6223 12540
rect 5977 12486 5979 12538
rect 6159 12486 6161 12538
rect 5915 12484 5921 12486
rect 5977 12484 6001 12486
rect 6057 12484 6081 12486
rect 6137 12484 6161 12486
rect 6217 12484 6223 12486
rect 5915 12464 6223 12484
rect 6288 12442 6316 13262
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 5915 11452 6223 11472
rect 5915 11450 5921 11452
rect 5977 11450 6001 11452
rect 6057 11450 6081 11452
rect 6137 11450 6161 11452
rect 6217 11450 6223 11452
rect 5977 11398 5979 11450
rect 6159 11398 6161 11450
rect 5915 11396 5921 11398
rect 5977 11396 6001 11398
rect 6057 11396 6081 11398
rect 6137 11396 6161 11398
rect 6217 11396 6223 11398
rect 5915 11376 6223 11396
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6288 10674 6316 11018
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 5915 10364 6223 10384
rect 5915 10362 5921 10364
rect 5977 10362 6001 10364
rect 6057 10362 6081 10364
rect 6137 10362 6161 10364
rect 6217 10362 6223 10364
rect 5977 10310 5979 10362
rect 6159 10310 6161 10362
rect 5915 10308 5921 10310
rect 5977 10308 6001 10310
rect 6057 10308 6081 10310
rect 6137 10308 6161 10310
rect 6217 10308 6223 10310
rect 5915 10288 6223 10308
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6288 10062 6316 10134
rect 6000 10056 6052 10062
rect 5920 10016 6000 10044
rect 5920 9625 5948 10016
rect 6276 10056 6328 10062
rect 6000 9998 6052 10004
rect 6196 10016 6276 10044
rect 5906 9616 5962 9625
rect 5906 9551 5962 9560
rect 6196 9489 6224 10016
rect 6276 9998 6328 10004
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6182 9480 6238 9489
rect 6182 9415 6238 9424
rect 5915 9276 6223 9296
rect 5915 9274 5921 9276
rect 5977 9274 6001 9276
rect 6057 9274 6081 9276
rect 6137 9274 6161 9276
rect 6217 9274 6223 9276
rect 5977 9222 5979 9274
rect 6159 9222 6161 9274
rect 5915 9220 5921 9222
rect 5977 9220 6001 9222
rect 6057 9220 6081 9222
rect 6137 9220 6161 9222
rect 6217 9220 6223 9222
rect 5915 9200 6223 9220
rect 6288 8906 6316 9862
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 5552 8486 5672 8514
rect 5736 8758 5856 8786
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4816 3942 4844 7686
rect 5092 6662 5120 7754
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5184 6730 5212 7346
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6186 5120 6598
rect 5276 6322 5304 6870
rect 5460 6866 5488 7822
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5092 4078 5120 6122
rect 5276 5370 5304 6258
rect 5368 6254 5396 6734
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5368 5710 5396 6190
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5184 4146 5212 4762
rect 5460 4690 5488 6666
rect 5552 5098 5580 8486
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5644 6798 5672 8366
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5356 4140 5408 4146
rect 5460 4128 5488 4626
rect 5644 4622 5672 6258
rect 5736 6186 5764 8758
rect 5915 8188 6223 8208
rect 5915 8186 5921 8188
rect 5977 8186 6001 8188
rect 6057 8186 6081 8188
rect 6137 8186 6161 8188
rect 6217 8186 6223 8188
rect 5977 8134 5979 8186
rect 6159 8134 6161 8186
rect 5915 8132 5921 8134
rect 5977 8132 6001 8134
rect 6057 8132 6081 8134
rect 6137 8132 6161 8134
rect 6217 8132 6223 8134
rect 5915 8112 6223 8132
rect 5816 8016 5868 8022
rect 5816 7958 5868 7964
rect 5828 7478 5856 7958
rect 6288 7886 6316 8842
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5828 6882 5856 7414
rect 5915 7100 6223 7120
rect 5915 7098 5921 7100
rect 5977 7098 6001 7100
rect 6057 7098 6081 7100
rect 6137 7098 6161 7100
rect 6217 7098 6223 7100
rect 5977 7046 5979 7098
rect 6159 7046 6161 7098
rect 5915 7044 5921 7046
rect 5977 7044 6001 7046
rect 6057 7044 6081 7046
rect 6137 7044 6161 7046
rect 6217 7044 6223 7046
rect 5915 7024 6223 7044
rect 5828 6854 5948 6882
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5828 6168 5856 6734
rect 5920 6730 5948 6854
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 6288 6662 6316 7822
rect 6380 7002 6408 13194
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6090 6352 6146 6361
rect 6288 6322 6316 6598
rect 6090 6287 6092 6296
rect 6144 6287 6146 6296
rect 6276 6316 6328 6322
rect 6092 6258 6144 6264
rect 6276 6258 6328 6264
rect 5908 6180 5960 6186
rect 5828 6140 5908 6168
rect 5828 5846 5856 6140
rect 5908 6122 5960 6128
rect 5915 6012 6223 6032
rect 5915 6010 5921 6012
rect 5977 6010 6001 6012
rect 6057 6010 6081 6012
rect 6137 6010 6161 6012
rect 6217 6010 6223 6012
rect 5977 5958 5979 6010
rect 6159 5958 6161 6010
rect 5915 5956 5921 5958
rect 5977 5956 6001 5958
rect 6057 5956 6081 5958
rect 6137 5956 6161 5958
rect 6217 5956 6223 5958
rect 5915 5936 6223 5956
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6012 5166 6040 5646
rect 6380 5370 6408 6598
rect 6472 5846 6500 13806
rect 6564 10810 6592 14826
rect 6656 13938 6684 14962
rect 6748 14958 6776 15370
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6748 14498 6776 14894
rect 6840 14618 6868 18924
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6932 15026 6960 15914
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6918 14512 6974 14521
rect 6748 14470 6868 14498
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6840 14362 6868 14470
rect 6918 14447 6920 14456
rect 6972 14447 6974 14456
rect 6920 14418 6972 14424
rect 7024 14414 7052 15846
rect 7116 15178 7144 20810
rect 7208 20058 7236 28086
rect 7300 26246 7328 28086
rect 7380 27872 7432 27878
rect 7380 27814 7432 27820
rect 7392 27674 7420 27814
rect 7380 27668 7432 27674
rect 7380 27610 7432 27616
rect 7392 26926 7420 27610
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7288 26240 7340 26246
rect 7288 26182 7340 26188
rect 7288 25492 7340 25498
rect 7288 25434 7340 25440
rect 7300 23866 7328 25434
rect 7392 24818 7420 26862
rect 7484 26432 7512 28562
rect 7564 26988 7616 26994
rect 7564 26930 7616 26936
rect 7576 26586 7604 26930
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 7564 26444 7616 26450
rect 7484 26404 7564 26432
rect 7564 26386 7616 26392
rect 7472 26036 7524 26042
rect 7472 25978 7524 25984
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7392 23866 7420 24142
rect 7288 23860 7340 23866
rect 7288 23802 7340 23808
rect 7380 23860 7432 23866
rect 7380 23802 7432 23808
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7300 23322 7328 23666
rect 7288 23316 7340 23322
rect 7288 23258 7340 23264
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7196 19916 7248 19922
rect 7196 19858 7248 19864
rect 7208 19718 7236 19858
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7300 18086 7328 23122
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 7392 21350 7420 22170
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7392 21010 7420 21286
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7484 18714 7512 25978
rect 7576 25838 7604 26386
rect 7564 25832 7616 25838
rect 7564 25774 7616 25780
rect 7564 25424 7616 25430
rect 7564 25366 7616 25372
rect 7576 24342 7604 25366
rect 7668 24954 7696 29446
rect 7852 29152 7880 31726
rect 8128 31142 8156 33798
rect 8220 33522 8248 34054
rect 8298 34031 8354 34040
rect 8300 33924 8352 33930
rect 8300 33866 8352 33872
rect 8208 33516 8260 33522
rect 8208 33458 8260 33464
rect 8312 33114 8340 33866
rect 8404 33658 8432 35142
rect 8760 35080 8812 35086
rect 8760 35022 8812 35028
rect 8668 34944 8720 34950
rect 8668 34886 8720 34892
rect 8680 34610 8708 34886
rect 8772 34746 8800 35022
rect 8760 34740 8812 34746
rect 8760 34682 8812 34688
rect 8668 34604 8720 34610
rect 8668 34546 8720 34552
rect 8484 34536 8536 34542
rect 8484 34478 8536 34484
rect 8496 33998 8524 34478
rect 8484 33992 8536 33998
rect 8484 33934 8536 33940
rect 8392 33652 8444 33658
rect 8392 33594 8444 33600
rect 8404 33454 8432 33594
rect 8496 33504 8524 33934
rect 8576 33516 8628 33522
rect 8496 33476 8576 33504
rect 8576 33458 8628 33464
rect 8392 33448 8444 33454
rect 8444 33396 8616 33402
rect 8392 33390 8616 33396
rect 8404 33374 8616 33390
rect 8300 33108 8352 33114
rect 8300 33050 8352 33056
rect 8116 31136 8168 31142
rect 8116 31078 8168 31084
rect 8312 30734 8340 33050
rect 8588 31414 8616 33374
rect 8760 33380 8812 33386
rect 8760 33322 8812 33328
rect 8772 32570 8800 33322
rect 8760 32564 8812 32570
rect 8760 32506 8812 32512
rect 8576 31408 8628 31414
rect 8576 31350 8628 31356
rect 8576 31136 8628 31142
rect 8576 31078 8628 31084
rect 8300 30728 8352 30734
rect 8300 30670 8352 30676
rect 8588 30054 8616 31078
rect 8772 30258 8800 32506
rect 8864 31686 8892 35158
rect 8942 34640 8998 34649
rect 8942 34575 8944 34584
rect 8996 34575 8998 34584
rect 8944 34546 8996 34552
rect 9048 34406 9076 38286
rect 9232 37330 9260 38354
rect 9324 38350 9352 38830
rect 9508 38350 9536 39782
rect 9692 38554 9720 39986
rect 9680 38548 9732 38554
rect 9680 38490 9732 38496
rect 9312 38344 9364 38350
rect 9312 38286 9364 38292
rect 9496 38344 9548 38350
rect 9496 38286 9548 38292
rect 9324 38214 9352 38286
rect 9312 38208 9364 38214
rect 9312 38150 9364 38156
rect 9220 37324 9272 37330
rect 9220 37266 9272 37272
rect 9324 37262 9352 38150
rect 9128 37256 9180 37262
rect 9128 37198 9180 37204
rect 9312 37256 9364 37262
rect 9312 37198 9364 37204
rect 9140 35766 9168 37198
rect 9324 36378 9352 37198
rect 9508 36718 9536 38286
rect 9680 38276 9732 38282
rect 9680 38218 9732 38224
rect 9588 37664 9640 37670
rect 9588 37606 9640 37612
rect 9600 37398 9628 37606
rect 9588 37392 9640 37398
rect 9588 37334 9640 37340
rect 9692 37262 9720 38218
rect 9784 37806 9812 42774
rect 9876 42770 9904 44338
rect 9956 44260 10008 44266
rect 9956 44202 10008 44208
rect 9968 43450 9996 44202
rect 15846 44092 16154 44112
rect 15846 44090 15852 44092
rect 15908 44090 15932 44092
rect 15988 44090 16012 44092
rect 16068 44090 16092 44092
rect 16148 44090 16154 44092
rect 15908 44038 15910 44090
rect 16090 44038 16092 44090
rect 15846 44036 15852 44038
rect 15908 44036 15932 44038
rect 15988 44036 16012 44038
rect 16068 44036 16092 44038
rect 16148 44036 16154 44038
rect 15846 44016 16154 44036
rect 20088 43994 20116 44338
rect 25776 44092 26084 44112
rect 25776 44090 25782 44092
rect 25838 44090 25862 44092
rect 25918 44090 25942 44092
rect 25998 44090 26022 44092
rect 26078 44090 26084 44092
rect 25838 44038 25840 44090
rect 26020 44038 26022 44090
rect 25776 44036 25782 44038
rect 25838 44036 25862 44038
rect 25918 44036 25942 44038
rect 25998 44036 26022 44038
rect 26078 44036 26084 44038
rect 25776 44016 26084 44036
rect 20076 43988 20128 43994
rect 20076 43930 20128 43936
rect 29012 43858 29040 45222
rect 30024 44878 30052 46951
rect 30104 45484 30156 45490
rect 30104 45426 30156 45432
rect 30116 44985 30144 45426
rect 30102 44976 30158 44985
rect 30102 44911 30158 44920
rect 30012 44872 30064 44878
rect 30012 44814 30064 44820
rect 29920 44736 29972 44742
rect 29920 44678 29972 44684
rect 29000 43852 29052 43858
rect 29000 43794 29052 43800
rect 29932 43790 29960 44678
rect 10416 43784 10468 43790
rect 10416 43726 10468 43732
rect 20168 43784 20220 43790
rect 20168 43726 20220 43732
rect 29920 43784 29972 43790
rect 29920 43726 29972 43732
rect 10428 43450 10456 43726
rect 10880 43548 11188 43568
rect 10880 43546 10886 43548
rect 10942 43546 10966 43548
rect 11022 43546 11046 43548
rect 11102 43546 11126 43548
rect 11182 43546 11188 43548
rect 10942 43494 10944 43546
rect 11124 43494 11126 43546
rect 10880 43492 10886 43494
rect 10942 43492 10966 43494
rect 11022 43492 11046 43494
rect 11102 43492 11126 43494
rect 11182 43492 11188 43494
rect 10880 43472 11188 43492
rect 9956 43444 10008 43450
rect 9956 43386 10008 43392
rect 10416 43444 10468 43450
rect 10416 43386 10468 43392
rect 15846 43004 16154 43024
rect 15846 43002 15852 43004
rect 15908 43002 15932 43004
rect 15988 43002 16012 43004
rect 16068 43002 16092 43004
rect 16148 43002 16154 43004
rect 15908 42950 15910 43002
rect 16090 42950 16092 43002
rect 15846 42948 15852 42950
rect 15908 42948 15932 42950
rect 15988 42948 16012 42950
rect 16068 42948 16092 42950
rect 16148 42948 16154 42950
rect 15846 42928 16154 42948
rect 9864 42764 9916 42770
rect 9864 42706 9916 42712
rect 9876 41414 9904 42706
rect 20180 42634 20208 43726
rect 20811 43548 21119 43568
rect 20811 43546 20817 43548
rect 20873 43546 20897 43548
rect 20953 43546 20977 43548
rect 21033 43546 21057 43548
rect 21113 43546 21119 43548
rect 20873 43494 20875 43546
rect 21055 43494 21057 43546
rect 20811 43492 20817 43494
rect 20873 43492 20897 43494
rect 20953 43492 20977 43494
rect 21033 43492 21057 43494
rect 21113 43492 21119 43494
rect 20811 43472 21119 43492
rect 30104 43308 30156 43314
rect 30104 43250 30156 43256
rect 29920 43104 29972 43110
rect 29920 43046 29972 43052
rect 25776 43004 26084 43024
rect 25776 43002 25782 43004
rect 25838 43002 25862 43004
rect 25918 43002 25942 43004
rect 25998 43002 26022 43004
rect 26078 43002 26084 43004
rect 25838 42950 25840 43002
rect 26020 42950 26022 43002
rect 25776 42948 25782 42950
rect 25838 42948 25862 42950
rect 25918 42948 25942 42950
rect 25998 42948 26022 42950
rect 26078 42948 26084 42950
rect 25776 42928 26084 42948
rect 29932 42702 29960 43046
rect 30116 42945 30144 43250
rect 30102 42936 30158 42945
rect 30102 42871 30158 42880
rect 29920 42696 29972 42702
rect 29920 42638 29972 42644
rect 20168 42628 20220 42634
rect 20168 42570 20220 42576
rect 10232 42560 10284 42566
rect 10232 42502 10284 42508
rect 10244 41546 10272 42502
rect 10880 42460 11188 42480
rect 10880 42458 10886 42460
rect 10942 42458 10966 42460
rect 11022 42458 11046 42460
rect 11102 42458 11126 42460
rect 11182 42458 11188 42460
rect 10942 42406 10944 42458
rect 11124 42406 11126 42458
rect 10880 42404 10886 42406
rect 10942 42404 10966 42406
rect 11022 42404 11046 42406
rect 11102 42404 11126 42406
rect 11182 42404 11188 42406
rect 10880 42384 11188 42404
rect 15846 41916 16154 41936
rect 15846 41914 15852 41916
rect 15908 41914 15932 41916
rect 15988 41914 16012 41916
rect 16068 41914 16092 41916
rect 16148 41914 16154 41916
rect 15908 41862 15910 41914
rect 16090 41862 16092 41914
rect 15846 41860 15852 41862
rect 15908 41860 15932 41862
rect 15988 41860 16012 41862
rect 16068 41860 16092 41862
rect 16148 41860 16154 41862
rect 15846 41840 16154 41860
rect 10232 41540 10284 41546
rect 10232 41482 10284 41488
rect 9876 41386 9996 41414
rect 9864 40112 9916 40118
rect 9864 40054 9916 40060
rect 9772 37800 9824 37806
rect 9772 37742 9824 37748
rect 9876 37652 9904 40054
rect 9784 37624 9904 37652
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 9784 36718 9812 37624
rect 9496 36712 9548 36718
rect 9496 36654 9548 36660
rect 9772 36712 9824 36718
rect 9772 36654 9824 36660
rect 9312 36372 9364 36378
rect 9312 36314 9364 36320
rect 9680 36304 9732 36310
rect 9680 36246 9732 36252
rect 9404 35828 9456 35834
rect 9404 35770 9456 35776
rect 9128 35760 9180 35766
rect 9128 35702 9180 35708
rect 9036 34400 9088 34406
rect 9036 34342 9088 34348
rect 8944 34196 8996 34202
rect 8944 34138 8996 34144
rect 8956 34066 8984 34138
rect 8944 34060 8996 34066
rect 8944 34002 8996 34008
rect 8956 33454 8984 34002
rect 9048 33862 9076 34342
rect 9312 33992 9364 33998
rect 9312 33934 9364 33940
rect 9036 33856 9088 33862
rect 9036 33798 9088 33804
rect 9324 33590 9352 33934
rect 9312 33584 9364 33590
rect 9312 33526 9364 33532
rect 8944 33448 8996 33454
rect 8944 33390 8996 33396
rect 9324 32910 9352 33526
rect 9312 32904 9364 32910
rect 9312 32846 9364 32852
rect 8852 31680 8904 31686
rect 8852 31622 8904 31628
rect 8864 30870 8892 31622
rect 9416 31346 9444 35770
rect 9692 33946 9720 36246
rect 9784 34134 9812 36654
rect 9968 35306 9996 41386
rect 10140 37868 10192 37874
rect 10140 37810 10192 37816
rect 10048 37732 10100 37738
rect 10048 37674 10100 37680
rect 10060 37126 10088 37674
rect 10048 37120 10100 37126
rect 10048 37062 10100 37068
rect 10060 36242 10088 37062
rect 10152 36786 10180 37810
rect 10140 36780 10192 36786
rect 10140 36722 10192 36728
rect 10048 36236 10100 36242
rect 10048 36178 10100 36184
rect 10048 35692 10100 35698
rect 10152 35680 10180 36722
rect 10244 35698 10272 41482
rect 10880 41372 11188 41392
rect 10880 41370 10886 41372
rect 10942 41370 10966 41372
rect 11022 41370 11046 41372
rect 11102 41370 11126 41372
rect 11182 41370 11188 41372
rect 10942 41318 10944 41370
rect 11124 41318 11126 41370
rect 10880 41316 10886 41318
rect 10942 41316 10966 41318
rect 11022 41316 11046 41318
rect 11102 41316 11126 41318
rect 11182 41316 11188 41318
rect 10880 41296 11188 41316
rect 16212 41132 16264 41138
rect 16212 41074 16264 41080
rect 16856 41132 16908 41138
rect 16856 41074 16908 41080
rect 15846 40828 16154 40848
rect 15846 40826 15852 40828
rect 15908 40826 15932 40828
rect 15988 40826 16012 40828
rect 16068 40826 16092 40828
rect 16148 40826 16154 40828
rect 15908 40774 15910 40826
rect 16090 40774 16092 40826
rect 15846 40772 15852 40774
rect 15908 40772 15932 40774
rect 15988 40772 16012 40774
rect 16068 40772 16092 40774
rect 16148 40772 16154 40774
rect 15846 40752 16154 40772
rect 15120 40594 15240 40610
rect 15108 40588 15240 40594
rect 15160 40582 15240 40588
rect 15108 40530 15160 40536
rect 12164 40520 12216 40526
rect 12164 40462 12216 40468
rect 12992 40520 13044 40526
rect 12992 40462 13044 40468
rect 14464 40520 14516 40526
rect 14464 40462 14516 40468
rect 14648 40520 14700 40526
rect 14648 40462 14700 40468
rect 10416 40384 10468 40390
rect 10416 40326 10468 40332
rect 10428 40050 10456 40326
rect 10880 40284 11188 40304
rect 10880 40282 10886 40284
rect 10942 40282 10966 40284
rect 11022 40282 11046 40284
rect 11102 40282 11126 40284
rect 11182 40282 11188 40284
rect 10942 40230 10944 40282
rect 11124 40230 11126 40282
rect 10880 40228 10886 40230
rect 10942 40228 10966 40230
rect 11022 40228 11046 40230
rect 11102 40228 11126 40230
rect 11182 40228 11188 40230
rect 10880 40208 11188 40228
rect 12176 40186 12204 40462
rect 12532 40384 12584 40390
rect 12532 40326 12584 40332
rect 12164 40180 12216 40186
rect 12164 40122 12216 40128
rect 12544 40050 12572 40326
rect 10416 40044 10468 40050
rect 10416 39986 10468 39992
rect 12532 40044 12584 40050
rect 12532 39986 12584 39992
rect 10880 39196 11188 39216
rect 10880 39194 10886 39196
rect 10942 39194 10966 39196
rect 11022 39194 11046 39196
rect 11102 39194 11126 39196
rect 11182 39194 11188 39196
rect 10942 39142 10944 39194
rect 11124 39142 11126 39194
rect 10880 39140 10886 39142
rect 10942 39140 10966 39142
rect 11022 39140 11046 39142
rect 11102 39140 11126 39142
rect 11182 39140 11188 39142
rect 10880 39120 11188 39140
rect 12544 38962 12572 39986
rect 12624 39908 12676 39914
rect 12624 39850 12676 39856
rect 12636 39370 12664 39850
rect 13004 39642 13032 40462
rect 13544 40384 13596 40390
rect 13544 40326 13596 40332
rect 13176 40180 13228 40186
rect 13176 40122 13228 40128
rect 12992 39636 13044 39642
rect 12992 39578 13044 39584
rect 12624 39364 12676 39370
rect 12624 39306 12676 39312
rect 11428 38956 11480 38962
rect 11428 38898 11480 38904
rect 12532 38956 12584 38962
rect 12532 38898 12584 38904
rect 10600 38752 10652 38758
rect 10600 38694 10652 38700
rect 10416 38344 10468 38350
rect 10416 38286 10468 38292
rect 10324 37936 10376 37942
rect 10324 37878 10376 37884
rect 10336 36786 10364 37878
rect 10324 36780 10376 36786
rect 10324 36722 10376 36728
rect 10336 36258 10364 36722
rect 10428 36582 10456 38286
rect 10508 37800 10560 37806
rect 10508 37742 10560 37748
rect 10520 36786 10548 37742
rect 10612 37262 10640 38694
rect 10880 38108 11188 38128
rect 10880 38106 10886 38108
rect 10942 38106 10966 38108
rect 11022 38106 11046 38108
rect 11102 38106 11126 38108
rect 11182 38106 11188 38108
rect 10942 38054 10944 38106
rect 11124 38054 11126 38106
rect 10880 38052 10886 38054
rect 10942 38052 10966 38054
rect 11022 38052 11046 38054
rect 11102 38052 11126 38054
rect 11182 38052 11188 38054
rect 10880 38032 11188 38052
rect 11244 37936 11296 37942
rect 11244 37878 11296 37884
rect 10876 37664 10928 37670
rect 10876 37606 10928 37612
rect 10888 37262 10916 37606
rect 10600 37256 10652 37262
rect 10600 37198 10652 37204
rect 10876 37256 10928 37262
rect 10876 37198 10928 37204
rect 10880 37020 11188 37040
rect 10880 37018 10886 37020
rect 10942 37018 10966 37020
rect 11022 37018 11046 37020
rect 11102 37018 11126 37020
rect 11182 37018 11188 37020
rect 10942 36966 10944 37018
rect 11124 36966 11126 37018
rect 10880 36964 10886 36966
rect 10942 36964 10966 36966
rect 11022 36964 11046 36966
rect 11102 36964 11126 36966
rect 11182 36964 11188 36966
rect 10880 36944 11188 36964
rect 11256 36922 11284 37878
rect 11336 37188 11388 37194
rect 11336 37130 11388 37136
rect 11244 36916 11296 36922
rect 11244 36858 11296 36864
rect 10508 36780 10560 36786
rect 10508 36722 10560 36728
rect 10784 36780 10836 36786
rect 10784 36722 10836 36728
rect 10416 36576 10468 36582
rect 10416 36518 10468 36524
rect 10336 36230 10456 36258
rect 10324 36168 10376 36174
rect 10324 36110 10376 36116
rect 10100 35652 10180 35680
rect 10048 35634 10100 35640
rect 10152 35494 10180 35652
rect 10232 35692 10284 35698
rect 10232 35634 10284 35640
rect 10140 35488 10192 35494
rect 10140 35430 10192 35436
rect 9968 35278 10272 35306
rect 10336 35290 10364 36110
rect 10428 35766 10456 36230
rect 10416 35760 10468 35766
rect 10416 35702 10468 35708
rect 9956 35148 10008 35154
rect 9956 35090 10008 35096
rect 9864 34536 9916 34542
rect 9864 34478 9916 34484
rect 9876 34202 9904 34478
rect 9864 34196 9916 34202
rect 9864 34138 9916 34144
rect 9772 34128 9824 34134
rect 9772 34070 9824 34076
rect 9588 33924 9640 33930
rect 9692 33918 9904 33946
rect 9588 33866 9640 33872
rect 9496 33856 9548 33862
rect 9496 33798 9548 33804
rect 9508 33590 9536 33798
rect 9496 33584 9548 33590
rect 9496 33526 9548 33532
rect 9600 32910 9628 33866
rect 9772 33516 9824 33522
rect 9772 33458 9824 33464
rect 9680 32972 9732 32978
rect 9680 32914 9732 32920
rect 9588 32904 9640 32910
rect 9588 32846 9640 32852
rect 9692 32042 9720 32914
rect 9784 32570 9812 33458
rect 9876 32756 9904 33918
rect 9968 33522 9996 35090
rect 10140 34536 10192 34542
rect 10140 34478 10192 34484
rect 10152 33522 10180 34478
rect 9956 33516 10008 33522
rect 9956 33458 10008 33464
rect 10140 33516 10192 33522
rect 10140 33458 10192 33464
rect 9968 33046 9996 33458
rect 10048 33448 10100 33454
rect 10046 33416 10048 33425
rect 10100 33416 10102 33425
rect 10046 33351 10102 33360
rect 10060 33114 10088 33351
rect 10048 33108 10100 33114
rect 10048 33050 10100 33056
rect 9956 33040 10008 33046
rect 9956 32982 10008 32988
rect 9956 32904 10008 32910
rect 10152 32892 10180 33458
rect 10008 32864 10180 32892
rect 9956 32846 10008 32852
rect 9876 32728 9996 32756
rect 9772 32564 9824 32570
rect 9772 32506 9824 32512
rect 9508 32014 9720 32042
rect 9508 31754 9536 32014
rect 9680 31884 9732 31890
rect 9680 31826 9732 31832
rect 9496 31748 9548 31754
rect 9496 31690 9548 31696
rect 9692 31634 9720 31826
rect 9784 31822 9812 32506
rect 9864 32020 9916 32026
rect 9864 31962 9916 31968
rect 9772 31816 9824 31822
rect 9772 31758 9824 31764
rect 9692 31606 9812 31634
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 9404 31340 9456 31346
rect 9404 31282 9456 31288
rect 9312 31272 9364 31278
rect 9312 31214 9364 31220
rect 8852 30864 8904 30870
rect 8852 30806 8904 30812
rect 8944 30592 8996 30598
rect 8944 30534 8996 30540
rect 8760 30252 8812 30258
rect 8760 30194 8812 30200
rect 8208 30048 8260 30054
rect 8208 29990 8260 29996
rect 8576 30048 8628 30054
rect 8576 29990 8628 29996
rect 8220 29170 8248 29990
rect 8852 29844 8904 29850
rect 8852 29786 8904 29792
rect 8576 29300 8628 29306
rect 8576 29242 8628 29248
rect 7760 29124 7880 29152
rect 8208 29164 8260 29170
rect 7760 25906 7788 29124
rect 8208 29106 8260 29112
rect 7840 29028 7892 29034
rect 7840 28970 7892 28976
rect 8392 29028 8444 29034
rect 8392 28970 8444 28976
rect 7852 26382 7880 28970
rect 8404 28558 8432 28970
rect 8392 28552 8444 28558
rect 8392 28494 8444 28500
rect 8024 28416 8076 28422
rect 8024 28358 8076 28364
rect 8036 28218 8064 28358
rect 8024 28212 8076 28218
rect 8024 28154 8076 28160
rect 7932 28076 7984 28082
rect 8116 28076 8168 28082
rect 7984 28036 8116 28064
rect 7932 28018 7984 28024
rect 8116 28018 8168 28024
rect 8484 28076 8536 28082
rect 8484 28018 8536 28024
rect 8208 28008 8260 28014
rect 8260 27968 8432 27996
rect 8208 27950 8260 27956
rect 8116 27940 8168 27946
rect 8116 27882 8168 27888
rect 7930 27704 7986 27713
rect 7930 27639 7986 27648
rect 7944 26994 7972 27639
rect 7932 26988 7984 26994
rect 7932 26930 7984 26936
rect 7944 26858 7972 26930
rect 8128 26926 8156 27882
rect 8404 27606 8432 27968
rect 8392 27600 8444 27606
rect 8392 27542 8444 27548
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8404 27130 8432 27270
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8116 26920 8168 26926
rect 8116 26862 8168 26868
rect 7932 26852 7984 26858
rect 7932 26794 7984 26800
rect 8024 26852 8076 26858
rect 8024 26794 8076 26800
rect 7932 26580 7984 26586
rect 7932 26522 7984 26528
rect 7944 26382 7972 26522
rect 7840 26376 7892 26382
rect 7840 26318 7892 26324
rect 7932 26376 7984 26382
rect 7932 26318 7984 26324
rect 7932 26240 7984 26246
rect 7932 26182 7984 26188
rect 7748 25900 7800 25906
rect 7944 25888 7972 26182
rect 8036 26042 8064 26794
rect 8024 26036 8076 26042
rect 8024 25978 8076 25984
rect 8024 25900 8076 25906
rect 7944 25860 8024 25888
rect 7748 25842 7800 25848
rect 8024 25842 8076 25848
rect 7840 25832 7892 25838
rect 7840 25774 7892 25780
rect 7852 25498 7880 25774
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 7840 25492 7892 25498
rect 7840 25434 7892 25440
rect 7656 24948 7708 24954
rect 7656 24890 7708 24896
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7564 24336 7616 24342
rect 7564 24278 7616 24284
rect 7668 24188 7696 24754
rect 7852 24750 7880 25434
rect 7944 25362 7972 25638
rect 7932 25356 7984 25362
rect 7932 25298 7984 25304
rect 7748 24744 7800 24750
rect 7748 24686 7800 24692
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7760 24410 7788 24686
rect 7748 24404 7800 24410
rect 7748 24346 7800 24352
rect 7748 24200 7800 24206
rect 7668 24160 7748 24188
rect 7748 24142 7800 24148
rect 7564 23792 7616 23798
rect 7564 23734 7616 23740
rect 7576 22166 7604 23734
rect 7656 23316 7708 23322
rect 7656 23258 7708 23264
rect 7564 22160 7616 22166
rect 7564 22102 7616 22108
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7576 21622 7604 21966
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7668 21350 7696 23258
rect 7760 21690 7788 24142
rect 7852 23186 7880 24686
rect 7944 23526 7972 25298
rect 8036 25226 8064 25842
rect 8024 25220 8076 25226
rect 8024 25162 8076 25168
rect 8036 23730 8064 25162
rect 8128 24614 8156 26862
rect 8220 25838 8248 27066
rect 8392 26512 8444 26518
rect 8392 26454 8444 26460
rect 8208 25832 8260 25838
rect 8208 25774 8260 25780
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8128 24274 8156 24550
rect 8116 24268 8168 24274
rect 8116 24210 8168 24216
rect 8024 23724 8076 23730
rect 8024 23666 8076 23672
rect 7932 23520 7984 23526
rect 7932 23462 7984 23468
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 7852 22642 7880 22918
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7944 22574 7972 23462
rect 8036 23338 8064 23666
rect 8128 23508 8156 24210
rect 8220 23730 8248 25094
rect 8208 23724 8260 23730
rect 8208 23666 8260 23672
rect 8128 23480 8340 23508
rect 8036 23310 8156 23338
rect 8024 22976 8076 22982
rect 8024 22918 8076 22924
rect 7932 22568 7984 22574
rect 7932 22510 7984 22516
rect 7930 21992 7986 22001
rect 7930 21927 7986 21936
rect 7840 21888 7892 21894
rect 7838 21856 7840 21865
rect 7892 21856 7894 21865
rect 7838 21791 7894 21800
rect 7838 21720 7894 21729
rect 7748 21684 7800 21690
rect 7838 21655 7894 21664
rect 7748 21626 7800 21632
rect 7852 21486 7880 21655
rect 7840 21480 7892 21486
rect 7840 21422 7892 21428
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7656 20324 7708 20330
rect 7656 20266 7708 20272
rect 7668 18766 7696 20266
rect 7852 19334 7880 21422
rect 7944 21078 7972 21927
rect 7932 21072 7984 21078
rect 7932 21014 7984 21020
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 7944 20330 7972 20878
rect 8036 20602 8064 22918
rect 8128 22273 8156 23310
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8114 22264 8170 22273
rect 8114 22199 8170 22208
rect 8116 22160 8168 22166
rect 8116 22102 8168 22108
rect 8024 20596 8076 20602
rect 8024 20538 8076 20544
rect 7932 20324 7984 20330
rect 7932 20266 7984 20272
rect 8036 19938 8064 20538
rect 7944 19910 8064 19938
rect 7944 19854 7972 19910
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 8036 19718 8064 19790
rect 8024 19712 8076 19718
rect 8024 19654 8076 19660
rect 7760 19306 7880 19334
rect 7392 18686 7512 18714
rect 7656 18760 7708 18766
rect 7656 18702 7708 18708
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7196 17196 7248 17202
rect 7248 17156 7328 17184
rect 7196 17138 7248 17144
rect 7194 16280 7250 16289
rect 7194 16215 7196 16224
rect 7248 16215 7250 16224
rect 7196 16186 7248 16192
rect 7208 15910 7236 16186
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7116 15150 7236 15178
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7116 14482 7144 14962
rect 7208 14618 7236 15150
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7012 14408 7064 14414
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6656 13394 6684 13874
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6656 12850 6684 13330
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6564 10470 6592 10610
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6656 10130 6684 10610
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6564 9586 6592 9930
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6564 8566 6592 9522
rect 6656 9178 6684 10066
rect 6748 9450 6776 14350
rect 6840 14334 6960 14362
rect 7116 14385 7144 14418
rect 7196 14408 7248 14414
rect 7012 14350 7064 14356
rect 7102 14376 7158 14385
rect 6826 13968 6882 13977
rect 6932 13954 6960 14334
rect 7196 14350 7248 14356
rect 7102 14311 7158 14320
rect 6932 13926 7052 13954
rect 6826 13903 6828 13912
rect 6880 13903 6882 13912
rect 6828 13874 6880 13880
rect 7024 13870 7052 13926
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7208 13376 7236 14350
rect 7116 13348 7236 13376
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6932 11898 6960 12786
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 7024 11218 7052 13126
rect 7116 12442 7144 13348
rect 7196 13252 7248 13258
rect 7196 13194 7248 13200
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7208 12306 7236 13194
rect 7300 12434 7328 17156
rect 7392 15434 7420 18686
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 7484 18358 7512 18566
rect 7668 18426 7696 18702
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 7564 18352 7616 18358
rect 7564 18294 7616 18300
rect 7472 17604 7524 17610
rect 7472 17546 7524 17552
rect 7484 17338 7512 17546
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7392 15162 7420 15370
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7392 14414 7420 14554
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7392 13394 7420 13670
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7300 12406 7420 12434
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 7300 11150 7328 11494
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6932 9908 6960 10746
rect 7208 10062 7236 11018
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6840 9880 6960 9908
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6840 9178 6868 9880
rect 7024 9586 7052 9930
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6840 8498 6868 9114
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6564 7886 6592 8366
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6748 7886 6776 8026
rect 6552 7880 6604 7886
rect 6736 7880 6788 7886
rect 6552 7822 6604 7828
rect 6656 7828 6736 7834
rect 6656 7822 6788 7828
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6564 7426 6592 7822
rect 6656 7806 6776 7822
rect 6656 7750 6684 7806
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6564 7410 6684 7426
rect 6564 7404 6696 7410
rect 6564 7398 6644 7404
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5915 4924 6223 4944
rect 5915 4922 5921 4924
rect 5977 4922 6001 4924
rect 6057 4922 6081 4924
rect 6137 4922 6161 4924
rect 6217 4922 6223 4924
rect 5977 4870 5979 4922
rect 6159 4870 6161 4922
rect 5915 4868 5921 4870
rect 5977 4868 6001 4870
rect 6057 4868 6081 4870
rect 6137 4868 6161 4870
rect 6217 4868 6223 4870
rect 5915 4848 6223 4868
rect 6472 4826 6500 5170
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 5920 4622 5948 4694
rect 6564 4622 6592 7398
rect 6644 7346 6696 7352
rect 6748 7018 6776 7686
rect 6840 7342 6868 7822
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6656 6990 6776 7018
rect 6656 6662 6684 6990
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6748 6322 6776 6802
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6840 5930 6868 7278
rect 6920 6792 6972 6798
rect 7024 6780 7052 9522
rect 7116 8838 7144 9590
rect 7392 9382 7420 12406
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 7886 7144 8774
rect 7300 8090 7328 8842
rect 7484 8106 7512 16118
rect 7576 15178 7604 18294
rect 7656 17672 7708 17678
rect 7760 17660 7788 19306
rect 8036 18850 8064 19654
rect 7944 18822 8064 18850
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7708 17632 7788 17660
rect 7656 17614 7708 17620
rect 7668 15638 7696 17614
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7668 15366 7696 15438
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7576 15150 7696 15178
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7576 14006 7604 14214
rect 7564 14000 7616 14006
rect 7564 13942 7616 13948
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7576 12714 7604 13806
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7576 12306 7604 12650
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7576 10470 7604 11630
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7576 8566 7604 9318
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7392 8078 7512 8106
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7208 7410 7236 7686
rect 7392 7478 7420 8078
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7472 7404 7524 7410
rect 7668 7392 7696 15150
rect 7760 12238 7788 16390
rect 7852 13870 7880 18022
rect 7944 17882 7972 18822
rect 8024 18760 8076 18766
rect 8128 18748 8156 22102
rect 8220 22098 8248 22578
rect 8312 22574 8340 23480
rect 8300 22568 8352 22574
rect 8300 22510 8352 22516
rect 8312 22098 8340 22510
rect 8404 22234 8432 26454
rect 8392 22228 8444 22234
rect 8392 22170 8444 22176
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 8300 21956 8352 21962
rect 8300 21898 8352 21904
rect 8206 21720 8262 21729
rect 8206 21655 8208 21664
rect 8260 21655 8262 21664
rect 8208 21626 8260 21632
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8220 21146 8248 21490
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8220 19990 8248 21082
rect 8312 20466 8340 21898
rect 8392 21412 8444 21418
rect 8392 21354 8444 21360
rect 8404 20602 8432 21354
rect 8496 21146 8524 28018
rect 8588 27402 8616 29242
rect 8864 28994 8892 29786
rect 8956 29646 8984 30534
rect 8944 29640 8996 29646
rect 8944 29582 8996 29588
rect 9128 29504 9180 29510
rect 9128 29446 9180 29452
rect 9140 29306 9168 29446
rect 9128 29300 9180 29306
rect 9128 29242 9180 29248
rect 9220 29096 9272 29102
rect 9220 29038 9272 29044
rect 8864 28966 8984 28994
rect 8760 28212 8812 28218
rect 8760 28154 8812 28160
rect 8666 27568 8722 27577
rect 8666 27503 8722 27512
rect 8680 27470 8708 27503
rect 8668 27464 8720 27470
rect 8668 27406 8720 27412
rect 8576 27396 8628 27402
rect 8576 27338 8628 27344
rect 8668 26444 8720 26450
rect 8668 26386 8720 26392
rect 8680 26353 8708 26386
rect 8666 26344 8722 26353
rect 8666 26279 8722 26288
rect 8576 25152 8628 25158
rect 8576 25094 8628 25100
rect 8588 24818 8616 25094
rect 8576 24812 8628 24818
rect 8576 24754 8628 24760
rect 8576 24064 8628 24070
rect 8576 24006 8628 24012
rect 8588 23798 8616 24006
rect 8576 23792 8628 23798
rect 8576 23734 8628 23740
rect 8588 22137 8616 23734
rect 8668 23588 8720 23594
rect 8668 23530 8720 23536
rect 8680 22166 8708 23530
rect 8668 22160 8720 22166
rect 8574 22128 8630 22137
rect 8668 22102 8720 22108
rect 8574 22063 8630 22072
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8392 20596 8444 20602
rect 8392 20538 8444 20544
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8208 19984 8260 19990
rect 8208 19926 8260 19932
rect 8076 18720 8156 18748
rect 8024 18702 8076 18708
rect 8036 18358 8064 18702
rect 8024 18352 8076 18358
rect 8024 18294 8076 18300
rect 7932 17876 7984 17882
rect 7932 17818 7984 17824
rect 7944 17202 7972 17818
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 7932 15428 7984 15434
rect 7932 15370 7984 15376
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7944 7886 7972 15370
rect 8128 15366 8156 16050
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 8036 14550 8064 14758
rect 8128 14618 8156 15302
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8024 14544 8076 14550
rect 8024 14486 8076 14492
rect 8128 14482 8156 14554
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8312 14346 8340 20402
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8404 19446 8432 19790
rect 8392 19440 8444 19446
rect 8392 19382 8444 19388
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8404 17202 8432 18702
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8496 14346 8524 20946
rect 8300 14340 8352 14346
rect 8484 14340 8536 14346
rect 8352 14300 8432 14328
rect 8300 14282 8352 14288
rect 8404 13870 8432 14300
rect 8484 14282 8536 14288
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8036 12782 8064 13738
rect 8220 13326 8248 13738
rect 8496 13410 8524 14282
rect 8312 13382 8524 13410
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8312 13002 8340 13382
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8220 12974 8340 13002
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 8036 11286 8064 12718
rect 8220 12306 8248 12974
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8128 9586 8156 10610
rect 8312 10538 8340 12854
rect 8404 12102 8432 13126
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8496 11762 8524 13262
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8496 11354 8524 11698
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 8312 9654 8340 10474
rect 8588 10266 8616 21830
rect 8668 21412 8720 21418
rect 8668 21354 8720 21360
rect 8680 20806 8708 21354
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8772 19854 8800 28154
rect 8852 27328 8904 27334
rect 8852 27270 8904 27276
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 8772 18426 8800 19314
rect 8864 18698 8892 27270
rect 8956 26994 8984 28966
rect 9036 28416 9088 28422
rect 9036 28358 9088 28364
rect 9048 28082 9076 28358
rect 9232 28218 9260 29038
rect 9324 28558 9352 31214
rect 9404 30592 9456 30598
rect 9404 30534 9456 30540
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 9416 28234 9444 30534
rect 9692 30258 9720 31418
rect 9680 30252 9732 30258
rect 9680 30194 9732 30200
rect 9692 28626 9720 30194
rect 9784 29646 9812 31606
rect 9876 31142 9904 31962
rect 9864 31136 9916 31142
rect 9864 31078 9916 31084
rect 9876 30938 9904 31078
rect 9864 30932 9916 30938
rect 9864 30874 9916 30880
rect 9968 30734 9996 32728
rect 10048 32224 10100 32230
rect 10048 32166 10100 32172
rect 10060 31822 10088 32166
rect 10244 31890 10272 35278
rect 10324 35284 10376 35290
rect 10324 35226 10376 35232
rect 10428 34542 10456 35702
rect 10520 35562 10548 36722
rect 10796 36582 10824 36722
rect 11348 36582 11376 37130
rect 11440 36922 11468 38898
rect 12636 38894 12664 39306
rect 12624 38888 12676 38894
rect 12624 38830 12676 38836
rect 13188 38826 13216 40122
rect 13556 39930 13584 40326
rect 13636 39976 13688 39982
rect 13556 39924 13636 39930
rect 13556 39918 13688 39924
rect 13820 39976 13872 39982
rect 13872 39924 13952 39930
rect 13820 39918 13952 39924
rect 13268 39908 13320 39914
rect 13268 39850 13320 39856
rect 13556 39902 13676 39918
rect 13832 39902 13952 39918
rect 13280 39574 13308 39850
rect 13360 39840 13412 39846
rect 13360 39782 13412 39788
rect 13268 39568 13320 39574
rect 13268 39510 13320 39516
rect 13372 38944 13400 39782
rect 13452 38956 13504 38962
rect 13372 38916 13452 38944
rect 13268 38888 13320 38894
rect 13268 38830 13320 38836
rect 13176 38820 13228 38826
rect 13176 38762 13228 38768
rect 13280 38486 13308 38830
rect 13372 38486 13400 38916
rect 13452 38898 13504 38904
rect 13556 38894 13584 39902
rect 13728 39432 13780 39438
rect 13728 39374 13780 39380
rect 13544 38888 13596 38894
rect 13544 38830 13596 38836
rect 13268 38480 13320 38486
rect 13268 38422 13320 38428
rect 13360 38480 13412 38486
rect 13360 38422 13412 38428
rect 12716 38344 12768 38350
rect 12716 38286 12768 38292
rect 11520 38208 11572 38214
rect 11520 38150 11572 38156
rect 11532 37874 11560 38150
rect 11520 37868 11572 37874
rect 11520 37810 11572 37816
rect 12440 37664 12492 37670
rect 12440 37606 12492 37612
rect 11428 36916 11480 36922
rect 11428 36858 11480 36864
rect 12452 36786 12480 37606
rect 12728 37466 12756 38286
rect 13280 38214 13308 38422
rect 13360 38344 13412 38350
rect 13360 38286 13412 38292
rect 13268 38208 13320 38214
rect 13268 38150 13320 38156
rect 13372 37806 13400 38286
rect 13556 38282 13584 38830
rect 13740 38554 13768 39374
rect 13924 38894 13952 39902
rect 14476 39438 14504 40462
rect 14660 39506 14688 40462
rect 15212 40390 15240 40582
rect 15476 40520 15528 40526
rect 15476 40462 15528 40468
rect 15200 40384 15252 40390
rect 15200 40326 15252 40332
rect 15212 40186 15240 40326
rect 15200 40180 15252 40186
rect 15200 40122 15252 40128
rect 15200 39976 15252 39982
rect 15200 39918 15252 39924
rect 14648 39500 14700 39506
rect 14648 39442 14700 39448
rect 14464 39432 14516 39438
rect 14464 39374 14516 39380
rect 13912 38888 13964 38894
rect 13912 38830 13964 38836
rect 13728 38548 13780 38554
rect 13728 38490 13780 38496
rect 14372 38412 14424 38418
rect 14372 38354 14424 38360
rect 14280 38344 14332 38350
rect 14280 38286 14332 38292
rect 13544 38276 13596 38282
rect 13544 38218 13596 38224
rect 14292 38010 14320 38286
rect 14280 38004 14332 38010
rect 14280 37946 14332 37952
rect 14384 37874 14412 38354
rect 14476 38010 14504 39374
rect 14832 39296 14884 39302
rect 14832 39238 14884 39244
rect 14844 38962 14872 39238
rect 15212 39098 15240 39918
rect 15488 39846 15516 40462
rect 15752 40384 15804 40390
rect 15752 40326 15804 40332
rect 15476 39840 15528 39846
rect 15476 39782 15528 39788
rect 15488 39506 15516 39782
rect 15660 39636 15712 39642
rect 15660 39578 15712 39584
rect 15476 39500 15528 39506
rect 15476 39442 15528 39448
rect 15200 39092 15252 39098
rect 15200 39034 15252 39040
rect 15672 38962 15700 39578
rect 14832 38956 14884 38962
rect 14832 38898 14884 38904
rect 15660 38956 15712 38962
rect 15660 38898 15712 38904
rect 14464 38004 14516 38010
rect 14464 37946 14516 37952
rect 13820 37868 13872 37874
rect 13820 37810 13872 37816
rect 14188 37868 14240 37874
rect 14188 37810 14240 37816
rect 14372 37868 14424 37874
rect 14372 37810 14424 37816
rect 12992 37800 13044 37806
rect 12992 37742 13044 37748
rect 13360 37800 13412 37806
rect 13360 37742 13412 37748
rect 12900 37664 12952 37670
rect 12900 37606 12952 37612
rect 12716 37460 12768 37466
rect 12716 37402 12768 37408
rect 12912 36854 12940 37606
rect 13004 37262 13032 37742
rect 13728 37664 13780 37670
rect 13728 37606 13780 37612
rect 12992 37256 13044 37262
rect 12992 37198 13044 37204
rect 13084 37256 13136 37262
rect 13084 37198 13136 37204
rect 12900 36848 12952 36854
rect 12900 36790 12952 36796
rect 12440 36780 12492 36786
rect 12440 36722 12492 36728
rect 11888 36712 11940 36718
rect 11888 36654 11940 36660
rect 10784 36576 10836 36582
rect 10784 36518 10836 36524
rect 11336 36576 11388 36582
rect 11336 36518 11388 36524
rect 10692 36100 10744 36106
rect 10692 36042 10744 36048
rect 10600 36032 10652 36038
rect 10600 35974 10652 35980
rect 10612 35766 10640 35974
rect 10704 35834 10732 36042
rect 10692 35828 10744 35834
rect 10692 35770 10744 35776
rect 10600 35760 10652 35766
rect 10600 35702 10652 35708
rect 10508 35556 10560 35562
rect 10508 35498 10560 35504
rect 10520 35154 10548 35498
rect 10508 35148 10560 35154
rect 10508 35090 10560 35096
rect 10796 35086 10824 36518
rect 10880 35932 11188 35952
rect 10880 35930 10886 35932
rect 10942 35930 10966 35932
rect 11022 35930 11046 35932
rect 11102 35930 11126 35932
rect 11182 35930 11188 35932
rect 10942 35878 10944 35930
rect 11124 35878 11126 35930
rect 10880 35876 10886 35878
rect 10942 35876 10966 35878
rect 11022 35876 11046 35878
rect 11102 35876 11126 35878
rect 11182 35876 11188 35878
rect 10880 35856 11188 35876
rect 10784 35080 10836 35086
rect 10784 35022 10836 35028
rect 11612 35080 11664 35086
rect 11612 35022 11664 35028
rect 10416 34536 10468 34542
rect 10416 34478 10468 34484
rect 10416 33924 10468 33930
rect 10416 33866 10468 33872
rect 10324 33856 10376 33862
rect 10324 33798 10376 33804
rect 10336 32910 10364 33798
rect 10428 33522 10456 33866
rect 10796 33862 10824 35022
rect 10880 34844 11188 34864
rect 10880 34842 10886 34844
rect 10942 34842 10966 34844
rect 11022 34842 11046 34844
rect 11102 34842 11126 34844
rect 11182 34842 11188 34844
rect 10942 34790 10944 34842
rect 11124 34790 11126 34842
rect 10880 34788 10886 34790
rect 10942 34788 10966 34790
rect 11022 34788 11046 34790
rect 11102 34788 11126 34790
rect 11182 34788 11188 34790
rect 10880 34768 11188 34788
rect 11624 34542 11652 35022
rect 11704 34604 11756 34610
rect 11704 34546 11756 34552
rect 11612 34536 11664 34542
rect 11612 34478 11664 34484
rect 11520 33992 11572 33998
rect 11520 33934 11572 33940
rect 11244 33924 11296 33930
rect 11244 33866 11296 33872
rect 11428 33924 11480 33930
rect 11428 33866 11480 33872
rect 10784 33856 10836 33862
rect 10784 33798 10836 33804
rect 10880 33756 11188 33776
rect 10880 33754 10886 33756
rect 10942 33754 10966 33756
rect 11022 33754 11046 33756
rect 11102 33754 11126 33756
rect 11182 33754 11188 33756
rect 10942 33702 10944 33754
rect 11124 33702 11126 33754
rect 10880 33700 10886 33702
rect 10942 33700 10966 33702
rect 11022 33700 11046 33702
rect 11102 33700 11126 33702
rect 11182 33700 11188 33702
rect 10880 33680 11188 33700
rect 10416 33516 10468 33522
rect 10416 33458 10468 33464
rect 10692 33312 10744 33318
rect 10692 33254 10744 33260
rect 10324 32904 10376 32910
rect 10324 32846 10376 32852
rect 10232 31884 10284 31890
rect 10232 31826 10284 31832
rect 10048 31816 10100 31822
rect 10048 31758 10100 31764
rect 10048 31204 10100 31210
rect 10048 31146 10100 31152
rect 9956 30728 10008 30734
rect 9956 30670 10008 30676
rect 9864 30252 9916 30258
rect 9864 30194 9916 30200
rect 9772 29640 9824 29646
rect 9772 29582 9824 29588
rect 9680 28620 9732 28626
rect 9680 28562 9732 28568
rect 9496 28552 9548 28558
rect 9496 28494 9548 28500
rect 9220 28212 9272 28218
rect 9220 28154 9272 28160
rect 9324 28206 9444 28234
rect 9324 28098 9352 28206
rect 9036 28076 9088 28082
rect 9036 28018 9088 28024
rect 9128 28076 9180 28082
rect 9128 28018 9180 28024
rect 9232 28070 9352 28098
rect 9140 27962 9168 28018
rect 9048 27934 9168 27962
rect 9048 27470 9076 27934
rect 9128 27872 9180 27878
rect 9128 27814 9180 27820
rect 9036 27464 9088 27470
rect 9036 27406 9088 27412
rect 8944 26988 8996 26994
rect 8944 26930 8996 26936
rect 8942 26480 8998 26489
rect 9048 26450 9076 27406
rect 8942 26415 8998 26424
rect 9036 26444 9088 26450
rect 8956 26382 8984 26415
rect 9036 26386 9088 26392
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 8956 23526 8984 26318
rect 9140 25294 9168 27814
rect 9232 26042 9260 28070
rect 9312 28008 9364 28014
rect 9312 27950 9364 27956
rect 9324 27470 9352 27950
rect 9508 27946 9536 28494
rect 9496 27940 9548 27946
rect 9496 27882 9548 27888
rect 9494 27704 9550 27713
rect 9494 27639 9550 27648
rect 9508 27606 9536 27639
rect 9876 27606 9904 30194
rect 9956 29640 10008 29646
rect 9956 29582 10008 29588
rect 9496 27600 9548 27606
rect 9496 27542 9548 27548
rect 9864 27600 9916 27606
rect 9864 27542 9916 27548
rect 9312 27464 9364 27470
rect 9680 27464 9732 27470
rect 9312 27406 9364 27412
rect 9508 27424 9680 27452
rect 9324 26382 9352 27406
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 8944 23520 8996 23526
rect 8944 23462 8996 23468
rect 9140 22778 9168 24142
rect 9220 23724 9272 23730
rect 9220 23666 9272 23672
rect 9232 23118 9260 23666
rect 9324 23644 9352 26318
rect 9404 25832 9456 25838
rect 9404 25774 9456 25780
rect 9416 25498 9444 25774
rect 9404 25492 9456 25498
rect 9404 25434 9456 25440
rect 9508 23730 9536 27424
rect 9680 27406 9732 27412
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9588 26512 9640 26518
rect 9588 26454 9640 26460
rect 9600 26314 9628 26454
rect 9588 26308 9640 26314
rect 9588 26250 9640 26256
rect 9588 26036 9640 26042
rect 9588 25978 9640 25984
rect 9600 24954 9628 25978
rect 9692 25294 9720 26726
rect 9784 26586 9812 26930
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 9968 26058 9996 29582
rect 10060 29170 10088 31146
rect 10140 30728 10192 30734
rect 10140 30670 10192 30676
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 10048 28076 10100 28082
rect 10048 28018 10100 28024
rect 10060 26518 10088 28018
rect 10048 26512 10100 26518
rect 10048 26454 10100 26460
rect 9968 26030 10088 26058
rect 9956 25900 10008 25906
rect 9956 25842 10008 25848
rect 9968 25702 9996 25842
rect 9956 25696 10008 25702
rect 9956 25638 10008 25644
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9588 24948 9640 24954
rect 9588 24890 9640 24896
rect 9864 24132 9916 24138
rect 9864 24074 9916 24080
rect 9876 23866 9904 24074
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9692 23746 9720 23802
rect 9496 23724 9548 23730
rect 9692 23718 9812 23746
rect 9496 23666 9548 23672
rect 9404 23656 9456 23662
rect 9324 23616 9404 23644
rect 9404 23598 9456 23604
rect 9508 23254 9536 23666
rect 9784 23662 9812 23718
rect 9588 23656 9640 23662
rect 9588 23598 9640 23604
rect 9772 23656 9824 23662
rect 9772 23598 9824 23604
rect 9496 23248 9548 23254
rect 9496 23190 9548 23196
rect 9220 23112 9272 23118
rect 9220 23054 9272 23060
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 9232 22710 9260 23054
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9220 22704 9272 22710
rect 9416 22681 9444 22714
rect 9220 22646 9272 22652
rect 9402 22672 9458 22681
rect 9128 22636 9180 22642
rect 9508 22642 9536 23190
rect 9600 23050 9628 23598
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9588 23044 9640 23050
rect 9588 22986 9640 22992
rect 9402 22607 9458 22616
rect 9496 22636 9548 22642
rect 9128 22578 9180 22584
rect 9496 22578 9548 22584
rect 8944 22500 8996 22506
rect 8944 22442 8996 22448
rect 8956 20466 8984 22442
rect 9034 22128 9090 22137
rect 9034 22063 9090 22072
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8956 20262 8984 20402
rect 8944 20256 8996 20262
rect 8944 20198 8996 20204
rect 8944 19780 8996 19786
rect 8944 19722 8996 19728
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 8864 17954 8892 18634
rect 8680 17926 8892 17954
rect 8680 12434 8708 17926
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8772 17270 8800 17478
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8772 16658 8800 17070
rect 8864 16726 8892 17138
rect 8852 16720 8904 16726
rect 8852 16662 8904 16668
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8864 16046 8892 16662
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8760 15564 8812 15570
rect 8812 15524 8892 15552
rect 8760 15506 8812 15512
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8772 15094 8800 15302
rect 8760 15088 8812 15094
rect 8760 15030 8812 15036
rect 8864 14396 8892 15524
rect 8956 15484 8984 19722
rect 9048 18952 9076 22063
rect 9140 20058 9168 22578
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9416 21865 9444 21966
rect 9402 21856 9458 21865
rect 9402 21791 9458 21800
rect 9416 21706 9444 21791
rect 9600 21729 9628 22986
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9324 21678 9444 21706
rect 9586 21720 9642 21729
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 9232 21146 9260 21490
rect 9324 21468 9352 21678
rect 9586 21655 9642 21664
rect 9494 21584 9550 21593
rect 9494 21519 9496 21528
rect 9548 21519 9550 21528
rect 9496 21490 9548 21496
rect 9404 21480 9456 21486
rect 9324 21440 9404 21468
rect 9404 21422 9456 21428
rect 9586 21448 9642 21457
rect 9586 21383 9642 21392
rect 9402 21176 9458 21185
rect 9220 21140 9272 21146
rect 9402 21111 9458 21120
rect 9220 21082 9272 21088
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9324 20602 9352 20878
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9324 19446 9352 19790
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9048 18924 9260 18952
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 9048 17134 9076 18770
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 9140 17338 9168 17546
rect 9232 17542 9260 18924
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 9128 15496 9180 15502
rect 8956 15464 9128 15484
rect 9180 15464 9182 15473
rect 8956 15456 9126 15464
rect 9126 15399 9182 15408
rect 8944 14408 8996 14414
rect 8864 14368 8944 14396
rect 8944 14350 8996 14356
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8772 12782 8800 13874
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8680 12406 8800 12434
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8128 8838 8156 9522
rect 8208 9512 8260 9518
rect 8484 9512 8536 9518
rect 8260 9460 8340 9466
rect 8208 9454 8340 9460
rect 8484 9454 8536 9460
rect 8220 9438 8340 9454
rect 8312 8974 8340 9438
rect 8496 9178 8524 9454
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8312 8634 8340 8910
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 7852 7546 7880 7754
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7472 7346 7524 7352
rect 7576 7364 7696 7392
rect 6972 6752 7052 6780
rect 6920 6734 6972 6740
rect 6932 6361 6960 6734
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6918 6352 6974 6361
rect 6918 6287 6974 6296
rect 6748 5902 6868 5930
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5408 4100 5488 4128
rect 5356 4082 5408 4088
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 3148 3120 3200 3126
rect 3148 3062 3200 3068
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2792 2502 2912 2530
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2792 1737 2820 2314
rect 2778 1728 2834 1737
rect 2778 1663 2834 1672
rect 2884 1057 2912 2502
rect 2870 1048 2926 1057
rect 2870 983 2926 992
rect 386 0 442 800
rect 1122 0 1178 800
rect 1858 0 1914 800
rect 2594 0 2650 800
rect 2976 377 3004 3062
rect 4172 3058 4200 3538
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 3436 800 3464 2994
rect 4264 2774 4292 3402
rect 5000 3126 5028 3878
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 5184 3058 5212 4082
rect 5552 3534 5580 4422
rect 5644 3738 5672 4558
rect 5920 4282 5948 4558
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 6380 4146 6408 4558
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6552 4140 6604 4146
rect 6656 4128 6684 4626
rect 6748 4554 6776 5902
rect 6932 5778 6960 6287
rect 6920 5772 6972 5778
rect 6840 5732 6920 5760
rect 6840 5302 6868 5732
rect 6920 5714 6972 5720
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6932 4826 6960 5578
rect 7024 5370 7052 6394
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 6748 4282 6776 4490
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6932 4146 6960 4762
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7116 4282 7144 4490
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7208 4162 7236 7346
rect 7484 7002 7512 7346
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 6736 4140 6788 4146
rect 6656 4100 6736 4128
rect 6552 4082 6604 4088
rect 6736 4082 6788 4088
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 7116 4134 7236 4162
rect 5816 4072 5868 4078
rect 5814 4040 5816 4049
rect 5868 4040 5870 4049
rect 5814 3975 5870 3984
rect 5915 3836 6223 3856
rect 5915 3834 5921 3836
rect 5977 3834 6001 3836
rect 6057 3834 6081 3836
rect 6137 3834 6161 3836
rect 6217 3834 6223 3836
rect 5977 3782 5979 3834
rect 6159 3782 6161 3834
rect 5915 3780 5921 3782
rect 5977 3780 6001 3782
rect 6057 3780 6081 3782
rect 6137 3780 6161 3782
rect 6217 3780 6223 3782
rect 5915 3760 6223 3780
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 6564 3670 6592 4082
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 4172 2746 4292 2774
rect 5915 2748 6223 2768
rect 5915 2746 5921 2748
rect 5977 2746 6001 2748
rect 6057 2746 6081 2748
rect 6137 2746 6161 2748
rect 6217 2746 6223 2748
rect 4172 800 4200 2746
rect 5977 2694 5979 2746
rect 6159 2694 6161 2746
rect 5915 2692 5921 2694
rect 5977 2692 6001 2694
rect 6057 2692 6081 2694
rect 6137 2692 6161 2694
rect 6217 2692 6223 2694
rect 5915 2672 6223 2692
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 4908 800 4936 2382
rect 5736 800 5764 2382
rect 6472 800 6500 2994
rect 6748 2922 6776 3878
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6840 2650 6868 3606
rect 7116 2854 7144 4134
rect 7576 4078 7604 7364
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7668 7002 7696 7210
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7760 6798 7788 7142
rect 8312 6798 8340 8570
rect 8404 8430 8432 8910
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8404 7410 8432 8366
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8312 6390 8340 6734
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8312 4690 8340 6326
rect 8404 5234 8432 7346
rect 8496 7274 8524 7754
rect 8680 7410 8708 11698
rect 8772 10198 8800 12406
rect 8864 11898 8892 13806
rect 8956 12696 8984 14350
rect 9232 12889 9260 17478
rect 9324 16658 9352 18702
rect 9416 17338 9444 21111
rect 9600 21010 9628 21383
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 9692 20874 9720 22034
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9784 20754 9812 23462
rect 9968 21962 9996 25638
rect 10060 23662 10088 26030
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 10060 22030 10088 22918
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9600 20726 9812 20754
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9508 18426 9536 18702
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9600 17490 9628 20726
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9680 19984 9732 19990
rect 9680 19926 9732 19932
rect 9692 19854 9720 19926
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9784 19378 9812 19994
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9692 17678 9720 18294
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9508 17462 9628 17490
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9416 15570 9444 16458
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9324 15026 9352 15302
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9416 14414 9444 15506
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9508 14346 9536 17462
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9600 16454 9628 17274
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9600 15502 9628 16186
rect 9692 16114 9720 17614
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9692 15502 9720 16050
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9692 15366 9720 15438
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9600 14618 9628 15030
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9586 14512 9642 14521
rect 9586 14447 9588 14456
rect 9640 14447 9642 14456
rect 9588 14418 9640 14424
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 13938 9720 14214
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9600 13530 9628 13806
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9218 12880 9274 12889
rect 9218 12815 9274 12824
rect 8956 12668 9168 12696
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8864 11150 8892 11698
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 8496 5846 8524 7210
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8312 4146 8340 4626
rect 8404 4622 8432 5170
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 8312 3602 8340 4082
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 7208 800 7236 2994
rect 8128 2854 8156 3334
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8588 2582 8616 5170
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 8680 2446 8708 7346
rect 8956 3670 8984 12242
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9048 11558 9076 12038
rect 9140 11801 9168 12668
rect 9126 11792 9182 11801
rect 9324 11762 9352 13466
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9126 11727 9182 11736
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9218 11656 9274 11665
rect 9218 11591 9274 11600
rect 9037 11552 9089 11558
rect 9037 11494 9089 11500
rect 9126 11384 9182 11393
rect 9126 11319 9182 11328
rect 9034 11248 9090 11257
rect 9034 11183 9090 11192
rect 9048 7750 9076 11183
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9048 6458 9076 7346
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9140 5574 9168 11319
rect 9232 8022 9260 11591
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9324 11150 9352 11494
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9324 8430 9352 8910
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 9324 7342 9352 8366
rect 9416 8294 9444 12718
rect 9508 9994 9536 13194
rect 9600 12850 9628 13194
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9586 12744 9642 12753
rect 9586 12679 9642 12688
rect 9600 12457 9628 12679
rect 9586 12448 9642 12457
rect 9586 12383 9642 12392
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9600 11218 9628 12106
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9508 7750 9536 9930
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 8974 9628 9318
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9692 8362 9720 13874
rect 9784 13172 9812 19314
rect 9876 18170 9904 19722
rect 9968 19258 9996 20198
rect 10048 19780 10100 19786
rect 10048 19722 10100 19728
rect 10060 19446 10088 19722
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 9968 19230 10088 19258
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9968 18290 9996 18566
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9876 18142 9996 18170
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9876 15706 9904 16050
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9876 13394 9904 15302
rect 9968 13870 9996 18142
rect 10060 17184 10088 19230
rect 10152 17377 10180 30670
rect 10244 28642 10272 31826
rect 10336 31346 10364 32846
rect 10704 32502 10732 33254
rect 11256 33114 11284 33866
rect 11440 33590 11468 33866
rect 11532 33658 11560 33934
rect 11520 33652 11572 33658
rect 11520 33594 11572 33600
rect 11428 33584 11480 33590
rect 11428 33526 11480 33532
rect 11336 33312 11388 33318
rect 11336 33254 11388 33260
rect 11244 33108 11296 33114
rect 11244 33050 11296 33056
rect 10784 32768 10836 32774
rect 10784 32710 10836 32716
rect 10796 32570 10824 32710
rect 10880 32668 11188 32688
rect 10880 32666 10886 32668
rect 10942 32666 10966 32668
rect 11022 32666 11046 32668
rect 11102 32666 11126 32668
rect 11182 32666 11188 32668
rect 10942 32614 10944 32666
rect 11124 32614 11126 32666
rect 10880 32612 10886 32614
rect 10942 32612 10966 32614
rect 11022 32612 11046 32614
rect 11102 32612 11126 32614
rect 11182 32612 11188 32614
rect 10880 32592 11188 32612
rect 10784 32564 10836 32570
rect 10784 32506 10836 32512
rect 10692 32496 10744 32502
rect 10692 32438 10744 32444
rect 11244 31884 11296 31890
rect 11244 31826 11296 31832
rect 10508 31816 10560 31822
rect 10508 31758 10560 31764
rect 10324 31340 10376 31346
rect 10324 31282 10376 31288
rect 10520 28744 10548 31758
rect 10880 31580 11188 31600
rect 10880 31578 10886 31580
rect 10942 31578 10966 31580
rect 11022 31578 11046 31580
rect 11102 31578 11126 31580
rect 11182 31578 11188 31580
rect 10942 31526 10944 31578
rect 11124 31526 11126 31578
rect 10880 31524 10886 31526
rect 10942 31524 10966 31526
rect 11022 31524 11046 31526
rect 11102 31524 11126 31526
rect 11182 31524 11188 31526
rect 10880 31504 11188 31524
rect 10876 31340 10928 31346
rect 10876 31282 10928 31288
rect 10692 31136 10744 31142
rect 10692 31078 10744 31084
rect 10704 30734 10732 31078
rect 10888 30938 10916 31282
rect 10876 30932 10928 30938
rect 10876 30874 10928 30880
rect 11256 30870 11284 31826
rect 11244 30864 11296 30870
rect 11244 30806 11296 30812
rect 10692 30728 10744 30734
rect 10692 30670 10744 30676
rect 10880 30492 11188 30512
rect 10880 30490 10886 30492
rect 10942 30490 10966 30492
rect 11022 30490 11046 30492
rect 11102 30490 11126 30492
rect 11182 30490 11188 30492
rect 10942 30438 10944 30490
rect 11124 30438 11126 30490
rect 10880 30436 10886 30438
rect 10942 30436 10966 30438
rect 11022 30436 11046 30438
rect 11102 30436 11126 30438
rect 11182 30436 11188 30438
rect 10880 30416 11188 30436
rect 10784 30388 10836 30394
rect 10784 30330 10836 30336
rect 10692 30116 10744 30122
rect 10692 30058 10744 30064
rect 10520 28716 10640 28744
rect 10244 28614 10548 28642
rect 10324 28484 10376 28490
rect 10324 28426 10376 28432
rect 10416 28484 10468 28490
rect 10416 28426 10468 28432
rect 10336 28218 10364 28426
rect 10324 28212 10376 28218
rect 10324 28154 10376 28160
rect 10232 28076 10284 28082
rect 10232 28018 10284 28024
rect 10244 27470 10272 28018
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 10324 27464 10376 27470
rect 10324 27406 10376 27412
rect 10244 26382 10272 27406
rect 10336 27130 10364 27406
rect 10324 27124 10376 27130
rect 10324 27066 10376 27072
rect 10428 27062 10456 28426
rect 10416 27056 10468 27062
rect 10416 26998 10468 27004
rect 10324 26988 10376 26994
rect 10324 26930 10376 26936
rect 10232 26376 10284 26382
rect 10232 26318 10284 26324
rect 10336 25430 10364 26930
rect 10428 26586 10456 26998
rect 10416 26580 10468 26586
rect 10416 26522 10468 26528
rect 10520 26466 10548 28614
rect 10428 26438 10548 26466
rect 10324 25424 10376 25430
rect 10324 25366 10376 25372
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 10244 23866 10272 24754
rect 10336 24750 10364 25366
rect 10324 24744 10376 24750
rect 10324 24686 10376 24692
rect 10232 23860 10284 23866
rect 10232 23802 10284 23808
rect 10428 23118 10456 26438
rect 10508 25356 10560 25362
rect 10508 25298 10560 25304
rect 10520 23730 10548 25298
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10416 23112 10468 23118
rect 10416 23054 10468 23060
rect 10324 22568 10376 22574
rect 10324 22510 10376 22516
rect 10336 21146 10364 22510
rect 10520 21554 10548 23666
rect 10612 22094 10640 28716
rect 10704 27577 10732 30058
rect 10796 29850 10824 30330
rect 11348 29850 11376 33254
rect 11624 32910 11652 34478
rect 11716 33522 11744 34546
rect 11900 33522 11928 36654
rect 12900 36236 12952 36242
rect 12900 36178 12952 36184
rect 12624 36032 12676 36038
rect 12624 35974 12676 35980
rect 11980 35692 12032 35698
rect 11980 35634 12032 35640
rect 11992 33998 12020 35634
rect 12072 35012 12124 35018
rect 12072 34954 12124 34960
rect 11980 33992 12032 33998
rect 11980 33934 12032 33940
rect 11992 33538 12020 33934
rect 12084 33658 12112 34954
rect 12636 34678 12664 35974
rect 12808 35692 12860 35698
rect 12912 35680 12940 36178
rect 12860 35652 12940 35680
rect 12808 35634 12860 35640
rect 12716 35488 12768 35494
rect 12716 35430 12768 35436
rect 12624 34672 12676 34678
rect 12624 34614 12676 34620
rect 12728 33674 12756 35430
rect 12072 33652 12124 33658
rect 12072 33594 12124 33600
rect 12636 33646 12756 33674
rect 11992 33522 12112 33538
rect 11704 33516 11756 33522
rect 11704 33458 11756 33464
rect 11888 33516 11940 33522
rect 11992 33516 12124 33522
rect 11992 33510 12072 33516
rect 11888 33458 11940 33464
rect 12072 33458 12124 33464
rect 11612 32904 11664 32910
rect 11612 32846 11664 32852
rect 11624 32366 11652 32846
rect 11612 32360 11664 32366
rect 11612 32302 11664 32308
rect 11520 31816 11572 31822
rect 11518 31784 11520 31793
rect 11572 31784 11574 31793
rect 11518 31719 11574 31728
rect 11624 31482 11652 32302
rect 11612 31476 11664 31482
rect 11612 31418 11664 31424
rect 11716 31362 11744 33458
rect 11980 32836 12032 32842
rect 11980 32778 12032 32784
rect 11520 31340 11572 31346
rect 11520 31282 11572 31288
rect 11624 31334 11744 31362
rect 11428 30728 11480 30734
rect 11428 30670 11480 30676
rect 10784 29844 10836 29850
rect 10784 29786 10836 29792
rect 11336 29844 11388 29850
rect 11336 29786 11388 29792
rect 10690 27568 10746 27577
rect 10690 27503 10746 27512
rect 10796 27130 10824 29786
rect 11440 29714 11468 30670
rect 11532 30666 11560 31282
rect 11520 30660 11572 30666
rect 11520 30602 11572 30608
rect 11624 30054 11652 31334
rect 11796 31272 11848 31278
rect 11796 31214 11848 31220
rect 11704 31204 11756 31210
rect 11704 31146 11756 31152
rect 11716 30734 11744 31146
rect 11704 30728 11756 30734
rect 11704 30670 11756 30676
rect 11612 30048 11664 30054
rect 11612 29990 11664 29996
rect 11428 29708 11480 29714
rect 11428 29650 11480 29656
rect 11612 29708 11664 29714
rect 11612 29650 11664 29656
rect 10880 29404 11188 29424
rect 10880 29402 10886 29404
rect 10942 29402 10966 29404
rect 11022 29402 11046 29404
rect 11102 29402 11126 29404
rect 11182 29402 11188 29404
rect 10942 29350 10944 29402
rect 11124 29350 11126 29402
rect 10880 29348 10886 29350
rect 10942 29348 10966 29350
rect 11022 29348 11046 29350
rect 11102 29348 11126 29350
rect 11182 29348 11188 29350
rect 10880 29328 11188 29348
rect 11336 28756 11388 28762
rect 11336 28698 11388 28704
rect 11244 28416 11296 28422
rect 11244 28358 11296 28364
rect 10880 28316 11188 28336
rect 10880 28314 10886 28316
rect 10942 28314 10966 28316
rect 11022 28314 11046 28316
rect 11102 28314 11126 28316
rect 11182 28314 11188 28316
rect 10942 28262 10944 28314
rect 11124 28262 11126 28314
rect 10880 28260 10886 28262
rect 10942 28260 10966 28262
rect 11022 28260 11046 28262
rect 11102 28260 11126 28262
rect 11182 28260 11188 28262
rect 10880 28240 11188 28260
rect 10968 27940 11020 27946
rect 10968 27882 11020 27888
rect 10980 27470 11008 27882
rect 11256 27606 11284 28358
rect 11348 28082 11376 28698
rect 11624 28082 11652 29650
rect 11716 29510 11744 30670
rect 11704 29504 11756 29510
rect 11704 29446 11756 29452
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11612 28076 11664 28082
rect 11612 28018 11664 28024
rect 11244 27600 11296 27606
rect 11244 27542 11296 27548
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 10880 27228 11188 27248
rect 10880 27226 10886 27228
rect 10942 27226 10966 27228
rect 11022 27226 11046 27228
rect 11102 27226 11126 27228
rect 11182 27226 11188 27228
rect 10942 27174 10944 27226
rect 11124 27174 11126 27226
rect 10880 27172 10886 27174
rect 10942 27172 10966 27174
rect 11022 27172 11046 27174
rect 11102 27172 11126 27174
rect 11182 27172 11188 27174
rect 10880 27152 11188 27172
rect 10692 27124 10744 27130
rect 10692 27066 10744 27072
rect 10784 27124 10836 27130
rect 10784 27066 10836 27072
rect 10704 25276 10732 27066
rect 10796 26450 10824 27066
rect 11440 26926 11468 27406
rect 11520 27396 11572 27402
rect 11520 27338 11572 27344
rect 11428 26920 11480 26926
rect 11428 26862 11480 26868
rect 11244 26512 11296 26518
rect 11244 26454 11296 26460
rect 10784 26444 10836 26450
rect 10784 26386 10836 26392
rect 10796 25906 10824 26386
rect 10880 26140 11188 26160
rect 10880 26138 10886 26140
rect 10942 26138 10966 26140
rect 11022 26138 11046 26140
rect 11102 26138 11126 26140
rect 11182 26138 11188 26140
rect 10942 26086 10944 26138
rect 11124 26086 11126 26138
rect 10880 26084 10886 26086
rect 10942 26084 10966 26086
rect 11022 26084 11046 26086
rect 11102 26084 11126 26086
rect 11182 26084 11188 26086
rect 10880 26064 11188 26084
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 10796 25430 10824 25842
rect 10784 25424 10836 25430
rect 10784 25366 10836 25372
rect 10704 25248 10824 25276
rect 10692 24948 10744 24954
rect 10692 24890 10744 24896
rect 10704 24818 10732 24890
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10704 24410 10732 24618
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 10796 24274 10824 25248
rect 10880 25052 11188 25072
rect 10880 25050 10886 25052
rect 10942 25050 10966 25052
rect 11022 25050 11046 25052
rect 11102 25050 11126 25052
rect 11182 25050 11188 25052
rect 10942 24998 10944 25050
rect 11124 24998 11126 25050
rect 10880 24996 10886 24998
rect 10942 24996 10966 24998
rect 11022 24996 11046 24998
rect 11102 24996 11126 24998
rect 11182 24996 11188 24998
rect 10880 24976 11188 24996
rect 11256 24818 11284 26454
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11348 25226 11376 26318
rect 11336 25220 11388 25226
rect 11336 25162 11388 25168
rect 11244 24812 11296 24818
rect 11244 24754 11296 24760
rect 11348 24698 11376 25162
rect 11440 24818 11468 26862
rect 11532 26042 11560 27338
rect 11520 26036 11572 26042
rect 11520 25978 11572 25984
rect 11624 25294 11652 28018
rect 11808 25498 11836 31214
rect 11992 30870 12020 32778
rect 12084 31822 12112 33458
rect 12256 32428 12308 32434
rect 12256 32370 12308 32376
rect 12072 31816 12124 31822
rect 12072 31758 12124 31764
rect 12268 31482 12296 32370
rect 12256 31476 12308 31482
rect 12256 31418 12308 31424
rect 11980 30864 12032 30870
rect 11980 30806 12032 30812
rect 12440 30864 12492 30870
rect 12440 30806 12492 30812
rect 11888 30796 11940 30802
rect 11888 30738 11940 30744
rect 12072 30796 12124 30802
rect 12072 30738 12124 30744
rect 11796 25492 11848 25498
rect 11796 25434 11848 25440
rect 11900 25362 11928 30738
rect 12084 30394 12112 30738
rect 12256 30660 12308 30666
rect 12256 30602 12308 30608
rect 12072 30388 12124 30394
rect 12072 30330 12124 30336
rect 12072 30252 12124 30258
rect 12072 30194 12124 30200
rect 12084 29578 12112 30194
rect 12072 29572 12124 29578
rect 12072 29514 12124 29520
rect 11980 29504 12032 29510
rect 11980 29446 12032 29452
rect 11888 25356 11940 25362
rect 11888 25298 11940 25304
rect 11612 25288 11664 25294
rect 11612 25230 11664 25236
rect 11520 25152 11572 25158
rect 11520 25094 11572 25100
rect 11428 24812 11480 24818
rect 11428 24754 11480 24760
rect 11256 24670 11376 24698
rect 10784 24268 10836 24274
rect 10784 24210 10836 24216
rect 10880 23964 11188 23984
rect 10880 23962 10886 23964
rect 10942 23962 10966 23964
rect 11022 23962 11046 23964
rect 11102 23962 11126 23964
rect 11182 23962 11188 23964
rect 10942 23910 10944 23962
rect 11124 23910 11126 23962
rect 10880 23908 10886 23910
rect 10942 23908 10966 23910
rect 11022 23908 11046 23910
rect 11102 23908 11126 23910
rect 11182 23908 11188 23910
rect 10880 23888 11188 23908
rect 10880 22876 11188 22896
rect 10880 22874 10886 22876
rect 10942 22874 10966 22876
rect 11022 22874 11046 22876
rect 11102 22874 11126 22876
rect 11182 22874 11188 22876
rect 10942 22822 10944 22874
rect 11124 22822 11126 22874
rect 10880 22820 10886 22822
rect 10942 22820 10966 22822
rect 11022 22820 11046 22822
rect 11102 22820 11126 22822
rect 11182 22820 11188 22822
rect 10880 22800 11188 22820
rect 10612 22066 10732 22094
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10324 21140 10376 21146
rect 10324 21082 10376 21088
rect 10232 20528 10284 20534
rect 10232 20470 10284 20476
rect 10244 19446 10272 20470
rect 10336 20398 10364 21082
rect 10416 20868 10468 20874
rect 10416 20810 10468 20816
rect 10600 20868 10652 20874
rect 10600 20810 10652 20816
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10232 19440 10284 19446
rect 10232 19382 10284 19388
rect 10138 17368 10194 17377
rect 10138 17303 10194 17312
rect 10060 17156 10272 17184
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 15638 10180 16526
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10060 15094 10088 15438
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 10060 13938 10088 14350
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 10060 13530 10088 13874
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9864 13184 9916 13190
rect 9784 13144 9864 13172
rect 9864 13126 9916 13132
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9784 11150 9812 12582
rect 9876 11626 9904 12786
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9862 11520 9918 11529
rect 9862 11455 9918 11464
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9876 10996 9904 11455
rect 9784 10968 9904 10996
rect 9784 9194 9812 10968
rect 9968 10674 9996 11766
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9876 9654 9904 10610
rect 9968 10198 9996 10610
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9968 9382 9996 9862
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9784 9166 9904 9194
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9232 6322 9260 7142
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9324 5914 9352 7278
rect 9692 6866 9720 7414
rect 9784 7274 9812 8978
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 9048 2922 9076 4558
rect 9140 4214 9168 4966
rect 9692 4690 9720 5238
rect 9876 4826 9904 9166
rect 9968 8498 9996 9318
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9968 7478 9996 8434
rect 10060 8090 10088 13126
rect 10152 12986 10180 14282
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10244 12322 10272 17156
rect 10336 15434 10364 19858
rect 10428 16590 10456 20810
rect 10612 20534 10640 20810
rect 10704 20534 10732 22066
rect 10880 21788 11188 21808
rect 10880 21786 10886 21788
rect 10942 21786 10966 21788
rect 11022 21786 11046 21788
rect 11102 21786 11126 21788
rect 11182 21786 11188 21788
rect 10942 21734 10944 21786
rect 11124 21734 11126 21786
rect 10880 21732 10886 21734
rect 10942 21732 10966 21734
rect 11022 21732 11046 21734
rect 11102 21732 11126 21734
rect 11182 21732 11188 21734
rect 10880 21712 11188 21732
rect 10880 20700 11188 20720
rect 10880 20698 10886 20700
rect 10942 20698 10966 20700
rect 11022 20698 11046 20700
rect 11102 20698 11126 20700
rect 11182 20698 11188 20700
rect 10942 20646 10944 20698
rect 11124 20646 11126 20698
rect 10880 20644 10886 20646
rect 10942 20644 10966 20646
rect 11022 20644 11046 20646
rect 11102 20644 11126 20646
rect 11182 20644 11188 20646
rect 10880 20624 11188 20644
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10692 20528 10744 20534
rect 10692 20470 10744 20476
rect 10600 19780 10652 19786
rect 10600 19722 10652 19728
rect 10612 19258 10640 19722
rect 10704 19378 10732 20470
rect 10880 19612 11188 19632
rect 10880 19610 10886 19612
rect 10942 19610 10966 19612
rect 11022 19610 11046 19612
rect 11102 19610 11126 19612
rect 11182 19610 11188 19612
rect 10942 19558 10944 19610
rect 11124 19558 11126 19610
rect 10880 19556 10886 19558
rect 10942 19556 10966 19558
rect 11022 19556 11046 19558
rect 11102 19556 11126 19558
rect 11182 19556 11188 19558
rect 10880 19536 11188 19556
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10612 19230 10732 19258
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10324 15428 10376 15434
rect 10324 15370 10376 15376
rect 10324 15088 10376 15094
rect 10324 15030 10376 15036
rect 10336 14346 10364 15030
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10336 13326 10364 14282
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10152 12294 10272 12322
rect 10152 10792 10180 12294
rect 10232 12232 10284 12238
rect 10336 12220 10364 13262
rect 10428 12764 10456 16526
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 13938 10548 15846
rect 10612 15366 10640 18090
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 14482 10640 14758
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10520 12918 10548 13874
rect 10612 13326 10640 14214
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10428 12736 10640 12764
rect 10506 12336 10562 12345
rect 10506 12271 10562 12280
rect 10284 12192 10364 12220
rect 10232 12174 10284 12180
rect 10244 11150 10272 12174
rect 10322 12064 10378 12073
rect 10322 11999 10378 12008
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10152 10764 10272 10792
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10152 9178 10180 10610
rect 10244 10266 10272 10764
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10244 9586 10272 9930
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10244 8838 10272 9522
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10152 8022 10180 8230
rect 10140 8016 10192 8022
rect 10046 7984 10102 7993
rect 10140 7958 10192 7964
rect 10046 7919 10102 7928
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9968 6798 9996 7210
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9968 5166 9996 6734
rect 10060 6474 10088 7919
rect 10152 7546 10180 7958
rect 10244 7886 10272 8774
rect 10336 7993 10364 11999
rect 10520 11762 10548 12271
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10322 7984 10378 7993
rect 10322 7919 10378 7928
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10060 6446 10180 6474
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 5234 10088 6258
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9312 4548 9364 4554
rect 9312 4490 9364 4496
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 9324 4078 9352 4490
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9232 3058 9260 3538
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9600 3194 9628 3402
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9692 3126 9720 4422
rect 9784 3194 9812 4558
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9876 4146 9904 4490
rect 9968 4486 9996 5102
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 10060 4282 10088 5170
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10152 3738 10180 6446
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8772 2650 8800 2790
rect 10244 2774 10272 7822
rect 10336 7546 10364 7822
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10428 5914 10456 11698
rect 10520 10538 10548 11698
rect 10612 11529 10640 12736
rect 10598 11520 10654 11529
rect 10598 11455 10654 11464
rect 10704 11234 10732 19230
rect 10796 18698 10824 19314
rect 11058 19136 11114 19145
rect 11058 19071 11114 19080
rect 11072 18902 11100 19071
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10796 18358 10824 18634
rect 10880 18524 11188 18544
rect 10880 18522 10886 18524
rect 10942 18522 10966 18524
rect 11022 18522 11046 18524
rect 11102 18522 11126 18524
rect 11182 18522 11188 18524
rect 10942 18470 10944 18522
rect 11124 18470 11126 18522
rect 10880 18468 10886 18470
rect 10942 18468 10966 18470
rect 11022 18468 11046 18470
rect 11102 18468 11126 18470
rect 11182 18468 11188 18470
rect 10880 18448 11188 18468
rect 10784 18352 10836 18358
rect 10784 18294 10836 18300
rect 11256 17882 11284 24670
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11348 23798 11376 24006
rect 11440 23798 11468 24754
rect 11336 23792 11388 23798
rect 11336 23734 11388 23740
rect 11428 23792 11480 23798
rect 11428 23734 11480 23740
rect 11532 23322 11560 25094
rect 11624 24070 11652 25230
rect 11704 24948 11756 24954
rect 11704 24890 11756 24896
rect 11612 24064 11664 24070
rect 11612 24006 11664 24012
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 11532 22234 11560 23258
rect 11520 22228 11572 22234
rect 11520 22170 11572 22176
rect 11532 22094 11560 22170
rect 11440 22066 11560 22094
rect 11440 19990 11468 22066
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 11428 19984 11480 19990
rect 11428 19926 11480 19932
rect 11532 19922 11560 21966
rect 11624 21554 11652 23802
rect 11716 23186 11744 24890
rect 11992 24410 12020 29446
rect 12084 29306 12112 29514
rect 12072 29300 12124 29306
rect 12072 29242 12124 29248
rect 12164 27940 12216 27946
rect 12164 27882 12216 27888
rect 12176 26518 12204 27882
rect 12072 26512 12124 26518
rect 12072 26454 12124 26460
rect 12164 26512 12216 26518
rect 12164 26454 12216 26460
rect 12084 25498 12112 26454
rect 12176 25906 12204 26454
rect 12164 25900 12216 25906
rect 12164 25842 12216 25848
rect 12072 25492 12124 25498
rect 12072 25434 12124 25440
rect 12084 25294 12112 25434
rect 12072 25288 12124 25294
rect 12072 25230 12124 25236
rect 11980 24404 12032 24410
rect 11980 24346 12032 24352
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11612 21548 11664 21554
rect 11716 21536 11744 23122
rect 11796 22976 11848 22982
rect 11796 22918 11848 22924
rect 11808 21978 11836 22918
rect 11808 21962 11928 21978
rect 11808 21956 11940 21962
rect 11808 21950 11888 21956
rect 11888 21898 11940 21904
rect 11992 21842 12020 24346
rect 12084 24206 12112 25230
rect 12176 24954 12204 25842
rect 12164 24948 12216 24954
rect 12164 24890 12216 24896
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 12084 23118 12112 24142
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 12176 23186 12204 24074
rect 12268 23866 12296 30602
rect 12452 28694 12480 30806
rect 12532 29640 12584 29646
rect 12532 29582 12584 29588
rect 12544 29170 12572 29582
rect 12532 29164 12584 29170
rect 12532 29106 12584 29112
rect 12532 29028 12584 29034
rect 12532 28970 12584 28976
rect 12440 28688 12492 28694
rect 12440 28630 12492 28636
rect 12440 26784 12492 26790
rect 12440 26726 12492 26732
rect 12452 26382 12480 26726
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12544 26314 12572 28970
rect 12636 28762 12664 33646
rect 12820 33454 12848 35634
rect 12900 35556 12952 35562
rect 12900 35498 12952 35504
rect 12912 35290 12940 35498
rect 12900 35284 12952 35290
rect 12900 35226 12952 35232
rect 12808 33448 12860 33454
rect 12808 33390 12860 33396
rect 12716 32224 12768 32230
rect 12716 32166 12768 32172
rect 12728 31346 12756 32166
rect 12820 31414 12848 33390
rect 12900 32768 12952 32774
rect 13004 32756 13032 37198
rect 13096 36786 13124 37198
rect 13740 37194 13768 37606
rect 13832 37466 13860 37810
rect 14004 37800 14056 37806
rect 14004 37742 14056 37748
rect 14016 37466 14044 37742
rect 13820 37460 13872 37466
rect 13820 37402 13872 37408
rect 14004 37460 14056 37466
rect 14004 37402 14056 37408
rect 13728 37188 13780 37194
rect 13728 37130 13780 37136
rect 13740 36786 13768 37130
rect 13832 36786 13860 37402
rect 14096 37256 14148 37262
rect 14096 37198 14148 37204
rect 14108 37126 14136 37198
rect 14096 37120 14148 37126
rect 14096 37062 14148 37068
rect 14200 36786 14228 37810
rect 14844 37126 14872 38898
rect 14924 38344 14976 38350
rect 14924 38286 14976 38292
rect 15108 38344 15160 38350
rect 15108 38286 15160 38292
rect 14936 37738 14964 38286
rect 15120 37806 15148 38286
rect 15108 37800 15160 37806
rect 15108 37742 15160 37748
rect 14924 37732 14976 37738
rect 14924 37674 14976 37680
rect 14936 37262 14964 37674
rect 15200 37392 15252 37398
rect 15200 37334 15252 37340
rect 14924 37256 14976 37262
rect 14924 37198 14976 37204
rect 14832 37120 14884 37126
rect 14832 37062 14884 37068
rect 13084 36780 13136 36786
rect 13084 36722 13136 36728
rect 13728 36780 13780 36786
rect 13728 36722 13780 36728
rect 13820 36780 13872 36786
rect 13820 36722 13872 36728
rect 14188 36780 14240 36786
rect 14844 36768 14872 37062
rect 14936 36922 14964 37198
rect 15212 37194 15240 37334
rect 15672 37330 15700 38898
rect 15384 37324 15436 37330
rect 15384 37266 15436 37272
rect 15660 37324 15712 37330
rect 15660 37266 15712 37272
rect 15292 37256 15344 37262
rect 15292 37198 15344 37204
rect 15200 37188 15252 37194
rect 15200 37130 15252 37136
rect 14924 36916 14976 36922
rect 14924 36858 14976 36864
rect 14924 36780 14976 36786
rect 14844 36740 14924 36768
rect 14188 36722 14240 36728
rect 14924 36722 14976 36728
rect 13740 36582 13768 36722
rect 13544 36576 13596 36582
rect 13544 36518 13596 36524
rect 13728 36576 13780 36582
rect 13728 36518 13780 36524
rect 13084 36168 13136 36174
rect 13084 36110 13136 36116
rect 13268 36168 13320 36174
rect 13268 36110 13320 36116
rect 13096 35698 13124 36110
rect 13176 36032 13228 36038
rect 13176 35974 13228 35980
rect 13084 35692 13136 35698
rect 13084 35634 13136 35640
rect 13096 34610 13124 35634
rect 13084 34604 13136 34610
rect 13084 34546 13136 34552
rect 12952 32728 13032 32756
rect 12900 32710 12952 32716
rect 12808 31408 12860 31414
rect 12808 31350 12860 31356
rect 12716 31340 12768 31346
rect 12716 31282 12768 31288
rect 12912 30734 12940 32710
rect 12992 32564 13044 32570
rect 12992 32506 13044 32512
rect 13004 31346 13032 32506
rect 12992 31340 13044 31346
rect 12992 31282 13044 31288
rect 13084 31340 13136 31346
rect 13084 31282 13136 31288
rect 13096 30734 13124 31282
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12716 30252 12768 30258
rect 12716 30194 12768 30200
rect 12728 29238 12756 30194
rect 12820 29646 12848 30330
rect 13188 30122 13216 35974
rect 13280 35834 13308 36110
rect 13360 36100 13412 36106
rect 13360 36042 13412 36048
rect 13268 35828 13320 35834
rect 13268 35770 13320 35776
rect 13280 32570 13308 35770
rect 13372 34746 13400 36042
rect 13360 34740 13412 34746
rect 13360 34682 13412 34688
rect 13268 32564 13320 32570
rect 13268 32506 13320 32512
rect 13268 30728 13320 30734
rect 13268 30670 13320 30676
rect 13176 30116 13228 30122
rect 13176 30058 13228 30064
rect 13084 30048 13136 30054
rect 13084 29990 13136 29996
rect 12808 29640 12860 29646
rect 12808 29582 12860 29588
rect 12716 29232 12768 29238
rect 12716 29174 12768 29180
rect 12820 29102 12848 29582
rect 12808 29096 12860 29102
rect 12808 29038 12860 29044
rect 12624 28756 12676 28762
rect 12624 28698 12676 28704
rect 12716 28688 12768 28694
rect 12716 28630 12768 28636
rect 12728 27418 12756 28630
rect 12820 28558 12848 29038
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 12820 28150 12848 28494
rect 13096 28490 13124 29990
rect 13176 29572 13228 29578
rect 13176 29514 13228 29520
rect 13188 29306 13216 29514
rect 13176 29300 13228 29306
rect 13176 29242 13228 29248
rect 13280 29050 13308 30670
rect 13452 29164 13504 29170
rect 13452 29106 13504 29112
rect 13188 29034 13308 29050
rect 13176 29028 13308 29034
rect 13228 29022 13308 29028
rect 13176 28970 13228 28976
rect 13084 28484 13136 28490
rect 13084 28426 13136 28432
rect 12808 28144 12860 28150
rect 12808 28086 12860 28092
rect 12728 27390 12848 27418
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12624 26988 12676 26994
rect 12624 26930 12676 26936
rect 12636 26518 12664 26930
rect 12728 26518 12756 27270
rect 12624 26512 12676 26518
rect 12624 26454 12676 26460
rect 12716 26512 12768 26518
rect 12716 26454 12768 26460
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 12360 25498 12388 25842
rect 12544 25838 12572 26250
rect 12728 25974 12756 26454
rect 12820 26382 12848 27390
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12808 26376 12860 26382
rect 12808 26318 12860 26324
rect 12716 25968 12768 25974
rect 12716 25910 12768 25916
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 12348 25492 12400 25498
rect 12348 25434 12400 25440
rect 12544 25362 12572 25774
rect 12624 25696 12676 25702
rect 12624 25638 12676 25644
rect 12348 25356 12400 25362
rect 12348 25298 12400 25304
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12360 24274 12388 25298
rect 12544 24274 12572 25298
rect 12636 25294 12664 25638
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 12532 24268 12584 24274
rect 12532 24210 12584 24216
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 11900 21814 12020 21842
rect 11796 21548 11848 21554
rect 11716 21508 11796 21536
rect 11612 21490 11664 21496
rect 11796 21490 11848 21496
rect 11624 20262 11652 21490
rect 11900 21486 11928 21814
rect 11888 21480 11940 21486
rect 11888 21422 11940 21428
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11348 19378 11376 19654
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11440 18834 11468 19382
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 10880 17436 11188 17456
rect 10880 17434 10886 17436
rect 10942 17434 10966 17436
rect 11022 17434 11046 17436
rect 11102 17434 11126 17436
rect 11182 17434 11188 17436
rect 10942 17382 10944 17434
rect 11124 17382 11126 17434
rect 10880 17380 10886 17382
rect 10942 17380 10966 17382
rect 11022 17380 11046 17382
rect 11102 17380 11126 17382
rect 11182 17380 11188 17382
rect 10880 17360 11188 17380
rect 11256 17270 11284 17818
rect 11244 17264 11296 17270
rect 11244 17206 11296 17212
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10888 16794 10916 17138
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 10880 16348 11188 16368
rect 10880 16346 10886 16348
rect 10942 16346 10966 16348
rect 11022 16346 11046 16348
rect 11102 16346 11126 16348
rect 11182 16346 11188 16348
rect 10942 16294 10944 16346
rect 11124 16294 11126 16346
rect 10880 16292 10886 16294
rect 10942 16292 10966 16294
rect 11022 16292 11046 16294
rect 11102 16292 11126 16294
rect 11182 16292 11188 16294
rect 10880 16272 11188 16292
rect 11256 16182 11284 16390
rect 11440 16250 11468 18770
rect 11624 18766 11652 20198
rect 11900 18834 11928 21422
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 10880 15260 11188 15280
rect 10880 15258 10886 15260
rect 10942 15258 10966 15260
rect 11022 15258 11046 15260
rect 11102 15258 11126 15260
rect 11182 15258 11188 15260
rect 10942 15206 10944 15258
rect 11124 15206 11126 15258
rect 10880 15204 10886 15206
rect 10942 15204 10966 15206
rect 11022 15204 11046 15206
rect 11102 15204 11126 15206
rect 11182 15204 11188 15206
rect 10880 15184 11188 15204
rect 10876 14408 10928 14414
rect 10796 14368 10876 14396
rect 10796 12646 10824 14368
rect 10876 14350 10928 14356
rect 10880 14172 11188 14192
rect 10880 14170 10886 14172
rect 10942 14170 10966 14172
rect 11022 14170 11046 14172
rect 11102 14170 11126 14172
rect 11182 14170 11188 14172
rect 10942 14118 10944 14170
rect 11124 14118 11126 14170
rect 10880 14116 10886 14118
rect 10942 14116 10966 14118
rect 11022 14116 11046 14118
rect 11102 14116 11126 14118
rect 11182 14116 11188 14118
rect 10880 14096 11188 14116
rect 11256 13734 11284 15370
rect 11716 14482 11744 17070
rect 11992 16590 12020 18838
rect 12084 18426 12112 23054
rect 12176 20534 12204 23122
rect 12256 23112 12308 23118
rect 12256 23054 12308 23060
rect 12268 22778 12296 23054
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 12360 22642 12388 23666
rect 12544 23186 12572 24210
rect 12532 23180 12584 23186
rect 12532 23122 12584 23128
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12820 22710 12848 22918
rect 12808 22704 12860 22710
rect 12808 22646 12860 22652
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12360 22030 12388 22578
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12544 21690 12572 22578
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 12176 18834 12204 20470
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12268 18970 12296 19722
rect 12452 18970 12480 20402
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12544 18766 12572 19994
rect 12912 19514 12940 26522
rect 12992 26308 13044 26314
rect 12992 26250 13044 26256
rect 13004 25226 13032 26250
rect 12992 25220 13044 25226
rect 12992 25162 13044 25168
rect 13004 23798 13032 25162
rect 12992 23792 13044 23798
rect 12992 23734 13044 23740
rect 13096 23322 13124 28426
rect 13188 24834 13216 28970
rect 13360 28416 13412 28422
rect 13360 28358 13412 28364
rect 13372 28082 13400 28358
rect 13360 28076 13412 28082
rect 13360 28018 13412 28024
rect 13464 26489 13492 29106
rect 13450 26480 13506 26489
rect 13450 26415 13506 26424
rect 13360 25900 13412 25906
rect 13360 25842 13412 25848
rect 13372 25498 13400 25842
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13556 25362 13584 36518
rect 13740 35018 13768 36518
rect 13728 35012 13780 35018
rect 13728 34954 13780 34960
rect 13832 33318 13860 36722
rect 14372 35488 14424 35494
rect 14372 35430 14424 35436
rect 14188 34536 14240 34542
rect 14188 34478 14240 34484
rect 14004 33924 14056 33930
rect 14004 33866 14056 33872
rect 14016 33590 14044 33866
rect 14004 33584 14056 33590
rect 14004 33526 14056 33532
rect 13820 33312 13872 33318
rect 13820 33254 13872 33260
rect 14200 32298 14228 34478
rect 14384 33930 14412 35430
rect 14648 35080 14700 35086
rect 14648 35022 14700 35028
rect 14464 35012 14516 35018
rect 14464 34954 14516 34960
rect 14476 34610 14504 34954
rect 14660 34950 14688 35022
rect 14936 34950 14964 36722
rect 15212 36310 15240 37130
rect 15304 36718 15332 37198
rect 15292 36712 15344 36718
rect 15292 36654 15344 36660
rect 15200 36304 15252 36310
rect 15200 36246 15252 36252
rect 15212 36174 15240 36246
rect 15304 36242 15332 36654
rect 15292 36236 15344 36242
rect 15292 36178 15344 36184
rect 15200 36168 15252 36174
rect 15200 36110 15252 36116
rect 15212 35222 15240 36110
rect 15200 35216 15252 35222
rect 15200 35158 15252 35164
rect 14648 34944 14700 34950
rect 14648 34886 14700 34892
rect 14924 34944 14976 34950
rect 14924 34886 14976 34892
rect 14464 34604 14516 34610
rect 14464 34546 14516 34552
rect 14660 34542 14688 34886
rect 15212 34626 15240 35158
rect 15396 35154 15424 37266
rect 15764 36242 15792 40326
rect 15846 39740 16154 39760
rect 15846 39738 15852 39740
rect 15908 39738 15932 39740
rect 15988 39738 16012 39740
rect 16068 39738 16092 39740
rect 16148 39738 16154 39740
rect 15908 39686 15910 39738
rect 16090 39686 16092 39738
rect 15846 39684 15852 39686
rect 15908 39684 15932 39686
rect 15988 39684 16012 39686
rect 16068 39684 16092 39686
rect 16148 39684 16154 39686
rect 15846 39664 16154 39684
rect 16224 39098 16252 41074
rect 16764 40928 16816 40934
rect 16764 40870 16816 40876
rect 16304 40588 16356 40594
rect 16304 40530 16356 40536
rect 16316 39982 16344 40530
rect 16580 40452 16632 40458
rect 16580 40394 16632 40400
rect 16304 39976 16356 39982
rect 16304 39918 16356 39924
rect 16316 39506 16344 39918
rect 16304 39500 16356 39506
rect 16304 39442 16356 39448
rect 16212 39092 16264 39098
rect 16212 39034 16264 39040
rect 16316 38894 16344 39442
rect 16592 39030 16620 40394
rect 16776 40050 16804 40870
rect 16868 40050 16896 41074
rect 17408 40520 17460 40526
rect 17408 40462 17460 40468
rect 17040 40384 17092 40390
rect 17040 40326 17092 40332
rect 17132 40384 17184 40390
rect 17132 40326 17184 40332
rect 16764 40044 16816 40050
rect 16764 39986 16816 39992
rect 16856 40044 16908 40050
rect 16856 39986 16908 39992
rect 16856 39908 16908 39914
rect 16856 39850 16908 39856
rect 16868 39642 16896 39850
rect 16856 39636 16908 39642
rect 16856 39578 16908 39584
rect 16868 39506 16896 39578
rect 17052 39506 17080 40326
rect 16856 39500 16908 39506
rect 16856 39442 16908 39448
rect 17040 39500 17092 39506
rect 17040 39442 17092 39448
rect 16580 39024 16632 39030
rect 16580 38966 16632 38972
rect 16304 38888 16356 38894
rect 16304 38830 16356 38836
rect 15846 38652 16154 38672
rect 15846 38650 15852 38652
rect 15908 38650 15932 38652
rect 15988 38650 16012 38652
rect 16068 38650 16092 38652
rect 16148 38650 16154 38652
rect 15908 38598 15910 38650
rect 16090 38598 16092 38650
rect 15846 38596 15852 38598
rect 15908 38596 15932 38598
rect 15988 38596 16012 38598
rect 16068 38596 16092 38598
rect 16148 38596 16154 38598
rect 15846 38576 16154 38596
rect 16212 38004 16264 38010
rect 16212 37946 16264 37952
rect 15846 37564 16154 37584
rect 15846 37562 15852 37564
rect 15908 37562 15932 37564
rect 15988 37562 16012 37564
rect 16068 37562 16092 37564
rect 16148 37562 16154 37564
rect 15908 37510 15910 37562
rect 16090 37510 16092 37562
rect 15846 37508 15852 37510
rect 15908 37508 15932 37510
rect 15988 37508 16012 37510
rect 16068 37508 16092 37510
rect 16148 37508 16154 37510
rect 15846 37488 16154 37508
rect 16120 37324 16172 37330
rect 16224 37312 16252 37946
rect 16316 37330 16344 38830
rect 16764 38752 16816 38758
rect 16764 38694 16816 38700
rect 16172 37284 16252 37312
rect 16120 37266 16172 37272
rect 15846 36476 16154 36496
rect 15846 36474 15852 36476
rect 15908 36474 15932 36476
rect 15988 36474 16012 36476
rect 16068 36474 16092 36476
rect 16148 36474 16154 36476
rect 15908 36422 15910 36474
rect 16090 36422 16092 36474
rect 15846 36420 15852 36422
rect 15908 36420 15932 36422
rect 15988 36420 16012 36422
rect 16068 36420 16092 36422
rect 16148 36420 16154 36422
rect 15846 36400 16154 36420
rect 15752 36236 15804 36242
rect 15752 36178 15804 36184
rect 16120 36236 16172 36242
rect 16224 36224 16252 37284
rect 16304 37324 16356 37330
rect 16304 37266 16356 37272
rect 16172 36196 16252 36224
rect 16120 36178 16172 36184
rect 15764 35766 15792 36178
rect 16316 36174 16344 37266
rect 16580 36712 16632 36718
rect 16580 36654 16632 36660
rect 16304 36168 16356 36174
rect 16304 36110 16356 36116
rect 15752 35760 15804 35766
rect 15752 35702 15804 35708
rect 15384 35148 15436 35154
rect 15384 35090 15436 35096
rect 15212 34610 15332 34626
rect 15212 34604 15344 34610
rect 15212 34598 15292 34604
rect 15292 34546 15344 34552
rect 14648 34536 14700 34542
rect 14648 34478 14700 34484
rect 15016 34468 15068 34474
rect 15068 34428 15240 34456
rect 15016 34410 15068 34416
rect 15212 34134 15240 34428
rect 15200 34128 15252 34134
rect 15200 34070 15252 34076
rect 15396 33946 15424 35090
rect 15660 35080 15712 35086
rect 15660 35022 15712 35028
rect 15672 34950 15700 35022
rect 15660 34944 15712 34950
rect 15660 34886 15712 34892
rect 15660 34536 15712 34542
rect 15660 34478 15712 34484
rect 14372 33924 14424 33930
rect 14372 33866 14424 33872
rect 14556 33924 14608 33930
rect 15396 33918 15516 33946
rect 14556 33866 14608 33872
rect 14568 33522 14596 33866
rect 15384 33856 15436 33862
rect 15384 33798 15436 33804
rect 15396 33522 15424 33798
rect 14280 33516 14332 33522
rect 14280 33458 14332 33464
rect 14556 33516 14608 33522
rect 14556 33458 14608 33464
rect 15384 33516 15436 33522
rect 15384 33458 15436 33464
rect 14188 32292 14240 32298
rect 14188 32234 14240 32240
rect 13820 32224 13872 32230
rect 13820 32166 13872 32172
rect 13832 32042 13860 32166
rect 13740 32014 13860 32042
rect 13740 31890 13768 32014
rect 13832 31890 13952 31906
rect 13728 31884 13780 31890
rect 13728 31826 13780 31832
rect 13820 31884 13952 31890
rect 13872 31878 13952 31884
rect 13820 31826 13872 31832
rect 13820 31748 13872 31754
rect 13820 31690 13872 31696
rect 13832 31482 13860 31690
rect 13924 31686 13952 31878
rect 14096 31884 14148 31890
rect 14096 31826 14148 31832
rect 13912 31680 13964 31686
rect 13912 31622 13964 31628
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 14004 31340 14056 31346
rect 14004 31282 14056 31288
rect 13728 31272 13780 31278
rect 13728 31214 13780 31220
rect 13740 30734 13768 31214
rect 13820 31136 13872 31142
rect 13820 31078 13872 31084
rect 13728 30728 13780 30734
rect 13728 30670 13780 30676
rect 13740 30258 13768 30670
rect 13728 30252 13780 30258
rect 13728 30194 13780 30200
rect 13636 27668 13688 27674
rect 13636 27610 13688 27616
rect 13544 25356 13596 25362
rect 13544 25298 13596 25304
rect 13268 25288 13320 25294
rect 13360 25288 13412 25294
rect 13268 25230 13320 25236
rect 13358 25256 13360 25265
rect 13412 25256 13414 25265
rect 13280 24954 13308 25230
rect 13358 25191 13414 25200
rect 13648 24954 13676 27610
rect 13832 25974 13860 31078
rect 14016 29102 14044 31282
rect 14108 30258 14136 31826
rect 14292 30870 14320 33458
rect 14372 33312 14424 33318
rect 14372 33254 14424 33260
rect 14280 30864 14332 30870
rect 14280 30806 14332 30812
rect 14384 30716 14412 33254
rect 14568 32416 14596 33458
rect 15396 33114 15424 33458
rect 15488 33114 15516 33918
rect 15384 33108 15436 33114
rect 15384 33050 15436 33056
rect 15476 33108 15528 33114
rect 15476 33050 15528 33056
rect 14648 32564 14700 32570
rect 14648 32506 14700 32512
rect 14660 32434 14688 32506
rect 15488 32502 15516 33050
rect 15476 32496 15528 32502
rect 15476 32438 15528 32444
rect 14476 32388 14596 32416
rect 14648 32428 14700 32434
rect 14476 32026 14504 32388
rect 14648 32370 14700 32376
rect 15384 32428 15436 32434
rect 15384 32370 15436 32376
rect 14464 32020 14516 32026
rect 14464 31962 14516 31968
rect 14556 31476 14608 31482
rect 14556 31418 14608 31424
rect 14464 31340 14516 31346
rect 14464 31282 14516 31288
rect 14476 31142 14504 31282
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14568 30734 14596 31418
rect 14464 30728 14516 30734
rect 14384 30688 14464 30716
rect 14464 30670 14516 30676
rect 14556 30728 14608 30734
rect 14556 30670 14608 30676
rect 14568 30394 14596 30670
rect 14556 30388 14608 30394
rect 14556 30330 14608 30336
rect 14096 30252 14148 30258
rect 14096 30194 14148 30200
rect 14108 29714 14136 30194
rect 14096 29708 14148 29714
rect 14096 29650 14148 29656
rect 14004 29096 14056 29102
rect 14004 29038 14056 29044
rect 14004 28484 14056 28490
rect 14004 28426 14056 28432
rect 13820 25968 13872 25974
rect 13820 25910 13872 25916
rect 13268 24948 13320 24954
rect 13268 24890 13320 24896
rect 13636 24948 13688 24954
rect 13636 24890 13688 24896
rect 13188 24806 13308 24834
rect 13176 24064 13228 24070
rect 13176 24006 13228 24012
rect 13188 23798 13216 24006
rect 13176 23792 13228 23798
rect 13176 23734 13228 23740
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 12992 23044 13044 23050
rect 12992 22986 13044 22992
rect 13004 22234 13032 22986
rect 12992 22228 13044 22234
rect 12992 22170 13044 22176
rect 13004 21622 13032 22170
rect 13280 22094 13308 24806
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13740 22778 13768 23054
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 13096 22066 13308 22094
rect 12992 21616 13044 21622
rect 12992 21558 13044 21564
rect 13096 20466 13124 22066
rect 13740 21554 13768 22714
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12728 18358 12756 18702
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 17270 12572 17478
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12070 15192 12126 15201
rect 12070 15127 12126 15136
rect 12084 14550 12112 15127
rect 12544 15026 12572 15302
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12360 14906 12388 14962
rect 12360 14878 12480 14906
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11532 14074 11560 14350
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11440 13977 11468 14010
rect 11426 13968 11482 13977
rect 11426 13903 11482 13912
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 10880 13084 11188 13104
rect 10880 13082 10886 13084
rect 10942 13082 10966 13084
rect 11022 13082 11046 13084
rect 11102 13082 11126 13084
rect 11182 13082 11188 13084
rect 10942 13030 10944 13082
rect 11124 13030 11126 13082
rect 10880 13028 10886 13030
rect 10942 13028 10966 13030
rect 11022 13028 11046 13030
rect 11102 13028 11126 13030
rect 11182 13028 11188 13030
rect 10880 13008 11188 13028
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 11256 12345 11284 13670
rect 12084 13530 12112 13806
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11348 12714 11376 13262
rect 12176 12918 12204 14418
rect 12452 14278 12480 14878
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12636 13190 12664 18226
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12820 16590 12848 16934
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12820 16114 12848 16526
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12820 14006 12848 14894
rect 13096 14346 13124 16458
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12820 13258 12848 13670
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12624 13184 12676 13190
rect 12820 13138 12848 13194
rect 12624 13126 12676 13132
rect 12728 13110 12848 13138
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11242 12336 11298 12345
rect 11242 12271 11298 12280
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 10880 11996 11188 12016
rect 10880 11994 10886 11996
rect 10942 11994 10966 11996
rect 11022 11994 11046 11996
rect 11102 11994 11126 11996
rect 11182 11994 11188 11996
rect 10942 11942 10944 11994
rect 11124 11942 11126 11994
rect 10880 11940 10886 11942
rect 10942 11940 10966 11942
rect 11022 11940 11046 11942
rect 11102 11940 11126 11942
rect 11182 11940 11188 11942
rect 10880 11920 11188 11940
rect 11256 11898 11284 12106
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11348 11898 11376 12038
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 10612 11206 10732 11234
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10612 7750 10640 11206
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10704 10810 10732 11018
rect 10880 10908 11188 10928
rect 10880 10906 10886 10908
rect 10942 10906 10966 10908
rect 11022 10906 11046 10908
rect 11102 10906 11126 10908
rect 11182 10906 11188 10908
rect 10942 10854 10944 10906
rect 11124 10854 11126 10906
rect 10880 10852 10886 10854
rect 10942 10852 10966 10854
rect 11022 10852 11046 10854
rect 11102 10852 11126 10854
rect 11182 10852 11188 10854
rect 10880 10832 11188 10852
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10796 10062 10824 10746
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 10980 10198 11008 10474
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10704 9654 10732 9862
rect 10880 9820 11188 9840
rect 10880 9818 10886 9820
rect 10942 9818 10966 9820
rect 11022 9818 11046 9820
rect 11102 9818 11126 9820
rect 11182 9818 11188 9820
rect 10942 9766 10944 9818
rect 11124 9766 11126 9818
rect 10880 9764 10886 9766
rect 10942 9764 10966 9766
rect 11022 9764 11046 9766
rect 11102 9764 11126 9766
rect 11182 9764 11188 9766
rect 10880 9744 11188 9764
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10880 8732 11188 8752
rect 10880 8730 10886 8732
rect 10942 8730 10966 8732
rect 11022 8730 11046 8732
rect 11102 8730 11126 8732
rect 11182 8730 11188 8732
rect 10942 8678 10944 8730
rect 11124 8678 11126 8730
rect 10880 8676 10886 8678
rect 10942 8676 10966 8678
rect 11022 8676 11046 8678
rect 11102 8676 11126 8678
rect 11182 8676 11188 8678
rect 10880 8656 11188 8676
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10704 7818 10732 8434
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10612 7342 10640 7686
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10598 6760 10654 6769
rect 10598 6695 10654 6704
rect 10612 6390 10640 6695
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10520 4622 10548 6258
rect 10600 5296 10652 5302
rect 10600 5238 10652 5244
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10428 4146 10456 4422
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10612 4078 10640 5238
rect 10704 4826 10732 7754
rect 10880 7644 11188 7664
rect 10880 7642 10886 7644
rect 10942 7642 10966 7644
rect 11022 7642 11046 7644
rect 11102 7642 11126 7644
rect 11182 7642 11188 7644
rect 10942 7590 10944 7642
rect 11124 7590 11126 7642
rect 10880 7588 10886 7590
rect 10942 7588 10966 7590
rect 11022 7588 11046 7590
rect 11102 7588 11126 7590
rect 11182 7588 11188 7590
rect 10880 7568 11188 7588
rect 10880 6556 11188 6576
rect 10880 6554 10886 6556
rect 10942 6554 10966 6556
rect 11022 6554 11046 6556
rect 11102 6554 11126 6556
rect 11182 6554 11188 6556
rect 10942 6502 10944 6554
rect 11124 6502 11126 6554
rect 10880 6500 10886 6502
rect 10942 6500 10966 6502
rect 11022 6500 11046 6502
rect 11102 6500 11126 6502
rect 11182 6500 11188 6502
rect 10880 6480 11188 6500
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10796 4146 10824 6326
rect 10980 6254 11008 6326
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 11256 5710 11284 11562
rect 11808 11218 11836 12786
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11900 11694 11928 12650
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11428 10668 11480 10674
rect 11532 10656 11560 10950
rect 11624 10742 11652 10950
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11480 10628 11560 10656
rect 11428 10610 11480 10616
rect 11532 10266 11560 10628
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11348 8566 11376 9046
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11440 7478 11468 8910
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11532 7954 11560 8774
rect 11716 8634 11744 10610
rect 11900 10606 11928 11630
rect 11992 10674 12020 12718
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11900 8362 11928 8978
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11992 8430 12020 8910
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11900 7954 11928 8298
rect 11992 8090 12020 8366
rect 12084 8090 12112 12786
rect 12176 12434 12204 12854
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12176 12406 12296 12434
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12176 11150 12204 12310
rect 12268 12238 12296 12406
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12268 11762 12296 12174
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11830 12388 12038
rect 12636 11830 12664 12582
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12360 10742 12388 11766
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12268 9994 12296 10406
rect 12452 10062 12480 11494
rect 12728 10810 12756 13110
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13004 12238 13032 12786
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 11898 12940 12038
rect 13004 11898 13032 12174
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 12900 11144 12952 11150
rect 12820 11104 12900 11132
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12636 10198 12664 10610
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8634 12204 8774
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11992 7970 12020 8026
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11888 7948 11940 7954
rect 11992 7942 12112 7970
rect 11888 7890 11940 7896
rect 11900 7834 11928 7890
rect 11704 7812 11756 7818
rect 11900 7806 12020 7834
rect 11704 7754 11756 7760
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11716 7410 11744 7754
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11808 6798 11836 7686
rect 11900 7002 11928 7686
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 10880 5468 11188 5488
rect 10880 5466 10886 5468
rect 10942 5466 10966 5468
rect 11022 5466 11046 5468
rect 11102 5466 11126 5468
rect 11182 5466 11188 5468
rect 10942 5414 10944 5466
rect 11124 5414 11126 5466
rect 10880 5412 10886 5414
rect 10942 5412 10966 5414
rect 11022 5412 11046 5414
rect 11102 5412 11126 5414
rect 11182 5412 11188 5414
rect 10880 5392 11188 5412
rect 11256 5234 11284 5510
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 10880 4380 11188 4400
rect 10880 4378 10886 4380
rect 10942 4378 10966 4380
rect 11022 4378 11046 4380
rect 11102 4378 11126 4380
rect 11182 4378 11188 4380
rect 10942 4326 10944 4378
rect 11124 4326 11126 4378
rect 10880 4324 10886 4326
rect 10942 4324 10966 4326
rect 11022 4324 11046 4326
rect 11102 4324 11126 4326
rect 11182 4324 11188 4326
rect 10880 4304 11188 4324
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10796 3738 10824 4082
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10796 3126 10824 3538
rect 10888 3534 10916 3878
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10880 3292 11188 3312
rect 10880 3290 10886 3292
rect 10942 3290 10966 3292
rect 11022 3290 11046 3292
rect 11102 3290 11126 3292
rect 11182 3290 11188 3292
rect 10942 3238 10944 3290
rect 11124 3238 11126 3290
rect 10880 3236 10886 3238
rect 10942 3236 10966 3238
rect 11022 3236 11046 3238
rect 11102 3236 11126 3238
rect 11182 3236 11188 3238
rect 10880 3216 11188 3236
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 9968 2746 10272 2774
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 9968 2514 9996 2746
rect 11440 2582 11468 6734
rect 11992 6254 12020 7806
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 12084 6066 12112 7942
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12452 7018 12480 7278
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12360 6990 12480 7018
rect 12360 6254 12388 6990
rect 12544 6730 12572 7142
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 11992 6038 12112 6066
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 11532 5370 11560 5578
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11532 3466 11560 5102
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11624 3194 11652 4490
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11716 3058 11744 5170
rect 11808 4010 11836 5646
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11900 4078 11928 4490
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 11900 3534 11928 4014
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11716 2650 11744 2994
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11428 2576 11480 2582
rect 11428 2518 11480 2524
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 7944 800 7972 2382
rect 8772 800 8800 2382
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 9416 1426 9444 2314
rect 9404 1420 9456 1426
rect 9404 1362 9456 1368
rect 9508 800 9536 2382
rect 10244 800 10272 2382
rect 10880 2204 11188 2224
rect 10880 2202 10886 2204
rect 10942 2202 10966 2204
rect 11022 2202 11046 2204
rect 11102 2202 11126 2204
rect 11182 2202 11188 2204
rect 10942 2150 10944 2202
rect 11124 2150 11126 2202
rect 10880 2148 10886 2150
rect 10942 2148 10966 2150
rect 11022 2148 11046 2150
rect 11102 2148 11126 2150
rect 11182 2148 11188 2150
rect 10880 2128 11188 2148
rect 11060 1420 11112 1426
rect 11060 1362 11112 1368
rect 11072 800 11100 1362
rect 11808 800 11836 2926
rect 11992 2514 12020 6038
rect 12452 5778 12480 6122
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12544 5098 12572 6666
rect 12636 6390 12664 9862
rect 12820 6934 12848 11104
rect 12900 11086 12952 11092
rect 13004 10674 13032 11222
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13004 10062 13032 10610
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13004 9518 13032 9998
rect 13096 9602 13124 13874
rect 13188 9722 13216 19450
rect 13280 19446 13308 20198
rect 13372 20058 13400 20878
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13464 19786 13492 20402
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13556 19514 13584 19790
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13268 19440 13320 19446
rect 13268 19382 13320 19388
rect 13280 17678 13308 19382
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13280 17338 13308 17614
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13372 16454 13400 16662
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 16046 13400 16390
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13280 15026 13308 15846
rect 13372 15502 13400 15982
rect 13464 15910 13492 16662
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13280 14414 13308 14758
rect 13372 14550 13400 15438
rect 13556 15026 13584 17546
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13280 10606 13308 11086
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13280 9722 13308 10542
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13096 9574 13216 9602
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 8634 12940 8774
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12912 8090 12940 8434
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12808 6928 12860 6934
rect 12808 6870 12860 6876
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12728 6474 12756 6734
rect 12728 6446 12848 6474
rect 12820 6390 12848 6446
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12084 4146 12112 4422
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 12084 2310 12112 4082
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12176 3398 12204 4014
rect 12452 3942 12480 4490
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12544 4146 12572 4422
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12636 4078 12664 6190
rect 12820 5166 12848 6326
rect 12912 5778 12940 7346
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 13004 6798 13032 7142
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13096 6186 13124 9386
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12912 5234 12940 5714
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 13096 5370 13124 5510
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12820 4078 12848 5102
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 3738 12480 3878
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12452 3534 12480 3674
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 12544 800 12572 3946
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 3058 13032 3470
rect 13096 3058 13124 4626
rect 13188 3602 13216 9574
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13280 8974 13308 9318
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13372 5642 13400 13806
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13464 5914 13492 10610
rect 13648 9586 13676 18566
rect 14016 18290 14044 28426
rect 14108 28150 14136 29650
rect 14660 29306 14688 32370
rect 15108 32224 15160 32230
rect 15108 32166 15160 32172
rect 15120 31958 15148 32166
rect 15108 31952 15160 31958
rect 15108 31894 15160 31900
rect 15120 31754 15148 31894
rect 15396 31822 15424 32370
rect 15384 31816 15436 31822
rect 15384 31758 15436 31764
rect 14936 31726 15148 31754
rect 14740 31136 14792 31142
rect 14740 31078 14792 31084
rect 14752 30258 14780 31078
rect 14740 30252 14792 30258
rect 14740 30194 14792 30200
rect 14648 29300 14700 29306
rect 14648 29242 14700 29248
rect 14660 28762 14688 29242
rect 14740 29164 14792 29170
rect 14740 29106 14792 29112
rect 14648 28756 14700 28762
rect 14648 28698 14700 28704
rect 14464 28620 14516 28626
rect 14464 28562 14516 28568
rect 14476 28218 14504 28562
rect 14752 28558 14780 29106
rect 14740 28552 14792 28558
rect 14740 28494 14792 28500
rect 14464 28212 14516 28218
rect 14464 28154 14516 28160
rect 14096 28144 14148 28150
rect 14096 28086 14148 28092
rect 14280 27600 14332 27606
rect 14280 27542 14332 27548
rect 14476 27554 14504 28154
rect 14648 28076 14700 28082
rect 14648 28018 14700 28024
rect 14292 26858 14320 27542
rect 14476 27526 14596 27554
rect 14568 27470 14596 27526
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14384 26926 14412 27406
rect 14372 26920 14424 26926
rect 14372 26862 14424 26868
rect 14280 26852 14332 26858
rect 14280 26794 14332 26800
rect 14292 26586 14320 26794
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14384 26314 14412 26862
rect 14568 26450 14596 27406
rect 14660 26586 14688 28018
rect 14648 26580 14700 26586
rect 14648 26522 14700 26528
rect 14556 26444 14608 26450
rect 14556 26386 14608 26392
rect 14372 26308 14424 26314
rect 14372 26250 14424 26256
rect 14384 25906 14412 26250
rect 14372 25900 14424 25906
rect 14372 25842 14424 25848
rect 14660 24206 14688 26522
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14752 24410 14780 24754
rect 14740 24404 14792 24410
rect 14740 24346 14792 24352
rect 14280 24200 14332 24206
rect 14648 24200 14700 24206
rect 14280 24142 14332 24148
rect 14568 24160 14648 24188
rect 14292 23866 14320 24142
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 14292 23186 14320 23666
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 14292 22778 14320 23122
rect 14568 23050 14596 24160
rect 14648 24142 14700 24148
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14752 23050 14780 23802
rect 14556 23044 14608 23050
rect 14556 22986 14608 22992
rect 14740 23044 14792 23050
rect 14740 22986 14792 22992
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14372 21888 14424 21894
rect 14372 21830 14424 21836
rect 14096 20324 14148 20330
rect 14096 20266 14148 20272
rect 14108 19854 14136 20266
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14200 18766 14228 19110
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13740 16998 13768 17274
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 13938 13768 16934
rect 13924 16590 13952 17206
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13912 16584 13964 16590
rect 13912 16526 13964 16532
rect 14016 16250 14044 17138
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 14108 16114 14136 17614
rect 14200 17134 14228 18702
rect 14384 17746 14412 21830
rect 14936 20924 14964 31726
rect 15396 31482 15424 31758
rect 15476 31680 15528 31686
rect 15476 31622 15528 31628
rect 15384 31476 15436 31482
rect 15384 31418 15436 31424
rect 15200 31340 15252 31346
rect 15200 31282 15252 31288
rect 15108 30728 15160 30734
rect 15108 30670 15160 30676
rect 15120 29782 15148 30670
rect 15108 29776 15160 29782
rect 15108 29718 15160 29724
rect 15120 29102 15148 29718
rect 15108 29096 15160 29102
rect 15108 29038 15160 29044
rect 15120 28694 15148 29038
rect 15108 28688 15160 28694
rect 15108 28630 15160 28636
rect 15212 28490 15240 31282
rect 15488 31210 15516 31622
rect 15568 31408 15620 31414
rect 15568 31350 15620 31356
rect 15476 31204 15528 31210
rect 15476 31146 15528 31152
rect 15488 29594 15516 31146
rect 15580 30122 15608 31350
rect 15568 30116 15620 30122
rect 15568 30058 15620 30064
rect 15396 29566 15516 29594
rect 15200 28484 15252 28490
rect 15200 28426 15252 28432
rect 15016 26988 15068 26994
rect 15016 26930 15068 26936
rect 15108 26988 15160 26994
rect 15108 26930 15160 26936
rect 15028 26586 15056 26930
rect 15016 26580 15068 26586
rect 15016 26522 15068 26528
rect 15120 26042 15148 26930
rect 15108 26036 15160 26042
rect 15108 25978 15160 25984
rect 15212 25922 15240 28426
rect 15292 27872 15344 27878
rect 15292 27814 15344 27820
rect 15304 27470 15332 27814
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 15120 25894 15240 25922
rect 15120 25276 15148 25894
rect 15200 25832 15252 25838
rect 15200 25774 15252 25780
rect 15212 25430 15240 25774
rect 15200 25424 15252 25430
rect 15200 25366 15252 25372
rect 15292 25288 15344 25294
rect 15120 25248 15240 25276
rect 15016 24676 15068 24682
rect 15016 24618 15068 24624
rect 15028 24070 15056 24618
rect 15108 24608 15160 24614
rect 15212 24596 15240 25248
rect 15292 25230 15344 25236
rect 15396 25242 15424 29566
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 15488 29238 15516 29446
rect 15476 29232 15528 29238
rect 15476 29174 15528 29180
rect 15672 27538 15700 34478
rect 15764 34134 15792 35702
rect 15846 35388 16154 35408
rect 15846 35386 15852 35388
rect 15908 35386 15932 35388
rect 15988 35386 16012 35388
rect 16068 35386 16092 35388
rect 16148 35386 16154 35388
rect 15908 35334 15910 35386
rect 16090 35334 16092 35386
rect 15846 35332 15852 35334
rect 15908 35332 15932 35334
rect 15988 35332 16012 35334
rect 16068 35332 16092 35334
rect 16148 35332 16154 35334
rect 15846 35312 16154 35332
rect 16316 35154 16344 36110
rect 16592 36038 16620 36654
rect 16580 36032 16632 36038
rect 16580 35974 16632 35980
rect 16592 35850 16620 35974
rect 16592 35822 16712 35850
rect 16580 35692 16632 35698
rect 16580 35634 16632 35640
rect 16592 35290 16620 35634
rect 16684 35630 16712 35822
rect 16672 35624 16724 35630
rect 16672 35566 16724 35572
rect 16580 35284 16632 35290
rect 16580 35226 16632 35232
rect 16304 35148 16356 35154
rect 16304 35090 16356 35096
rect 15936 35080 15988 35086
rect 15856 35040 15936 35068
rect 15856 34542 15884 35040
rect 15936 35022 15988 35028
rect 15844 34536 15896 34542
rect 15844 34478 15896 34484
rect 15846 34300 16154 34320
rect 15846 34298 15852 34300
rect 15908 34298 15932 34300
rect 15988 34298 16012 34300
rect 16068 34298 16092 34300
rect 16148 34298 16154 34300
rect 15908 34246 15910 34298
rect 16090 34246 16092 34298
rect 15846 34244 15852 34246
rect 15908 34244 15932 34246
rect 15988 34244 16012 34246
rect 16068 34244 16092 34246
rect 16148 34244 16154 34246
rect 15846 34224 16154 34244
rect 15752 34128 15804 34134
rect 15752 34070 15804 34076
rect 15846 33212 16154 33232
rect 15846 33210 15852 33212
rect 15908 33210 15932 33212
rect 15988 33210 16012 33212
rect 16068 33210 16092 33212
rect 16148 33210 16154 33212
rect 15908 33158 15910 33210
rect 16090 33158 16092 33210
rect 15846 33156 15852 33158
rect 15908 33156 15932 33158
rect 15988 33156 16012 33158
rect 16068 33156 16092 33158
rect 16148 33156 16154 33158
rect 15846 33136 16154 33156
rect 15752 32836 15804 32842
rect 15752 32778 15804 32784
rect 15764 32570 15792 32778
rect 15752 32564 15804 32570
rect 15752 32506 15804 32512
rect 15752 32428 15804 32434
rect 15752 32370 15804 32376
rect 16580 32428 16632 32434
rect 16580 32370 16632 32376
rect 15764 32026 15792 32370
rect 15846 32124 16154 32144
rect 15846 32122 15852 32124
rect 15908 32122 15932 32124
rect 15988 32122 16012 32124
rect 16068 32122 16092 32124
rect 16148 32122 16154 32124
rect 15908 32070 15910 32122
rect 16090 32070 16092 32122
rect 15846 32068 15852 32070
rect 15908 32068 15932 32070
rect 15988 32068 16012 32070
rect 16068 32068 16092 32070
rect 16148 32068 16154 32070
rect 15846 32048 16154 32068
rect 15752 32020 15804 32026
rect 15752 31962 15804 31968
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 15846 31036 16154 31056
rect 15846 31034 15852 31036
rect 15908 31034 15932 31036
rect 15988 31034 16012 31036
rect 16068 31034 16092 31036
rect 16148 31034 16154 31036
rect 15908 30982 15910 31034
rect 16090 30982 16092 31034
rect 15846 30980 15852 30982
rect 15908 30980 15932 30982
rect 15988 30980 16012 30982
rect 16068 30980 16092 30982
rect 16148 30980 16154 30982
rect 15846 30960 16154 30980
rect 16212 30660 16264 30666
rect 16212 30602 16264 30608
rect 16224 30394 16252 30602
rect 16212 30388 16264 30394
rect 16212 30330 16264 30336
rect 15846 29948 16154 29968
rect 15846 29946 15852 29948
rect 15908 29946 15932 29948
rect 15988 29946 16012 29948
rect 16068 29946 16092 29948
rect 16148 29946 16154 29948
rect 15908 29894 15910 29946
rect 16090 29894 16092 29946
rect 15846 29892 15852 29894
rect 15908 29892 15932 29894
rect 15988 29892 16012 29894
rect 16068 29892 16092 29894
rect 16148 29892 16154 29894
rect 15846 29872 16154 29892
rect 15846 28860 16154 28880
rect 15846 28858 15852 28860
rect 15908 28858 15932 28860
rect 15988 28858 16012 28860
rect 16068 28858 16092 28860
rect 16148 28858 16154 28860
rect 15908 28806 15910 28858
rect 16090 28806 16092 28858
rect 15846 28804 15852 28806
rect 15908 28804 15932 28806
rect 15988 28804 16012 28806
rect 16068 28804 16092 28806
rect 16148 28804 16154 28806
rect 15846 28784 16154 28804
rect 16224 28694 16252 30330
rect 16212 28688 16264 28694
rect 16212 28630 16264 28636
rect 15752 28076 15804 28082
rect 15752 28018 15804 28024
rect 16212 28076 16264 28082
rect 16212 28018 16264 28024
rect 15660 27532 15712 27538
rect 15660 27474 15712 27480
rect 15568 27328 15620 27334
rect 15566 27296 15568 27305
rect 15620 27296 15622 27305
rect 15566 27231 15622 27240
rect 15568 27056 15620 27062
rect 15568 26998 15620 27004
rect 15580 26450 15608 26998
rect 15672 26926 15700 27474
rect 15660 26920 15712 26926
rect 15660 26862 15712 26868
rect 15568 26444 15620 26450
rect 15568 26386 15620 26392
rect 15304 24750 15332 25230
rect 15396 25214 15516 25242
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15292 24744 15344 24750
rect 15292 24686 15344 24692
rect 15212 24568 15332 24596
rect 15108 24550 15160 24556
rect 15120 24138 15148 24550
rect 15108 24132 15160 24138
rect 15108 24074 15160 24080
rect 15016 24064 15068 24070
rect 15016 24006 15068 24012
rect 15028 23322 15056 24006
rect 15108 23792 15160 23798
rect 15108 23734 15160 23740
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 15120 21418 15148 23734
rect 15304 22080 15332 24568
rect 15396 24342 15424 25094
rect 15488 24750 15516 25214
rect 15580 24818 15608 26386
rect 15764 25974 15792 28018
rect 15846 27772 16154 27792
rect 15846 27770 15852 27772
rect 15908 27770 15932 27772
rect 15988 27770 16012 27772
rect 16068 27770 16092 27772
rect 16148 27770 16154 27772
rect 15908 27718 15910 27770
rect 16090 27718 16092 27770
rect 15846 27716 15852 27718
rect 15908 27716 15932 27718
rect 15988 27716 16012 27718
rect 16068 27716 16092 27718
rect 16148 27716 16154 27718
rect 15846 27696 16154 27716
rect 16224 27674 16252 28018
rect 16212 27668 16264 27674
rect 16212 27610 16264 27616
rect 15846 26684 16154 26704
rect 15846 26682 15852 26684
rect 15908 26682 15932 26684
rect 15988 26682 16012 26684
rect 16068 26682 16092 26684
rect 16148 26682 16154 26684
rect 15908 26630 15910 26682
rect 16090 26630 16092 26682
rect 15846 26628 15852 26630
rect 15908 26628 15932 26630
rect 15988 26628 16012 26630
rect 16068 26628 16092 26630
rect 16148 26628 16154 26630
rect 15846 26608 16154 26628
rect 15752 25968 15804 25974
rect 15752 25910 15804 25916
rect 15752 25696 15804 25702
rect 15752 25638 15804 25644
rect 15660 25424 15712 25430
rect 15660 25366 15712 25372
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 15476 24744 15528 24750
rect 15476 24686 15528 24692
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15384 24336 15436 24342
rect 15384 24278 15436 24284
rect 15488 24274 15516 24550
rect 15580 24342 15608 24754
rect 15568 24336 15620 24342
rect 15568 24278 15620 24284
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 15568 24200 15620 24206
rect 15488 24148 15568 24154
rect 15488 24142 15620 24148
rect 15488 24126 15608 24142
rect 15488 23662 15516 24126
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 15488 22166 15516 23598
rect 15580 23322 15608 23598
rect 15568 23316 15620 23322
rect 15568 23258 15620 23264
rect 15672 22642 15700 25366
rect 15764 23118 15792 25638
rect 15846 25596 16154 25616
rect 15846 25594 15852 25596
rect 15908 25594 15932 25596
rect 15988 25594 16012 25596
rect 16068 25594 16092 25596
rect 16148 25594 16154 25596
rect 15908 25542 15910 25594
rect 16090 25542 16092 25594
rect 15846 25540 15852 25542
rect 15908 25540 15932 25542
rect 15988 25540 16012 25542
rect 16068 25540 16092 25542
rect 16148 25540 16154 25542
rect 15846 25520 16154 25540
rect 15846 24508 16154 24528
rect 15846 24506 15852 24508
rect 15908 24506 15932 24508
rect 15988 24506 16012 24508
rect 16068 24506 16092 24508
rect 16148 24506 16154 24508
rect 15908 24454 15910 24506
rect 16090 24454 16092 24506
rect 15846 24452 15852 24454
rect 15908 24452 15932 24454
rect 15988 24452 16012 24454
rect 16068 24452 16092 24454
rect 16148 24452 16154 24454
rect 15846 24432 16154 24452
rect 16120 24064 16172 24070
rect 16120 24006 16172 24012
rect 16132 23662 16160 24006
rect 16316 23798 16344 31282
rect 16396 28008 16448 28014
rect 16396 27950 16448 27956
rect 16408 27538 16436 27950
rect 16396 27532 16448 27538
rect 16396 27474 16448 27480
rect 16408 25498 16436 27474
rect 16488 25900 16540 25906
rect 16488 25842 16540 25848
rect 16396 25492 16448 25498
rect 16396 25434 16448 25440
rect 16408 24274 16436 25434
rect 16500 25158 16528 25842
rect 16488 25152 16540 25158
rect 16488 25094 16540 25100
rect 16592 25106 16620 32370
rect 16672 31340 16724 31346
rect 16672 31282 16724 31288
rect 16684 30394 16712 31282
rect 16672 30388 16724 30394
rect 16672 30330 16724 30336
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16684 28218 16712 29106
rect 16672 28212 16724 28218
rect 16672 28154 16724 28160
rect 16672 27328 16724 27334
rect 16672 27270 16724 27276
rect 16684 27130 16712 27270
rect 16672 27124 16724 27130
rect 16672 27066 16724 27072
rect 16776 25498 16804 38694
rect 16868 36718 16896 39442
rect 17144 38962 17172 40326
rect 17420 39982 17448 40462
rect 17592 40452 17644 40458
rect 17592 40394 17644 40400
rect 17604 40050 17632 40394
rect 17868 40180 17920 40186
rect 17868 40122 17920 40128
rect 17592 40044 17644 40050
rect 17592 39986 17644 39992
rect 17408 39976 17460 39982
rect 17408 39918 17460 39924
rect 17420 39098 17448 39918
rect 17776 39840 17828 39846
rect 17776 39782 17828 39788
rect 17684 39296 17736 39302
rect 17684 39238 17736 39244
rect 17696 39098 17724 39238
rect 17788 39098 17816 39782
rect 17880 39370 17908 40122
rect 19340 40044 19392 40050
rect 19340 39986 19392 39992
rect 18052 39976 18104 39982
rect 18052 39918 18104 39924
rect 18064 39642 18092 39918
rect 18972 39840 19024 39846
rect 18972 39782 19024 39788
rect 18052 39636 18104 39642
rect 18052 39578 18104 39584
rect 18788 39568 18840 39574
rect 18788 39510 18840 39516
rect 18144 39432 18196 39438
rect 18144 39374 18196 39380
rect 17868 39364 17920 39370
rect 17868 39306 17920 39312
rect 17408 39092 17460 39098
rect 17408 39034 17460 39040
rect 17684 39092 17736 39098
rect 17684 39034 17736 39040
rect 17776 39092 17828 39098
rect 17776 39034 17828 39040
rect 17132 38956 17184 38962
rect 17132 38898 17184 38904
rect 17788 38350 17816 39034
rect 17960 38888 18012 38894
rect 17960 38830 18012 38836
rect 17776 38344 17828 38350
rect 17776 38286 17828 38292
rect 17684 37868 17736 37874
rect 17684 37810 17736 37816
rect 17696 37262 17724 37810
rect 17972 37330 18000 38830
rect 18156 38554 18184 39374
rect 18800 39098 18828 39510
rect 18984 39098 19012 39782
rect 18788 39092 18840 39098
rect 18788 39034 18840 39040
rect 18972 39092 19024 39098
rect 18972 39034 19024 39040
rect 18144 38548 18196 38554
rect 18144 38490 18196 38496
rect 18800 38350 18828 39034
rect 19156 38752 19208 38758
rect 19156 38694 19208 38700
rect 18788 38344 18840 38350
rect 18788 38286 18840 38292
rect 18512 37664 18564 37670
rect 18512 37606 18564 37612
rect 17960 37324 18012 37330
rect 17960 37266 18012 37272
rect 18524 37262 18552 37606
rect 17684 37256 17736 37262
rect 17684 37198 17736 37204
rect 18512 37256 18564 37262
rect 18512 37198 18564 37204
rect 18788 37256 18840 37262
rect 18788 37198 18840 37204
rect 16948 37120 17000 37126
rect 16948 37062 17000 37068
rect 16960 36922 16988 37062
rect 17696 36922 17724 37198
rect 18144 37120 18196 37126
rect 18144 37062 18196 37068
rect 16948 36916 17000 36922
rect 16948 36858 17000 36864
rect 17684 36916 17736 36922
rect 17684 36858 17736 36864
rect 16856 36712 16908 36718
rect 16856 36654 16908 36660
rect 17132 36712 17184 36718
rect 17132 36654 17184 36660
rect 17144 36378 17172 36654
rect 17132 36372 17184 36378
rect 17132 36314 17184 36320
rect 16948 35624 17000 35630
rect 16948 35566 17000 35572
rect 16960 34746 16988 35566
rect 17316 35488 17368 35494
rect 17316 35430 17368 35436
rect 17224 35216 17276 35222
rect 17224 35158 17276 35164
rect 16948 34740 17000 34746
rect 16948 34682 17000 34688
rect 16946 33416 17002 33425
rect 16946 33351 17002 33360
rect 16960 33318 16988 33351
rect 16856 33312 16908 33318
rect 16856 33254 16908 33260
rect 16948 33312 17000 33318
rect 16948 33254 17000 33260
rect 16868 32978 16896 33254
rect 16856 32972 16908 32978
rect 16856 32914 16908 32920
rect 17236 32434 17264 35158
rect 17328 35154 17356 35430
rect 17316 35148 17368 35154
rect 17316 35090 17368 35096
rect 17408 34944 17460 34950
rect 17408 34886 17460 34892
rect 17420 34746 17448 34886
rect 17408 34740 17460 34746
rect 17408 34682 17460 34688
rect 18052 34604 18104 34610
rect 18052 34546 18104 34552
rect 17500 34536 17552 34542
rect 17500 34478 17552 34484
rect 17224 32428 17276 32434
rect 17224 32370 17276 32376
rect 17132 32360 17184 32366
rect 17132 32302 17184 32308
rect 17144 32026 17172 32302
rect 17408 32292 17460 32298
rect 17408 32234 17460 32240
rect 17132 32020 17184 32026
rect 17132 31962 17184 31968
rect 17420 31822 17448 32234
rect 17512 31890 17540 34478
rect 18064 34202 18092 34546
rect 18052 34196 18104 34202
rect 18052 34138 18104 34144
rect 17960 32836 18012 32842
rect 17960 32778 18012 32784
rect 17972 32570 18000 32778
rect 17960 32564 18012 32570
rect 17960 32506 18012 32512
rect 18052 32496 18104 32502
rect 18052 32438 18104 32444
rect 18064 32366 18092 32438
rect 17868 32360 17920 32366
rect 17868 32302 17920 32308
rect 18052 32360 18104 32366
rect 18052 32302 18104 32308
rect 17880 32230 17908 32302
rect 17868 32224 17920 32230
rect 17868 32166 17920 32172
rect 17500 31884 17552 31890
rect 17500 31826 17552 31832
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 17592 31748 17644 31754
rect 17592 31690 17644 31696
rect 17224 31136 17276 31142
rect 17224 31078 17276 31084
rect 17132 30728 17184 30734
rect 17132 30670 17184 30676
rect 17040 30660 17092 30666
rect 17040 30602 17092 30608
rect 16948 29504 17000 29510
rect 16948 29446 17000 29452
rect 16960 29238 16988 29446
rect 16948 29232 17000 29238
rect 16948 29174 17000 29180
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16868 28762 16896 29106
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 16960 28626 16988 29174
rect 16948 28620 17000 28626
rect 16948 28562 17000 28568
rect 16856 28416 16908 28422
rect 16856 28358 16908 28364
rect 16868 28218 16896 28358
rect 16856 28212 16908 28218
rect 16856 28154 16908 28160
rect 16868 27470 16896 28154
rect 16856 27464 16908 27470
rect 16856 27406 16908 27412
rect 17052 26432 17080 30602
rect 17144 29850 17172 30670
rect 17132 29844 17184 29850
rect 17132 29786 17184 29792
rect 17132 29300 17184 29306
rect 17132 29242 17184 29248
rect 17144 26994 17172 29242
rect 17236 29170 17264 31078
rect 17604 30870 17632 31690
rect 17880 31482 17908 32166
rect 17868 31476 17920 31482
rect 17868 31418 17920 31424
rect 17592 30864 17644 30870
rect 17592 30806 17644 30812
rect 17500 30728 17552 30734
rect 17500 30670 17552 30676
rect 17512 30394 17540 30670
rect 18052 30592 18104 30598
rect 18052 30534 18104 30540
rect 17500 30388 17552 30394
rect 17500 30330 17552 30336
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 17408 30252 17460 30258
rect 17408 30194 17460 30200
rect 17328 29646 17356 30194
rect 17316 29640 17368 29646
rect 17316 29582 17368 29588
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17328 29050 17356 29582
rect 17420 29510 17448 30194
rect 17776 30116 17828 30122
rect 17776 30058 17828 30064
rect 17408 29504 17460 29510
rect 17408 29446 17460 29452
rect 17420 29238 17448 29446
rect 17408 29232 17460 29238
rect 17408 29174 17460 29180
rect 17236 29022 17356 29050
rect 17132 26988 17184 26994
rect 17132 26930 17184 26936
rect 16868 26404 17080 26432
rect 16672 25492 16724 25498
rect 16672 25434 16724 25440
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16684 25362 16712 25434
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16396 24132 16448 24138
rect 16396 24074 16448 24080
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16408 23594 16436 24074
rect 16500 24070 16528 25094
rect 16592 25078 16804 25106
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16500 23730 16528 24006
rect 16488 23724 16540 23730
rect 16488 23666 16540 23672
rect 16396 23588 16448 23594
rect 16396 23530 16448 23536
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 16304 23520 16356 23526
rect 16304 23462 16356 23468
rect 15846 23420 16154 23440
rect 15846 23418 15852 23420
rect 15908 23418 15932 23420
rect 15988 23418 16012 23420
rect 16068 23418 16092 23420
rect 16148 23418 16154 23420
rect 15908 23366 15910 23418
rect 16090 23366 16092 23418
rect 15846 23364 15852 23366
rect 15908 23364 15932 23366
rect 15988 23364 16012 23366
rect 16068 23364 16092 23366
rect 16148 23364 16154 23366
rect 15846 23344 16154 23364
rect 16224 23118 16252 23462
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 16212 23112 16264 23118
rect 16212 23054 16264 23060
rect 16316 22778 16344 23462
rect 16408 22778 16436 23530
rect 15752 22772 15804 22778
rect 15752 22714 15804 22720
rect 16304 22772 16356 22778
rect 16304 22714 16356 22720
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15476 22160 15528 22166
rect 15476 22102 15528 22108
rect 15221 22052 15332 22080
rect 15568 22092 15620 22098
rect 15221 21876 15249 22052
rect 15568 22034 15620 22040
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15212 21848 15249 21876
rect 15108 21412 15160 21418
rect 15108 21354 15160 21360
rect 14752 20896 14964 20924
rect 14556 20324 14608 20330
rect 14556 20266 14608 20272
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14476 19990 14504 20198
rect 14464 19984 14516 19990
rect 14464 19926 14516 19932
rect 14476 17814 14504 19926
rect 14568 19854 14596 20266
rect 14752 19922 14780 20896
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14752 19446 14780 19654
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14476 16794 14504 17750
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14568 16590 14596 17274
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14108 15570 14136 16050
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13832 14006 13860 15030
rect 14476 15026 14504 16050
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 14476 13462 14504 14962
rect 14568 14618 14596 14962
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14660 14414 14688 18022
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14752 15706 14780 15982
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14740 15496 14792 15502
rect 14844 15484 14872 20742
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14936 18902 14964 20334
rect 14924 18896 14976 18902
rect 14924 18838 14976 18844
rect 15212 17338 15240 21848
rect 15304 21690 15332 21898
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15396 21570 15424 21898
rect 15304 21554 15424 21570
rect 15292 21548 15424 21554
rect 15344 21542 15424 21548
rect 15292 21490 15344 21496
rect 15292 20800 15344 20806
rect 15292 20742 15344 20748
rect 15304 20602 15332 20742
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15304 18358 15332 19654
rect 15396 18714 15424 21542
rect 15488 19961 15516 21966
rect 15580 21554 15608 22034
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15568 21412 15620 21418
rect 15568 21354 15620 21360
rect 15474 19952 15530 19961
rect 15474 19887 15530 19896
rect 15396 18686 15516 18714
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15396 18426 15424 18566
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15488 17746 15516 18686
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15120 16726 15148 16934
rect 15108 16720 15160 16726
rect 15108 16662 15160 16668
rect 15304 16590 15332 17206
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14792 15456 14872 15484
rect 14740 15438 14792 15444
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14844 15162 14872 15302
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14844 14414 14872 15098
rect 14924 14476 14976 14482
rect 15028 14464 15056 15506
rect 15120 15366 15148 15846
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 14976 14436 15056 14464
rect 14924 14418 14976 14424
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 14464 13456 14516 13462
rect 14464 13398 14516 13404
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13740 10606 13768 11154
rect 13832 11014 13860 13330
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14292 12850 14320 13194
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14292 12442 14320 12786
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14108 11218 14136 11698
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13740 10130 13768 10542
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13740 9654 13768 10066
rect 14200 9994 14228 12106
rect 14476 11830 14504 13398
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14384 10810 14412 11698
rect 14568 11082 14596 13942
rect 15120 13938 15148 15302
rect 15212 14414 15240 15506
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15488 14006 15516 17682
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 13728 9648 13780 9654
rect 13726 9616 13728 9625
rect 13780 9616 13782 9625
rect 13636 9580 13688 9586
rect 13726 9551 13782 9560
rect 13636 9522 13688 9528
rect 13740 9525 13768 9551
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13556 8974 13584 9114
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13556 8498 13584 8910
rect 13648 8566 13676 9522
rect 14094 8936 14150 8945
rect 14094 8871 14096 8880
rect 14148 8871 14150 8880
rect 14096 8842 14148 8848
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14016 7818 14044 8366
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14004 7812 14056 7818
rect 14004 7754 14056 7760
rect 14016 7410 14044 7754
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13556 6390 13584 7278
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 6798 13676 7142
rect 14004 6928 14056 6934
rect 14004 6870 14056 6876
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13648 6118 13676 6734
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13648 5778 13676 6054
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13372 4622 13400 5578
rect 13556 4842 13584 5646
rect 13648 5030 13676 5714
rect 13740 5710 13768 6802
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 14016 5302 14044 6870
rect 14108 5710 14136 7822
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13556 4814 13676 4842
rect 13648 4622 13676 4814
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13372 4214 13400 4558
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13648 3738 13676 4558
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13268 3460 13320 3466
rect 13268 3402 13320 3408
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 13004 2854 13032 2994
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 13096 1970 13124 2994
rect 13084 1964 13136 1970
rect 13084 1906 13136 1912
rect 13280 800 13308 3402
rect 13648 2990 13676 3674
rect 13740 3602 13768 4082
rect 13924 4010 13952 5170
rect 14108 4690 14136 5646
rect 14200 4826 14228 7346
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13740 2446 13768 3538
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 14016 2446 14044 2926
rect 14108 2650 14136 2994
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14200 2530 14228 3946
rect 14292 3194 14320 9998
rect 14568 7954 14596 9998
rect 14660 9926 14688 13194
rect 15028 12850 15056 13262
rect 15120 13258 15148 13874
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15488 13190 15516 13942
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15488 12646 15516 13126
rect 15580 12918 15608 21354
rect 15672 19378 15700 22578
rect 15764 20040 15792 22714
rect 16500 22658 16528 23666
rect 16592 23118 16620 24006
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16684 23322 16712 23666
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16670 23216 16726 23225
rect 16670 23151 16672 23160
rect 16724 23151 16726 23160
rect 16672 23122 16724 23128
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 16316 22630 16528 22658
rect 15846 22332 16154 22352
rect 15846 22330 15852 22332
rect 15908 22330 15932 22332
rect 15988 22330 16012 22332
rect 16068 22330 16092 22332
rect 16148 22330 16154 22332
rect 15908 22278 15910 22330
rect 16090 22278 16092 22330
rect 15846 22276 15852 22278
rect 15908 22276 15932 22278
rect 15988 22276 16012 22278
rect 16068 22276 16092 22278
rect 16148 22276 16154 22278
rect 15846 22256 16154 22276
rect 15844 22160 15896 22166
rect 15844 22102 15896 22108
rect 15856 21486 15884 22102
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15846 21244 16154 21264
rect 15846 21242 15852 21244
rect 15908 21242 15932 21244
rect 15988 21242 16012 21244
rect 16068 21242 16092 21244
rect 16148 21242 16154 21244
rect 15908 21190 15910 21242
rect 16090 21190 16092 21242
rect 15846 21188 15852 21190
rect 15908 21188 15932 21190
rect 15988 21188 16012 21190
rect 16068 21188 16092 21190
rect 16148 21188 16154 21190
rect 15846 21168 16154 21188
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 16224 20466 16252 20810
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 15846 20156 16154 20176
rect 15846 20154 15852 20156
rect 15908 20154 15932 20156
rect 15988 20154 16012 20156
rect 16068 20154 16092 20156
rect 16148 20154 16154 20156
rect 15908 20102 15910 20154
rect 16090 20102 16092 20154
rect 15846 20100 15852 20102
rect 15908 20100 15932 20102
rect 15988 20100 16012 20102
rect 16068 20100 16092 20102
rect 16148 20100 16154 20102
rect 15846 20080 16154 20100
rect 16224 20058 16252 20402
rect 16212 20052 16264 20058
rect 15764 20012 16068 20040
rect 15842 19952 15898 19961
rect 15752 19916 15804 19922
rect 16040 19922 16068 20012
rect 16212 19994 16264 20000
rect 15842 19887 15898 19896
rect 16028 19916 16080 19922
rect 15752 19858 15804 19864
rect 15764 19378 15792 19858
rect 15856 19854 15884 19887
rect 16028 19858 16080 19864
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15948 19514 15976 19790
rect 16316 19514 16344 22630
rect 16684 22556 16712 23122
rect 16408 22528 16712 22556
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15764 17882 15792 19314
rect 15846 19068 16154 19088
rect 15846 19066 15852 19068
rect 15908 19066 15932 19068
rect 15988 19066 16012 19068
rect 16068 19066 16092 19068
rect 16148 19066 16154 19068
rect 15908 19014 15910 19066
rect 16090 19014 16092 19066
rect 15846 19012 15852 19014
rect 15908 19012 15932 19014
rect 15988 19012 16012 19014
rect 16068 19012 16092 19014
rect 16148 19012 16154 19014
rect 15846 18992 16154 19012
rect 16212 18148 16264 18154
rect 16212 18090 16264 18096
rect 15846 17980 16154 18000
rect 15846 17978 15852 17980
rect 15908 17978 15932 17980
rect 15988 17978 16012 17980
rect 16068 17978 16092 17980
rect 16148 17978 16154 17980
rect 15908 17926 15910 17978
rect 16090 17926 16092 17978
rect 15846 17924 15852 17926
rect 15908 17924 15932 17926
rect 15988 17924 16012 17926
rect 16068 17924 16092 17926
rect 16148 17924 16154 17926
rect 15846 17904 16154 17924
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15846 16892 16154 16912
rect 15846 16890 15852 16892
rect 15908 16890 15932 16892
rect 15988 16890 16012 16892
rect 16068 16890 16092 16892
rect 16148 16890 16154 16892
rect 15908 16838 15910 16890
rect 16090 16838 16092 16890
rect 15846 16836 15852 16838
rect 15908 16836 15932 16838
rect 15988 16836 16012 16838
rect 16068 16836 16092 16838
rect 16148 16836 16154 16838
rect 15846 16816 16154 16836
rect 16224 15910 16252 18090
rect 16316 17678 16344 19450
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 15846 15804 16154 15824
rect 15846 15802 15852 15804
rect 15908 15802 15932 15804
rect 15988 15802 16012 15804
rect 16068 15802 16092 15804
rect 16148 15802 16154 15804
rect 15908 15750 15910 15802
rect 16090 15750 16092 15802
rect 15846 15748 15852 15750
rect 15908 15748 15932 15750
rect 15988 15748 16012 15750
rect 16068 15748 16092 15750
rect 16148 15748 16154 15750
rect 15846 15728 16154 15748
rect 16316 15706 16344 16390
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16316 14958 16344 15642
rect 16408 15473 16436 22528
rect 16580 22092 16632 22098
rect 16776 22094 16804 25078
rect 16580 22034 16632 22040
rect 16684 22066 16804 22094
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16500 21690 16528 21966
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16500 20874 16528 21422
rect 16488 20868 16540 20874
rect 16488 20810 16540 20816
rect 16592 20806 16620 22034
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16684 20618 16712 22066
rect 16868 22030 16896 26404
rect 17040 26308 17092 26314
rect 17040 26250 17092 26256
rect 16948 26240 17000 26246
rect 16948 26182 17000 26188
rect 16960 24834 16988 26182
rect 17052 26042 17080 26250
rect 17040 26036 17092 26042
rect 17040 25978 17092 25984
rect 17040 25492 17092 25498
rect 17040 25434 17092 25440
rect 17052 25158 17080 25434
rect 17236 25242 17264 29022
rect 17420 28082 17448 29174
rect 17788 29170 17816 30058
rect 17960 29504 18012 29510
rect 17960 29446 18012 29452
rect 17776 29164 17828 29170
rect 17776 29106 17828 29112
rect 17684 28620 17736 28626
rect 17684 28562 17736 28568
rect 17592 28144 17644 28150
rect 17592 28086 17644 28092
rect 17408 28076 17460 28082
rect 17408 28018 17460 28024
rect 17420 27538 17448 28018
rect 17408 27532 17460 27538
rect 17408 27474 17460 27480
rect 17500 27464 17552 27470
rect 17500 27406 17552 27412
rect 17408 27328 17460 27334
rect 17408 27270 17460 27276
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 17328 26450 17356 26930
rect 17316 26444 17368 26450
rect 17316 26386 17368 26392
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17328 25498 17356 26250
rect 17316 25492 17368 25498
rect 17316 25434 17368 25440
rect 17236 25214 17356 25242
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 17224 25152 17276 25158
rect 17224 25094 17276 25100
rect 17132 24948 17184 24954
rect 17132 24890 17184 24896
rect 16960 24806 17080 24834
rect 16948 24744 17000 24750
rect 16948 24686 17000 24692
rect 16960 24138 16988 24686
rect 16948 24132 17000 24138
rect 16948 24074 17000 24080
rect 16960 22409 16988 24074
rect 17052 23186 17080 24806
rect 17144 24070 17172 24890
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 16946 22400 17002 22409
rect 16946 22335 17002 22344
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16764 21548 16816 21554
rect 16764 21490 16816 21496
rect 16776 21146 16804 21490
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16592 20590 16712 20618
rect 16592 15502 16620 20590
rect 16776 20466 16804 20742
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 16684 18222 16712 19858
rect 16776 19514 16804 20402
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16776 18970 16804 19110
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16776 17746 16804 18158
rect 16764 17740 16816 17746
rect 16764 17682 16816 17688
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16580 15496 16632 15502
rect 16394 15464 16450 15473
rect 16580 15438 16632 15444
rect 16394 15399 16396 15408
rect 16448 15399 16450 15408
rect 16396 15370 16448 15376
rect 16408 15339 16436 15370
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 15846 14716 16154 14736
rect 15846 14714 15852 14716
rect 15908 14714 15932 14716
rect 15988 14714 16012 14716
rect 16068 14714 16092 14716
rect 16148 14714 16154 14716
rect 15908 14662 15910 14714
rect 16090 14662 16092 14714
rect 15846 14660 15852 14662
rect 15908 14660 15932 14662
rect 15988 14660 16012 14662
rect 16068 14660 16092 14662
rect 16148 14660 16154 14662
rect 15846 14640 16154 14660
rect 16120 14476 16172 14482
rect 16224 14464 16252 14758
rect 16316 14634 16344 14894
rect 16316 14606 16436 14634
rect 16684 14618 16712 17478
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16776 15910 16804 16526
rect 16868 16454 16896 21966
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16960 20806 16988 21286
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16960 19854 16988 20198
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 17052 18834 17080 22578
rect 17144 22386 17172 23666
rect 17236 23662 17264 25094
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 17144 22358 17264 22386
rect 17236 22098 17264 22358
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 17144 21146 17172 21898
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17236 20602 17264 21490
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16960 17338 16988 18702
rect 17052 17882 17080 18770
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 17052 17202 17080 17546
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16856 15632 16908 15638
rect 16960 15620 16988 16594
rect 17052 16590 17080 17138
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 16908 15592 16988 15620
rect 16856 15574 16908 15580
rect 16172 14436 16252 14464
rect 16120 14418 16172 14424
rect 16224 14278 16252 14436
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 15752 13796 15804 13802
rect 15752 13738 15804 13744
rect 15764 13462 15792 13738
rect 15846 13628 16154 13648
rect 15846 13626 15852 13628
rect 15908 13626 15932 13628
rect 15988 13626 16012 13628
rect 16068 13626 16092 13628
rect 16148 13626 16154 13628
rect 15908 13574 15910 13626
rect 16090 13574 16092 13626
rect 15846 13572 15852 13574
rect 15908 13572 15932 13574
rect 15988 13572 16012 13574
rect 16068 13572 16092 13574
rect 16148 13572 16154 13574
rect 15846 13552 16154 13572
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15764 12434 15792 13398
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16040 12986 16068 13330
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16224 12850 16252 14214
rect 16316 13530 16344 14418
rect 16408 14414 16436 14606
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16684 14464 16712 14554
rect 16592 14436 16712 14464
rect 16764 14476 16816 14482
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16592 13870 16620 14436
rect 16764 14418 16816 14424
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16672 13728 16724 13734
rect 16672 13670 16724 13676
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16684 13326 16712 13670
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 15846 12540 16154 12560
rect 15846 12538 15852 12540
rect 15908 12538 15932 12540
rect 15988 12538 16012 12540
rect 16068 12538 16092 12540
rect 16148 12538 16154 12540
rect 15908 12486 15910 12538
rect 16090 12486 16092 12538
rect 15846 12484 15852 12486
rect 15908 12484 15932 12486
rect 15988 12484 16012 12486
rect 16068 12484 16092 12486
rect 16148 12484 16154 12486
rect 15846 12464 16154 12484
rect 15672 12406 15792 12434
rect 15672 12306 15700 12406
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14844 10674 14872 11494
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15028 10674 15056 10950
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14844 8906 14872 9862
rect 15106 9616 15162 9625
rect 15304 9586 15332 11698
rect 15672 11218 15700 12038
rect 15846 11452 16154 11472
rect 15846 11450 15852 11452
rect 15908 11450 15932 11452
rect 15988 11450 16012 11452
rect 16068 11450 16092 11452
rect 16148 11450 16154 11452
rect 15908 11398 15910 11450
rect 16090 11398 16092 11450
rect 15846 11396 15852 11398
rect 15908 11396 15932 11398
rect 15988 11396 16012 11398
rect 16068 11396 16092 11398
rect 16148 11396 16154 11398
rect 15846 11376 16154 11396
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15672 9994 15700 10610
rect 15764 10606 15792 11086
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15846 10364 16154 10384
rect 15846 10362 15852 10364
rect 15908 10362 15932 10364
rect 15988 10362 16012 10364
rect 16068 10362 16092 10364
rect 16148 10362 16154 10364
rect 15908 10310 15910 10362
rect 16090 10310 16092 10362
rect 15846 10308 15852 10310
rect 15908 10308 15932 10310
rect 15988 10308 16012 10310
rect 16068 10308 16092 10310
rect 16148 10308 16154 10310
rect 15846 10288 16154 10308
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15764 10062 15792 10202
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15568 9988 15620 9994
rect 15568 9930 15620 9936
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15106 9551 15108 9560
rect 15160 9551 15162 9560
rect 15292 9580 15344 9586
rect 15108 9522 15160 9528
rect 15292 9522 15344 9528
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14108 2502 14228 2530
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 14108 800 14136 2502
rect 14384 2378 14412 7822
rect 14568 7426 14596 7890
rect 14660 7546 14688 8434
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14476 7410 14596 7426
rect 14844 7410 14872 7822
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 14464 7404 14596 7410
rect 14516 7398 14596 7404
rect 14832 7404 14884 7410
rect 14464 7346 14516 7352
rect 14832 7346 14884 7352
rect 15028 6866 15056 7414
rect 15120 7274 15148 9522
rect 15304 8838 15332 9522
rect 15580 8974 15608 9930
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15212 7546 15240 7822
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 15212 6866 15240 7346
rect 15304 7342 15332 8230
rect 15476 7812 15528 7818
rect 15476 7754 15528 7760
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 4690 14596 6598
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14568 3058 14596 4626
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 14844 800 14872 6666
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 14936 5370 14964 6258
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15028 5166 15056 6802
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15304 6118 15332 6734
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15016 4548 15068 4554
rect 15016 4490 15068 4496
rect 15028 2650 15056 4490
rect 15120 3210 15148 4966
rect 15396 4826 15424 7346
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15120 3182 15240 3210
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15016 2644 15068 2650
rect 15016 2586 15068 2592
rect 15120 2446 15148 2994
rect 15212 2990 15240 3182
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15212 2854 15240 2926
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15304 2582 15332 4014
rect 15396 3058 15424 4082
rect 15488 3738 15516 7754
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15580 5234 15608 6802
rect 15672 6186 15700 9522
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15764 8362 15792 9454
rect 15846 9276 16154 9296
rect 15846 9274 15852 9276
rect 15908 9274 15932 9276
rect 15988 9274 16012 9276
rect 16068 9274 16092 9276
rect 16148 9274 16154 9276
rect 15908 9222 15910 9274
rect 16090 9222 16092 9274
rect 15846 9220 15852 9222
rect 15908 9220 15932 9222
rect 15988 9220 16012 9222
rect 16068 9220 16092 9222
rect 16148 9220 16154 9222
rect 15846 9200 16154 9220
rect 15752 8356 15804 8362
rect 15752 8298 15804 8304
rect 15846 8188 16154 8208
rect 15846 8186 15852 8188
rect 15908 8186 15932 8188
rect 15988 8186 16012 8188
rect 16068 8186 16092 8188
rect 16148 8186 16154 8188
rect 15908 8134 15910 8186
rect 16090 8134 16092 8186
rect 15846 8132 15852 8134
rect 15908 8132 15932 8134
rect 15988 8132 16012 8134
rect 16068 8132 16092 8134
rect 16148 8132 16154 8134
rect 15846 8112 16154 8132
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15672 5386 15700 6122
rect 15764 5642 15792 7142
rect 15846 7100 16154 7120
rect 15846 7098 15852 7100
rect 15908 7098 15932 7100
rect 15988 7098 16012 7100
rect 16068 7098 16092 7100
rect 16148 7098 16154 7100
rect 15908 7046 15910 7098
rect 16090 7046 16092 7098
rect 15846 7044 15852 7046
rect 15908 7044 15932 7046
rect 15988 7044 16012 7046
rect 16068 7044 16092 7046
rect 16148 7044 16154 7046
rect 15846 7024 16154 7044
rect 16224 6769 16252 12786
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16500 12646 16528 12718
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16316 11218 16344 12174
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16408 10130 16436 12174
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 8945 16344 9318
rect 16408 9110 16436 10066
rect 16500 9654 16528 11086
rect 16592 10810 16620 13194
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16684 12442 16712 12718
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16776 11150 16804 14418
rect 16868 13938 16896 15574
rect 17040 15496 17092 15502
rect 16960 15456 17040 15484
rect 16960 15366 16988 15456
rect 17144 15484 17172 19654
rect 17236 19378 17264 19994
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17236 17270 17264 19314
rect 17328 18834 17356 25214
rect 17420 24206 17448 27270
rect 17512 26586 17540 27406
rect 17500 26580 17552 26586
rect 17500 26522 17552 26528
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17512 25770 17540 26318
rect 17500 25764 17552 25770
rect 17500 25706 17552 25712
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 17408 23656 17460 23662
rect 17408 23598 17460 23604
rect 17420 22778 17448 23598
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17408 22568 17460 22574
rect 17512 22556 17540 24822
rect 17460 22528 17540 22556
rect 17408 22510 17460 22516
rect 17420 21010 17448 22510
rect 17604 22080 17632 28086
rect 17696 28014 17724 28562
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 17684 27532 17736 27538
rect 17684 27474 17736 27480
rect 17696 27441 17724 27474
rect 17682 27432 17738 27441
rect 17682 27367 17738 27376
rect 17684 26784 17736 26790
rect 17684 26726 17736 26732
rect 17512 22052 17632 22080
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 17408 20868 17460 20874
rect 17408 20810 17460 20816
rect 17420 20398 17448 20810
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17420 18222 17448 20334
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17236 16794 17264 17070
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17236 15706 17264 16050
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17224 15496 17276 15502
rect 17144 15456 17224 15484
rect 17040 15438 17092 15444
rect 17224 15438 17276 15444
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 17130 15328 17186 15337
rect 16960 15162 16988 15302
rect 17130 15263 17186 15272
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 17040 15088 17092 15094
rect 17038 15056 17040 15065
rect 17092 15056 17094 15065
rect 17144 15026 17172 15263
rect 17222 15192 17278 15201
rect 17222 15127 17278 15136
rect 17236 15026 17264 15127
rect 17038 14991 17094 15000
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17328 14906 17356 15846
rect 17408 15496 17460 15502
rect 17406 15464 17408 15473
rect 17460 15464 17462 15473
rect 17406 15399 17462 15408
rect 17406 15328 17462 15337
rect 17406 15263 17462 15272
rect 17052 14878 17356 14906
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16868 13190 16896 13874
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16960 12442 16988 14758
rect 17052 13938 17080 14878
rect 17316 14816 17368 14822
rect 17236 14764 17316 14770
rect 17236 14758 17368 14764
rect 17236 14742 17356 14758
rect 17236 14482 17264 14742
rect 17420 14634 17448 15263
rect 17512 14770 17540 22052
rect 17590 21992 17646 22001
rect 17590 21927 17646 21936
rect 17604 21078 17632 21927
rect 17592 21072 17644 21078
rect 17592 21014 17644 21020
rect 17604 19922 17632 21014
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 17696 19854 17724 26726
rect 17788 23730 17816 29106
rect 17868 29028 17920 29034
rect 17868 28970 17920 28976
rect 17880 24954 17908 28970
rect 17868 24948 17920 24954
rect 17868 24890 17920 24896
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17880 24410 17908 24686
rect 17868 24404 17920 24410
rect 17868 24346 17920 24352
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 17788 21622 17816 23666
rect 17880 22166 17908 23666
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17880 21690 17908 21966
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17776 21616 17828 21622
rect 17776 21558 17828 21564
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 17880 21350 17908 21490
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17592 19712 17644 19718
rect 17788 19666 17816 20402
rect 17880 20058 17908 21082
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17592 19654 17644 19660
rect 17604 19514 17632 19654
rect 17696 19638 17816 19666
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17604 18154 17632 19314
rect 17696 18290 17724 19638
rect 17972 19530 18000 29446
rect 18064 29170 18092 30534
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 18156 28626 18184 37062
rect 18800 36922 18828 37198
rect 18788 36916 18840 36922
rect 18788 36858 18840 36864
rect 18512 36100 18564 36106
rect 18512 36042 18564 36048
rect 18236 36032 18288 36038
rect 18236 35974 18288 35980
rect 18248 35698 18276 35974
rect 18236 35692 18288 35698
rect 18236 35634 18288 35640
rect 18420 35692 18472 35698
rect 18420 35634 18472 35640
rect 18328 34944 18380 34950
rect 18328 34886 18380 34892
rect 18236 33924 18288 33930
rect 18236 33866 18288 33872
rect 18248 33522 18276 33866
rect 18236 33516 18288 33522
rect 18236 33458 18288 33464
rect 18248 29510 18276 33458
rect 18340 30326 18368 34886
rect 18432 33658 18460 35634
rect 18524 35018 18552 36042
rect 19168 35306 19196 38694
rect 19352 38554 19380 39986
rect 19432 39432 19484 39438
rect 19432 39374 19484 39380
rect 19340 38548 19392 38554
rect 19340 38490 19392 38496
rect 19444 38282 19472 39374
rect 19616 39364 19668 39370
rect 19616 39306 19668 39312
rect 19628 39098 19656 39306
rect 19616 39092 19668 39098
rect 19616 39034 19668 39040
rect 20076 38956 20128 38962
rect 20076 38898 20128 38904
rect 20088 38554 20116 38898
rect 20076 38548 20128 38554
rect 20076 38490 20128 38496
rect 19432 38276 19484 38282
rect 19432 38218 19484 38224
rect 19444 37942 19472 38218
rect 19432 37936 19484 37942
rect 19432 37878 19484 37884
rect 19248 37120 19300 37126
rect 19248 37062 19300 37068
rect 19260 36786 19288 37062
rect 19340 36848 19392 36854
rect 19340 36790 19392 36796
rect 19248 36780 19300 36786
rect 19248 36722 19300 36728
rect 19352 36242 19380 36790
rect 19340 36236 19392 36242
rect 19340 36178 19392 36184
rect 19444 36106 19472 37878
rect 20180 36938 20208 42570
rect 20811 42460 21119 42480
rect 20811 42458 20817 42460
rect 20873 42458 20897 42460
rect 20953 42458 20977 42460
rect 21033 42458 21057 42460
rect 21113 42458 21119 42460
rect 20873 42406 20875 42458
rect 21055 42406 21057 42458
rect 20811 42404 20817 42406
rect 20873 42404 20897 42406
rect 20953 42404 20977 42406
rect 21033 42404 21057 42406
rect 21113 42404 21119 42406
rect 20811 42384 21119 42404
rect 21916 42220 21968 42226
rect 21916 42162 21968 42168
rect 20811 41372 21119 41392
rect 20811 41370 20817 41372
rect 20873 41370 20897 41372
rect 20953 41370 20977 41372
rect 21033 41370 21057 41372
rect 21113 41370 21119 41372
rect 20873 41318 20875 41370
rect 21055 41318 21057 41370
rect 20811 41316 20817 41318
rect 20873 41316 20897 41318
rect 20953 41316 20977 41318
rect 21033 41316 21057 41318
rect 21113 41316 21119 41318
rect 20811 41296 21119 41316
rect 20811 40284 21119 40304
rect 20811 40282 20817 40284
rect 20873 40282 20897 40284
rect 20953 40282 20977 40284
rect 21033 40282 21057 40284
rect 21113 40282 21119 40284
rect 20873 40230 20875 40282
rect 21055 40230 21057 40282
rect 20811 40228 20817 40230
rect 20873 40228 20897 40230
rect 20953 40228 20977 40230
rect 21033 40228 21057 40230
rect 21113 40228 21119 40230
rect 20811 40208 21119 40228
rect 21824 39976 21876 39982
rect 21824 39918 21876 39924
rect 20260 39296 20312 39302
rect 20260 39238 20312 39244
rect 20272 38350 20300 39238
rect 20811 39196 21119 39216
rect 20811 39194 20817 39196
rect 20873 39194 20897 39196
rect 20953 39194 20977 39196
rect 21033 39194 21057 39196
rect 21113 39194 21119 39196
rect 20873 39142 20875 39194
rect 21055 39142 21057 39194
rect 20811 39140 20817 39142
rect 20873 39140 20897 39142
rect 20953 39140 20977 39142
rect 21033 39140 21057 39142
rect 21113 39140 21119 39142
rect 20811 39120 21119 39140
rect 21364 38752 21416 38758
rect 21364 38694 21416 38700
rect 20260 38344 20312 38350
rect 20260 38286 20312 38292
rect 20811 38108 21119 38128
rect 20811 38106 20817 38108
rect 20873 38106 20897 38108
rect 20953 38106 20977 38108
rect 21033 38106 21057 38108
rect 21113 38106 21119 38108
rect 20873 38054 20875 38106
rect 21055 38054 21057 38106
rect 20811 38052 20817 38054
rect 20873 38052 20897 38054
rect 20953 38052 20977 38054
rect 21033 38052 21057 38054
rect 21113 38052 21119 38054
rect 20811 38032 21119 38052
rect 20352 37460 20404 37466
rect 20352 37402 20404 37408
rect 20180 36910 20300 36938
rect 20168 36848 20220 36854
rect 20168 36790 20220 36796
rect 19524 36780 19576 36786
rect 19524 36722 19576 36728
rect 19432 36100 19484 36106
rect 19432 36042 19484 36048
rect 19432 35828 19484 35834
rect 19432 35770 19484 35776
rect 19168 35278 19288 35306
rect 18512 35012 18564 35018
rect 18512 34954 18564 34960
rect 18420 33652 18472 33658
rect 18420 33594 18472 33600
rect 18420 32768 18472 32774
rect 18420 32710 18472 32716
rect 18432 32570 18460 32710
rect 18420 32564 18472 32570
rect 18420 32506 18472 32512
rect 18524 32450 18552 34954
rect 18604 34944 18656 34950
rect 18604 34886 18656 34892
rect 18616 34678 18644 34886
rect 19156 34740 19208 34746
rect 19156 34682 19208 34688
rect 18604 34672 18656 34678
rect 18604 34614 18656 34620
rect 18604 33992 18656 33998
rect 18604 33934 18656 33940
rect 18616 33658 18644 33934
rect 19064 33856 19116 33862
rect 19064 33798 19116 33804
rect 18604 33652 18656 33658
rect 18604 33594 18656 33600
rect 19076 33522 19104 33798
rect 19168 33658 19196 34682
rect 19156 33652 19208 33658
rect 19156 33594 19208 33600
rect 19064 33516 19116 33522
rect 19064 33458 19116 33464
rect 18880 32904 18932 32910
rect 18880 32846 18932 32852
rect 18788 32496 18840 32502
rect 18524 32422 18644 32450
rect 18788 32438 18840 32444
rect 18512 31816 18564 31822
rect 18512 31758 18564 31764
rect 18524 31414 18552 31758
rect 18512 31408 18564 31414
rect 18512 31350 18564 31356
rect 18420 31136 18472 31142
rect 18420 31078 18472 31084
rect 18432 30802 18460 31078
rect 18524 30938 18552 31350
rect 18512 30932 18564 30938
rect 18512 30874 18564 30880
rect 18420 30796 18472 30802
rect 18420 30738 18472 30744
rect 18328 30320 18380 30326
rect 18328 30262 18380 30268
rect 18328 30184 18380 30190
rect 18328 30126 18380 30132
rect 18340 29782 18368 30126
rect 18420 29844 18472 29850
rect 18420 29786 18472 29792
rect 18328 29776 18380 29782
rect 18328 29718 18380 29724
rect 18340 29578 18368 29718
rect 18328 29572 18380 29578
rect 18328 29514 18380 29520
rect 18236 29504 18288 29510
rect 18236 29446 18288 29452
rect 18340 29322 18368 29514
rect 18248 29294 18368 29322
rect 18052 28620 18104 28626
rect 18052 28562 18104 28568
rect 18144 28620 18196 28626
rect 18144 28562 18196 28568
rect 18064 28506 18092 28562
rect 18248 28506 18276 29294
rect 18328 29164 18380 29170
rect 18328 29106 18380 29112
rect 18340 28626 18368 29106
rect 18328 28620 18380 28626
rect 18328 28562 18380 28568
rect 18064 28478 18276 28506
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 18064 26858 18092 28358
rect 18340 28234 18368 28562
rect 18432 28558 18460 29786
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 18512 28416 18564 28422
rect 18512 28358 18564 28364
rect 18248 28206 18368 28234
rect 18144 27464 18196 27470
rect 18144 27406 18196 27412
rect 18052 26852 18104 26858
rect 18052 26794 18104 26800
rect 18156 26586 18184 27406
rect 18248 26994 18276 28206
rect 18328 28076 18380 28082
rect 18328 28018 18380 28024
rect 18236 26988 18288 26994
rect 18236 26930 18288 26936
rect 18236 26852 18288 26858
rect 18236 26794 18288 26800
rect 18144 26580 18196 26586
rect 18144 26522 18196 26528
rect 18052 26444 18104 26450
rect 18052 26386 18104 26392
rect 18064 25838 18092 26386
rect 18248 26246 18276 26794
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 18052 25832 18104 25838
rect 18052 25774 18104 25780
rect 18064 25362 18092 25774
rect 18052 25356 18104 25362
rect 18052 25298 18104 25304
rect 18050 25256 18106 25265
rect 18050 25191 18052 25200
rect 18104 25191 18106 25200
rect 18052 25162 18104 25168
rect 18144 25152 18196 25158
rect 18248 25106 18276 26182
rect 18340 26042 18368 28018
rect 18420 27872 18472 27878
rect 18420 27814 18472 27820
rect 18432 26994 18460 27814
rect 18524 27470 18552 28358
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18616 27418 18644 32422
rect 18696 31952 18748 31958
rect 18696 31894 18748 31900
rect 18708 31346 18736 31894
rect 18696 31340 18748 31346
rect 18696 31282 18748 31288
rect 18800 30920 18828 32438
rect 18892 32434 18920 32846
rect 18880 32428 18932 32434
rect 18880 32370 18932 32376
rect 18892 31346 18920 32370
rect 19064 32224 19116 32230
rect 19064 32166 19116 32172
rect 18972 31748 19024 31754
rect 18972 31690 19024 31696
rect 18880 31340 18932 31346
rect 18880 31282 18932 31288
rect 18800 30892 18920 30920
rect 18788 30796 18840 30802
rect 18788 30738 18840 30744
rect 18696 30252 18748 30258
rect 18696 30194 18748 30200
rect 18708 28082 18736 30194
rect 18696 28076 18748 28082
rect 18696 28018 18748 28024
rect 18708 27606 18736 28018
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 18616 27390 18736 27418
rect 18800 27402 18828 30738
rect 18892 30122 18920 30892
rect 18984 30258 19012 31690
rect 19076 31482 19104 32166
rect 19168 32026 19196 33594
rect 19156 32020 19208 32026
rect 19156 31962 19208 31968
rect 19064 31476 19116 31482
rect 19064 31418 19116 31424
rect 19076 30734 19104 31418
rect 19168 31346 19196 31962
rect 19156 31340 19208 31346
rect 19156 31282 19208 31288
rect 19156 31204 19208 31210
rect 19156 31146 19208 31152
rect 19064 30728 19116 30734
rect 19064 30670 19116 30676
rect 19168 30666 19196 31146
rect 19156 30660 19208 30666
rect 19156 30602 19208 30608
rect 18972 30252 19024 30258
rect 18972 30194 19024 30200
rect 18880 30116 18932 30122
rect 18880 30058 18932 30064
rect 18880 28552 18932 28558
rect 18880 28494 18932 28500
rect 18512 27328 18564 27334
rect 18512 27270 18564 27276
rect 18604 27328 18656 27334
rect 18604 27270 18656 27276
rect 18420 26988 18472 26994
rect 18420 26930 18472 26936
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18196 25100 18276 25106
rect 18144 25094 18276 25100
rect 18156 25078 18276 25094
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 18064 22098 18092 24754
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18052 22092 18104 22098
rect 18052 22034 18104 22040
rect 18156 21690 18184 23462
rect 18144 21684 18196 21690
rect 18144 21626 18196 21632
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 17880 19502 18000 19530
rect 17880 18850 17908 19502
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17972 18970 18000 19314
rect 18156 19310 18184 20878
rect 18248 19446 18276 25078
rect 18328 24268 18380 24274
rect 18380 24228 18460 24256
rect 18328 24210 18380 24216
rect 18328 24064 18380 24070
rect 18328 24006 18380 24012
rect 18340 23866 18368 24006
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18340 22234 18368 22578
rect 18432 22574 18460 24228
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18328 22228 18380 22234
rect 18328 22170 18380 22176
rect 18432 22094 18460 22510
rect 18340 22066 18460 22094
rect 18340 21010 18368 22066
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 18432 21078 18460 21422
rect 18420 21072 18472 21078
rect 18420 21014 18472 21020
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18524 20924 18552 27270
rect 18616 26994 18644 27270
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 18708 26432 18736 27390
rect 18788 27396 18840 27402
rect 18788 27338 18840 27344
rect 18788 26988 18840 26994
rect 18788 26930 18840 26936
rect 18800 26450 18828 26930
rect 18616 26404 18736 26432
rect 18788 26444 18840 26450
rect 18616 24342 18644 26404
rect 18788 26386 18840 26392
rect 18696 26308 18748 26314
rect 18696 26250 18748 26256
rect 18708 25838 18736 26250
rect 18788 25968 18840 25974
rect 18788 25910 18840 25916
rect 18696 25832 18748 25838
rect 18696 25774 18748 25780
rect 18604 24336 18656 24342
rect 18656 24284 18736 24290
rect 18604 24278 18736 24284
rect 18616 24262 18736 24278
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18616 22778 18644 23598
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18616 21486 18644 22034
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18432 20896 18552 20924
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 18052 18896 18104 18902
rect 17880 18822 18000 18850
rect 18052 18838 18104 18844
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17592 18148 17644 18154
rect 17592 18090 17644 18096
rect 17512 14742 17632 14770
rect 17328 14606 17448 14634
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 17328 14414 17356 14606
rect 17604 14498 17632 14742
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17512 14470 17632 14498
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17052 13258 17080 13874
rect 17224 13728 17276 13734
rect 17144 13676 17224 13682
rect 17144 13670 17276 13676
rect 17144 13654 17264 13670
rect 17144 13326 17172 13654
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17052 12714 17080 13194
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17328 12850 17356 13126
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17420 11898 17448 14418
rect 17512 13530 17540 14470
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17604 14074 17632 14350
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17512 13326 17540 13466
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16580 10804 16632 10810
rect 16632 10764 16712 10792
rect 16580 10746 16632 10752
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16592 10130 16620 10610
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16684 10062 16712 10764
rect 16868 10674 16896 11562
rect 16960 11286 16988 11698
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16960 10674 16988 11018
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 17052 10606 17080 11154
rect 17328 11150 17356 11494
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 17144 10130 17172 11086
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 17236 9722 17264 10610
rect 17696 10266 17724 18226
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17880 17270 17908 17614
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17788 13734 17816 17138
rect 17866 15056 17922 15065
rect 17972 15042 18000 18822
rect 18064 17814 18092 18838
rect 18156 18834 18184 19246
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18144 18692 18196 18698
rect 18144 18634 18196 18640
rect 18052 17808 18104 17814
rect 18052 17750 18104 17756
rect 18156 17678 18184 18634
rect 18248 17814 18276 19382
rect 18432 19334 18460 20896
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18524 20602 18552 20742
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18340 19306 18460 19334
rect 18236 17808 18288 17814
rect 18236 17750 18288 17756
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18156 16590 18184 17614
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18156 16250 18184 16526
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18248 15434 18276 16050
rect 18236 15428 18288 15434
rect 17922 15014 18000 15042
rect 18156 15388 18236 15416
rect 17866 14991 17868 15000
rect 17920 14991 17922 15000
rect 17868 14962 17920 14968
rect 17880 14931 17908 14962
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17972 14414 18000 14894
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17880 11354 17908 13806
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18064 12102 18092 12582
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 18064 11898 18092 12038
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18064 10810 18092 11086
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17696 10062 17724 10202
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17420 9722 17448 9930
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 16302 8936 16358 8945
rect 16302 8871 16358 8880
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 7818 16528 8774
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 16210 6760 16266 6769
rect 16210 6695 16266 6704
rect 16500 6390 16528 7754
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16868 6866 16896 7142
rect 16960 6866 16988 7346
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 15846 6012 16154 6032
rect 15846 6010 15852 6012
rect 15908 6010 15932 6012
rect 15988 6010 16012 6012
rect 16068 6010 16092 6012
rect 16148 6010 16154 6012
rect 15908 5958 15910 6010
rect 16090 5958 16092 6010
rect 15846 5956 15852 5958
rect 15908 5956 15932 5958
rect 15988 5956 16012 5958
rect 16068 5956 16092 5958
rect 16148 5956 16154 5958
rect 15846 5936 16154 5956
rect 16500 5794 16528 6326
rect 16408 5766 16528 5794
rect 16408 5710 16436 5766
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15672 5358 15792 5386
rect 15764 5302 15792 5358
rect 15752 5296 15804 5302
rect 15752 5238 15804 5244
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 15846 4924 16154 4944
rect 15846 4922 15852 4924
rect 15908 4922 15932 4924
rect 15988 4922 16012 4924
rect 16068 4922 16092 4924
rect 16148 4922 16154 4924
rect 15908 4870 15910 4922
rect 16090 4870 16092 4922
rect 15846 4868 15852 4870
rect 15908 4868 15932 4870
rect 15988 4868 16012 4870
rect 16068 4868 16092 4870
rect 16148 4868 16154 4870
rect 15846 4848 16154 4868
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15580 4282 15608 4422
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15764 4146 15792 4422
rect 15948 4146 15976 4626
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 16040 4146 16068 4490
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 16028 4140 16080 4146
rect 16080 4100 16252 4128
rect 16028 4082 16080 4088
rect 15846 3836 16154 3856
rect 15846 3834 15852 3836
rect 15908 3834 15932 3836
rect 15988 3834 16012 3836
rect 16068 3834 16092 3836
rect 16148 3834 16154 3836
rect 15908 3782 15910 3834
rect 16090 3782 16092 3834
rect 15846 3780 15852 3782
rect 15908 3780 15932 3782
rect 15988 3780 16012 3782
rect 16068 3780 16092 3782
rect 16148 3780 16154 3782
rect 15846 3760 16154 3780
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 16224 3670 16252 4100
rect 16316 4010 16344 5170
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16408 4078 16436 4558
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15396 2650 15424 2994
rect 15846 2748 16154 2768
rect 15846 2746 15852 2748
rect 15908 2746 15932 2748
rect 15988 2746 16012 2748
rect 16068 2746 16092 2748
rect 16148 2746 16154 2748
rect 15908 2694 15910 2746
rect 16090 2694 16092 2746
rect 15846 2692 15852 2694
rect 15908 2692 15932 2694
rect 15988 2692 16012 2694
rect 16068 2692 16092 2694
rect 16148 2692 16154 2694
rect 15846 2672 16154 2692
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15304 2446 15332 2518
rect 16224 2514 16252 3606
rect 16500 3534 16528 4422
rect 16592 4282 16620 5102
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16684 3738 16712 6734
rect 16960 5914 16988 6802
rect 17236 6798 17264 9522
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17880 9178 17908 9454
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17774 9072 17830 9081
rect 17774 9007 17830 9016
rect 17788 8974 17816 9007
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17788 8498 17816 8910
rect 17880 8498 17908 9114
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17328 7478 17356 8434
rect 17972 7546 18000 10610
rect 18156 10062 18184 15388
rect 18236 15370 18288 15376
rect 18340 15337 18368 19306
rect 18616 17202 18644 19722
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18326 15328 18382 15337
rect 18382 15286 18460 15314
rect 18326 15263 18382 15272
rect 18328 14408 18380 14414
rect 18328 14350 18380 14356
rect 18340 14278 18368 14350
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18340 13938 18368 14214
rect 18432 14074 18460 15286
rect 18524 15026 18552 17070
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18616 15502 18644 16390
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18616 15026 18644 15438
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18524 13938 18552 14962
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18616 14618 18644 14758
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18602 13968 18658 13977
rect 18328 13932 18380 13938
rect 18512 13932 18564 13938
rect 18328 13874 18380 13880
rect 18432 13892 18512 13920
rect 18432 13802 18460 13892
rect 18602 13903 18658 13912
rect 18512 13874 18564 13880
rect 18616 13802 18644 13903
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18248 12918 18276 13262
rect 18432 12986 18460 13738
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18524 13530 18552 13670
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18328 12368 18380 12374
rect 18328 12310 18380 12316
rect 18340 11762 18368 12310
rect 18616 12238 18644 13126
rect 18708 12986 18736 24262
rect 18800 19514 18828 25910
rect 18892 25838 18920 28494
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 18984 27674 19012 28018
rect 18972 27668 19024 27674
rect 18972 27610 19024 27616
rect 18972 27532 19024 27538
rect 18972 27474 19024 27480
rect 18984 27062 19012 27474
rect 19064 27464 19116 27470
rect 19062 27432 19064 27441
rect 19116 27432 19118 27441
rect 19062 27367 19118 27376
rect 19156 27396 19208 27402
rect 19156 27338 19208 27344
rect 19064 27328 19116 27334
rect 19168 27305 19196 27338
rect 19064 27270 19116 27276
rect 19154 27296 19210 27305
rect 18972 27056 19024 27062
rect 18972 26998 19024 27004
rect 19076 26858 19104 27270
rect 19154 27231 19210 27240
rect 19156 26920 19208 26926
rect 19156 26862 19208 26868
rect 19064 26852 19116 26858
rect 19064 26794 19116 26800
rect 18880 25832 18932 25838
rect 18880 25774 18932 25780
rect 18892 24886 18920 25774
rect 18880 24880 18932 24886
rect 18880 24822 18932 24828
rect 19168 24750 19196 26862
rect 19156 24744 19208 24750
rect 19156 24686 19208 24692
rect 18880 24608 18932 24614
rect 18880 24550 18932 24556
rect 18972 24608 19024 24614
rect 18972 24550 19024 24556
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18800 18766 18828 19450
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18892 15094 18920 24550
rect 18984 24410 19012 24550
rect 18972 24404 19024 24410
rect 18972 24346 19024 24352
rect 19168 23662 19196 24686
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 19168 23118 19196 23598
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 19156 23112 19208 23118
rect 19156 23054 19208 23060
rect 18984 21026 19012 23054
rect 19156 22976 19208 22982
rect 19156 22918 19208 22924
rect 19168 22642 19196 22918
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 19064 22432 19116 22438
rect 19064 22374 19116 22380
rect 19076 21554 19104 22374
rect 19156 22160 19208 22166
rect 19156 22102 19208 22108
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 19168 21418 19196 22102
rect 19260 22098 19288 35278
rect 19340 34400 19392 34406
rect 19340 34342 19392 34348
rect 19352 33590 19380 34342
rect 19444 33998 19472 35770
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 19340 33584 19392 33590
rect 19340 33526 19392 33532
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 19444 31822 19472 33458
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19536 31482 19564 36722
rect 19800 36236 19852 36242
rect 19800 36178 19852 36184
rect 19616 36032 19668 36038
rect 19616 35974 19668 35980
rect 19628 34610 19656 35974
rect 19616 34604 19668 34610
rect 19616 34546 19668 34552
rect 19812 33998 19840 36178
rect 19984 34944 20036 34950
rect 19984 34886 20036 34892
rect 19892 34400 19944 34406
rect 19892 34342 19944 34348
rect 19616 33992 19668 33998
rect 19616 33934 19668 33940
rect 19800 33992 19852 33998
rect 19800 33934 19852 33940
rect 19628 33114 19656 33934
rect 19708 33584 19760 33590
rect 19708 33526 19760 33532
rect 19616 33108 19668 33114
rect 19616 33050 19668 33056
rect 19616 32224 19668 32230
rect 19616 32166 19668 32172
rect 19524 31476 19576 31482
rect 19524 31418 19576 31424
rect 19628 31278 19656 32166
rect 19616 31272 19668 31278
rect 19616 31214 19668 31220
rect 19616 31136 19668 31142
rect 19616 31078 19668 31084
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19352 28082 19380 29582
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 19432 27872 19484 27878
rect 19432 27814 19484 27820
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 19352 26518 19380 26930
rect 19444 26790 19472 27814
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19340 26512 19392 26518
rect 19340 26454 19392 26460
rect 19352 26042 19380 26454
rect 19340 26036 19392 26042
rect 19340 25978 19392 25984
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19352 24818 19380 25842
rect 19444 25702 19472 26726
rect 19524 26036 19576 26042
rect 19524 25978 19576 25984
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19352 23798 19380 24754
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 19340 22704 19392 22710
rect 19444 22692 19472 25638
rect 19536 25294 19564 25978
rect 19628 25498 19656 31078
rect 19720 28422 19748 33526
rect 19904 33522 19932 34342
rect 19996 34066 20024 34886
rect 20076 34536 20128 34542
rect 20076 34478 20128 34484
rect 20088 34202 20116 34478
rect 20076 34196 20128 34202
rect 20076 34138 20128 34144
rect 19984 34060 20036 34066
rect 19984 34002 20036 34008
rect 20088 33946 20116 34138
rect 20180 34066 20208 36790
rect 20272 36242 20300 36910
rect 20260 36236 20312 36242
rect 20260 36178 20312 36184
rect 20260 36032 20312 36038
rect 20260 35974 20312 35980
rect 20272 35834 20300 35974
rect 20260 35828 20312 35834
rect 20260 35770 20312 35776
rect 20272 35698 20300 35770
rect 20260 35692 20312 35698
rect 20260 35634 20312 35640
rect 20364 34746 20392 37402
rect 20811 37020 21119 37040
rect 20811 37018 20817 37020
rect 20873 37018 20897 37020
rect 20953 37018 20977 37020
rect 21033 37018 21057 37020
rect 21113 37018 21119 37020
rect 20873 36966 20875 37018
rect 21055 36966 21057 37018
rect 20811 36964 20817 36966
rect 20873 36964 20897 36966
rect 20953 36964 20977 36966
rect 21033 36964 21057 36966
rect 21113 36964 21119 36966
rect 20811 36944 21119 36964
rect 20628 36576 20680 36582
rect 20628 36518 20680 36524
rect 21272 36576 21324 36582
rect 21272 36518 21324 36524
rect 20640 36174 20668 36518
rect 20628 36168 20680 36174
rect 20628 36110 20680 36116
rect 21180 36168 21232 36174
rect 21180 36110 21232 36116
rect 20640 35698 20668 36110
rect 20811 35932 21119 35952
rect 20811 35930 20817 35932
rect 20873 35930 20897 35932
rect 20953 35930 20977 35932
rect 21033 35930 21057 35932
rect 21113 35930 21119 35932
rect 20873 35878 20875 35930
rect 21055 35878 21057 35930
rect 20811 35876 20817 35878
rect 20873 35876 20897 35878
rect 20953 35876 20977 35878
rect 21033 35876 21057 35878
rect 21113 35876 21119 35878
rect 20811 35856 21119 35876
rect 21192 35834 21220 36110
rect 20720 35828 20772 35834
rect 20720 35770 20772 35776
rect 21180 35828 21232 35834
rect 21180 35770 21232 35776
rect 20628 35692 20680 35698
rect 20548 35652 20628 35680
rect 20444 35080 20496 35086
rect 20444 35022 20496 35028
rect 20352 34740 20404 34746
rect 20352 34682 20404 34688
rect 20456 34678 20484 35022
rect 20444 34672 20496 34678
rect 20444 34614 20496 34620
rect 20168 34060 20220 34066
rect 20168 34002 20220 34008
rect 20352 33992 20404 33998
rect 20088 33918 20208 33946
rect 20352 33934 20404 33940
rect 20076 33856 20128 33862
rect 20076 33798 20128 33804
rect 19892 33516 19944 33522
rect 19892 33458 19944 33464
rect 19800 32904 19852 32910
rect 19800 32846 19852 32852
rect 19812 32434 19840 32846
rect 19892 32768 19944 32774
rect 19892 32710 19944 32716
rect 19800 32428 19852 32434
rect 19800 32370 19852 32376
rect 19800 32020 19852 32026
rect 19800 31962 19852 31968
rect 19812 30938 19840 31962
rect 19800 30932 19852 30938
rect 19800 30874 19852 30880
rect 19904 30666 19932 32710
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 19996 31958 20024 32370
rect 19984 31952 20036 31958
rect 19984 31894 20036 31900
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 19892 30660 19944 30666
rect 19892 30602 19944 30608
rect 19904 29714 19932 30602
rect 19996 30258 20024 31078
rect 19984 30252 20036 30258
rect 19984 30194 20036 30200
rect 19892 29708 19944 29714
rect 19892 29650 19944 29656
rect 19904 29510 19932 29650
rect 19996 29646 20024 30194
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19892 29504 19944 29510
rect 19892 29446 19944 29452
rect 19708 28416 19760 28422
rect 19708 28358 19760 28364
rect 20088 27062 20116 33798
rect 20180 29510 20208 33918
rect 20364 33522 20392 33934
rect 20352 33516 20404 33522
rect 20272 33476 20352 33504
rect 20272 32298 20300 33476
rect 20352 33458 20404 33464
rect 20352 33108 20404 33114
rect 20352 33050 20404 33056
rect 20364 32502 20392 33050
rect 20456 32978 20484 34614
rect 20548 33538 20576 35652
rect 20628 35634 20680 35640
rect 20732 35290 20760 35770
rect 20720 35284 20772 35290
rect 20720 35226 20772 35232
rect 20628 35012 20680 35018
rect 20628 34954 20680 34960
rect 20640 34678 20668 34954
rect 20811 34844 21119 34864
rect 20811 34842 20817 34844
rect 20873 34842 20897 34844
rect 20953 34842 20977 34844
rect 21033 34842 21057 34844
rect 21113 34842 21119 34844
rect 20873 34790 20875 34842
rect 21055 34790 21057 34842
rect 20811 34788 20817 34790
rect 20873 34788 20897 34790
rect 20953 34788 20977 34790
rect 21033 34788 21057 34790
rect 21113 34788 21119 34790
rect 20811 34768 21119 34788
rect 20720 34740 20772 34746
rect 20720 34682 20772 34688
rect 21180 34740 21232 34746
rect 21180 34682 21232 34688
rect 20628 34672 20680 34678
rect 20628 34614 20680 34620
rect 20732 34082 20760 34682
rect 20996 34604 21048 34610
rect 20996 34546 21048 34552
rect 20824 34134 20852 34165
rect 20812 34128 20864 34134
rect 20732 34076 20812 34082
rect 20732 34070 20864 34076
rect 20732 34054 20852 34070
rect 20824 33998 20852 34054
rect 21008 33998 21036 34546
rect 20812 33992 20864 33998
rect 20812 33934 20864 33940
rect 20996 33992 21048 33998
rect 20996 33934 21048 33940
rect 20720 33924 20772 33930
rect 20720 33866 20772 33872
rect 20548 33510 20668 33538
rect 20536 33448 20588 33454
rect 20536 33390 20588 33396
rect 20444 32972 20496 32978
rect 20444 32914 20496 32920
rect 20352 32496 20404 32502
rect 20352 32438 20404 32444
rect 20260 32292 20312 32298
rect 20260 32234 20312 32240
rect 20272 31958 20300 32234
rect 20364 32026 20392 32438
rect 20352 32020 20404 32026
rect 20352 31962 20404 31968
rect 20260 31952 20312 31958
rect 20260 31894 20312 31900
rect 20352 31816 20404 31822
rect 20456 31804 20484 32914
rect 20548 32570 20576 33390
rect 20536 32564 20588 32570
rect 20536 32506 20588 32512
rect 20404 31776 20484 31804
rect 20352 31758 20404 31764
rect 20364 31346 20392 31758
rect 20352 31340 20404 31346
rect 20352 31282 20404 31288
rect 20548 30598 20576 32506
rect 20640 32434 20668 33510
rect 20732 33114 20760 33866
rect 21192 33862 21220 34682
rect 21180 33856 21232 33862
rect 21180 33798 21232 33804
rect 20811 33756 21119 33776
rect 20811 33754 20817 33756
rect 20873 33754 20897 33756
rect 20953 33754 20977 33756
rect 21033 33754 21057 33756
rect 21113 33754 21119 33756
rect 20873 33702 20875 33754
rect 21055 33702 21057 33754
rect 20811 33700 20817 33702
rect 20873 33700 20897 33702
rect 20953 33700 20977 33702
rect 21033 33700 21057 33702
rect 21113 33700 21119 33702
rect 20811 33680 21119 33700
rect 21192 33454 21220 33798
rect 20812 33448 20864 33454
rect 20812 33390 20864 33396
rect 21180 33448 21232 33454
rect 21180 33390 21232 33396
rect 20720 33108 20772 33114
rect 20720 33050 20772 33056
rect 20824 32756 20852 33390
rect 21284 33386 21312 36518
rect 21272 33380 21324 33386
rect 21272 33322 21324 33328
rect 20732 32728 20852 32756
rect 20628 32428 20680 32434
rect 20628 32370 20680 32376
rect 20640 32230 20668 32370
rect 20628 32224 20680 32230
rect 20628 32166 20680 32172
rect 20732 31346 20760 32728
rect 20811 32668 21119 32688
rect 20811 32666 20817 32668
rect 20873 32666 20897 32668
rect 20953 32666 20977 32668
rect 21033 32666 21057 32668
rect 21113 32666 21119 32668
rect 20873 32614 20875 32666
rect 21055 32614 21057 32666
rect 20811 32612 20817 32614
rect 20873 32612 20897 32614
rect 20953 32612 20977 32614
rect 21033 32612 21057 32614
rect 21113 32612 21119 32614
rect 20811 32592 21119 32612
rect 21180 31816 21232 31822
rect 21180 31758 21232 31764
rect 20811 31580 21119 31600
rect 20811 31578 20817 31580
rect 20873 31578 20897 31580
rect 20953 31578 20977 31580
rect 21033 31578 21057 31580
rect 21113 31578 21119 31580
rect 20873 31526 20875 31578
rect 21055 31526 21057 31578
rect 20811 31524 20817 31526
rect 20873 31524 20897 31526
rect 20953 31524 20977 31526
rect 21033 31524 21057 31526
rect 21113 31524 21119 31526
rect 20811 31504 21119 31524
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20732 30802 20760 31282
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20996 31272 21048 31278
rect 20996 31214 21048 31220
rect 20824 30870 20852 31214
rect 21008 30938 21036 31214
rect 21192 31210 21220 31758
rect 21180 31204 21232 31210
rect 21180 31146 21232 31152
rect 20996 30932 21048 30938
rect 20996 30874 21048 30880
rect 20812 30864 20864 30870
rect 20812 30806 20864 30812
rect 20720 30796 20772 30802
rect 20720 30738 20772 30744
rect 20824 30648 20852 30806
rect 21272 30728 21324 30734
rect 21272 30670 21324 30676
rect 20732 30620 20852 30648
rect 20536 30592 20588 30598
rect 20536 30534 20588 30540
rect 20548 30258 20576 30534
rect 20732 30326 20760 30620
rect 20811 30492 21119 30512
rect 20811 30490 20817 30492
rect 20873 30490 20897 30492
rect 20953 30490 20977 30492
rect 21033 30490 21057 30492
rect 21113 30490 21119 30492
rect 20873 30438 20875 30490
rect 21055 30438 21057 30490
rect 20811 30436 20817 30438
rect 20873 30436 20897 30438
rect 20953 30436 20977 30438
rect 21033 30436 21057 30438
rect 21113 30436 21119 30438
rect 20811 30416 21119 30436
rect 21284 30394 21312 30670
rect 21272 30388 21324 30394
rect 21272 30330 21324 30336
rect 20720 30320 20772 30326
rect 20720 30262 20772 30268
rect 20536 30252 20588 30258
rect 20588 30212 20668 30240
rect 20536 30194 20588 30200
rect 20640 29782 20668 30212
rect 20536 29776 20588 29782
rect 20536 29718 20588 29724
rect 20628 29776 20680 29782
rect 20628 29718 20680 29724
rect 20548 29578 20576 29718
rect 20260 29572 20312 29578
rect 20260 29514 20312 29520
rect 20536 29572 20588 29578
rect 20536 29514 20588 29520
rect 20168 29504 20220 29510
rect 20168 29446 20220 29452
rect 20180 29170 20208 29446
rect 20168 29164 20220 29170
rect 20168 29106 20220 29112
rect 20076 27056 20128 27062
rect 20076 26998 20128 27004
rect 19892 25832 19944 25838
rect 19892 25774 19944 25780
rect 19616 25492 19668 25498
rect 19616 25434 19668 25440
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19628 24682 19656 25434
rect 19904 24954 19932 25774
rect 20088 25514 20116 26998
rect 19996 25486 20116 25514
rect 19892 24948 19944 24954
rect 19892 24890 19944 24896
rect 19996 24818 20024 25486
rect 20076 25356 20128 25362
rect 20076 25298 20128 25304
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19616 24676 19668 24682
rect 19616 24618 19668 24624
rect 19628 24410 19656 24618
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 20088 23866 20116 25298
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20076 23860 20128 23866
rect 19996 23820 20076 23848
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 19536 23322 19564 23462
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19392 22664 19472 22692
rect 19340 22646 19392 22652
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19352 21690 19380 22646
rect 19536 22094 19564 23258
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19616 22704 19668 22710
rect 19616 22646 19668 22652
rect 19444 22066 19564 22094
rect 19444 22030 19472 22066
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19524 21888 19576 21894
rect 19524 21830 19576 21836
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19536 21554 19564 21830
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19524 21548 19576 21554
rect 19524 21490 19576 21496
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 18984 20998 19104 21026
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18984 18426 19012 20878
rect 19076 20534 19104 20998
rect 19260 20602 19288 21286
rect 19352 21146 19380 21490
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19064 20528 19116 20534
rect 19064 20470 19116 20476
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19076 19922 19104 20334
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 19076 18834 19104 19858
rect 19352 19530 19380 20946
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19260 19502 19380 19530
rect 19260 19394 19288 19502
rect 19168 19366 19288 19394
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 19168 18290 19196 19366
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 19260 18222 19288 19246
rect 19352 18970 19380 19382
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19260 17338 19288 17818
rect 19352 17746 19380 18362
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19156 17060 19208 17066
rect 19156 17002 19208 17008
rect 19168 16402 19196 17002
rect 19260 16522 19288 17274
rect 19340 17264 19392 17270
rect 19338 17232 19340 17241
rect 19392 17232 19394 17241
rect 19338 17167 19394 17176
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19248 16516 19300 16522
rect 19248 16458 19300 16464
rect 19168 16374 19288 16402
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19076 16114 19104 16186
rect 19260 16114 19288 16374
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19260 15366 19288 16050
rect 19352 16046 19380 17070
rect 19444 16114 19472 20198
rect 19536 19174 19564 21286
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19524 18352 19576 18358
rect 19524 18294 19576 18300
rect 19536 17814 19564 18294
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19628 16658 19656 22646
rect 19720 22506 19748 23054
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 19708 22500 19760 22506
rect 19708 22442 19760 22448
rect 19708 21956 19760 21962
rect 19708 21898 19760 21904
rect 19720 21146 19748 21898
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19720 18426 19748 21082
rect 19812 20942 19840 22714
rect 19996 22642 20024 23820
rect 20076 23802 20128 23808
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 20088 22778 20116 23054
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 20180 22658 20208 24754
rect 20272 23118 20300 29514
rect 20640 29102 20668 29718
rect 20732 29646 20760 30262
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20811 29404 21119 29424
rect 20811 29402 20817 29404
rect 20873 29402 20897 29404
rect 20953 29402 20977 29404
rect 21033 29402 21057 29404
rect 21113 29402 21119 29404
rect 20873 29350 20875 29402
rect 21055 29350 21057 29402
rect 20811 29348 20817 29350
rect 20873 29348 20897 29350
rect 20953 29348 20977 29350
rect 21033 29348 21057 29350
rect 21113 29348 21119 29350
rect 20811 29328 21119 29348
rect 20536 29096 20588 29102
rect 20536 29038 20588 29044
rect 20628 29096 20680 29102
rect 20628 29038 20680 29044
rect 20548 28642 20576 29038
rect 20548 28614 20668 28642
rect 20536 28484 20588 28490
rect 20536 28426 20588 28432
rect 20444 28416 20496 28422
rect 20444 28358 20496 28364
rect 20352 25832 20404 25838
rect 20352 25774 20404 25780
rect 20364 25158 20392 25774
rect 20352 25152 20404 25158
rect 20352 25094 20404 25100
rect 20364 24206 20392 25094
rect 20456 24698 20484 28358
rect 20548 28218 20576 28426
rect 20640 28422 20668 28614
rect 20628 28416 20680 28422
rect 20628 28358 20680 28364
rect 20811 28316 21119 28336
rect 20811 28314 20817 28316
rect 20873 28314 20897 28316
rect 20953 28314 20977 28316
rect 21033 28314 21057 28316
rect 21113 28314 21119 28316
rect 20873 28262 20875 28314
rect 21055 28262 21057 28314
rect 20811 28260 20817 28262
rect 20873 28260 20897 28262
rect 20953 28260 20977 28262
rect 21033 28260 21057 28262
rect 21113 28260 21119 28262
rect 20811 28240 21119 28260
rect 20536 28212 20588 28218
rect 20536 28154 20588 28160
rect 21272 28144 21324 28150
rect 21272 28086 21324 28092
rect 20720 28076 20772 28082
rect 20720 28018 20772 28024
rect 20812 28076 20864 28082
rect 20812 28018 20864 28024
rect 20732 27606 20760 28018
rect 20824 27674 20852 28018
rect 20812 27668 20864 27674
rect 20812 27610 20864 27616
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 21180 27600 21232 27606
rect 21180 27542 21232 27548
rect 20812 27532 20864 27538
rect 20812 27474 20864 27480
rect 20824 27418 20852 27474
rect 20536 27396 20588 27402
rect 20536 27338 20588 27344
rect 20732 27390 20852 27418
rect 20548 27130 20576 27338
rect 20536 27124 20588 27130
rect 20536 27066 20588 27072
rect 20732 26586 20760 27390
rect 20811 27228 21119 27248
rect 20811 27226 20817 27228
rect 20873 27226 20897 27228
rect 20953 27226 20977 27228
rect 21033 27226 21057 27228
rect 21113 27226 21119 27228
rect 20873 27174 20875 27226
rect 21055 27174 21057 27226
rect 20811 27172 20817 27174
rect 20873 27172 20897 27174
rect 20953 27172 20977 27174
rect 21033 27172 21057 27174
rect 21113 27172 21119 27174
rect 20811 27152 21119 27172
rect 20720 26580 20772 26586
rect 20720 26522 20772 26528
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20640 25294 20668 25842
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 20548 24886 20576 25230
rect 20536 24880 20588 24886
rect 20536 24822 20588 24828
rect 20536 24744 20588 24750
rect 20456 24692 20536 24698
rect 20456 24686 20588 24692
rect 20456 24670 20576 24686
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20260 23112 20312 23118
rect 20260 23054 20312 23060
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 20088 22630 20208 22658
rect 19892 22092 19944 22098
rect 19892 22034 19944 22040
rect 19904 21486 19932 22034
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 19996 21010 20024 21966
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19812 19854 19840 20878
rect 19984 20800 20036 20806
rect 19984 20742 20036 20748
rect 19892 20528 19944 20534
rect 19892 20470 19944 20476
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19536 16182 19564 16526
rect 19524 16176 19576 16182
rect 19524 16118 19576 16124
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19352 15570 19380 15982
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 18880 15088 18932 15094
rect 19352 15076 19380 15506
rect 19536 15502 19564 16118
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19432 15088 19484 15094
rect 19352 15048 19432 15076
rect 18880 15030 18932 15036
rect 19432 15030 19484 15036
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18340 11218 18368 11698
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18432 11354 18460 11630
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18156 9654 18184 9862
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18236 9104 18288 9110
rect 18234 9072 18236 9081
rect 18288 9072 18290 9081
rect 18234 9007 18290 9016
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18052 7812 18104 7818
rect 18052 7754 18104 7760
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 17500 7268 17552 7274
rect 17500 7210 17552 7216
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17052 6186 17080 6734
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6322 17264 6598
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17512 5710 17540 7210
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17604 5778 17632 7142
rect 17776 6724 17828 6730
rect 17776 6666 17828 6672
rect 17788 5846 17816 6666
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17512 4622 17540 5646
rect 17604 5098 17632 5714
rect 17788 5710 17816 5782
rect 17972 5778 18000 7482
rect 18064 7478 18092 7754
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 18064 6730 18092 7414
rect 18052 6724 18104 6730
rect 18052 6666 18104 6672
rect 18064 5914 18092 6666
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17592 5092 17644 5098
rect 17592 5034 17644 5040
rect 17788 4690 17816 5646
rect 17960 5636 18012 5642
rect 17960 5578 18012 5584
rect 17776 4684 17828 4690
rect 17776 4626 17828 4632
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16776 3466 16804 4558
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 16776 3194 16804 3402
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15580 800 15608 2382
rect 16408 800 16436 2994
rect 17052 2514 17080 4150
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17236 3602 17264 4014
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17144 2650 17172 3334
rect 17236 3058 17264 3334
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17236 2582 17264 2994
rect 17328 2854 17356 4082
rect 17972 3738 18000 5578
rect 18156 5352 18184 8910
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18248 5914 18276 7346
rect 18340 6984 18368 8910
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18432 8634 18460 8774
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18420 6996 18472 7002
rect 18340 6956 18420 6984
rect 18420 6938 18472 6944
rect 18432 6254 18460 6938
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18156 5324 18276 5352
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 4758 18092 4966
rect 18052 4752 18104 4758
rect 18052 4694 18104 4700
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 17972 3126 18000 3402
rect 18064 3194 18092 4558
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 18156 3058 18184 5170
rect 18248 5166 18276 5324
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 3194 18276 4966
rect 18524 4622 18552 11086
rect 18984 10742 19012 13194
rect 19352 12918 19380 14758
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 19076 11830 19104 12174
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 18972 10736 19024 10742
rect 18972 10678 19024 10684
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18616 7546 18644 10406
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18708 10010 18736 10066
rect 18892 10062 18920 10610
rect 19076 10470 19104 11766
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 18880 10056 18932 10062
rect 18708 9982 18828 10010
rect 18880 9998 18932 10004
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 18800 8906 18828 9982
rect 19260 9722 19288 9998
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 19248 9716 19300 9722
rect 19248 9658 19300 9664
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 18880 8900 18932 8906
rect 18880 8842 18932 8848
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8498 18736 8774
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18800 6934 18828 8842
rect 18892 8090 18920 8842
rect 19076 8838 19104 9658
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18788 6928 18840 6934
rect 18788 6870 18840 6876
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18524 4282 18552 4558
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18340 3194 18368 3334
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18524 2990 18552 3538
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18708 2854 18736 4762
rect 18984 2990 19012 5102
rect 19352 4826 19380 12242
rect 19444 9382 19472 13262
rect 19536 12832 19564 15438
rect 19628 15026 19656 16594
rect 19720 15994 19748 18226
rect 19812 17066 19840 18566
rect 19800 17060 19852 17066
rect 19800 17002 19852 17008
rect 19720 15966 19840 15994
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 19720 15502 19748 15846
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19812 15178 19840 15966
rect 19720 15150 19840 15178
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19720 13682 19748 15150
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19812 14414 19840 14962
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 19812 13938 19840 14350
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19628 13654 19748 13682
rect 19628 13462 19656 13654
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19616 13456 19668 13462
rect 19616 13398 19668 13404
rect 19616 12844 19668 12850
rect 19536 12804 19616 12832
rect 19616 12786 19668 12792
rect 19720 12238 19748 13466
rect 19904 13326 19932 20470
rect 19996 19378 20024 20742
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 19996 18970 20024 19110
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19996 16726 20024 17614
rect 19984 16720 20036 16726
rect 19984 16662 20036 16668
rect 20088 15722 20116 22630
rect 20272 22094 20300 23054
rect 20180 22066 20300 22094
rect 20180 20874 20208 22066
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20180 20058 20208 20810
rect 20272 20602 20300 21490
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20260 19848 20312 19854
rect 20180 19808 20260 19836
rect 20180 17746 20208 19808
rect 20260 19790 20312 19796
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20272 19378 20300 19654
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20364 19258 20392 23734
rect 20456 23730 20484 24550
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 20456 21690 20484 23666
rect 20548 23662 20576 24670
rect 20732 23662 20760 26522
rect 20811 26140 21119 26160
rect 20811 26138 20817 26140
rect 20873 26138 20897 26140
rect 20953 26138 20977 26140
rect 21033 26138 21057 26140
rect 21113 26138 21119 26140
rect 20873 26086 20875 26138
rect 21055 26086 21057 26138
rect 20811 26084 20817 26086
rect 20873 26084 20897 26086
rect 20953 26084 20977 26086
rect 21033 26084 21057 26086
rect 21113 26084 21119 26086
rect 20811 26064 21119 26084
rect 21192 25974 21220 27542
rect 21284 27470 21312 28086
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21284 26314 21312 27406
rect 21272 26308 21324 26314
rect 21272 26250 21324 26256
rect 20904 25968 20956 25974
rect 20904 25910 20956 25916
rect 21180 25968 21232 25974
rect 21180 25910 21232 25916
rect 20916 25294 20944 25910
rect 21088 25900 21140 25906
rect 21088 25842 21140 25848
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21008 25362 21036 25638
rect 20996 25356 21048 25362
rect 20996 25298 21048 25304
rect 21100 25294 21128 25842
rect 21180 25832 21232 25838
rect 21180 25774 21232 25780
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 21088 25288 21140 25294
rect 21088 25230 21140 25236
rect 20811 25052 21119 25072
rect 20811 25050 20817 25052
rect 20873 25050 20897 25052
rect 20953 25050 20977 25052
rect 21033 25050 21057 25052
rect 21113 25050 21119 25052
rect 20873 24998 20875 25050
rect 21055 24998 21057 25050
rect 20811 24996 20817 24998
rect 20873 24996 20897 24998
rect 20953 24996 20977 24998
rect 21033 24996 21057 24998
rect 21113 24996 21119 24998
rect 20811 24976 21119 24996
rect 21192 24954 21220 25774
rect 21272 25696 21324 25702
rect 21272 25638 21324 25644
rect 21284 25294 21312 25638
rect 21272 25288 21324 25294
rect 21272 25230 21324 25236
rect 21180 24948 21232 24954
rect 21180 24890 21232 24896
rect 20811 23964 21119 23984
rect 20811 23962 20817 23964
rect 20873 23962 20897 23964
rect 20953 23962 20977 23964
rect 21033 23962 21057 23964
rect 21113 23962 21119 23964
rect 20873 23910 20875 23962
rect 21055 23910 21057 23962
rect 20811 23908 20817 23910
rect 20873 23908 20897 23910
rect 20953 23908 20977 23910
rect 21033 23908 21057 23910
rect 21113 23908 21119 23910
rect 20811 23888 21119 23908
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 20720 23656 20772 23662
rect 20720 23598 20772 23604
rect 20628 23588 20680 23594
rect 20628 23530 20680 23536
rect 20536 23044 20588 23050
rect 20536 22986 20588 22992
rect 20548 22710 20576 22986
rect 20536 22704 20588 22710
rect 20536 22646 20588 22652
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20456 20398 20484 20946
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 20456 19446 20484 20334
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20548 19378 20576 21286
rect 20640 20602 20668 23530
rect 20732 23186 20760 23598
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20732 22760 20760 22918
rect 20811 22876 21119 22896
rect 20811 22874 20817 22876
rect 20873 22874 20897 22876
rect 20953 22874 20977 22876
rect 21033 22874 21057 22876
rect 21113 22874 21119 22876
rect 20873 22822 20875 22874
rect 21055 22822 21057 22874
rect 20811 22820 20817 22822
rect 20873 22820 20897 22822
rect 20953 22820 20977 22822
rect 21033 22820 21057 22822
rect 21113 22820 21119 22822
rect 20811 22800 21119 22820
rect 21192 22778 21220 23054
rect 21180 22772 21232 22778
rect 20732 22732 20852 22760
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20732 22234 20760 22578
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20824 22098 20852 22732
rect 21180 22714 21232 22720
rect 21284 22642 21312 23122
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20732 21078 20760 21966
rect 20811 21788 21119 21808
rect 20811 21786 20817 21788
rect 20873 21786 20897 21788
rect 20953 21786 20977 21788
rect 21033 21786 21057 21788
rect 21113 21786 21119 21788
rect 20873 21734 20875 21786
rect 21055 21734 21057 21786
rect 20811 21732 20817 21734
rect 20873 21732 20897 21734
rect 20953 21732 20977 21734
rect 21033 21732 21057 21734
rect 21113 21732 21119 21734
rect 20811 21712 21119 21732
rect 20720 21072 20772 21078
rect 20720 21014 20772 21020
rect 21376 20942 21404 38694
rect 21548 36304 21600 36310
rect 21548 36246 21600 36252
rect 21456 31680 21508 31686
rect 21456 31622 21508 31628
rect 21468 31414 21496 31622
rect 21456 31408 21508 31414
rect 21456 31350 21508 31356
rect 21456 31204 21508 31210
rect 21456 31146 21508 31152
rect 21468 29102 21496 31146
rect 21560 30870 21588 36246
rect 21732 33992 21784 33998
rect 21732 33934 21784 33940
rect 21744 33658 21772 33934
rect 21732 33652 21784 33658
rect 21732 33594 21784 33600
rect 21836 33318 21864 39918
rect 21928 39098 21956 42162
rect 25776 41916 26084 41936
rect 25776 41914 25782 41916
rect 25838 41914 25862 41916
rect 25918 41914 25942 41916
rect 25998 41914 26022 41916
rect 26078 41914 26084 41916
rect 25838 41862 25840 41914
rect 26020 41862 26022 41914
rect 25776 41860 25782 41862
rect 25838 41860 25862 41862
rect 25918 41860 25942 41862
rect 25998 41860 26022 41862
rect 26078 41860 26084 41862
rect 25776 41840 26084 41860
rect 30104 41132 30156 41138
rect 30104 41074 30156 41080
rect 30116 41041 30144 41074
rect 30102 41032 30158 41041
rect 30102 40967 30158 40976
rect 29920 40928 29972 40934
rect 29920 40870 29972 40876
rect 25776 40828 26084 40848
rect 25776 40826 25782 40828
rect 25838 40826 25862 40828
rect 25918 40826 25942 40828
rect 25998 40826 26022 40828
rect 26078 40826 26084 40828
rect 25838 40774 25840 40826
rect 26020 40774 26022 40826
rect 25776 40772 25782 40774
rect 25838 40772 25862 40774
rect 25918 40772 25942 40774
rect 25998 40772 26022 40774
rect 26078 40772 26084 40774
rect 25776 40752 26084 40772
rect 22100 40044 22152 40050
rect 22100 39986 22152 39992
rect 21916 39092 21968 39098
rect 21916 39034 21968 39040
rect 22112 38962 22140 39986
rect 29932 39982 29960 40870
rect 29920 39976 29972 39982
rect 29920 39918 29972 39924
rect 25776 39740 26084 39760
rect 25776 39738 25782 39740
rect 25838 39738 25862 39740
rect 25918 39738 25942 39740
rect 25998 39738 26022 39740
rect 26078 39738 26084 39740
rect 25838 39686 25840 39738
rect 26020 39686 26022 39738
rect 25776 39684 25782 39686
rect 25838 39684 25862 39686
rect 25918 39684 25942 39686
rect 25998 39684 26022 39686
rect 26078 39684 26084 39686
rect 25776 39664 26084 39684
rect 30104 39432 30156 39438
rect 30104 39374 30156 39380
rect 29920 39296 29972 39302
rect 29920 39238 29972 39244
rect 22100 38956 22152 38962
rect 22100 38898 22152 38904
rect 22112 36786 22140 38898
rect 29932 38894 29960 39238
rect 30116 39001 30144 39374
rect 30102 38992 30158 39001
rect 30102 38927 30158 38936
rect 29920 38888 29972 38894
rect 29920 38830 29972 38836
rect 25776 38652 26084 38672
rect 25776 38650 25782 38652
rect 25838 38650 25862 38652
rect 25918 38650 25942 38652
rect 25998 38650 26022 38652
rect 26078 38650 26084 38652
rect 25838 38598 25840 38650
rect 26020 38598 26022 38650
rect 25776 38596 25782 38598
rect 25838 38596 25862 38598
rect 25918 38596 25942 38598
rect 25998 38596 26022 38598
rect 26078 38596 26084 38598
rect 25776 38576 26084 38596
rect 25776 37564 26084 37584
rect 25776 37562 25782 37564
rect 25838 37562 25862 37564
rect 25918 37562 25942 37564
rect 25998 37562 26022 37564
rect 26078 37562 26084 37564
rect 25838 37510 25840 37562
rect 26020 37510 26022 37562
rect 25776 37508 25782 37510
rect 25838 37508 25862 37510
rect 25918 37508 25942 37510
rect 25998 37508 26022 37510
rect 26078 37508 26084 37510
rect 25776 37488 26084 37508
rect 30104 37256 30156 37262
rect 30104 37198 30156 37204
rect 29920 37120 29972 37126
rect 29920 37062 29972 37068
rect 22100 36780 22152 36786
rect 22100 36722 22152 36728
rect 22112 35894 22140 36722
rect 29932 36718 29960 37062
rect 30116 36961 30144 37198
rect 30102 36952 30158 36961
rect 30102 36887 30158 36896
rect 29920 36712 29972 36718
rect 29920 36654 29972 36660
rect 25776 36476 26084 36496
rect 25776 36474 25782 36476
rect 25838 36474 25862 36476
rect 25918 36474 25942 36476
rect 25998 36474 26022 36476
rect 26078 36474 26084 36476
rect 25838 36422 25840 36474
rect 26020 36422 26022 36474
rect 25776 36420 25782 36422
rect 25838 36420 25862 36422
rect 25918 36420 25942 36422
rect 25998 36420 26022 36422
rect 26078 36420 26084 36422
rect 25776 36400 26084 36420
rect 22112 35866 22232 35894
rect 22204 35086 22232 35866
rect 25776 35388 26084 35408
rect 25776 35386 25782 35388
rect 25838 35386 25862 35388
rect 25918 35386 25942 35388
rect 25998 35386 26022 35388
rect 26078 35386 26084 35388
rect 25838 35334 25840 35386
rect 26020 35334 26022 35386
rect 25776 35332 25782 35334
rect 25838 35332 25862 35334
rect 25918 35332 25942 35334
rect 25998 35332 26022 35334
rect 26078 35332 26084 35334
rect 25776 35312 26084 35332
rect 22192 35080 22244 35086
rect 30104 35080 30156 35086
rect 30102 35048 30104 35057
rect 30156 35048 30158 35057
rect 22244 35028 22324 35034
rect 22192 35022 22324 35028
rect 22204 35006 22324 35022
rect 21916 34944 21968 34950
rect 21916 34886 21968 34892
rect 21928 34406 21956 34886
rect 21916 34400 21968 34406
rect 21916 34342 21968 34348
rect 22008 34128 22060 34134
rect 22008 34070 22060 34076
rect 21824 33312 21876 33318
rect 21824 33254 21876 33260
rect 21640 32224 21692 32230
rect 21640 32166 21692 32172
rect 21548 30864 21600 30870
rect 21548 30806 21600 30812
rect 21652 30734 21680 32166
rect 22020 31890 22048 34070
rect 22296 32910 22324 35006
rect 30102 34983 30158 34992
rect 25776 34300 26084 34320
rect 25776 34298 25782 34300
rect 25838 34298 25862 34300
rect 25918 34298 25942 34300
rect 25998 34298 26022 34300
rect 26078 34298 26084 34300
rect 25838 34246 25840 34298
rect 26020 34246 26022 34298
rect 25776 34244 25782 34246
rect 25838 34244 25862 34246
rect 25918 34244 25942 34246
rect 25998 34244 26022 34246
rect 26078 34244 26084 34246
rect 25776 34224 26084 34244
rect 22376 33856 22428 33862
rect 22376 33798 22428 33804
rect 22388 33522 22416 33798
rect 22376 33516 22428 33522
rect 22376 33458 22428 33464
rect 30104 33516 30156 33522
rect 30104 33458 30156 33464
rect 22560 33312 22612 33318
rect 22560 33254 22612 33260
rect 29920 33312 29972 33318
rect 29920 33254 29972 33260
rect 22284 32904 22336 32910
rect 22284 32846 22336 32852
rect 22100 32768 22152 32774
rect 22100 32710 22152 32716
rect 22008 31884 22060 31890
rect 22008 31826 22060 31832
rect 22020 31754 22048 31826
rect 21928 31726 22048 31754
rect 21732 31272 21784 31278
rect 21732 31214 21784 31220
rect 21640 30728 21692 30734
rect 21744 30716 21772 31214
rect 21824 30728 21876 30734
rect 21744 30688 21824 30716
rect 21640 30670 21692 30676
rect 21824 30670 21876 30676
rect 21836 30190 21864 30670
rect 21824 30184 21876 30190
rect 21824 30126 21876 30132
rect 21836 29866 21864 30126
rect 21928 30036 21956 31726
rect 22112 31414 22140 32710
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 22020 30734 22048 31282
rect 22296 31278 22324 32846
rect 22284 31272 22336 31278
rect 22284 31214 22336 31220
rect 22008 30728 22060 30734
rect 22008 30670 22060 30676
rect 22376 30728 22428 30734
rect 22376 30670 22428 30676
rect 22388 30258 22416 30670
rect 22376 30252 22428 30258
rect 22376 30194 22428 30200
rect 22008 30048 22060 30054
rect 21928 30008 22008 30036
rect 22008 29990 22060 29996
rect 22192 30048 22244 30054
rect 22192 29990 22244 29996
rect 21548 29844 21600 29850
rect 21836 29838 21956 29866
rect 21548 29786 21600 29792
rect 21560 29238 21588 29786
rect 21824 29640 21876 29646
rect 21824 29582 21876 29588
rect 21836 29306 21864 29582
rect 21824 29300 21876 29306
rect 21824 29242 21876 29248
rect 21548 29232 21600 29238
rect 21548 29174 21600 29180
rect 21456 29096 21508 29102
rect 21456 29038 21508 29044
rect 21732 29096 21784 29102
rect 21732 29038 21784 29044
rect 21548 28008 21600 28014
rect 21548 27950 21600 27956
rect 21560 27470 21588 27950
rect 21548 27464 21600 27470
rect 21548 27406 21600 27412
rect 21456 25900 21508 25906
rect 21456 25842 21508 25848
rect 21468 25498 21496 25842
rect 21456 25492 21508 25498
rect 21456 25434 21508 25440
rect 21560 25226 21588 27406
rect 21640 26784 21692 26790
rect 21640 26726 21692 26732
rect 21652 26450 21680 26726
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21548 25220 21600 25226
rect 21548 25162 21600 25168
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21468 23186 21496 24006
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 21560 22506 21588 25162
rect 21744 24886 21772 29038
rect 21928 28218 21956 29838
rect 22100 29572 22152 29578
rect 22100 29514 22152 29520
rect 22008 28756 22060 28762
rect 22008 28698 22060 28704
rect 21916 28212 21968 28218
rect 21916 28154 21968 28160
rect 21824 25832 21876 25838
rect 21824 25774 21876 25780
rect 21836 25362 21864 25774
rect 21824 25356 21876 25362
rect 21824 25298 21876 25304
rect 21732 24880 21784 24886
rect 21732 24822 21784 24828
rect 21928 24274 21956 28154
rect 22020 28150 22048 28698
rect 22112 28558 22140 29514
rect 22100 28552 22152 28558
rect 22100 28494 22152 28500
rect 22008 28144 22060 28150
rect 22008 28086 22060 28092
rect 22112 28082 22140 28494
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22112 26518 22140 26862
rect 22100 26512 22152 26518
rect 22100 26454 22152 26460
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 22008 26308 22060 26314
rect 22008 26250 22060 26256
rect 21916 24268 21968 24274
rect 21916 24210 21968 24216
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21548 22500 21600 22506
rect 21548 22442 21600 22448
rect 21456 21956 21508 21962
rect 21456 21898 21508 21904
rect 21468 21554 21496 21898
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20732 20466 20760 20742
rect 20811 20700 21119 20720
rect 20811 20698 20817 20700
rect 20873 20698 20897 20700
rect 20953 20698 20977 20700
rect 21033 20698 21057 20700
rect 21113 20698 21119 20700
rect 20873 20646 20875 20698
rect 21055 20646 21057 20698
rect 20811 20644 20817 20646
rect 20873 20644 20897 20646
rect 20953 20644 20977 20646
rect 21033 20644 21057 20646
rect 21113 20644 21119 20646
rect 20811 20624 21119 20644
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20640 19446 20668 19790
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20272 19230 20392 19258
rect 20168 17740 20220 17746
rect 20168 17682 20220 17688
rect 20180 17338 20208 17682
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 19996 15694 20116 15722
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19996 12918 20024 15694
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19904 11762 19932 12038
rect 19996 11830 20024 12854
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 20088 11354 20116 14350
rect 20272 13530 20300 19230
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20364 18766 20392 19110
rect 20456 18834 20484 19110
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20364 16794 20392 17070
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20364 16182 20392 16730
rect 20456 16590 20484 16934
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20548 15994 20576 18906
rect 20640 18426 20668 19382
rect 20732 18426 20760 20402
rect 20811 19612 21119 19632
rect 20811 19610 20817 19612
rect 20873 19610 20897 19612
rect 20953 19610 20977 19612
rect 21033 19610 21057 19612
rect 21113 19610 21119 19612
rect 20873 19558 20875 19610
rect 21055 19558 21057 19610
rect 20811 19556 20817 19558
rect 20873 19556 20897 19558
rect 20953 19556 20977 19558
rect 21033 19556 21057 19558
rect 21113 19556 21119 19558
rect 20811 19536 21119 19556
rect 20811 18524 21119 18544
rect 20811 18522 20817 18524
rect 20873 18522 20897 18524
rect 20953 18522 20977 18524
rect 21033 18522 21057 18524
rect 21113 18522 21119 18524
rect 20873 18470 20875 18522
rect 21055 18470 21057 18522
rect 20811 18468 20817 18470
rect 20873 18468 20897 18470
rect 20953 18468 20977 18470
rect 21033 18468 21057 18470
rect 21113 18468 21119 18470
rect 20811 18448 21119 18468
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 20640 17241 20668 17614
rect 21284 17542 21312 17614
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 20811 17436 21119 17456
rect 20811 17434 20817 17436
rect 20873 17434 20897 17436
rect 20953 17434 20977 17436
rect 21033 17434 21057 17436
rect 21113 17434 21119 17436
rect 20873 17382 20875 17434
rect 21055 17382 21057 17434
rect 20811 17380 20817 17382
rect 20873 17380 20897 17382
rect 20953 17380 20977 17382
rect 21033 17380 21057 17382
rect 21113 17380 21119 17382
rect 20811 17360 21119 17380
rect 20626 17232 20682 17241
rect 21284 17202 21312 17478
rect 20626 17167 20682 17176
rect 21272 17196 21324 17202
rect 20640 17134 20668 17167
rect 21272 17138 21324 17144
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 20811 16348 21119 16368
rect 20811 16346 20817 16348
rect 20873 16346 20897 16348
rect 20953 16346 20977 16348
rect 21033 16346 21057 16348
rect 21113 16346 21119 16348
rect 20873 16294 20875 16346
rect 21055 16294 21057 16346
rect 20811 16292 20817 16294
rect 20873 16292 20897 16294
rect 20953 16292 20977 16294
rect 21033 16292 21057 16294
rect 21113 16292 21119 16294
rect 20811 16272 21119 16292
rect 21284 16182 21312 17138
rect 21272 16176 21324 16182
rect 21272 16118 21324 16124
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 20548 15966 20760 15994
rect 20732 15910 20760 15966
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20364 13326 20392 13874
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20364 12238 20392 13262
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 20180 11234 20208 11630
rect 20088 11218 20208 11234
rect 20088 11212 20220 11218
rect 20088 11206 20168 11212
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19444 8022 19472 8366
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19536 6866 19564 11086
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19996 10266 20024 10610
rect 20088 10606 20116 11206
rect 20168 11154 20220 11160
rect 20180 11123 20208 11154
rect 20272 11150 20300 11630
rect 20364 11354 20392 11698
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20272 10606 20300 11086
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19812 8634 19840 8842
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19720 7342 19748 7822
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19720 6390 19748 7278
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19444 5710 19472 6258
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19352 4214 19380 4558
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 19352 3738 19380 4150
rect 19444 4146 19472 4422
rect 19720 4146 19748 6326
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19812 4622 19840 5646
rect 19904 5370 19932 9998
rect 20364 9722 20392 10610
rect 20352 9716 20404 9722
rect 20352 9658 20404 9664
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20272 9042 20300 9318
rect 20456 9178 20484 11698
rect 20548 10810 20576 14962
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20640 14414 20668 14894
rect 20732 14618 20760 15846
rect 20824 15706 20852 16050
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20811 15260 21119 15280
rect 20811 15258 20817 15260
rect 20873 15258 20897 15260
rect 20953 15258 20977 15260
rect 21033 15258 21057 15260
rect 21113 15258 21119 15260
rect 20873 15206 20875 15258
rect 21055 15206 21057 15258
rect 20811 15204 20817 15206
rect 20873 15204 20897 15206
rect 20953 15204 20977 15206
rect 21033 15204 21057 15206
rect 21113 15204 21119 15206
rect 20811 15184 21119 15204
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 21192 14414 21220 16050
rect 21468 15502 21496 21490
rect 21652 19990 21680 24074
rect 21928 23798 21956 24210
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 22020 22778 22048 26250
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 22020 22098 22048 22714
rect 22112 22658 22140 26318
rect 22204 23254 22232 29990
rect 22388 28082 22416 30194
rect 22468 29504 22520 29510
rect 22468 29446 22520 29452
rect 22480 29170 22508 29446
rect 22572 29170 22600 33254
rect 25776 33212 26084 33232
rect 25776 33210 25782 33212
rect 25838 33210 25862 33212
rect 25918 33210 25942 33212
rect 25998 33210 26022 33212
rect 26078 33210 26084 33212
rect 25838 33158 25840 33210
rect 26020 33158 26022 33210
rect 25776 33156 25782 33158
rect 25838 33156 25862 33158
rect 25918 33156 25942 33158
rect 25998 33156 26022 33158
rect 26078 33156 26084 33158
rect 25776 33136 26084 33156
rect 29932 32910 29960 33254
rect 30116 33017 30144 33458
rect 30102 33008 30158 33017
rect 30102 32943 30158 32952
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 29828 32360 29880 32366
rect 29828 32302 29880 32308
rect 25776 32124 26084 32144
rect 25776 32122 25782 32124
rect 25838 32122 25862 32124
rect 25918 32122 25942 32124
rect 25998 32122 26022 32124
rect 26078 32122 26084 32124
rect 25838 32070 25840 32122
rect 26020 32070 26022 32122
rect 25776 32068 25782 32070
rect 25838 32068 25862 32070
rect 25918 32068 25942 32070
rect 25998 32068 26022 32070
rect 26078 32068 26084 32070
rect 25776 32048 26084 32068
rect 29840 31346 29868 32302
rect 29828 31340 29880 31346
rect 29828 31282 29880 31288
rect 30104 31272 30156 31278
rect 30104 31214 30156 31220
rect 25776 31036 26084 31056
rect 25776 31034 25782 31036
rect 25838 31034 25862 31036
rect 25918 31034 25942 31036
rect 25998 31034 26022 31036
rect 26078 31034 26084 31036
rect 25838 30982 25840 31034
rect 26020 30982 26022 31034
rect 25776 30980 25782 30982
rect 25838 30980 25862 30982
rect 25918 30980 25942 30982
rect 25998 30980 26022 30982
rect 26078 30980 26084 30982
rect 25776 30960 26084 30980
rect 30116 30977 30144 31214
rect 30102 30968 30158 30977
rect 30102 30903 30158 30912
rect 22652 30660 22704 30666
rect 22652 30602 22704 30608
rect 22664 30258 22692 30602
rect 22652 30252 22704 30258
rect 22652 30194 22704 30200
rect 25776 29948 26084 29968
rect 25776 29946 25782 29948
rect 25838 29946 25862 29948
rect 25918 29946 25942 29948
rect 25998 29946 26022 29948
rect 26078 29946 26084 29948
rect 25838 29894 25840 29946
rect 26020 29894 26022 29946
rect 25776 29892 25782 29894
rect 25838 29892 25862 29894
rect 25918 29892 25942 29894
rect 25998 29892 26022 29894
rect 26078 29892 26084 29894
rect 25776 29872 26084 29892
rect 29736 29640 29788 29646
rect 29736 29582 29788 29588
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 25776 28860 26084 28880
rect 25776 28858 25782 28860
rect 25838 28858 25862 28860
rect 25918 28858 25942 28860
rect 25998 28858 26022 28860
rect 26078 28858 26084 28860
rect 25838 28806 25840 28858
rect 26020 28806 26022 28858
rect 25776 28804 25782 28806
rect 25838 28804 25862 28806
rect 25918 28804 25942 28806
rect 25998 28804 26022 28806
rect 26078 28804 26084 28806
rect 25776 28784 26084 28804
rect 29092 28416 29144 28422
rect 29092 28358 29144 28364
rect 22376 28076 22428 28082
rect 22376 28018 22428 28024
rect 22284 27056 22336 27062
rect 22284 26998 22336 27004
rect 22296 26042 22324 26998
rect 22388 26450 22416 28018
rect 25776 27772 26084 27792
rect 25776 27770 25782 27772
rect 25838 27770 25862 27772
rect 25918 27770 25942 27772
rect 25998 27770 26022 27772
rect 26078 27770 26084 27772
rect 25838 27718 25840 27770
rect 26020 27718 26022 27770
rect 25776 27716 25782 27718
rect 25838 27716 25862 27718
rect 25918 27716 25942 27718
rect 25998 27716 26022 27718
rect 26078 27716 26084 27718
rect 25776 27696 26084 27716
rect 25776 26684 26084 26704
rect 25776 26682 25782 26684
rect 25838 26682 25862 26684
rect 25918 26682 25942 26684
rect 25998 26682 26022 26684
rect 26078 26682 26084 26684
rect 25838 26630 25840 26682
rect 26020 26630 26022 26682
rect 25776 26628 25782 26630
rect 25838 26628 25862 26630
rect 25918 26628 25942 26630
rect 25998 26628 26022 26630
rect 26078 26628 26084 26630
rect 25776 26608 26084 26628
rect 22376 26444 22428 26450
rect 22376 26386 22428 26392
rect 23112 26376 23164 26382
rect 23112 26318 23164 26324
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 22296 24138 22324 25978
rect 23124 25702 23152 26318
rect 23204 26036 23256 26042
rect 23204 25978 23256 25984
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 23112 25696 23164 25702
rect 23112 25638 23164 25644
rect 22480 25158 22508 25638
rect 23216 25498 23244 25978
rect 25776 25596 26084 25616
rect 25776 25594 25782 25596
rect 25838 25594 25862 25596
rect 25918 25594 25942 25596
rect 25998 25594 26022 25596
rect 26078 25594 26084 25596
rect 25838 25542 25840 25594
rect 26020 25542 26022 25594
rect 25776 25540 25782 25542
rect 25838 25540 25862 25542
rect 25918 25540 25942 25542
rect 25998 25540 26022 25542
rect 26078 25540 26084 25542
rect 25776 25520 26084 25540
rect 23204 25492 23256 25498
rect 23204 25434 23256 25440
rect 22468 25152 22520 25158
rect 22468 25094 22520 25100
rect 22480 24274 22508 25094
rect 25776 24508 26084 24528
rect 25776 24506 25782 24508
rect 25838 24506 25862 24508
rect 25918 24506 25942 24508
rect 25998 24506 26022 24508
rect 26078 24506 26084 24508
rect 25838 24454 25840 24506
rect 26020 24454 26022 24506
rect 25776 24452 25782 24454
rect 25838 24452 25862 24454
rect 25918 24452 25942 24454
rect 25998 24452 26022 24454
rect 26078 24452 26084 24454
rect 25776 24432 26084 24452
rect 22468 24268 22520 24274
rect 22468 24210 22520 24216
rect 22284 24132 22336 24138
rect 22284 24074 22336 24080
rect 22296 23866 22324 24074
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22192 23248 22244 23254
rect 22192 23190 22244 23196
rect 22192 23112 22244 23118
rect 22192 23054 22244 23060
rect 22204 22778 22232 23054
rect 22296 23050 22324 23802
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22284 23044 22336 23050
rect 22284 22986 22336 22992
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22112 22630 22324 22658
rect 22100 22228 22152 22234
rect 22100 22170 22152 22176
rect 22008 22092 22060 22098
rect 22008 22034 22060 22040
rect 22020 20942 22048 22034
rect 22112 22030 22140 22170
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22008 20936 22060 20942
rect 21928 20896 22008 20924
rect 21928 20398 21956 20896
rect 22008 20878 22060 20884
rect 22296 20602 22324 22630
rect 22388 21962 22416 23122
rect 22480 22710 22508 24210
rect 22836 23724 22888 23730
rect 22836 23666 22888 23672
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22664 23322 22692 23598
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22848 22710 22876 23666
rect 22928 23656 22980 23662
rect 22928 23598 22980 23604
rect 22940 23186 22968 23598
rect 25776 23420 26084 23440
rect 25776 23418 25782 23420
rect 25838 23418 25862 23420
rect 25918 23418 25942 23420
rect 25998 23418 26022 23420
rect 26078 23418 26084 23420
rect 25838 23366 25840 23418
rect 26020 23366 26022 23418
rect 25776 23364 25782 23366
rect 25838 23364 25862 23366
rect 25918 23364 25942 23366
rect 25998 23364 26022 23366
rect 26078 23364 26084 23366
rect 25776 23344 26084 23364
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 22928 23044 22980 23050
rect 22928 22986 22980 22992
rect 22940 22778 22968 22986
rect 23388 22976 23440 22982
rect 23388 22918 23440 22924
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 23400 22710 23428 22918
rect 22468 22704 22520 22710
rect 22468 22646 22520 22652
rect 22836 22704 22888 22710
rect 22836 22646 22888 22652
rect 23020 22704 23072 22710
rect 23020 22646 23072 22652
rect 23388 22704 23440 22710
rect 23388 22646 23440 22652
rect 22848 22234 22876 22646
rect 22836 22228 22888 22234
rect 22836 22170 22888 22176
rect 22376 21956 22428 21962
rect 22376 21898 22428 21904
rect 22388 20942 22416 21898
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 22388 20534 22416 20878
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 22376 20528 22428 20534
rect 22376 20470 22428 20476
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 21640 19984 21692 19990
rect 21640 19926 21692 19932
rect 21652 16114 21680 19926
rect 21928 19854 21956 20334
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 21928 19514 21956 19790
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 21928 18834 21956 19450
rect 22020 19446 22048 20470
rect 23032 19854 23060 22646
rect 25776 22332 26084 22352
rect 25776 22330 25782 22332
rect 25838 22330 25862 22332
rect 25918 22330 25942 22332
rect 25998 22330 26022 22332
rect 26078 22330 26084 22332
rect 25838 22278 25840 22330
rect 26020 22278 26022 22330
rect 25776 22276 25782 22278
rect 25838 22276 25862 22278
rect 25918 22276 25942 22278
rect 25998 22276 26022 22278
rect 26078 22276 26084 22278
rect 25776 22256 26084 22276
rect 25776 21244 26084 21264
rect 25776 21242 25782 21244
rect 25838 21242 25862 21244
rect 25918 21242 25942 21244
rect 25998 21242 26022 21244
rect 26078 21242 26084 21244
rect 25838 21190 25840 21242
rect 26020 21190 26022 21242
rect 25776 21188 25782 21190
rect 25838 21188 25862 21190
rect 25918 21188 25942 21190
rect 25998 21188 26022 21190
rect 26078 21188 26084 21190
rect 25776 21168 26084 21188
rect 25776 20156 26084 20176
rect 25776 20154 25782 20156
rect 25838 20154 25862 20156
rect 25918 20154 25942 20156
rect 25998 20154 26022 20156
rect 26078 20154 26084 20156
rect 25838 20102 25840 20154
rect 26020 20102 26022 20154
rect 25776 20100 25782 20102
rect 25838 20100 25862 20102
rect 25918 20100 25942 20102
rect 25998 20100 26022 20102
rect 26078 20100 26084 20102
rect 25776 20080 26084 20100
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 22008 19440 22060 19446
rect 22008 19382 22060 19388
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 22020 18766 22048 19382
rect 22480 19378 22508 19790
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22480 18766 22508 19314
rect 25776 19068 26084 19088
rect 25776 19066 25782 19068
rect 25838 19066 25862 19068
rect 25918 19066 25942 19068
rect 25998 19066 26022 19068
rect 26078 19066 26084 19068
rect 25838 19014 25840 19066
rect 26020 19014 26022 19066
rect 25776 19012 25782 19014
rect 25838 19012 25862 19014
rect 25918 19012 25942 19014
rect 25998 19012 26022 19014
rect 26078 19012 26084 19014
rect 25776 18992 26084 19012
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21836 17338 21864 18226
rect 22020 17882 22048 18226
rect 25776 17980 26084 18000
rect 25776 17978 25782 17980
rect 25838 17978 25862 17980
rect 25918 17978 25942 17980
rect 25998 17978 26022 17980
rect 26078 17978 26084 17980
rect 25838 17926 25840 17978
rect 26020 17926 26022 17978
rect 25776 17924 25782 17926
rect 25838 17924 25862 17926
rect 25918 17924 25942 17926
rect 25998 17924 26022 17926
rect 26078 17924 26084 17926
rect 25776 17904 26084 17924
rect 22008 17876 22060 17882
rect 22008 17818 22060 17824
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21836 16794 21864 17138
rect 25776 16892 26084 16912
rect 25776 16890 25782 16892
rect 25838 16890 25862 16892
rect 25918 16890 25942 16892
rect 25998 16890 26022 16892
rect 26078 16890 26084 16892
rect 25838 16838 25840 16890
rect 26020 16838 26022 16890
rect 25776 16836 25782 16838
rect 25838 16836 25862 16838
rect 25918 16836 25942 16838
rect 25998 16836 26022 16838
rect 26078 16836 26084 16838
rect 25776 16816 26084 16836
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 25776 15804 26084 15824
rect 25776 15802 25782 15804
rect 25838 15802 25862 15804
rect 25918 15802 25942 15804
rect 25998 15802 26022 15804
rect 26078 15802 26084 15804
rect 25838 15750 25840 15802
rect 26020 15750 26022 15802
rect 25776 15748 25782 15750
rect 25838 15748 25862 15750
rect 25918 15748 25942 15750
rect 25998 15748 26022 15750
rect 26078 15748 26084 15750
rect 25776 15728 26084 15748
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 20640 14260 20668 14350
rect 20720 14272 20772 14278
rect 20640 14232 20720 14260
rect 20720 14214 20772 14220
rect 20732 13938 20760 14214
rect 20811 14172 21119 14192
rect 20811 14170 20817 14172
rect 20873 14170 20897 14172
rect 20953 14170 20977 14172
rect 21033 14170 21057 14172
rect 21113 14170 21119 14172
rect 20873 14118 20875 14170
rect 21055 14118 21057 14170
rect 20811 14116 20817 14118
rect 20873 14116 20897 14118
rect 20953 14116 20977 14118
rect 21033 14116 21057 14118
rect 21113 14116 21119 14118
rect 20811 14096 21119 14116
rect 21192 14006 21220 14350
rect 21180 14000 21232 14006
rect 21180 13942 21232 13948
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20732 13326 20760 13874
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20628 12232 20680 12238
rect 20732 12220 20760 13262
rect 20811 13084 21119 13104
rect 20811 13082 20817 13084
rect 20873 13082 20897 13084
rect 20953 13082 20977 13084
rect 21033 13082 21057 13084
rect 21113 13082 21119 13084
rect 20873 13030 20875 13082
rect 21055 13030 21057 13082
rect 20811 13028 20817 13030
rect 20873 13028 20897 13030
rect 20953 13028 20977 13030
rect 21033 13028 21057 13030
rect 21113 13028 21119 13030
rect 20811 13008 21119 13028
rect 21468 12238 21496 15438
rect 21824 15360 21876 15366
rect 21824 15302 21876 15308
rect 21836 15026 21864 15302
rect 21824 15020 21876 15026
rect 21824 14962 21876 14968
rect 25776 14716 26084 14736
rect 25776 14714 25782 14716
rect 25838 14714 25862 14716
rect 25918 14714 25942 14716
rect 25998 14714 26022 14716
rect 26078 14714 26084 14716
rect 25838 14662 25840 14714
rect 26020 14662 26022 14714
rect 25776 14660 25782 14662
rect 25838 14660 25862 14662
rect 25918 14660 25942 14662
rect 25998 14660 26022 14662
rect 26078 14660 26084 14662
rect 25776 14640 26084 14660
rect 29012 14550 29040 16050
rect 29000 14544 29052 14550
rect 29000 14486 29052 14492
rect 25776 13628 26084 13648
rect 25776 13626 25782 13628
rect 25838 13626 25862 13628
rect 25918 13626 25942 13628
rect 25998 13626 26022 13628
rect 26078 13626 26084 13628
rect 25838 13574 25840 13626
rect 26020 13574 26022 13626
rect 25776 13572 25782 13574
rect 25838 13572 25862 13574
rect 25918 13572 25942 13574
rect 25998 13572 26022 13574
rect 26078 13572 26084 13574
rect 25776 13552 26084 13572
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 20812 12232 20864 12238
rect 20732 12192 20812 12220
rect 20628 12174 20680 12180
rect 20812 12174 20864 12180
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 20640 11898 20668 12174
rect 21652 12170 21680 12786
rect 25776 12540 26084 12560
rect 25776 12538 25782 12540
rect 25838 12538 25862 12540
rect 25918 12538 25942 12540
rect 25998 12538 26022 12540
rect 26078 12538 26084 12540
rect 25838 12486 25840 12538
rect 26020 12486 26022 12538
rect 25776 12484 25782 12486
rect 25838 12484 25862 12486
rect 25918 12484 25942 12486
rect 25998 12484 26022 12486
rect 26078 12484 26084 12486
rect 25776 12464 26084 12484
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 20811 11996 21119 12016
rect 20811 11994 20817 11996
rect 20873 11994 20897 11996
rect 20953 11994 20977 11996
rect 21033 11994 21057 11996
rect 21113 11994 21119 11996
rect 20873 11942 20875 11994
rect 21055 11942 21057 11994
rect 20811 11940 20817 11942
rect 20873 11940 20897 11942
rect 20953 11940 20977 11942
rect 21033 11940 21057 11942
rect 21113 11940 21119 11942
rect 20811 11920 21119 11940
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20640 11150 20668 11494
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20732 10810 20760 11018
rect 20811 10908 21119 10928
rect 20811 10906 20817 10908
rect 20873 10906 20897 10908
rect 20953 10906 20977 10908
rect 21033 10906 21057 10908
rect 21113 10906 21119 10908
rect 20873 10854 20875 10906
rect 21055 10854 21057 10906
rect 20811 10852 20817 10854
rect 20873 10852 20897 10854
rect 20953 10852 20977 10854
rect 21033 10852 21057 10854
rect 21113 10852 21119 10854
rect 20811 10832 21119 10852
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 20732 9602 20760 9930
rect 20811 9820 21119 9840
rect 20811 9818 20817 9820
rect 20873 9818 20897 9820
rect 20953 9818 20977 9820
rect 21033 9818 21057 9820
rect 21113 9818 21119 9820
rect 20873 9766 20875 9818
rect 21055 9766 21057 9818
rect 20811 9764 20817 9766
rect 20873 9764 20897 9766
rect 20953 9764 20977 9766
rect 21033 9764 21057 9766
rect 21113 9764 21119 9766
rect 20811 9744 21119 9764
rect 20732 9574 20944 9602
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 20916 8974 20944 9574
rect 21192 9178 21220 9930
rect 21284 9382 21312 9998
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20364 8634 20392 8910
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20364 7410 20392 8570
rect 20444 8424 20496 8430
rect 20548 8401 20576 8910
rect 20444 8366 20496 8372
rect 20534 8392 20590 8401
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19904 4758 19932 5306
rect 19892 4752 19944 4758
rect 19892 4694 19944 4700
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19812 4146 19840 4558
rect 19996 4554 20024 5782
rect 20272 5778 20300 6258
rect 20456 5794 20484 8366
rect 20732 8362 20760 8910
rect 20811 8732 21119 8752
rect 20811 8730 20817 8732
rect 20873 8730 20897 8732
rect 20953 8730 20977 8732
rect 21033 8730 21057 8732
rect 21113 8730 21119 8732
rect 20873 8678 20875 8730
rect 21055 8678 21057 8730
rect 20811 8676 20817 8678
rect 20873 8676 20897 8678
rect 20953 8676 20977 8678
rect 21033 8676 21057 8678
rect 21113 8676 21119 8678
rect 20811 8656 21119 8676
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 20534 8327 20590 8336
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20536 8288 20588 8294
rect 20536 8230 20588 8236
rect 20548 7886 20576 8230
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20732 7426 20760 8298
rect 20811 7644 21119 7664
rect 20811 7642 20817 7644
rect 20873 7642 20897 7644
rect 20953 7642 20977 7644
rect 21033 7642 21057 7644
rect 21113 7642 21119 7644
rect 20873 7590 20875 7642
rect 21055 7590 21057 7642
rect 20811 7588 20817 7590
rect 20873 7588 20897 7590
rect 20953 7588 20977 7590
rect 21033 7588 21057 7590
rect 21113 7588 21119 7590
rect 20811 7568 21119 7588
rect 20732 7410 20944 7426
rect 20732 7404 20956 7410
rect 20732 7398 20904 7404
rect 20904 7346 20956 7352
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 20824 7206 20852 7278
rect 20812 7200 20864 7206
rect 20640 7160 20812 7188
rect 20640 6322 20668 7160
rect 20812 7142 20864 7148
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20732 5914 20760 6666
rect 20811 6556 21119 6576
rect 20811 6554 20817 6556
rect 20873 6554 20897 6556
rect 20953 6554 20977 6556
rect 21033 6554 21057 6556
rect 21113 6554 21119 6556
rect 20873 6502 20875 6554
rect 21055 6502 21057 6554
rect 20811 6500 20817 6502
rect 20873 6500 20897 6502
rect 20953 6500 20977 6502
rect 21033 6500 21057 6502
rect 21113 6500 21119 6502
rect 20811 6480 21119 6500
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20364 5778 20484 5794
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20364 5772 20496 5778
rect 20364 5766 20444 5772
rect 20364 5658 20392 5766
rect 20444 5714 20496 5720
rect 20272 5630 20392 5658
rect 20444 5636 20496 5642
rect 20272 4826 20300 5630
rect 20444 5578 20496 5584
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20272 4622 20300 4762
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 19996 4078 20024 4490
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 20088 4010 20116 4558
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20076 4004 20128 4010
rect 20076 3946 20128 3952
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19248 3460 19300 3466
rect 19248 3402 19300 3408
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19260 3058 19288 3402
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 17696 2650 17724 2790
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17696 2446 17724 2586
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16868 2106 16896 2246
rect 16856 2100 16908 2106
rect 16856 2042 16908 2048
rect 17132 1420 17184 1426
rect 17132 1362 17184 1368
rect 17144 800 17172 1362
rect 17880 800 17908 2450
rect 17960 2440 18012 2446
rect 18156 2428 18184 2790
rect 18012 2400 18184 2428
rect 18696 2440 18748 2446
rect 17960 2382 18012 2388
rect 18696 2382 18748 2388
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18340 2106 18368 2246
rect 18328 2100 18380 2106
rect 18328 2042 18380 2048
rect 18604 2100 18656 2106
rect 18604 2042 18656 2048
rect 18616 800 18644 2042
rect 18708 1426 18736 2382
rect 18984 2378 19012 2926
rect 18972 2372 19024 2378
rect 18972 2314 19024 2320
rect 18696 1420 18748 1426
rect 18696 1362 18748 1368
rect 19444 800 19472 3402
rect 20364 3126 20392 4082
rect 20456 3738 20484 5578
rect 20811 5468 21119 5488
rect 20811 5466 20817 5468
rect 20873 5466 20897 5468
rect 20953 5466 20977 5468
rect 21033 5466 21057 5468
rect 21113 5466 21119 5468
rect 20873 5414 20875 5466
rect 21055 5414 21057 5466
rect 20811 5412 20817 5414
rect 20873 5412 20897 5414
rect 20953 5412 20977 5414
rect 21033 5412 21057 5414
rect 21113 5412 21119 5414
rect 20811 5392 21119 5412
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20640 4826 20668 5170
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 20548 4078 20576 4490
rect 20811 4380 21119 4400
rect 20811 4378 20817 4380
rect 20873 4378 20897 4380
rect 20953 4378 20977 4380
rect 21033 4378 21057 4380
rect 21113 4378 21119 4380
rect 20873 4326 20875 4378
rect 21055 4326 21057 4378
rect 20811 4324 20817 4326
rect 20873 4324 20897 4326
rect 20953 4324 20977 4326
rect 21033 4324 21057 4326
rect 21113 4324 21119 4326
rect 20811 4304 21119 4324
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20628 4004 20680 4010
rect 20628 3946 20680 3952
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20352 3120 20404 3126
rect 20352 3062 20404 3068
rect 20456 2854 20484 3674
rect 20640 3058 20668 3946
rect 21192 3942 21220 8434
rect 21284 8362 21312 8978
rect 21376 8566 21404 11086
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 21284 7206 21312 8298
rect 21376 8090 21404 8502
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21284 5234 21312 6734
rect 21468 6662 21496 10610
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21560 9042 21588 9318
rect 21548 9036 21600 9042
rect 21548 8978 21600 8984
rect 21560 8480 21588 8978
rect 21652 8906 21680 12106
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22204 11762 22232 12038
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 25776 11452 26084 11472
rect 25776 11450 25782 11452
rect 25838 11450 25862 11452
rect 25918 11450 25942 11452
rect 25998 11450 26022 11452
rect 26078 11450 26084 11452
rect 25838 11398 25840 11450
rect 26020 11398 26022 11450
rect 25776 11396 25782 11398
rect 25838 11396 25862 11398
rect 25918 11396 25942 11398
rect 25998 11396 26022 11398
rect 26078 11396 26084 11398
rect 25776 11376 26084 11396
rect 25776 10364 26084 10384
rect 25776 10362 25782 10364
rect 25838 10362 25862 10364
rect 25918 10362 25942 10364
rect 25998 10362 26022 10364
rect 26078 10362 26084 10364
rect 25838 10310 25840 10362
rect 26020 10310 26022 10362
rect 25776 10308 25782 10310
rect 25838 10308 25862 10310
rect 25918 10308 25942 10310
rect 25998 10308 26022 10310
rect 26078 10308 26084 10310
rect 25776 10288 26084 10308
rect 28724 10260 28776 10266
rect 28724 10202 28776 10208
rect 25776 9276 26084 9296
rect 25776 9274 25782 9276
rect 25838 9274 25862 9276
rect 25918 9274 25942 9276
rect 25998 9274 26022 9276
rect 26078 9274 26084 9276
rect 25838 9222 25840 9274
rect 26020 9222 26022 9274
rect 25776 9220 25782 9222
rect 25838 9220 25862 9222
rect 25918 9220 25942 9222
rect 25998 9220 26022 9222
rect 26078 9220 26084 9222
rect 25776 9200 26084 9220
rect 21640 8900 21692 8906
rect 21640 8842 21692 8848
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21836 8634 21864 8842
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 22020 8498 22048 8774
rect 22008 8492 22060 8498
rect 21560 8452 21680 8480
rect 21652 7410 21680 8452
rect 22008 8434 22060 8440
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22204 8294 22232 8434
rect 22282 8392 22338 8401
rect 22282 8327 22338 8336
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21652 6798 21680 7346
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21468 5710 21496 6598
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 20916 3534 20944 3878
rect 21192 3754 21220 3878
rect 21100 3726 21220 3754
rect 21100 3534 21128 3726
rect 21284 3618 21312 5170
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 21192 3602 21312 3618
rect 21180 3596 21312 3602
rect 21232 3590 21312 3596
rect 21180 3538 21232 3544
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 21088 3528 21140 3534
rect 21140 3476 21220 3482
rect 21088 3470 21220 3476
rect 21100 3454 21220 3470
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 20732 2650 20760 3334
rect 20811 3292 21119 3312
rect 20811 3290 20817 3292
rect 20873 3290 20897 3292
rect 20953 3290 20977 3292
rect 21033 3290 21057 3292
rect 21113 3290 21119 3292
rect 20873 3238 20875 3290
rect 21055 3238 21057 3290
rect 20811 3236 20817 3238
rect 20873 3236 20897 3238
rect 20953 3236 20977 3238
rect 21033 3236 21057 3238
rect 21113 3236 21119 3238
rect 20811 3216 21119 3236
rect 21192 3058 21220 3454
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21284 3194 21312 3334
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21100 2650 21128 2790
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 21088 2644 21140 2650
rect 21088 2586 21140 2592
rect 20260 2576 20312 2582
rect 20260 2518 20312 2524
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 20180 1970 20208 2246
rect 20168 1964 20220 1970
rect 20168 1906 20220 1912
rect 20272 1306 20300 2518
rect 21192 2514 21220 2790
rect 21376 2774 21404 4082
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 21468 3602 21496 3946
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21560 3738 21588 3878
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 21456 3596 21508 3602
rect 21456 3538 21508 3544
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21836 3126 21864 3402
rect 22112 3194 22140 7142
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 21824 3120 21876 3126
rect 21824 3062 21876 3068
rect 21732 2984 21784 2990
rect 21732 2926 21784 2932
rect 21284 2746 21404 2774
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 20811 2204 21119 2224
rect 20811 2202 20817 2204
rect 20873 2202 20897 2204
rect 20953 2202 20977 2204
rect 21033 2202 21057 2204
rect 21113 2202 21119 2204
rect 20873 2150 20875 2202
rect 21055 2150 21057 2202
rect 20811 2148 20817 2150
rect 20873 2148 20897 2150
rect 20953 2148 20977 2150
rect 21033 2148 21057 2150
rect 21113 2148 21119 2150
rect 20811 2128 21119 2148
rect 20180 1278 20300 1306
rect 20180 800 20208 1278
rect 20916 870 21036 898
rect 20916 800 20944 870
rect 2962 368 3018 377
rect 2962 303 3018 312
rect 3422 0 3478 800
rect 4158 0 4214 800
rect 4894 0 4950 800
rect 5722 0 5778 800
rect 6458 0 6514 800
rect 7194 0 7250 800
rect 7930 0 7986 800
rect 8758 0 8814 800
rect 9494 0 9550 800
rect 10230 0 10286 800
rect 11058 0 11114 800
rect 11794 0 11850 800
rect 12530 0 12586 800
rect 13266 0 13322 800
rect 14094 0 14150 800
rect 14830 0 14886 800
rect 15566 0 15622 800
rect 16394 0 16450 800
rect 17130 0 17186 800
rect 17866 0 17922 800
rect 18602 0 18658 800
rect 19430 0 19486 800
rect 20166 0 20222 800
rect 20902 0 20958 800
rect 21008 762 21036 870
rect 21284 762 21312 2746
rect 21744 800 21772 2926
rect 21836 2514 21864 3062
rect 22112 3058 22140 3130
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 21928 2650 21956 2994
rect 22020 2922 22232 2938
rect 22008 2916 22232 2922
rect 22060 2910 22232 2916
rect 22008 2858 22060 2864
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 21824 2508 21876 2514
rect 21824 2450 21876 2456
rect 22204 2428 22232 2910
rect 22296 2854 22324 8327
rect 22388 3126 22416 8434
rect 25776 8188 26084 8208
rect 25776 8186 25782 8188
rect 25838 8186 25862 8188
rect 25918 8186 25942 8188
rect 25998 8186 26022 8188
rect 26078 8186 26084 8188
rect 25838 8134 25840 8186
rect 26020 8134 26022 8186
rect 25776 8132 25782 8134
rect 25838 8132 25862 8134
rect 25918 8132 25942 8134
rect 25998 8132 26022 8134
rect 26078 8132 26084 8134
rect 25776 8112 26084 8132
rect 25776 7100 26084 7120
rect 25776 7098 25782 7100
rect 25838 7098 25862 7100
rect 25918 7098 25942 7100
rect 25998 7098 26022 7100
rect 26078 7098 26084 7100
rect 25838 7046 25840 7098
rect 26020 7046 26022 7098
rect 25776 7044 25782 7046
rect 25838 7044 25862 7046
rect 25918 7044 25942 7046
rect 25998 7044 26022 7046
rect 26078 7044 26084 7046
rect 25776 7024 26084 7044
rect 25776 6012 26084 6032
rect 25776 6010 25782 6012
rect 25838 6010 25862 6012
rect 25918 6010 25942 6012
rect 25998 6010 26022 6012
rect 26078 6010 26084 6012
rect 25838 5958 25840 6010
rect 26020 5958 26022 6010
rect 25776 5956 25782 5958
rect 25838 5956 25862 5958
rect 25918 5956 25942 5958
rect 25998 5956 26022 5958
rect 26078 5956 26084 5958
rect 25776 5936 26084 5956
rect 25776 4924 26084 4944
rect 25776 4922 25782 4924
rect 25838 4922 25862 4924
rect 25918 4922 25942 4924
rect 25998 4922 26022 4924
rect 26078 4922 26084 4924
rect 25838 4870 25840 4922
rect 26020 4870 26022 4922
rect 25776 4868 25782 4870
rect 25838 4868 25862 4870
rect 25918 4868 25942 4870
rect 25998 4868 26022 4870
rect 26078 4868 26084 4870
rect 25776 4848 26084 4868
rect 25776 3836 26084 3856
rect 25776 3834 25782 3836
rect 25838 3834 25862 3836
rect 25918 3834 25942 3836
rect 25998 3834 26022 3836
rect 26078 3834 26084 3836
rect 25838 3782 25840 3834
rect 26020 3782 26022 3834
rect 25776 3780 25782 3782
rect 25838 3780 25862 3782
rect 25918 3780 25942 3782
rect 25998 3780 26022 3782
rect 26078 3780 26084 3782
rect 25776 3760 26084 3780
rect 22928 3664 22980 3670
rect 22928 3606 22980 3612
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22376 3120 22428 3126
rect 22376 3062 22428 3068
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 22284 2440 22336 2446
rect 22204 2400 22284 2428
rect 22284 2382 22336 2388
rect 22480 800 22508 3470
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22572 2650 22600 2994
rect 22940 2854 22968 3606
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 27804 3392 27856 3398
rect 27804 3334 27856 3340
rect 25044 3120 25096 3126
rect 25044 3062 25096 3068
rect 23204 3052 23256 3058
rect 23204 2994 23256 3000
rect 22928 2848 22980 2854
rect 22928 2790 22980 2796
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 22572 2310 22600 2586
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 22664 2310 22692 2382
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 22848 2106 22876 2382
rect 22836 2100 22888 2106
rect 22836 2042 22888 2048
rect 23216 800 23244 2994
rect 24400 2916 24452 2922
rect 24400 2858 24452 2864
rect 24412 2582 24440 2858
rect 25056 2582 25084 3062
rect 27160 3052 27212 3058
rect 27160 2994 27212 3000
rect 25776 2748 26084 2768
rect 25776 2746 25782 2748
rect 25838 2746 25862 2748
rect 25918 2746 25942 2748
rect 25998 2746 26022 2748
rect 26078 2746 26084 2748
rect 25838 2694 25840 2746
rect 26020 2694 26022 2746
rect 25776 2692 25782 2694
rect 25838 2692 25862 2694
rect 25918 2692 25942 2694
rect 25998 2692 26022 2694
rect 26078 2692 26084 2694
rect 25776 2672 26084 2692
rect 27172 2650 27200 2994
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 27632 2650 27660 2926
rect 27816 2854 27844 3334
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 27160 2644 27212 2650
rect 27160 2586 27212 2592
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 24400 2576 24452 2582
rect 24400 2518 24452 2524
rect 25044 2576 25096 2582
rect 25044 2518 25096 2524
rect 23296 2508 23348 2514
rect 23296 2450 23348 2456
rect 23308 2310 23336 2450
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 23952 800 23980 2382
rect 24780 800 24808 2382
rect 25516 800 25544 2382
rect 26252 800 26280 2382
rect 27080 800 27108 2382
rect 27908 1850 27936 3470
rect 27988 3392 28040 3398
rect 27988 3334 28040 3340
rect 28000 3126 28028 3334
rect 27988 3120 28040 3126
rect 27988 3062 28040 3068
rect 27816 1822 27936 1850
rect 27816 800 27844 1822
rect 28552 800 28580 3470
rect 28632 2848 28684 2854
rect 28632 2790 28684 2796
rect 28644 2378 28672 2790
rect 28736 2446 28764 10202
rect 29104 2446 29132 28358
rect 29748 28218 29776 29582
rect 30196 29164 30248 29170
rect 30196 29106 30248 29112
rect 29828 29028 29880 29034
rect 29828 28970 29880 28976
rect 30012 29028 30064 29034
rect 30012 28970 30064 28976
rect 29736 28212 29788 28218
rect 29564 28172 29736 28200
rect 29368 27464 29420 27470
rect 29368 27406 29420 27412
rect 29184 25288 29236 25294
rect 29184 25230 29236 25236
rect 29196 14890 29224 25230
rect 29276 18284 29328 18290
rect 29276 18226 29328 18232
rect 29184 14884 29236 14890
rect 29184 14826 29236 14832
rect 29288 13870 29316 18226
rect 29380 16250 29408 27406
rect 29460 23112 29512 23118
rect 29460 23054 29512 23060
rect 29368 16244 29420 16250
rect 29368 16186 29420 16192
rect 29472 15706 29500 23054
rect 29460 15700 29512 15706
rect 29460 15642 29512 15648
rect 29276 13864 29328 13870
rect 29276 13806 29328 13812
rect 29564 7410 29592 28172
rect 29736 28154 29788 28160
rect 29840 28082 29868 28970
rect 30024 28937 30052 28970
rect 30010 28928 30066 28937
rect 30010 28863 30066 28872
rect 29828 28076 29880 28082
rect 29828 28018 29880 28024
rect 29840 22094 29868 28018
rect 30012 27328 30064 27334
rect 30012 27270 30064 27276
rect 30024 27033 30052 27270
rect 30010 27024 30066 27033
rect 30010 26959 30066 26968
rect 30012 25152 30064 25158
rect 30012 25094 30064 25100
rect 30024 24993 30052 25094
rect 30010 24984 30066 24993
rect 30010 24919 30066 24928
rect 30012 22976 30064 22982
rect 30010 22944 30012 22953
rect 30064 22944 30066 22953
rect 30010 22879 30066 22888
rect 29748 22066 29868 22094
rect 29644 18760 29696 18766
rect 29644 18702 29696 18708
rect 29656 14482 29684 18702
rect 29644 14476 29696 14482
rect 29644 14418 29696 14424
rect 29552 7404 29604 7410
rect 29552 7346 29604 7352
rect 29748 5234 29776 22066
rect 29920 21548 29972 21554
rect 29920 21490 29972 21496
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 29840 18426 29868 19314
rect 29932 18970 29960 21490
rect 30012 21344 30064 21350
rect 30012 21286 30064 21292
rect 30024 21049 30052 21286
rect 30010 21040 30066 21049
rect 30010 20975 30066 20984
rect 30104 19440 30156 19446
rect 30104 19382 30156 19388
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 30024 19009 30052 19110
rect 30010 19000 30066 19009
rect 29920 18964 29972 18970
rect 30010 18935 30066 18944
rect 29920 18906 29972 18912
rect 30116 18766 30144 19382
rect 30104 18760 30156 18766
rect 30104 18702 30156 18708
rect 29828 18420 29880 18426
rect 29828 18362 29880 18368
rect 30116 18290 30144 18702
rect 30104 18284 30156 18290
rect 30104 18226 30156 18232
rect 29920 17196 29972 17202
rect 29920 17138 29972 17144
rect 29932 16574 29960 17138
rect 30012 16992 30064 16998
rect 30010 16960 30012 16969
rect 30064 16960 30066 16969
rect 30010 16895 30066 16904
rect 29840 16546 29960 16574
rect 29840 14074 29868 16546
rect 30116 16114 30144 18226
rect 30104 16108 30156 16114
rect 30104 16050 30156 16056
rect 30116 15502 30144 16050
rect 29920 15496 29972 15502
rect 29920 15438 29972 15444
rect 30104 15496 30156 15502
rect 30104 15438 30156 15444
rect 29932 15162 29960 15438
rect 29920 15156 29972 15162
rect 29920 15098 29972 15104
rect 29920 15020 29972 15026
rect 29920 14962 29972 14968
rect 29932 14618 29960 14962
rect 30116 14958 30144 15438
rect 30104 14952 30156 14958
rect 30010 14920 30066 14929
rect 30104 14894 30156 14900
rect 30010 14855 30012 14864
rect 30064 14855 30066 14864
rect 30012 14826 30064 14832
rect 29920 14612 29972 14618
rect 29920 14554 29972 14560
rect 30116 14414 30144 14894
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 29828 14068 29880 14074
rect 29828 14010 29880 14016
rect 30116 13938 30144 14350
rect 29920 13932 29972 13938
rect 29920 13874 29972 13880
rect 30104 13932 30156 13938
rect 30104 13874 30156 13880
rect 29932 13258 29960 13874
rect 30116 13326 30144 13874
rect 30104 13320 30156 13326
rect 30104 13262 30156 13268
rect 29920 13252 29972 13258
rect 29920 13194 29972 13200
rect 30012 13184 30064 13190
rect 30012 13126 30064 13132
rect 30024 13025 30052 13126
rect 30010 13016 30066 13025
rect 30010 12951 30066 12960
rect 30116 12850 30144 13262
rect 30208 12986 30236 29106
rect 30196 12980 30248 12986
rect 30196 12922 30248 12928
rect 29920 12844 29972 12850
rect 29920 12786 29972 12792
rect 30104 12844 30156 12850
rect 30104 12786 30156 12792
rect 29932 12306 29960 12786
rect 29920 12300 29972 12306
rect 29920 12242 29972 12248
rect 29828 11688 29880 11694
rect 29828 11630 29880 11636
rect 29840 11150 29868 11630
rect 29828 11144 29880 11150
rect 29828 11086 29880 11092
rect 29840 10418 29868 11086
rect 30012 11008 30064 11014
rect 30010 10976 30012 10985
rect 30064 10976 30066 10985
rect 30010 10911 30066 10920
rect 29840 10390 29960 10418
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 29840 8634 29868 8910
rect 29828 8628 29880 8634
rect 29828 8570 29880 8576
rect 29932 8498 29960 10390
rect 30010 8936 30066 8945
rect 30010 8871 30066 8880
rect 30024 8838 30052 8871
rect 30012 8832 30064 8838
rect 30012 8774 30064 8780
rect 29920 8492 29972 8498
rect 29920 8434 29972 8440
rect 30104 8492 30156 8498
rect 30104 8434 30156 8440
rect 30012 7200 30064 7206
rect 30012 7142 30064 7148
rect 30024 7041 30052 7142
rect 30010 7032 30066 7041
rect 30010 6967 30066 6976
rect 30116 6458 30144 8434
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 29736 5228 29788 5234
rect 29736 5170 29788 5176
rect 30012 5024 30064 5030
rect 30010 4992 30012 5001
rect 30064 4992 30066 5001
rect 30010 4927 30066 4936
rect 29644 4480 29696 4486
rect 29644 4422 29696 4428
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29276 3528 29328 3534
rect 29276 3470 29328 3476
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 29092 2440 29144 2446
rect 29092 2382 29144 2388
rect 28632 2372 28684 2378
rect 28632 2314 28684 2320
rect 28908 2304 28960 2310
rect 28908 2246 28960 2252
rect 28920 1057 28948 2246
rect 28906 1048 28962 1057
rect 28906 983 28962 992
rect 29288 800 29316 3470
rect 29564 3058 29592 3878
rect 29552 3052 29604 3058
rect 29552 2994 29604 3000
rect 29656 2854 29684 4422
rect 30104 4140 30156 4146
rect 30104 4082 30156 4088
rect 30012 3936 30064 3942
rect 30012 3878 30064 3884
rect 29920 3392 29972 3398
rect 29920 3334 29972 3340
rect 29932 3058 29960 3334
rect 30024 3058 30052 3878
rect 29920 3052 29972 3058
rect 29920 2994 29972 3000
rect 30012 3052 30064 3058
rect 30012 2994 30064 3000
rect 30010 2952 30066 2961
rect 30010 2887 30066 2896
rect 29644 2848 29696 2854
rect 29644 2790 29696 2796
rect 30024 2650 30052 2887
rect 30012 2644 30064 2650
rect 30012 2586 30064 2592
rect 30116 800 30144 4082
rect 31576 4072 31628 4078
rect 31576 4014 31628 4020
rect 30840 2848 30892 2854
rect 30840 2790 30892 2796
rect 30852 800 30880 2790
rect 31588 800 31616 4014
rect 21008 734 21312 762
rect 21730 0 21786 800
rect 22466 0 22522 800
rect 23202 0 23258 800
rect 23938 0 23994 800
rect 24766 0 24822 800
rect 25502 0 25558 800
rect 26238 0 26294 800
rect 27066 0 27122 800
rect 27802 0 27858 800
rect 28538 0 28594 800
rect 29274 0 29330 800
rect 30102 0 30158 800
rect 30838 0 30894 800
rect 31574 0 31630 800
<< via2 >>
rect 2778 47504 2834 47560
rect 1490 44512 1546 44568
rect 1490 43832 1546 43888
rect 1490 43016 1546 43072
rect 1398 42336 1454 42392
rect 1490 41656 1546 41712
rect 1398 40840 1454 40896
rect 1306 40160 1362 40216
rect 1490 39344 1546 39400
rect 1398 38664 1454 38720
rect 1490 36488 1546 36544
rect 1490 34992 1546 35048
rect 1490 32680 1546 32736
rect 1582 32000 1638 32056
rect 1490 31320 1546 31376
rect 1490 29028 1546 29064
rect 1490 29008 1492 29028
rect 1492 29008 1544 29028
rect 1544 29008 1546 29028
rect 2226 45348 2282 45384
rect 2226 45328 2228 45348
rect 2228 45328 2280 45348
rect 2280 45328 2282 45348
rect 30010 46960 30066 47016
rect 2870 46824 2926 46880
rect 2962 46008 3018 46064
rect 10886 45722 10942 45724
rect 10966 45722 11022 45724
rect 11046 45722 11102 45724
rect 11126 45722 11182 45724
rect 10886 45670 10932 45722
rect 10932 45670 10942 45722
rect 10966 45670 10996 45722
rect 10996 45670 11008 45722
rect 11008 45670 11022 45722
rect 11046 45670 11060 45722
rect 11060 45670 11072 45722
rect 11072 45670 11102 45722
rect 11126 45670 11136 45722
rect 11136 45670 11182 45722
rect 10886 45668 10942 45670
rect 10966 45668 11022 45670
rect 11046 45668 11102 45670
rect 11126 45668 11182 45670
rect 20817 45722 20873 45724
rect 20897 45722 20953 45724
rect 20977 45722 21033 45724
rect 21057 45722 21113 45724
rect 20817 45670 20863 45722
rect 20863 45670 20873 45722
rect 20897 45670 20927 45722
rect 20927 45670 20939 45722
rect 20939 45670 20953 45722
rect 20977 45670 20991 45722
rect 20991 45670 21003 45722
rect 21003 45670 21033 45722
rect 21057 45670 21067 45722
rect 21067 45670 21113 45722
rect 20817 45668 20873 45670
rect 20897 45668 20953 45670
rect 20977 45668 21033 45670
rect 21057 45668 21113 45670
rect 2410 44820 2412 44840
rect 2412 44820 2464 44840
rect 2464 44820 2466 44840
rect 2410 44784 2466 44820
rect 2226 35672 2282 35728
rect 4434 44532 4490 44568
rect 4434 44512 4436 44532
rect 4436 44512 4488 44532
rect 4488 44512 4490 44532
rect 3146 37848 3202 37904
rect 3146 37168 3202 37224
rect 3514 40568 3570 40624
rect 4250 40568 4306 40624
rect 4802 40588 4858 40624
rect 4802 40568 4804 40588
rect 4804 40568 4856 40588
rect 4856 40568 4858 40588
rect 5921 45178 5977 45180
rect 6001 45178 6057 45180
rect 6081 45178 6137 45180
rect 6161 45178 6217 45180
rect 5921 45126 5967 45178
rect 5967 45126 5977 45178
rect 6001 45126 6031 45178
rect 6031 45126 6043 45178
rect 6043 45126 6057 45178
rect 6081 45126 6095 45178
rect 6095 45126 6107 45178
rect 6107 45126 6137 45178
rect 6161 45126 6171 45178
rect 6171 45126 6217 45178
rect 5921 45124 5977 45126
rect 6001 45124 6057 45126
rect 6081 45124 6137 45126
rect 6161 45124 6217 45126
rect 3054 34176 3110 34232
rect 2962 33496 3018 33552
rect 5921 44090 5977 44092
rect 6001 44090 6057 44092
rect 6081 44090 6137 44092
rect 6161 44090 6217 44092
rect 5921 44038 5967 44090
rect 5967 44038 5977 44090
rect 6001 44038 6031 44090
rect 6031 44038 6043 44090
rect 6043 44038 6057 44090
rect 6081 44038 6095 44090
rect 6095 44038 6107 44090
rect 6107 44038 6137 44090
rect 6161 44038 6171 44090
rect 6171 44038 6217 44090
rect 5921 44036 5977 44038
rect 6001 44036 6057 44038
rect 6081 44036 6137 44038
rect 6161 44036 6217 44038
rect 15852 45178 15908 45180
rect 15932 45178 15988 45180
rect 16012 45178 16068 45180
rect 16092 45178 16148 45180
rect 15852 45126 15898 45178
rect 15898 45126 15908 45178
rect 15932 45126 15962 45178
rect 15962 45126 15974 45178
rect 15974 45126 15988 45178
rect 16012 45126 16026 45178
rect 16026 45126 16038 45178
rect 16038 45126 16068 45178
rect 16092 45126 16102 45178
rect 16102 45126 16148 45178
rect 15852 45124 15908 45126
rect 15932 45124 15988 45126
rect 16012 45124 16068 45126
rect 16092 45124 16148 45126
rect 25782 45178 25838 45180
rect 25862 45178 25918 45180
rect 25942 45178 25998 45180
rect 26022 45178 26078 45180
rect 25782 45126 25828 45178
rect 25828 45126 25838 45178
rect 25862 45126 25892 45178
rect 25892 45126 25904 45178
rect 25904 45126 25918 45178
rect 25942 45126 25956 45178
rect 25956 45126 25968 45178
rect 25968 45126 25998 45178
rect 26022 45126 26032 45178
rect 26032 45126 26078 45178
rect 25782 45124 25838 45126
rect 25862 45124 25918 45126
rect 25942 45124 25998 45126
rect 26022 45124 26078 45126
rect 5921 43002 5977 43004
rect 6001 43002 6057 43004
rect 6081 43002 6137 43004
rect 6161 43002 6217 43004
rect 5921 42950 5967 43002
rect 5967 42950 5977 43002
rect 6001 42950 6031 43002
rect 6031 42950 6043 43002
rect 6043 42950 6057 43002
rect 6081 42950 6095 43002
rect 6095 42950 6107 43002
rect 6107 42950 6137 43002
rect 6161 42950 6171 43002
rect 6171 42950 6217 43002
rect 5921 42948 5977 42950
rect 6001 42948 6057 42950
rect 6081 42948 6137 42950
rect 6161 42948 6217 42950
rect 5921 41914 5977 41916
rect 6001 41914 6057 41916
rect 6081 41914 6137 41916
rect 6161 41914 6217 41916
rect 5921 41862 5967 41914
rect 5967 41862 5977 41914
rect 6001 41862 6031 41914
rect 6031 41862 6043 41914
rect 6043 41862 6057 41914
rect 6081 41862 6095 41914
rect 6095 41862 6107 41914
rect 6107 41862 6137 41914
rect 6161 41862 6171 41914
rect 6171 41862 6217 41914
rect 5921 41860 5977 41862
rect 6001 41860 6057 41862
rect 6081 41860 6137 41862
rect 6161 41860 6217 41862
rect 5921 40826 5977 40828
rect 6001 40826 6057 40828
rect 6081 40826 6137 40828
rect 6161 40826 6217 40828
rect 5921 40774 5967 40826
rect 5967 40774 5977 40826
rect 6001 40774 6031 40826
rect 6031 40774 6043 40826
rect 6043 40774 6057 40826
rect 6081 40774 6095 40826
rect 6095 40774 6107 40826
rect 6107 40774 6137 40826
rect 6161 40774 6171 40826
rect 6171 40774 6217 40826
rect 5921 40772 5977 40774
rect 6001 40772 6057 40774
rect 6081 40772 6137 40774
rect 6161 40772 6217 40774
rect 2778 29824 2834 29880
rect 1490 28364 1492 28384
rect 1492 28364 1544 28384
rect 1544 28364 1546 28384
rect 1490 28328 1546 28364
rect 1490 27512 1546 27568
rect 1490 26852 1546 26888
rect 1490 26832 1492 26852
rect 1492 26832 1544 26852
rect 1544 26832 1546 26852
rect 1490 26188 1492 26208
rect 1492 26188 1544 26208
rect 1544 26188 1546 26208
rect 1490 26152 1546 26188
rect 1490 25336 1546 25392
rect 1490 24676 1546 24712
rect 1490 24656 1492 24676
rect 1492 24656 1544 24676
rect 1544 24656 1546 24676
rect 1490 23840 1546 23896
rect 1398 23160 1454 23216
rect 3974 30540 3976 30560
rect 3976 30540 4028 30560
rect 4028 30540 4030 30560
rect 3974 30504 4030 30540
rect 5921 39738 5977 39740
rect 6001 39738 6057 39740
rect 6081 39738 6137 39740
rect 6161 39738 6217 39740
rect 5921 39686 5967 39738
rect 5967 39686 5977 39738
rect 6001 39686 6031 39738
rect 6031 39686 6043 39738
rect 6043 39686 6057 39738
rect 6081 39686 6095 39738
rect 6095 39686 6107 39738
rect 6107 39686 6137 39738
rect 6161 39686 6171 39738
rect 6171 39686 6217 39738
rect 5921 39684 5977 39686
rect 6001 39684 6057 39686
rect 6081 39684 6137 39686
rect 6161 39684 6217 39686
rect 5921 38650 5977 38652
rect 6001 38650 6057 38652
rect 6081 38650 6137 38652
rect 6161 38650 6217 38652
rect 5921 38598 5967 38650
rect 5967 38598 5977 38650
rect 6001 38598 6031 38650
rect 6031 38598 6043 38650
rect 6043 38598 6057 38650
rect 6081 38598 6095 38650
rect 6095 38598 6107 38650
rect 6107 38598 6137 38650
rect 6161 38598 6171 38650
rect 6171 38598 6217 38650
rect 5921 38596 5977 38598
rect 6001 38596 6057 38598
rect 6081 38596 6137 38598
rect 6161 38596 6217 38598
rect 5921 37562 5977 37564
rect 6001 37562 6057 37564
rect 6081 37562 6137 37564
rect 6161 37562 6217 37564
rect 5921 37510 5967 37562
rect 5967 37510 5977 37562
rect 6001 37510 6031 37562
rect 6031 37510 6043 37562
rect 6043 37510 6057 37562
rect 6081 37510 6095 37562
rect 6095 37510 6107 37562
rect 6107 37510 6137 37562
rect 6161 37510 6171 37562
rect 6171 37510 6217 37562
rect 5921 37508 5977 37510
rect 6001 37508 6057 37510
rect 6081 37508 6137 37510
rect 6161 37508 6217 37510
rect 5921 36474 5977 36476
rect 6001 36474 6057 36476
rect 6081 36474 6137 36476
rect 6161 36474 6217 36476
rect 5921 36422 5967 36474
rect 5967 36422 5977 36474
rect 6001 36422 6031 36474
rect 6031 36422 6043 36474
rect 6043 36422 6057 36474
rect 6081 36422 6095 36474
rect 6095 36422 6107 36474
rect 6107 36422 6137 36474
rect 6161 36422 6171 36474
rect 6171 36422 6217 36474
rect 5921 36420 5977 36422
rect 6001 36420 6057 36422
rect 6081 36420 6137 36422
rect 6161 36420 6217 36422
rect 5921 35386 5977 35388
rect 6001 35386 6057 35388
rect 6081 35386 6137 35388
rect 6161 35386 6217 35388
rect 5921 35334 5967 35386
rect 5967 35334 5977 35386
rect 6001 35334 6031 35386
rect 6031 35334 6043 35386
rect 6043 35334 6057 35386
rect 6081 35334 6095 35386
rect 6095 35334 6107 35386
rect 6107 35334 6137 35386
rect 6161 35334 6171 35386
rect 6171 35334 6217 35386
rect 5921 35332 5977 35334
rect 6001 35332 6057 35334
rect 6081 35332 6137 35334
rect 6161 35332 6217 35334
rect 1214 14320 1270 14376
rect 1214 11328 1270 11384
rect 1214 5480 1270 5536
rect 1398 15816 1454 15872
rect 2042 22344 2098 22400
rect 1858 20984 1914 21040
rect 2962 21664 3018 21720
rect 2778 20168 2834 20224
rect 1398 13504 1454 13560
rect 1398 12824 1454 12880
rect 1398 12008 1454 12064
rect 3146 19488 3202 19544
rect 2962 18672 3018 18728
rect 2778 16496 2834 16552
rect 3238 16224 3294 16280
rect 3146 15000 3202 15056
rect 1398 10648 1454 10704
rect 1398 9152 1454 9208
rect 1398 8336 1454 8392
rect 1398 7656 1454 7712
rect 2318 9424 2374 9480
rect 2042 6840 2098 6896
rect 1398 4664 1454 4720
rect 1398 3984 1454 4040
rect 3054 9832 3110 9888
rect 4250 26324 4252 26344
rect 4252 26324 4304 26344
rect 4304 26324 4306 26344
rect 4250 26288 4306 26324
rect 4526 26288 4582 26344
rect 4158 24112 4214 24168
rect 4526 24148 4528 24168
rect 4528 24148 4580 24168
rect 4580 24148 4582 24168
rect 4526 24112 4582 24148
rect 3882 17992 3938 18048
rect 3974 17176 4030 17232
rect 2778 6160 2834 6216
rect 1858 2488 1914 2544
rect 3054 4004 3110 4040
rect 3054 3984 3056 4004
rect 3056 3984 3108 4004
rect 3108 3984 3110 4004
rect 2778 3168 2834 3224
rect 5078 15544 5134 15600
rect 4986 13932 5042 13968
rect 4986 13912 4988 13932
rect 4988 13912 5040 13932
rect 5040 13912 5042 13932
rect 6642 34584 6698 34640
rect 5921 34298 5977 34300
rect 6001 34298 6057 34300
rect 6081 34298 6137 34300
rect 6161 34298 6217 34300
rect 5921 34246 5967 34298
rect 5967 34246 5977 34298
rect 6001 34246 6031 34298
rect 6031 34246 6043 34298
rect 6043 34246 6057 34298
rect 6081 34246 6095 34298
rect 6095 34246 6107 34298
rect 6107 34246 6137 34298
rect 6161 34246 6171 34298
rect 6171 34246 6217 34298
rect 5921 34244 5977 34246
rect 6001 34244 6057 34246
rect 6081 34244 6137 34246
rect 6161 34244 6217 34246
rect 6182 34040 6238 34096
rect 5921 33210 5977 33212
rect 6001 33210 6057 33212
rect 6081 33210 6137 33212
rect 6161 33210 6217 33212
rect 5921 33158 5967 33210
rect 5967 33158 5977 33210
rect 6001 33158 6031 33210
rect 6031 33158 6043 33210
rect 6043 33158 6057 33210
rect 6081 33158 6095 33210
rect 6095 33158 6107 33210
rect 6107 33158 6137 33210
rect 6161 33158 6171 33210
rect 6171 33158 6217 33210
rect 5921 33156 5977 33158
rect 6001 33156 6057 33158
rect 6081 33156 6137 33158
rect 6161 33156 6217 33158
rect 5921 32122 5977 32124
rect 6001 32122 6057 32124
rect 6081 32122 6137 32124
rect 6161 32122 6217 32124
rect 5921 32070 5967 32122
rect 5967 32070 5977 32122
rect 6001 32070 6031 32122
rect 6031 32070 6043 32122
rect 6043 32070 6057 32122
rect 6081 32070 6095 32122
rect 6095 32070 6107 32122
rect 6107 32070 6137 32122
rect 6161 32070 6171 32122
rect 6171 32070 6217 32122
rect 5921 32068 5977 32070
rect 6001 32068 6057 32070
rect 6081 32068 6137 32070
rect 6161 32068 6217 32070
rect 5921 31034 5977 31036
rect 6001 31034 6057 31036
rect 6081 31034 6137 31036
rect 6161 31034 6217 31036
rect 5921 30982 5967 31034
rect 5967 30982 5977 31034
rect 6001 30982 6031 31034
rect 6031 30982 6043 31034
rect 6043 30982 6057 31034
rect 6081 30982 6095 31034
rect 6095 30982 6107 31034
rect 6107 30982 6137 31034
rect 6161 30982 6171 31034
rect 6171 30982 6217 31034
rect 5921 30980 5977 30982
rect 6001 30980 6057 30982
rect 6081 30980 6137 30982
rect 6161 30980 6217 30982
rect 5921 29946 5977 29948
rect 6001 29946 6057 29948
rect 6081 29946 6137 29948
rect 6161 29946 6217 29948
rect 5921 29894 5967 29946
rect 5967 29894 5977 29946
rect 6001 29894 6031 29946
rect 6031 29894 6043 29946
rect 6043 29894 6057 29946
rect 6081 29894 6095 29946
rect 6095 29894 6107 29946
rect 6107 29894 6137 29946
rect 6161 29894 6171 29946
rect 6171 29894 6217 29946
rect 5921 29892 5977 29894
rect 6001 29892 6057 29894
rect 6081 29892 6137 29894
rect 6161 29892 6217 29894
rect 8022 44784 8078 44840
rect 10886 44634 10942 44636
rect 10966 44634 11022 44636
rect 11046 44634 11102 44636
rect 11126 44634 11182 44636
rect 10886 44582 10932 44634
rect 10932 44582 10942 44634
rect 10966 44582 10996 44634
rect 10996 44582 11008 44634
rect 11008 44582 11022 44634
rect 11046 44582 11060 44634
rect 11060 44582 11072 44634
rect 11072 44582 11102 44634
rect 11126 44582 11136 44634
rect 11136 44582 11182 44634
rect 10886 44580 10942 44582
rect 10966 44580 11022 44582
rect 11046 44580 11102 44582
rect 11126 44580 11182 44582
rect 8206 44512 8262 44568
rect 20817 44634 20873 44636
rect 20897 44634 20953 44636
rect 20977 44634 21033 44636
rect 21057 44634 21113 44636
rect 20817 44582 20863 44634
rect 20863 44582 20873 44634
rect 20897 44582 20927 44634
rect 20927 44582 20939 44634
rect 20939 44582 20953 44634
rect 20977 44582 20991 44634
rect 20991 44582 21003 44634
rect 21003 44582 21033 44634
rect 21057 44582 21067 44634
rect 21067 44582 21113 44634
rect 20817 44580 20873 44582
rect 20897 44580 20953 44582
rect 20977 44580 21033 44582
rect 21057 44580 21113 44582
rect 5921 28858 5977 28860
rect 6001 28858 6057 28860
rect 6081 28858 6137 28860
rect 6161 28858 6217 28860
rect 5921 28806 5967 28858
rect 5967 28806 5977 28858
rect 6001 28806 6031 28858
rect 6031 28806 6043 28858
rect 6043 28806 6057 28858
rect 6081 28806 6095 28858
rect 6095 28806 6107 28858
rect 6107 28806 6137 28858
rect 6161 28806 6171 28858
rect 6171 28806 6217 28858
rect 5921 28804 5977 28806
rect 6001 28804 6057 28806
rect 6081 28804 6137 28806
rect 6161 28804 6217 28806
rect 5538 24148 5540 24168
rect 5540 24148 5592 24168
rect 5592 24148 5594 24168
rect 5538 24112 5594 24148
rect 5921 27770 5977 27772
rect 6001 27770 6057 27772
rect 6081 27770 6137 27772
rect 6161 27770 6217 27772
rect 5921 27718 5967 27770
rect 5967 27718 5977 27770
rect 6001 27718 6031 27770
rect 6031 27718 6043 27770
rect 6043 27718 6057 27770
rect 6081 27718 6095 27770
rect 6095 27718 6107 27770
rect 6107 27718 6137 27770
rect 6161 27718 6171 27770
rect 6171 27718 6217 27770
rect 5921 27716 5977 27718
rect 6001 27716 6057 27718
rect 6081 27716 6137 27718
rect 6161 27716 6217 27718
rect 5921 26682 5977 26684
rect 6001 26682 6057 26684
rect 6081 26682 6137 26684
rect 6161 26682 6217 26684
rect 5921 26630 5967 26682
rect 5967 26630 5977 26682
rect 6001 26630 6031 26682
rect 6031 26630 6043 26682
rect 6043 26630 6057 26682
rect 6081 26630 6095 26682
rect 6095 26630 6107 26682
rect 6107 26630 6137 26682
rect 6161 26630 6171 26682
rect 6171 26630 6217 26682
rect 5921 26628 5977 26630
rect 6001 26628 6057 26630
rect 6081 26628 6137 26630
rect 6161 26628 6217 26630
rect 5921 25594 5977 25596
rect 6001 25594 6057 25596
rect 6081 25594 6137 25596
rect 6161 25594 6217 25596
rect 5921 25542 5967 25594
rect 5967 25542 5977 25594
rect 6001 25542 6031 25594
rect 6031 25542 6043 25594
rect 6043 25542 6057 25594
rect 6081 25542 6095 25594
rect 6095 25542 6107 25594
rect 6107 25542 6137 25594
rect 6161 25542 6171 25594
rect 6171 25542 6217 25594
rect 5921 25540 5977 25542
rect 6001 25540 6057 25542
rect 6081 25540 6137 25542
rect 6161 25540 6217 25542
rect 5921 24506 5977 24508
rect 6001 24506 6057 24508
rect 6081 24506 6137 24508
rect 6161 24506 6217 24508
rect 5921 24454 5967 24506
rect 5967 24454 5977 24506
rect 6001 24454 6031 24506
rect 6031 24454 6043 24506
rect 6043 24454 6057 24506
rect 6081 24454 6095 24506
rect 6095 24454 6107 24506
rect 6107 24454 6137 24506
rect 6161 24454 6171 24506
rect 6171 24454 6217 24506
rect 5921 24452 5977 24454
rect 6001 24452 6057 24454
rect 6081 24452 6137 24454
rect 6161 24452 6217 24454
rect 5921 23418 5977 23420
rect 6001 23418 6057 23420
rect 6081 23418 6137 23420
rect 6161 23418 6217 23420
rect 5921 23366 5967 23418
rect 5967 23366 5977 23418
rect 6001 23366 6031 23418
rect 6031 23366 6043 23418
rect 6043 23366 6057 23418
rect 6081 23366 6095 23418
rect 6095 23366 6107 23418
rect 6107 23366 6137 23418
rect 6161 23366 6171 23418
rect 6171 23366 6217 23418
rect 5921 23364 5977 23366
rect 6001 23364 6057 23366
rect 6081 23364 6137 23366
rect 6161 23364 6217 23366
rect 5921 22330 5977 22332
rect 6001 22330 6057 22332
rect 6081 22330 6137 22332
rect 6161 22330 6217 22332
rect 5921 22278 5967 22330
rect 5967 22278 5977 22330
rect 6001 22278 6031 22330
rect 6031 22278 6043 22330
rect 6043 22278 6057 22330
rect 6081 22278 6095 22330
rect 6095 22278 6107 22330
rect 6107 22278 6137 22330
rect 6161 22278 6171 22330
rect 6171 22278 6217 22330
rect 5921 22276 5977 22278
rect 6001 22276 6057 22278
rect 6081 22276 6137 22278
rect 6161 22276 6217 22278
rect 5921 21242 5977 21244
rect 6001 21242 6057 21244
rect 6081 21242 6137 21244
rect 6161 21242 6217 21244
rect 5921 21190 5967 21242
rect 5967 21190 5977 21242
rect 6001 21190 6031 21242
rect 6031 21190 6043 21242
rect 6043 21190 6057 21242
rect 6081 21190 6095 21242
rect 6095 21190 6107 21242
rect 6107 21190 6137 21242
rect 6161 21190 6171 21242
rect 6171 21190 6217 21242
rect 5921 21188 5977 21190
rect 6001 21188 6057 21190
rect 6081 21188 6137 21190
rect 6161 21188 6217 21190
rect 5921 20154 5977 20156
rect 6001 20154 6057 20156
rect 6081 20154 6137 20156
rect 6161 20154 6217 20156
rect 5921 20102 5967 20154
rect 5967 20102 5977 20154
rect 6001 20102 6031 20154
rect 6031 20102 6043 20154
rect 6043 20102 6057 20154
rect 6081 20102 6095 20154
rect 6095 20102 6107 20154
rect 6107 20102 6137 20154
rect 6161 20102 6171 20154
rect 6171 20102 6217 20154
rect 5921 20100 5977 20102
rect 6001 20100 6057 20102
rect 6081 20100 6137 20102
rect 6161 20100 6217 20102
rect 5921 19066 5977 19068
rect 6001 19066 6057 19068
rect 6081 19066 6137 19068
rect 6161 19066 6217 19068
rect 5921 19014 5967 19066
rect 5967 19014 5977 19066
rect 6001 19014 6031 19066
rect 6031 19014 6043 19066
rect 6043 19014 6057 19066
rect 6081 19014 6095 19066
rect 6095 19014 6107 19066
rect 6107 19014 6137 19066
rect 6161 19014 6171 19066
rect 6171 19014 6217 19066
rect 5921 19012 5977 19014
rect 6001 19012 6057 19014
rect 6081 19012 6137 19014
rect 6161 19012 6217 19014
rect 5921 17978 5977 17980
rect 6001 17978 6057 17980
rect 6081 17978 6137 17980
rect 6161 17978 6217 17980
rect 5921 17926 5967 17978
rect 5967 17926 5977 17978
rect 6001 17926 6031 17978
rect 6031 17926 6043 17978
rect 6043 17926 6057 17978
rect 6081 17926 6095 17978
rect 6095 17926 6107 17978
rect 6107 17926 6137 17978
rect 6161 17926 6171 17978
rect 6171 17926 6217 17978
rect 5921 17924 5977 17926
rect 6001 17924 6057 17926
rect 6081 17924 6137 17926
rect 6161 17924 6217 17926
rect 5921 16890 5977 16892
rect 6001 16890 6057 16892
rect 6081 16890 6137 16892
rect 6161 16890 6217 16892
rect 5921 16838 5967 16890
rect 5967 16838 5977 16890
rect 6001 16838 6031 16890
rect 6031 16838 6043 16890
rect 6043 16838 6057 16890
rect 6081 16838 6095 16890
rect 6095 16838 6107 16890
rect 6107 16838 6137 16890
rect 6161 16838 6171 16890
rect 6171 16838 6217 16890
rect 5921 16836 5977 16838
rect 6001 16836 6057 16838
rect 6081 16836 6137 16838
rect 6161 16836 6217 16838
rect 5921 15802 5977 15804
rect 6001 15802 6057 15804
rect 6081 15802 6137 15804
rect 6161 15802 6217 15804
rect 5921 15750 5967 15802
rect 5967 15750 5977 15802
rect 6001 15750 6031 15802
rect 6031 15750 6043 15802
rect 6043 15750 6057 15802
rect 6081 15750 6095 15802
rect 6095 15750 6107 15802
rect 6107 15750 6137 15802
rect 6161 15750 6171 15802
rect 6171 15750 6217 15802
rect 5921 15748 5977 15750
rect 6001 15748 6057 15750
rect 6081 15748 6137 15750
rect 6161 15748 6217 15750
rect 5446 9560 5502 9616
rect 6182 15544 6238 15600
rect 5921 14714 5977 14716
rect 6001 14714 6057 14716
rect 6081 14714 6137 14716
rect 6161 14714 6217 14716
rect 5921 14662 5967 14714
rect 5967 14662 5977 14714
rect 6001 14662 6031 14714
rect 6031 14662 6043 14714
rect 6043 14662 6057 14714
rect 6081 14662 6095 14714
rect 6095 14662 6107 14714
rect 6107 14662 6137 14714
rect 6161 14662 6171 14714
rect 6171 14662 6217 14714
rect 5921 14660 5977 14662
rect 6001 14660 6057 14662
rect 6081 14660 6137 14662
rect 6161 14660 6217 14662
rect 5906 14320 5962 14376
rect 5921 13626 5977 13628
rect 6001 13626 6057 13628
rect 6081 13626 6137 13628
rect 6161 13626 6217 13628
rect 5921 13574 5967 13626
rect 5967 13574 5977 13626
rect 6001 13574 6031 13626
rect 6031 13574 6043 13626
rect 6043 13574 6057 13626
rect 6081 13574 6095 13626
rect 6095 13574 6107 13626
rect 6107 13574 6137 13626
rect 6161 13574 6171 13626
rect 6171 13574 6217 13626
rect 5921 13572 5977 13574
rect 6001 13572 6057 13574
rect 6081 13572 6137 13574
rect 6161 13572 6217 13574
rect 5921 12538 5977 12540
rect 6001 12538 6057 12540
rect 6081 12538 6137 12540
rect 6161 12538 6217 12540
rect 5921 12486 5967 12538
rect 5967 12486 5977 12538
rect 6001 12486 6031 12538
rect 6031 12486 6043 12538
rect 6043 12486 6057 12538
rect 6081 12486 6095 12538
rect 6095 12486 6107 12538
rect 6107 12486 6137 12538
rect 6161 12486 6171 12538
rect 6171 12486 6217 12538
rect 5921 12484 5977 12486
rect 6001 12484 6057 12486
rect 6081 12484 6137 12486
rect 6161 12484 6217 12486
rect 5921 11450 5977 11452
rect 6001 11450 6057 11452
rect 6081 11450 6137 11452
rect 6161 11450 6217 11452
rect 5921 11398 5967 11450
rect 5967 11398 5977 11450
rect 6001 11398 6031 11450
rect 6031 11398 6043 11450
rect 6043 11398 6057 11450
rect 6081 11398 6095 11450
rect 6095 11398 6107 11450
rect 6107 11398 6137 11450
rect 6161 11398 6171 11450
rect 6171 11398 6217 11450
rect 5921 11396 5977 11398
rect 6001 11396 6057 11398
rect 6081 11396 6137 11398
rect 6161 11396 6217 11398
rect 5921 10362 5977 10364
rect 6001 10362 6057 10364
rect 6081 10362 6137 10364
rect 6161 10362 6217 10364
rect 5921 10310 5967 10362
rect 5967 10310 5977 10362
rect 6001 10310 6031 10362
rect 6031 10310 6043 10362
rect 6043 10310 6057 10362
rect 6081 10310 6095 10362
rect 6095 10310 6107 10362
rect 6107 10310 6137 10362
rect 6161 10310 6171 10362
rect 6171 10310 6217 10362
rect 5921 10308 5977 10310
rect 6001 10308 6057 10310
rect 6081 10308 6137 10310
rect 6161 10308 6217 10310
rect 5906 9560 5962 9616
rect 6182 9424 6238 9480
rect 5921 9274 5977 9276
rect 6001 9274 6057 9276
rect 6081 9274 6137 9276
rect 6161 9274 6217 9276
rect 5921 9222 5967 9274
rect 5967 9222 5977 9274
rect 6001 9222 6031 9274
rect 6031 9222 6043 9274
rect 6043 9222 6057 9274
rect 6081 9222 6095 9274
rect 6095 9222 6107 9274
rect 6107 9222 6137 9274
rect 6161 9222 6171 9274
rect 6171 9222 6217 9274
rect 5921 9220 5977 9222
rect 6001 9220 6057 9222
rect 6081 9220 6137 9222
rect 6161 9220 6217 9222
rect 5921 8186 5977 8188
rect 6001 8186 6057 8188
rect 6081 8186 6137 8188
rect 6161 8186 6217 8188
rect 5921 8134 5967 8186
rect 5967 8134 5977 8186
rect 6001 8134 6031 8186
rect 6031 8134 6043 8186
rect 6043 8134 6057 8186
rect 6081 8134 6095 8186
rect 6095 8134 6107 8186
rect 6107 8134 6137 8186
rect 6161 8134 6171 8186
rect 6171 8134 6217 8186
rect 5921 8132 5977 8134
rect 6001 8132 6057 8134
rect 6081 8132 6137 8134
rect 6161 8132 6217 8134
rect 5921 7098 5977 7100
rect 6001 7098 6057 7100
rect 6081 7098 6137 7100
rect 6161 7098 6217 7100
rect 5921 7046 5967 7098
rect 5967 7046 5977 7098
rect 6001 7046 6031 7098
rect 6031 7046 6043 7098
rect 6043 7046 6057 7098
rect 6081 7046 6095 7098
rect 6095 7046 6107 7098
rect 6107 7046 6137 7098
rect 6161 7046 6171 7098
rect 6171 7046 6217 7098
rect 5921 7044 5977 7046
rect 6001 7044 6057 7046
rect 6081 7044 6137 7046
rect 6161 7044 6217 7046
rect 6090 6316 6146 6352
rect 6090 6296 6092 6316
rect 6092 6296 6144 6316
rect 6144 6296 6146 6316
rect 5921 6010 5977 6012
rect 6001 6010 6057 6012
rect 6081 6010 6137 6012
rect 6161 6010 6217 6012
rect 5921 5958 5967 6010
rect 5967 5958 5977 6010
rect 6001 5958 6031 6010
rect 6031 5958 6043 6010
rect 6043 5958 6057 6010
rect 6081 5958 6095 6010
rect 6095 5958 6107 6010
rect 6107 5958 6137 6010
rect 6161 5958 6171 6010
rect 6171 5958 6217 6010
rect 5921 5956 5977 5958
rect 6001 5956 6057 5958
rect 6081 5956 6137 5958
rect 6161 5956 6217 5958
rect 6918 14476 6974 14512
rect 6918 14456 6920 14476
rect 6920 14456 6972 14476
rect 6972 14456 6974 14476
rect 8298 34076 8300 34096
rect 8300 34076 8352 34096
rect 8352 34076 8354 34096
rect 8298 34040 8354 34076
rect 8942 34604 8998 34640
rect 8942 34584 8944 34604
rect 8944 34584 8996 34604
rect 8996 34584 8998 34604
rect 15852 44090 15908 44092
rect 15932 44090 15988 44092
rect 16012 44090 16068 44092
rect 16092 44090 16148 44092
rect 15852 44038 15898 44090
rect 15898 44038 15908 44090
rect 15932 44038 15962 44090
rect 15962 44038 15974 44090
rect 15974 44038 15988 44090
rect 16012 44038 16026 44090
rect 16026 44038 16038 44090
rect 16038 44038 16068 44090
rect 16092 44038 16102 44090
rect 16102 44038 16148 44090
rect 15852 44036 15908 44038
rect 15932 44036 15988 44038
rect 16012 44036 16068 44038
rect 16092 44036 16148 44038
rect 25782 44090 25838 44092
rect 25862 44090 25918 44092
rect 25942 44090 25998 44092
rect 26022 44090 26078 44092
rect 25782 44038 25828 44090
rect 25828 44038 25838 44090
rect 25862 44038 25892 44090
rect 25892 44038 25904 44090
rect 25904 44038 25918 44090
rect 25942 44038 25956 44090
rect 25956 44038 25968 44090
rect 25968 44038 25998 44090
rect 26022 44038 26032 44090
rect 26032 44038 26078 44090
rect 25782 44036 25838 44038
rect 25862 44036 25918 44038
rect 25942 44036 25998 44038
rect 26022 44036 26078 44038
rect 30102 44920 30158 44976
rect 10886 43546 10942 43548
rect 10966 43546 11022 43548
rect 11046 43546 11102 43548
rect 11126 43546 11182 43548
rect 10886 43494 10932 43546
rect 10932 43494 10942 43546
rect 10966 43494 10996 43546
rect 10996 43494 11008 43546
rect 11008 43494 11022 43546
rect 11046 43494 11060 43546
rect 11060 43494 11072 43546
rect 11072 43494 11102 43546
rect 11126 43494 11136 43546
rect 11136 43494 11182 43546
rect 10886 43492 10942 43494
rect 10966 43492 11022 43494
rect 11046 43492 11102 43494
rect 11126 43492 11182 43494
rect 15852 43002 15908 43004
rect 15932 43002 15988 43004
rect 16012 43002 16068 43004
rect 16092 43002 16148 43004
rect 15852 42950 15898 43002
rect 15898 42950 15908 43002
rect 15932 42950 15962 43002
rect 15962 42950 15974 43002
rect 15974 42950 15988 43002
rect 16012 42950 16026 43002
rect 16026 42950 16038 43002
rect 16038 42950 16068 43002
rect 16092 42950 16102 43002
rect 16102 42950 16148 43002
rect 15852 42948 15908 42950
rect 15932 42948 15988 42950
rect 16012 42948 16068 42950
rect 16092 42948 16148 42950
rect 20817 43546 20873 43548
rect 20897 43546 20953 43548
rect 20977 43546 21033 43548
rect 21057 43546 21113 43548
rect 20817 43494 20863 43546
rect 20863 43494 20873 43546
rect 20897 43494 20927 43546
rect 20927 43494 20939 43546
rect 20939 43494 20953 43546
rect 20977 43494 20991 43546
rect 20991 43494 21003 43546
rect 21003 43494 21033 43546
rect 21057 43494 21067 43546
rect 21067 43494 21113 43546
rect 20817 43492 20873 43494
rect 20897 43492 20953 43494
rect 20977 43492 21033 43494
rect 21057 43492 21113 43494
rect 25782 43002 25838 43004
rect 25862 43002 25918 43004
rect 25942 43002 25998 43004
rect 26022 43002 26078 43004
rect 25782 42950 25828 43002
rect 25828 42950 25838 43002
rect 25862 42950 25892 43002
rect 25892 42950 25904 43002
rect 25904 42950 25918 43002
rect 25942 42950 25956 43002
rect 25956 42950 25968 43002
rect 25968 42950 25998 43002
rect 26022 42950 26032 43002
rect 26032 42950 26078 43002
rect 25782 42948 25838 42950
rect 25862 42948 25918 42950
rect 25942 42948 25998 42950
rect 26022 42948 26078 42950
rect 30102 42880 30158 42936
rect 10886 42458 10942 42460
rect 10966 42458 11022 42460
rect 11046 42458 11102 42460
rect 11126 42458 11182 42460
rect 10886 42406 10932 42458
rect 10932 42406 10942 42458
rect 10966 42406 10996 42458
rect 10996 42406 11008 42458
rect 11008 42406 11022 42458
rect 11046 42406 11060 42458
rect 11060 42406 11072 42458
rect 11072 42406 11102 42458
rect 11126 42406 11136 42458
rect 11136 42406 11182 42458
rect 10886 42404 10942 42406
rect 10966 42404 11022 42406
rect 11046 42404 11102 42406
rect 11126 42404 11182 42406
rect 15852 41914 15908 41916
rect 15932 41914 15988 41916
rect 16012 41914 16068 41916
rect 16092 41914 16148 41916
rect 15852 41862 15898 41914
rect 15898 41862 15908 41914
rect 15932 41862 15962 41914
rect 15962 41862 15974 41914
rect 15974 41862 15988 41914
rect 16012 41862 16026 41914
rect 16026 41862 16038 41914
rect 16038 41862 16068 41914
rect 16092 41862 16102 41914
rect 16102 41862 16148 41914
rect 15852 41860 15908 41862
rect 15932 41860 15988 41862
rect 16012 41860 16068 41862
rect 16092 41860 16148 41862
rect 10886 41370 10942 41372
rect 10966 41370 11022 41372
rect 11046 41370 11102 41372
rect 11126 41370 11182 41372
rect 10886 41318 10932 41370
rect 10932 41318 10942 41370
rect 10966 41318 10996 41370
rect 10996 41318 11008 41370
rect 11008 41318 11022 41370
rect 11046 41318 11060 41370
rect 11060 41318 11072 41370
rect 11072 41318 11102 41370
rect 11126 41318 11136 41370
rect 11136 41318 11182 41370
rect 10886 41316 10942 41318
rect 10966 41316 11022 41318
rect 11046 41316 11102 41318
rect 11126 41316 11182 41318
rect 15852 40826 15908 40828
rect 15932 40826 15988 40828
rect 16012 40826 16068 40828
rect 16092 40826 16148 40828
rect 15852 40774 15898 40826
rect 15898 40774 15908 40826
rect 15932 40774 15962 40826
rect 15962 40774 15974 40826
rect 15974 40774 15988 40826
rect 16012 40774 16026 40826
rect 16026 40774 16038 40826
rect 16038 40774 16068 40826
rect 16092 40774 16102 40826
rect 16102 40774 16148 40826
rect 15852 40772 15908 40774
rect 15932 40772 15988 40774
rect 16012 40772 16068 40774
rect 16092 40772 16148 40774
rect 10886 40282 10942 40284
rect 10966 40282 11022 40284
rect 11046 40282 11102 40284
rect 11126 40282 11182 40284
rect 10886 40230 10932 40282
rect 10932 40230 10942 40282
rect 10966 40230 10996 40282
rect 10996 40230 11008 40282
rect 11008 40230 11022 40282
rect 11046 40230 11060 40282
rect 11060 40230 11072 40282
rect 11072 40230 11102 40282
rect 11126 40230 11136 40282
rect 11136 40230 11182 40282
rect 10886 40228 10942 40230
rect 10966 40228 11022 40230
rect 11046 40228 11102 40230
rect 11126 40228 11182 40230
rect 10886 39194 10942 39196
rect 10966 39194 11022 39196
rect 11046 39194 11102 39196
rect 11126 39194 11182 39196
rect 10886 39142 10932 39194
rect 10932 39142 10942 39194
rect 10966 39142 10996 39194
rect 10996 39142 11008 39194
rect 11008 39142 11022 39194
rect 11046 39142 11060 39194
rect 11060 39142 11072 39194
rect 11072 39142 11102 39194
rect 11126 39142 11136 39194
rect 11136 39142 11182 39194
rect 10886 39140 10942 39142
rect 10966 39140 11022 39142
rect 11046 39140 11102 39142
rect 11126 39140 11182 39142
rect 10886 38106 10942 38108
rect 10966 38106 11022 38108
rect 11046 38106 11102 38108
rect 11126 38106 11182 38108
rect 10886 38054 10932 38106
rect 10932 38054 10942 38106
rect 10966 38054 10996 38106
rect 10996 38054 11008 38106
rect 11008 38054 11022 38106
rect 11046 38054 11060 38106
rect 11060 38054 11072 38106
rect 11072 38054 11102 38106
rect 11126 38054 11136 38106
rect 11136 38054 11182 38106
rect 10886 38052 10942 38054
rect 10966 38052 11022 38054
rect 11046 38052 11102 38054
rect 11126 38052 11182 38054
rect 10886 37018 10942 37020
rect 10966 37018 11022 37020
rect 11046 37018 11102 37020
rect 11126 37018 11182 37020
rect 10886 36966 10932 37018
rect 10932 36966 10942 37018
rect 10966 36966 10996 37018
rect 10996 36966 11008 37018
rect 11008 36966 11022 37018
rect 11046 36966 11060 37018
rect 11060 36966 11072 37018
rect 11072 36966 11102 37018
rect 11126 36966 11136 37018
rect 11136 36966 11182 37018
rect 10886 36964 10942 36966
rect 10966 36964 11022 36966
rect 11046 36964 11102 36966
rect 11126 36964 11182 36966
rect 10046 33396 10048 33416
rect 10048 33396 10100 33416
rect 10100 33396 10102 33416
rect 10046 33360 10102 33396
rect 7930 27648 7986 27704
rect 7930 21936 7986 21992
rect 7838 21836 7840 21856
rect 7840 21836 7892 21856
rect 7892 21836 7894 21856
rect 7838 21800 7894 21836
rect 7838 21664 7894 21720
rect 8114 22208 8170 22264
rect 7194 16244 7250 16280
rect 7194 16224 7196 16244
rect 7196 16224 7248 16244
rect 7248 16224 7250 16244
rect 6826 13932 6882 13968
rect 6826 13912 6828 13932
rect 6828 13912 6880 13932
rect 6880 13912 6882 13932
rect 7102 14320 7158 14376
rect 5921 4922 5977 4924
rect 6001 4922 6057 4924
rect 6081 4922 6137 4924
rect 6161 4922 6217 4924
rect 5921 4870 5967 4922
rect 5967 4870 5977 4922
rect 6001 4870 6031 4922
rect 6031 4870 6043 4922
rect 6043 4870 6057 4922
rect 6081 4870 6095 4922
rect 6095 4870 6107 4922
rect 6107 4870 6137 4922
rect 6161 4870 6171 4922
rect 6171 4870 6217 4922
rect 5921 4868 5977 4870
rect 6001 4868 6057 4870
rect 6081 4868 6137 4870
rect 6161 4868 6217 4870
rect 8206 21684 8262 21720
rect 8206 21664 8208 21684
rect 8208 21664 8260 21684
rect 8260 21664 8262 21684
rect 8666 27512 8722 27568
rect 8666 26288 8722 26344
rect 8574 22072 8630 22128
rect 10886 35930 10942 35932
rect 10966 35930 11022 35932
rect 11046 35930 11102 35932
rect 11126 35930 11182 35932
rect 10886 35878 10932 35930
rect 10932 35878 10942 35930
rect 10966 35878 10996 35930
rect 10996 35878 11008 35930
rect 11008 35878 11022 35930
rect 11046 35878 11060 35930
rect 11060 35878 11072 35930
rect 11072 35878 11102 35930
rect 11126 35878 11136 35930
rect 11136 35878 11182 35930
rect 10886 35876 10942 35878
rect 10966 35876 11022 35878
rect 11046 35876 11102 35878
rect 11126 35876 11182 35878
rect 10886 34842 10942 34844
rect 10966 34842 11022 34844
rect 11046 34842 11102 34844
rect 11126 34842 11182 34844
rect 10886 34790 10932 34842
rect 10932 34790 10942 34842
rect 10966 34790 10996 34842
rect 10996 34790 11008 34842
rect 11008 34790 11022 34842
rect 11046 34790 11060 34842
rect 11060 34790 11072 34842
rect 11072 34790 11102 34842
rect 11126 34790 11136 34842
rect 11136 34790 11182 34842
rect 10886 34788 10942 34790
rect 10966 34788 11022 34790
rect 11046 34788 11102 34790
rect 11126 34788 11182 34790
rect 10886 33754 10942 33756
rect 10966 33754 11022 33756
rect 11046 33754 11102 33756
rect 11126 33754 11182 33756
rect 10886 33702 10932 33754
rect 10932 33702 10942 33754
rect 10966 33702 10996 33754
rect 10996 33702 11008 33754
rect 11008 33702 11022 33754
rect 11046 33702 11060 33754
rect 11060 33702 11072 33754
rect 11072 33702 11102 33754
rect 11126 33702 11136 33754
rect 11136 33702 11182 33754
rect 10886 33700 10942 33702
rect 10966 33700 11022 33702
rect 11046 33700 11102 33702
rect 11126 33700 11182 33702
rect 8942 26424 8998 26480
rect 9494 27648 9550 27704
rect 9402 22616 9458 22672
rect 9034 22072 9090 22128
rect 9402 21800 9458 21856
rect 9586 21664 9642 21720
rect 9494 21548 9550 21584
rect 9494 21528 9496 21548
rect 9496 21528 9548 21548
rect 9548 21528 9550 21548
rect 9586 21392 9642 21448
rect 9402 21120 9458 21176
rect 9126 15444 9128 15464
rect 9128 15444 9180 15464
rect 9180 15444 9182 15464
rect 9126 15408 9182 15444
rect 6918 6296 6974 6352
rect 2778 1672 2834 1728
rect 2870 992 2926 1048
rect 5814 4020 5816 4040
rect 5816 4020 5868 4040
rect 5868 4020 5870 4040
rect 5814 3984 5870 4020
rect 5921 3834 5977 3836
rect 6001 3834 6057 3836
rect 6081 3834 6137 3836
rect 6161 3834 6217 3836
rect 5921 3782 5967 3834
rect 5967 3782 5977 3834
rect 6001 3782 6031 3834
rect 6031 3782 6043 3834
rect 6043 3782 6057 3834
rect 6081 3782 6095 3834
rect 6095 3782 6107 3834
rect 6107 3782 6137 3834
rect 6161 3782 6171 3834
rect 6171 3782 6217 3834
rect 5921 3780 5977 3782
rect 6001 3780 6057 3782
rect 6081 3780 6137 3782
rect 6161 3780 6217 3782
rect 5921 2746 5977 2748
rect 6001 2746 6057 2748
rect 6081 2746 6137 2748
rect 6161 2746 6217 2748
rect 5921 2694 5967 2746
rect 5967 2694 5977 2746
rect 6001 2694 6031 2746
rect 6031 2694 6043 2746
rect 6043 2694 6057 2746
rect 6081 2694 6095 2746
rect 6095 2694 6107 2746
rect 6107 2694 6137 2746
rect 6161 2694 6171 2746
rect 6171 2694 6217 2746
rect 5921 2692 5977 2694
rect 6001 2692 6057 2694
rect 6081 2692 6137 2694
rect 6161 2692 6217 2694
rect 9586 14476 9642 14512
rect 9586 14456 9588 14476
rect 9588 14456 9640 14476
rect 9640 14456 9642 14476
rect 9218 12824 9274 12880
rect 9126 11736 9182 11792
rect 9218 11600 9274 11656
rect 9126 11328 9182 11384
rect 9034 11192 9090 11248
rect 9586 12688 9642 12744
rect 9586 12392 9642 12448
rect 10886 32666 10942 32668
rect 10966 32666 11022 32668
rect 11046 32666 11102 32668
rect 11126 32666 11182 32668
rect 10886 32614 10932 32666
rect 10932 32614 10942 32666
rect 10966 32614 10996 32666
rect 10996 32614 11008 32666
rect 11008 32614 11022 32666
rect 11046 32614 11060 32666
rect 11060 32614 11072 32666
rect 11072 32614 11102 32666
rect 11126 32614 11136 32666
rect 11136 32614 11182 32666
rect 10886 32612 10942 32614
rect 10966 32612 11022 32614
rect 11046 32612 11102 32614
rect 11126 32612 11182 32614
rect 10886 31578 10942 31580
rect 10966 31578 11022 31580
rect 11046 31578 11102 31580
rect 11126 31578 11182 31580
rect 10886 31526 10932 31578
rect 10932 31526 10942 31578
rect 10966 31526 10996 31578
rect 10996 31526 11008 31578
rect 11008 31526 11022 31578
rect 11046 31526 11060 31578
rect 11060 31526 11072 31578
rect 11072 31526 11102 31578
rect 11126 31526 11136 31578
rect 11136 31526 11182 31578
rect 10886 31524 10942 31526
rect 10966 31524 11022 31526
rect 11046 31524 11102 31526
rect 11126 31524 11182 31526
rect 10886 30490 10942 30492
rect 10966 30490 11022 30492
rect 11046 30490 11102 30492
rect 11126 30490 11182 30492
rect 10886 30438 10932 30490
rect 10932 30438 10942 30490
rect 10966 30438 10996 30490
rect 10996 30438 11008 30490
rect 11008 30438 11022 30490
rect 11046 30438 11060 30490
rect 11060 30438 11072 30490
rect 11072 30438 11102 30490
rect 11126 30438 11136 30490
rect 11136 30438 11182 30490
rect 10886 30436 10942 30438
rect 10966 30436 11022 30438
rect 11046 30436 11102 30438
rect 11126 30436 11182 30438
rect 11518 31764 11520 31784
rect 11520 31764 11572 31784
rect 11572 31764 11574 31784
rect 11518 31728 11574 31764
rect 10690 27512 10746 27568
rect 10886 29402 10942 29404
rect 10966 29402 11022 29404
rect 11046 29402 11102 29404
rect 11126 29402 11182 29404
rect 10886 29350 10932 29402
rect 10932 29350 10942 29402
rect 10966 29350 10996 29402
rect 10996 29350 11008 29402
rect 11008 29350 11022 29402
rect 11046 29350 11060 29402
rect 11060 29350 11072 29402
rect 11072 29350 11102 29402
rect 11126 29350 11136 29402
rect 11136 29350 11182 29402
rect 10886 29348 10942 29350
rect 10966 29348 11022 29350
rect 11046 29348 11102 29350
rect 11126 29348 11182 29350
rect 10886 28314 10942 28316
rect 10966 28314 11022 28316
rect 11046 28314 11102 28316
rect 11126 28314 11182 28316
rect 10886 28262 10932 28314
rect 10932 28262 10942 28314
rect 10966 28262 10996 28314
rect 10996 28262 11008 28314
rect 11008 28262 11022 28314
rect 11046 28262 11060 28314
rect 11060 28262 11072 28314
rect 11072 28262 11102 28314
rect 11126 28262 11136 28314
rect 11136 28262 11182 28314
rect 10886 28260 10942 28262
rect 10966 28260 11022 28262
rect 11046 28260 11102 28262
rect 11126 28260 11182 28262
rect 10886 27226 10942 27228
rect 10966 27226 11022 27228
rect 11046 27226 11102 27228
rect 11126 27226 11182 27228
rect 10886 27174 10932 27226
rect 10932 27174 10942 27226
rect 10966 27174 10996 27226
rect 10996 27174 11008 27226
rect 11008 27174 11022 27226
rect 11046 27174 11060 27226
rect 11060 27174 11072 27226
rect 11072 27174 11102 27226
rect 11126 27174 11136 27226
rect 11136 27174 11182 27226
rect 10886 27172 10942 27174
rect 10966 27172 11022 27174
rect 11046 27172 11102 27174
rect 11126 27172 11182 27174
rect 10886 26138 10942 26140
rect 10966 26138 11022 26140
rect 11046 26138 11102 26140
rect 11126 26138 11182 26140
rect 10886 26086 10932 26138
rect 10932 26086 10942 26138
rect 10966 26086 10996 26138
rect 10996 26086 11008 26138
rect 11008 26086 11022 26138
rect 11046 26086 11060 26138
rect 11060 26086 11072 26138
rect 11072 26086 11102 26138
rect 11126 26086 11136 26138
rect 11136 26086 11182 26138
rect 10886 26084 10942 26086
rect 10966 26084 11022 26086
rect 11046 26084 11102 26086
rect 11126 26084 11182 26086
rect 10886 25050 10942 25052
rect 10966 25050 11022 25052
rect 11046 25050 11102 25052
rect 11126 25050 11182 25052
rect 10886 24998 10932 25050
rect 10932 24998 10942 25050
rect 10966 24998 10996 25050
rect 10996 24998 11008 25050
rect 11008 24998 11022 25050
rect 11046 24998 11060 25050
rect 11060 24998 11072 25050
rect 11072 24998 11102 25050
rect 11126 24998 11136 25050
rect 11136 24998 11182 25050
rect 10886 24996 10942 24998
rect 10966 24996 11022 24998
rect 11046 24996 11102 24998
rect 11126 24996 11182 24998
rect 10886 23962 10942 23964
rect 10966 23962 11022 23964
rect 11046 23962 11102 23964
rect 11126 23962 11182 23964
rect 10886 23910 10932 23962
rect 10932 23910 10942 23962
rect 10966 23910 10996 23962
rect 10996 23910 11008 23962
rect 11008 23910 11022 23962
rect 11046 23910 11060 23962
rect 11060 23910 11072 23962
rect 11072 23910 11102 23962
rect 11126 23910 11136 23962
rect 11136 23910 11182 23962
rect 10886 23908 10942 23910
rect 10966 23908 11022 23910
rect 11046 23908 11102 23910
rect 11126 23908 11182 23910
rect 10886 22874 10942 22876
rect 10966 22874 11022 22876
rect 11046 22874 11102 22876
rect 11126 22874 11182 22876
rect 10886 22822 10932 22874
rect 10932 22822 10942 22874
rect 10966 22822 10996 22874
rect 10996 22822 11008 22874
rect 11008 22822 11022 22874
rect 11046 22822 11060 22874
rect 11060 22822 11072 22874
rect 11072 22822 11102 22874
rect 11126 22822 11136 22874
rect 11136 22822 11182 22874
rect 10886 22820 10942 22822
rect 10966 22820 11022 22822
rect 11046 22820 11102 22822
rect 11126 22820 11182 22822
rect 10138 17312 10194 17368
rect 9862 11464 9918 11520
rect 10886 21786 10942 21788
rect 10966 21786 11022 21788
rect 11046 21786 11102 21788
rect 11126 21786 11182 21788
rect 10886 21734 10932 21786
rect 10932 21734 10942 21786
rect 10966 21734 10996 21786
rect 10996 21734 11008 21786
rect 11008 21734 11022 21786
rect 11046 21734 11060 21786
rect 11060 21734 11072 21786
rect 11072 21734 11102 21786
rect 11126 21734 11136 21786
rect 11136 21734 11182 21786
rect 10886 21732 10942 21734
rect 10966 21732 11022 21734
rect 11046 21732 11102 21734
rect 11126 21732 11182 21734
rect 10886 20698 10942 20700
rect 10966 20698 11022 20700
rect 11046 20698 11102 20700
rect 11126 20698 11182 20700
rect 10886 20646 10932 20698
rect 10932 20646 10942 20698
rect 10966 20646 10996 20698
rect 10996 20646 11008 20698
rect 11008 20646 11022 20698
rect 11046 20646 11060 20698
rect 11060 20646 11072 20698
rect 11072 20646 11102 20698
rect 11126 20646 11136 20698
rect 11136 20646 11182 20698
rect 10886 20644 10942 20646
rect 10966 20644 11022 20646
rect 11046 20644 11102 20646
rect 11126 20644 11182 20646
rect 10886 19610 10942 19612
rect 10966 19610 11022 19612
rect 11046 19610 11102 19612
rect 11126 19610 11182 19612
rect 10886 19558 10932 19610
rect 10932 19558 10942 19610
rect 10966 19558 10996 19610
rect 10996 19558 11008 19610
rect 11008 19558 11022 19610
rect 11046 19558 11060 19610
rect 11060 19558 11072 19610
rect 11072 19558 11102 19610
rect 11126 19558 11136 19610
rect 11136 19558 11182 19610
rect 10886 19556 10942 19558
rect 10966 19556 11022 19558
rect 11046 19556 11102 19558
rect 11126 19556 11182 19558
rect 10506 12280 10562 12336
rect 10322 12008 10378 12064
rect 10046 7928 10102 7984
rect 10322 7928 10378 7984
rect 10598 11464 10654 11520
rect 11058 19080 11114 19136
rect 10886 18522 10942 18524
rect 10966 18522 11022 18524
rect 11046 18522 11102 18524
rect 11126 18522 11182 18524
rect 10886 18470 10932 18522
rect 10932 18470 10942 18522
rect 10966 18470 10996 18522
rect 10996 18470 11008 18522
rect 11008 18470 11022 18522
rect 11046 18470 11060 18522
rect 11060 18470 11072 18522
rect 11072 18470 11102 18522
rect 11126 18470 11136 18522
rect 11136 18470 11182 18522
rect 10886 18468 10942 18470
rect 10966 18468 11022 18470
rect 11046 18468 11102 18470
rect 11126 18468 11182 18470
rect 10886 17434 10942 17436
rect 10966 17434 11022 17436
rect 11046 17434 11102 17436
rect 11126 17434 11182 17436
rect 10886 17382 10932 17434
rect 10932 17382 10942 17434
rect 10966 17382 10996 17434
rect 10996 17382 11008 17434
rect 11008 17382 11022 17434
rect 11046 17382 11060 17434
rect 11060 17382 11072 17434
rect 11072 17382 11102 17434
rect 11126 17382 11136 17434
rect 11136 17382 11182 17434
rect 10886 17380 10942 17382
rect 10966 17380 11022 17382
rect 11046 17380 11102 17382
rect 11126 17380 11182 17382
rect 10886 16346 10942 16348
rect 10966 16346 11022 16348
rect 11046 16346 11102 16348
rect 11126 16346 11182 16348
rect 10886 16294 10932 16346
rect 10932 16294 10942 16346
rect 10966 16294 10996 16346
rect 10996 16294 11008 16346
rect 11008 16294 11022 16346
rect 11046 16294 11060 16346
rect 11060 16294 11072 16346
rect 11072 16294 11102 16346
rect 11126 16294 11136 16346
rect 11136 16294 11182 16346
rect 10886 16292 10942 16294
rect 10966 16292 11022 16294
rect 11046 16292 11102 16294
rect 11126 16292 11182 16294
rect 10886 15258 10942 15260
rect 10966 15258 11022 15260
rect 11046 15258 11102 15260
rect 11126 15258 11182 15260
rect 10886 15206 10932 15258
rect 10932 15206 10942 15258
rect 10966 15206 10996 15258
rect 10996 15206 11008 15258
rect 11008 15206 11022 15258
rect 11046 15206 11060 15258
rect 11060 15206 11072 15258
rect 11072 15206 11102 15258
rect 11126 15206 11136 15258
rect 11136 15206 11182 15258
rect 10886 15204 10942 15206
rect 10966 15204 11022 15206
rect 11046 15204 11102 15206
rect 11126 15204 11182 15206
rect 10886 14170 10942 14172
rect 10966 14170 11022 14172
rect 11046 14170 11102 14172
rect 11126 14170 11182 14172
rect 10886 14118 10932 14170
rect 10932 14118 10942 14170
rect 10966 14118 10996 14170
rect 10996 14118 11008 14170
rect 11008 14118 11022 14170
rect 11046 14118 11060 14170
rect 11060 14118 11072 14170
rect 11072 14118 11102 14170
rect 11126 14118 11136 14170
rect 11136 14118 11182 14170
rect 10886 14116 10942 14118
rect 10966 14116 11022 14118
rect 11046 14116 11102 14118
rect 11126 14116 11182 14118
rect 13450 26424 13506 26480
rect 15852 39738 15908 39740
rect 15932 39738 15988 39740
rect 16012 39738 16068 39740
rect 16092 39738 16148 39740
rect 15852 39686 15898 39738
rect 15898 39686 15908 39738
rect 15932 39686 15962 39738
rect 15962 39686 15974 39738
rect 15974 39686 15988 39738
rect 16012 39686 16026 39738
rect 16026 39686 16038 39738
rect 16038 39686 16068 39738
rect 16092 39686 16102 39738
rect 16102 39686 16148 39738
rect 15852 39684 15908 39686
rect 15932 39684 15988 39686
rect 16012 39684 16068 39686
rect 16092 39684 16148 39686
rect 15852 38650 15908 38652
rect 15932 38650 15988 38652
rect 16012 38650 16068 38652
rect 16092 38650 16148 38652
rect 15852 38598 15898 38650
rect 15898 38598 15908 38650
rect 15932 38598 15962 38650
rect 15962 38598 15974 38650
rect 15974 38598 15988 38650
rect 16012 38598 16026 38650
rect 16026 38598 16038 38650
rect 16038 38598 16068 38650
rect 16092 38598 16102 38650
rect 16102 38598 16148 38650
rect 15852 38596 15908 38598
rect 15932 38596 15988 38598
rect 16012 38596 16068 38598
rect 16092 38596 16148 38598
rect 15852 37562 15908 37564
rect 15932 37562 15988 37564
rect 16012 37562 16068 37564
rect 16092 37562 16148 37564
rect 15852 37510 15898 37562
rect 15898 37510 15908 37562
rect 15932 37510 15962 37562
rect 15962 37510 15974 37562
rect 15974 37510 15988 37562
rect 16012 37510 16026 37562
rect 16026 37510 16038 37562
rect 16038 37510 16068 37562
rect 16092 37510 16102 37562
rect 16102 37510 16148 37562
rect 15852 37508 15908 37510
rect 15932 37508 15988 37510
rect 16012 37508 16068 37510
rect 16092 37508 16148 37510
rect 15852 36474 15908 36476
rect 15932 36474 15988 36476
rect 16012 36474 16068 36476
rect 16092 36474 16148 36476
rect 15852 36422 15898 36474
rect 15898 36422 15908 36474
rect 15932 36422 15962 36474
rect 15962 36422 15974 36474
rect 15974 36422 15988 36474
rect 16012 36422 16026 36474
rect 16026 36422 16038 36474
rect 16038 36422 16068 36474
rect 16092 36422 16102 36474
rect 16102 36422 16148 36474
rect 15852 36420 15908 36422
rect 15932 36420 15988 36422
rect 16012 36420 16068 36422
rect 16092 36420 16148 36422
rect 13358 25236 13360 25256
rect 13360 25236 13412 25256
rect 13412 25236 13414 25256
rect 13358 25200 13414 25236
rect 12070 15136 12126 15192
rect 11426 13912 11482 13968
rect 10886 13082 10942 13084
rect 10966 13082 11022 13084
rect 11046 13082 11102 13084
rect 11126 13082 11182 13084
rect 10886 13030 10932 13082
rect 10932 13030 10942 13082
rect 10966 13030 10996 13082
rect 10996 13030 11008 13082
rect 11008 13030 11022 13082
rect 11046 13030 11060 13082
rect 11060 13030 11072 13082
rect 11072 13030 11102 13082
rect 11126 13030 11136 13082
rect 11136 13030 11182 13082
rect 10886 13028 10942 13030
rect 10966 13028 11022 13030
rect 11046 13028 11102 13030
rect 11126 13028 11182 13030
rect 11242 12280 11298 12336
rect 10886 11994 10942 11996
rect 10966 11994 11022 11996
rect 11046 11994 11102 11996
rect 11126 11994 11182 11996
rect 10886 11942 10932 11994
rect 10932 11942 10942 11994
rect 10966 11942 10996 11994
rect 10996 11942 11008 11994
rect 11008 11942 11022 11994
rect 11046 11942 11060 11994
rect 11060 11942 11072 11994
rect 11072 11942 11102 11994
rect 11126 11942 11136 11994
rect 11136 11942 11182 11994
rect 10886 11940 10942 11942
rect 10966 11940 11022 11942
rect 11046 11940 11102 11942
rect 11126 11940 11182 11942
rect 10886 10906 10942 10908
rect 10966 10906 11022 10908
rect 11046 10906 11102 10908
rect 11126 10906 11182 10908
rect 10886 10854 10932 10906
rect 10932 10854 10942 10906
rect 10966 10854 10996 10906
rect 10996 10854 11008 10906
rect 11008 10854 11022 10906
rect 11046 10854 11060 10906
rect 11060 10854 11072 10906
rect 11072 10854 11102 10906
rect 11126 10854 11136 10906
rect 11136 10854 11182 10906
rect 10886 10852 10942 10854
rect 10966 10852 11022 10854
rect 11046 10852 11102 10854
rect 11126 10852 11182 10854
rect 10886 9818 10942 9820
rect 10966 9818 11022 9820
rect 11046 9818 11102 9820
rect 11126 9818 11182 9820
rect 10886 9766 10932 9818
rect 10932 9766 10942 9818
rect 10966 9766 10996 9818
rect 10996 9766 11008 9818
rect 11008 9766 11022 9818
rect 11046 9766 11060 9818
rect 11060 9766 11072 9818
rect 11072 9766 11102 9818
rect 11126 9766 11136 9818
rect 11136 9766 11182 9818
rect 10886 9764 10942 9766
rect 10966 9764 11022 9766
rect 11046 9764 11102 9766
rect 11126 9764 11182 9766
rect 10886 8730 10942 8732
rect 10966 8730 11022 8732
rect 11046 8730 11102 8732
rect 11126 8730 11182 8732
rect 10886 8678 10932 8730
rect 10932 8678 10942 8730
rect 10966 8678 10996 8730
rect 10996 8678 11008 8730
rect 11008 8678 11022 8730
rect 11046 8678 11060 8730
rect 11060 8678 11072 8730
rect 11072 8678 11102 8730
rect 11126 8678 11136 8730
rect 11136 8678 11182 8730
rect 10886 8676 10942 8678
rect 10966 8676 11022 8678
rect 11046 8676 11102 8678
rect 11126 8676 11182 8678
rect 10598 6704 10654 6760
rect 10886 7642 10942 7644
rect 10966 7642 11022 7644
rect 11046 7642 11102 7644
rect 11126 7642 11182 7644
rect 10886 7590 10932 7642
rect 10932 7590 10942 7642
rect 10966 7590 10996 7642
rect 10996 7590 11008 7642
rect 11008 7590 11022 7642
rect 11046 7590 11060 7642
rect 11060 7590 11072 7642
rect 11072 7590 11102 7642
rect 11126 7590 11136 7642
rect 11136 7590 11182 7642
rect 10886 7588 10942 7590
rect 10966 7588 11022 7590
rect 11046 7588 11102 7590
rect 11126 7588 11182 7590
rect 10886 6554 10942 6556
rect 10966 6554 11022 6556
rect 11046 6554 11102 6556
rect 11126 6554 11182 6556
rect 10886 6502 10932 6554
rect 10932 6502 10942 6554
rect 10966 6502 10996 6554
rect 10996 6502 11008 6554
rect 11008 6502 11022 6554
rect 11046 6502 11060 6554
rect 11060 6502 11072 6554
rect 11072 6502 11102 6554
rect 11126 6502 11136 6554
rect 11136 6502 11182 6554
rect 10886 6500 10942 6502
rect 10966 6500 11022 6502
rect 11046 6500 11102 6502
rect 11126 6500 11182 6502
rect 10886 5466 10942 5468
rect 10966 5466 11022 5468
rect 11046 5466 11102 5468
rect 11126 5466 11182 5468
rect 10886 5414 10932 5466
rect 10932 5414 10942 5466
rect 10966 5414 10996 5466
rect 10996 5414 11008 5466
rect 11008 5414 11022 5466
rect 11046 5414 11060 5466
rect 11060 5414 11072 5466
rect 11072 5414 11102 5466
rect 11126 5414 11136 5466
rect 11136 5414 11182 5466
rect 10886 5412 10942 5414
rect 10966 5412 11022 5414
rect 11046 5412 11102 5414
rect 11126 5412 11182 5414
rect 10886 4378 10942 4380
rect 10966 4378 11022 4380
rect 11046 4378 11102 4380
rect 11126 4378 11182 4380
rect 10886 4326 10932 4378
rect 10932 4326 10942 4378
rect 10966 4326 10996 4378
rect 10996 4326 11008 4378
rect 11008 4326 11022 4378
rect 11046 4326 11060 4378
rect 11060 4326 11072 4378
rect 11072 4326 11102 4378
rect 11126 4326 11136 4378
rect 11136 4326 11182 4378
rect 10886 4324 10942 4326
rect 10966 4324 11022 4326
rect 11046 4324 11102 4326
rect 11126 4324 11182 4326
rect 10886 3290 10942 3292
rect 10966 3290 11022 3292
rect 11046 3290 11102 3292
rect 11126 3290 11182 3292
rect 10886 3238 10932 3290
rect 10932 3238 10942 3290
rect 10966 3238 10996 3290
rect 10996 3238 11008 3290
rect 11008 3238 11022 3290
rect 11046 3238 11060 3290
rect 11060 3238 11072 3290
rect 11072 3238 11102 3290
rect 11126 3238 11136 3290
rect 11136 3238 11182 3290
rect 10886 3236 10942 3238
rect 10966 3236 11022 3238
rect 11046 3236 11102 3238
rect 11126 3236 11182 3238
rect 10886 2202 10942 2204
rect 10966 2202 11022 2204
rect 11046 2202 11102 2204
rect 11126 2202 11182 2204
rect 10886 2150 10932 2202
rect 10932 2150 10942 2202
rect 10966 2150 10996 2202
rect 10996 2150 11008 2202
rect 11008 2150 11022 2202
rect 11046 2150 11060 2202
rect 11060 2150 11072 2202
rect 11072 2150 11102 2202
rect 11126 2150 11136 2202
rect 11136 2150 11182 2202
rect 10886 2148 10942 2150
rect 10966 2148 11022 2150
rect 11046 2148 11102 2150
rect 11126 2148 11182 2150
rect 15852 35386 15908 35388
rect 15932 35386 15988 35388
rect 16012 35386 16068 35388
rect 16092 35386 16148 35388
rect 15852 35334 15898 35386
rect 15898 35334 15908 35386
rect 15932 35334 15962 35386
rect 15962 35334 15974 35386
rect 15974 35334 15988 35386
rect 16012 35334 16026 35386
rect 16026 35334 16038 35386
rect 16038 35334 16068 35386
rect 16092 35334 16102 35386
rect 16102 35334 16148 35386
rect 15852 35332 15908 35334
rect 15932 35332 15988 35334
rect 16012 35332 16068 35334
rect 16092 35332 16148 35334
rect 15852 34298 15908 34300
rect 15932 34298 15988 34300
rect 16012 34298 16068 34300
rect 16092 34298 16148 34300
rect 15852 34246 15898 34298
rect 15898 34246 15908 34298
rect 15932 34246 15962 34298
rect 15962 34246 15974 34298
rect 15974 34246 15988 34298
rect 16012 34246 16026 34298
rect 16026 34246 16038 34298
rect 16038 34246 16068 34298
rect 16092 34246 16102 34298
rect 16102 34246 16148 34298
rect 15852 34244 15908 34246
rect 15932 34244 15988 34246
rect 16012 34244 16068 34246
rect 16092 34244 16148 34246
rect 15852 33210 15908 33212
rect 15932 33210 15988 33212
rect 16012 33210 16068 33212
rect 16092 33210 16148 33212
rect 15852 33158 15898 33210
rect 15898 33158 15908 33210
rect 15932 33158 15962 33210
rect 15962 33158 15974 33210
rect 15974 33158 15988 33210
rect 16012 33158 16026 33210
rect 16026 33158 16038 33210
rect 16038 33158 16068 33210
rect 16092 33158 16102 33210
rect 16102 33158 16148 33210
rect 15852 33156 15908 33158
rect 15932 33156 15988 33158
rect 16012 33156 16068 33158
rect 16092 33156 16148 33158
rect 15852 32122 15908 32124
rect 15932 32122 15988 32124
rect 16012 32122 16068 32124
rect 16092 32122 16148 32124
rect 15852 32070 15898 32122
rect 15898 32070 15908 32122
rect 15932 32070 15962 32122
rect 15962 32070 15974 32122
rect 15974 32070 15988 32122
rect 16012 32070 16026 32122
rect 16026 32070 16038 32122
rect 16038 32070 16068 32122
rect 16092 32070 16102 32122
rect 16102 32070 16148 32122
rect 15852 32068 15908 32070
rect 15932 32068 15988 32070
rect 16012 32068 16068 32070
rect 16092 32068 16148 32070
rect 15852 31034 15908 31036
rect 15932 31034 15988 31036
rect 16012 31034 16068 31036
rect 16092 31034 16148 31036
rect 15852 30982 15898 31034
rect 15898 30982 15908 31034
rect 15932 30982 15962 31034
rect 15962 30982 15974 31034
rect 15974 30982 15988 31034
rect 16012 30982 16026 31034
rect 16026 30982 16038 31034
rect 16038 30982 16068 31034
rect 16092 30982 16102 31034
rect 16102 30982 16148 31034
rect 15852 30980 15908 30982
rect 15932 30980 15988 30982
rect 16012 30980 16068 30982
rect 16092 30980 16148 30982
rect 15852 29946 15908 29948
rect 15932 29946 15988 29948
rect 16012 29946 16068 29948
rect 16092 29946 16148 29948
rect 15852 29894 15898 29946
rect 15898 29894 15908 29946
rect 15932 29894 15962 29946
rect 15962 29894 15974 29946
rect 15974 29894 15988 29946
rect 16012 29894 16026 29946
rect 16026 29894 16038 29946
rect 16038 29894 16068 29946
rect 16092 29894 16102 29946
rect 16102 29894 16148 29946
rect 15852 29892 15908 29894
rect 15932 29892 15988 29894
rect 16012 29892 16068 29894
rect 16092 29892 16148 29894
rect 15852 28858 15908 28860
rect 15932 28858 15988 28860
rect 16012 28858 16068 28860
rect 16092 28858 16148 28860
rect 15852 28806 15898 28858
rect 15898 28806 15908 28858
rect 15932 28806 15962 28858
rect 15962 28806 15974 28858
rect 15974 28806 15988 28858
rect 16012 28806 16026 28858
rect 16026 28806 16038 28858
rect 16038 28806 16068 28858
rect 16092 28806 16102 28858
rect 16102 28806 16148 28858
rect 15852 28804 15908 28806
rect 15932 28804 15988 28806
rect 16012 28804 16068 28806
rect 16092 28804 16148 28806
rect 15566 27276 15568 27296
rect 15568 27276 15620 27296
rect 15620 27276 15622 27296
rect 15566 27240 15622 27276
rect 15852 27770 15908 27772
rect 15932 27770 15988 27772
rect 16012 27770 16068 27772
rect 16092 27770 16148 27772
rect 15852 27718 15898 27770
rect 15898 27718 15908 27770
rect 15932 27718 15962 27770
rect 15962 27718 15974 27770
rect 15974 27718 15988 27770
rect 16012 27718 16026 27770
rect 16026 27718 16038 27770
rect 16038 27718 16068 27770
rect 16092 27718 16102 27770
rect 16102 27718 16148 27770
rect 15852 27716 15908 27718
rect 15932 27716 15988 27718
rect 16012 27716 16068 27718
rect 16092 27716 16148 27718
rect 15852 26682 15908 26684
rect 15932 26682 15988 26684
rect 16012 26682 16068 26684
rect 16092 26682 16148 26684
rect 15852 26630 15898 26682
rect 15898 26630 15908 26682
rect 15932 26630 15962 26682
rect 15962 26630 15974 26682
rect 15974 26630 15988 26682
rect 16012 26630 16026 26682
rect 16026 26630 16038 26682
rect 16038 26630 16068 26682
rect 16092 26630 16102 26682
rect 16102 26630 16148 26682
rect 15852 26628 15908 26630
rect 15932 26628 15988 26630
rect 16012 26628 16068 26630
rect 16092 26628 16148 26630
rect 15852 25594 15908 25596
rect 15932 25594 15988 25596
rect 16012 25594 16068 25596
rect 16092 25594 16148 25596
rect 15852 25542 15898 25594
rect 15898 25542 15908 25594
rect 15932 25542 15962 25594
rect 15962 25542 15974 25594
rect 15974 25542 15988 25594
rect 16012 25542 16026 25594
rect 16026 25542 16038 25594
rect 16038 25542 16068 25594
rect 16092 25542 16102 25594
rect 16102 25542 16148 25594
rect 15852 25540 15908 25542
rect 15932 25540 15988 25542
rect 16012 25540 16068 25542
rect 16092 25540 16148 25542
rect 15852 24506 15908 24508
rect 15932 24506 15988 24508
rect 16012 24506 16068 24508
rect 16092 24506 16148 24508
rect 15852 24454 15898 24506
rect 15898 24454 15908 24506
rect 15932 24454 15962 24506
rect 15962 24454 15974 24506
rect 15974 24454 15988 24506
rect 16012 24454 16026 24506
rect 16026 24454 16038 24506
rect 16038 24454 16068 24506
rect 16092 24454 16102 24506
rect 16102 24454 16148 24506
rect 15852 24452 15908 24454
rect 15932 24452 15988 24454
rect 16012 24452 16068 24454
rect 16092 24452 16148 24454
rect 16946 33360 17002 33416
rect 15852 23418 15908 23420
rect 15932 23418 15988 23420
rect 16012 23418 16068 23420
rect 16092 23418 16148 23420
rect 15852 23366 15898 23418
rect 15898 23366 15908 23418
rect 15932 23366 15962 23418
rect 15962 23366 15974 23418
rect 15974 23366 15988 23418
rect 16012 23366 16026 23418
rect 16026 23366 16038 23418
rect 16038 23366 16068 23418
rect 16092 23366 16102 23418
rect 16102 23366 16148 23418
rect 15852 23364 15908 23366
rect 15932 23364 15988 23366
rect 16012 23364 16068 23366
rect 16092 23364 16148 23366
rect 15474 19896 15530 19952
rect 13726 9596 13728 9616
rect 13728 9596 13780 9616
rect 13780 9596 13782 9616
rect 13726 9560 13782 9596
rect 14094 8900 14150 8936
rect 14094 8880 14096 8900
rect 14096 8880 14148 8900
rect 14148 8880 14150 8900
rect 16670 23180 16726 23216
rect 16670 23160 16672 23180
rect 16672 23160 16724 23180
rect 16724 23160 16726 23180
rect 15852 22330 15908 22332
rect 15932 22330 15988 22332
rect 16012 22330 16068 22332
rect 16092 22330 16148 22332
rect 15852 22278 15898 22330
rect 15898 22278 15908 22330
rect 15932 22278 15962 22330
rect 15962 22278 15974 22330
rect 15974 22278 15988 22330
rect 16012 22278 16026 22330
rect 16026 22278 16038 22330
rect 16038 22278 16068 22330
rect 16092 22278 16102 22330
rect 16102 22278 16148 22330
rect 15852 22276 15908 22278
rect 15932 22276 15988 22278
rect 16012 22276 16068 22278
rect 16092 22276 16148 22278
rect 15852 21242 15908 21244
rect 15932 21242 15988 21244
rect 16012 21242 16068 21244
rect 16092 21242 16148 21244
rect 15852 21190 15898 21242
rect 15898 21190 15908 21242
rect 15932 21190 15962 21242
rect 15962 21190 15974 21242
rect 15974 21190 15988 21242
rect 16012 21190 16026 21242
rect 16026 21190 16038 21242
rect 16038 21190 16068 21242
rect 16092 21190 16102 21242
rect 16102 21190 16148 21242
rect 15852 21188 15908 21190
rect 15932 21188 15988 21190
rect 16012 21188 16068 21190
rect 16092 21188 16148 21190
rect 15852 20154 15908 20156
rect 15932 20154 15988 20156
rect 16012 20154 16068 20156
rect 16092 20154 16148 20156
rect 15852 20102 15898 20154
rect 15898 20102 15908 20154
rect 15932 20102 15962 20154
rect 15962 20102 15974 20154
rect 15974 20102 15988 20154
rect 16012 20102 16026 20154
rect 16026 20102 16038 20154
rect 16038 20102 16068 20154
rect 16092 20102 16102 20154
rect 16102 20102 16148 20154
rect 15852 20100 15908 20102
rect 15932 20100 15988 20102
rect 16012 20100 16068 20102
rect 16092 20100 16148 20102
rect 15842 19896 15898 19952
rect 15852 19066 15908 19068
rect 15932 19066 15988 19068
rect 16012 19066 16068 19068
rect 16092 19066 16148 19068
rect 15852 19014 15898 19066
rect 15898 19014 15908 19066
rect 15932 19014 15962 19066
rect 15962 19014 15974 19066
rect 15974 19014 15988 19066
rect 16012 19014 16026 19066
rect 16026 19014 16038 19066
rect 16038 19014 16068 19066
rect 16092 19014 16102 19066
rect 16102 19014 16148 19066
rect 15852 19012 15908 19014
rect 15932 19012 15988 19014
rect 16012 19012 16068 19014
rect 16092 19012 16148 19014
rect 15852 17978 15908 17980
rect 15932 17978 15988 17980
rect 16012 17978 16068 17980
rect 16092 17978 16148 17980
rect 15852 17926 15898 17978
rect 15898 17926 15908 17978
rect 15932 17926 15962 17978
rect 15962 17926 15974 17978
rect 15974 17926 15988 17978
rect 16012 17926 16026 17978
rect 16026 17926 16038 17978
rect 16038 17926 16068 17978
rect 16092 17926 16102 17978
rect 16102 17926 16148 17978
rect 15852 17924 15908 17926
rect 15932 17924 15988 17926
rect 16012 17924 16068 17926
rect 16092 17924 16148 17926
rect 15852 16890 15908 16892
rect 15932 16890 15988 16892
rect 16012 16890 16068 16892
rect 16092 16890 16148 16892
rect 15852 16838 15898 16890
rect 15898 16838 15908 16890
rect 15932 16838 15962 16890
rect 15962 16838 15974 16890
rect 15974 16838 15988 16890
rect 16012 16838 16026 16890
rect 16026 16838 16038 16890
rect 16038 16838 16068 16890
rect 16092 16838 16102 16890
rect 16102 16838 16148 16890
rect 15852 16836 15908 16838
rect 15932 16836 15988 16838
rect 16012 16836 16068 16838
rect 16092 16836 16148 16838
rect 15852 15802 15908 15804
rect 15932 15802 15988 15804
rect 16012 15802 16068 15804
rect 16092 15802 16148 15804
rect 15852 15750 15898 15802
rect 15898 15750 15908 15802
rect 15932 15750 15962 15802
rect 15962 15750 15974 15802
rect 15974 15750 15988 15802
rect 16012 15750 16026 15802
rect 16026 15750 16038 15802
rect 16038 15750 16068 15802
rect 16092 15750 16102 15802
rect 16102 15750 16148 15802
rect 15852 15748 15908 15750
rect 15932 15748 15988 15750
rect 16012 15748 16068 15750
rect 16092 15748 16148 15750
rect 16946 22344 17002 22400
rect 16394 15428 16450 15464
rect 16394 15408 16396 15428
rect 16396 15408 16448 15428
rect 16448 15408 16450 15428
rect 15852 14714 15908 14716
rect 15932 14714 15988 14716
rect 16012 14714 16068 14716
rect 16092 14714 16148 14716
rect 15852 14662 15898 14714
rect 15898 14662 15908 14714
rect 15932 14662 15962 14714
rect 15962 14662 15974 14714
rect 15974 14662 15988 14714
rect 16012 14662 16026 14714
rect 16026 14662 16038 14714
rect 16038 14662 16068 14714
rect 16092 14662 16102 14714
rect 16102 14662 16148 14714
rect 15852 14660 15908 14662
rect 15932 14660 15988 14662
rect 16012 14660 16068 14662
rect 16092 14660 16148 14662
rect 15852 13626 15908 13628
rect 15932 13626 15988 13628
rect 16012 13626 16068 13628
rect 16092 13626 16148 13628
rect 15852 13574 15898 13626
rect 15898 13574 15908 13626
rect 15932 13574 15962 13626
rect 15962 13574 15974 13626
rect 15974 13574 15988 13626
rect 16012 13574 16026 13626
rect 16026 13574 16038 13626
rect 16038 13574 16068 13626
rect 16092 13574 16102 13626
rect 16102 13574 16148 13626
rect 15852 13572 15908 13574
rect 15932 13572 15988 13574
rect 16012 13572 16068 13574
rect 16092 13572 16148 13574
rect 15852 12538 15908 12540
rect 15932 12538 15988 12540
rect 16012 12538 16068 12540
rect 16092 12538 16148 12540
rect 15852 12486 15898 12538
rect 15898 12486 15908 12538
rect 15932 12486 15962 12538
rect 15962 12486 15974 12538
rect 15974 12486 15988 12538
rect 16012 12486 16026 12538
rect 16026 12486 16038 12538
rect 16038 12486 16068 12538
rect 16092 12486 16102 12538
rect 16102 12486 16148 12538
rect 15852 12484 15908 12486
rect 15932 12484 15988 12486
rect 16012 12484 16068 12486
rect 16092 12484 16148 12486
rect 15106 9580 15162 9616
rect 15852 11450 15908 11452
rect 15932 11450 15988 11452
rect 16012 11450 16068 11452
rect 16092 11450 16148 11452
rect 15852 11398 15898 11450
rect 15898 11398 15908 11450
rect 15932 11398 15962 11450
rect 15962 11398 15974 11450
rect 15974 11398 15988 11450
rect 16012 11398 16026 11450
rect 16026 11398 16038 11450
rect 16038 11398 16068 11450
rect 16092 11398 16102 11450
rect 16102 11398 16148 11450
rect 15852 11396 15908 11398
rect 15932 11396 15988 11398
rect 16012 11396 16068 11398
rect 16092 11396 16148 11398
rect 15852 10362 15908 10364
rect 15932 10362 15988 10364
rect 16012 10362 16068 10364
rect 16092 10362 16148 10364
rect 15852 10310 15898 10362
rect 15898 10310 15908 10362
rect 15932 10310 15962 10362
rect 15962 10310 15974 10362
rect 15974 10310 15988 10362
rect 16012 10310 16026 10362
rect 16026 10310 16038 10362
rect 16038 10310 16068 10362
rect 16092 10310 16102 10362
rect 16102 10310 16148 10362
rect 15852 10308 15908 10310
rect 15932 10308 15988 10310
rect 16012 10308 16068 10310
rect 16092 10308 16148 10310
rect 15106 9560 15108 9580
rect 15108 9560 15160 9580
rect 15160 9560 15162 9580
rect 15852 9274 15908 9276
rect 15932 9274 15988 9276
rect 16012 9274 16068 9276
rect 16092 9274 16148 9276
rect 15852 9222 15898 9274
rect 15898 9222 15908 9274
rect 15932 9222 15962 9274
rect 15962 9222 15974 9274
rect 15974 9222 15988 9274
rect 16012 9222 16026 9274
rect 16026 9222 16038 9274
rect 16038 9222 16068 9274
rect 16092 9222 16102 9274
rect 16102 9222 16148 9274
rect 15852 9220 15908 9222
rect 15932 9220 15988 9222
rect 16012 9220 16068 9222
rect 16092 9220 16148 9222
rect 15852 8186 15908 8188
rect 15932 8186 15988 8188
rect 16012 8186 16068 8188
rect 16092 8186 16148 8188
rect 15852 8134 15898 8186
rect 15898 8134 15908 8186
rect 15932 8134 15962 8186
rect 15962 8134 15974 8186
rect 15974 8134 15988 8186
rect 16012 8134 16026 8186
rect 16026 8134 16038 8186
rect 16038 8134 16068 8186
rect 16092 8134 16102 8186
rect 16102 8134 16148 8186
rect 15852 8132 15908 8134
rect 15932 8132 15988 8134
rect 16012 8132 16068 8134
rect 16092 8132 16148 8134
rect 15852 7098 15908 7100
rect 15932 7098 15988 7100
rect 16012 7098 16068 7100
rect 16092 7098 16148 7100
rect 15852 7046 15898 7098
rect 15898 7046 15908 7098
rect 15932 7046 15962 7098
rect 15962 7046 15974 7098
rect 15974 7046 15988 7098
rect 16012 7046 16026 7098
rect 16026 7046 16038 7098
rect 16038 7046 16068 7098
rect 16092 7046 16102 7098
rect 16102 7046 16148 7098
rect 15852 7044 15908 7046
rect 15932 7044 15988 7046
rect 16012 7044 16068 7046
rect 16092 7044 16148 7046
rect 17682 27376 17738 27432
rect 17130 15272 17186 15328
rect 17038 15036 17040 15056
rect 17040 15036 17092 15056
rect 17092 15036 17094 15056
rect 17038 15000 17094 15036
rect 17222 15136 17278 15192
rect 17406 15444 17408 15464
rect 17408 15444 17460 15464
rect 17460 15444 17462 15464
rect 17406 15408 17462 15444
rect 17406 15272 17462 15328
rect 17590 21936 17646 21992
rect 20817 42458 20873 42460
rect 20897 42458 20953 42460
rect 20977 42458 21033 42460
rect 21057 42458 21113 42460
rect 20817 42406 20863 42458
rect 20863 42406 20873 42458
rect 20897 42406 20927 42458
rect 20927 42406 20939 42458
rect 20939 42406 20953 42458
rect 20977 42406 20991 42458
rect 20991 42406 21003 42458
rect 21003 42406 21033 42458
rect 21057 42406 21067 42458
rect 21067 42406 21113 42458
rect 20817 42404 20873 42406
rect 20897 42404 20953 42406
rect 20977 42404 21033 42406
rect 21057 42404 21113 42406
rect 20817 41370 20873 41372
rect 20897 41370 20953 41372
rect 20977 41370 21033 41372
rect 21057 41370 21113 41372
rect 20817 41318 20863 41370
rect 20863 41318 20873 41370
rect 20897 41318 20927 41370
rect 20927 41318 20939 41370
rect 20939 41318 20953 41370
rect 20977 41318 20991 41370
rect 20991 41318 21003 41370
rect 21003 41318 21033 41370
rect 21057 41318 21067 41370
rect 21067 41318 21113 41370
rect 20817 41316 20873 41318
rect 20897 41316 20953 41318
rect 20977 41316 21033 41318
rect 21057 41316 21113 41318
rect 20817 40282 20873 40284
rect 20897 40282 20953 40284
rect 20977 40282 21033 40284
rect 21057 40282 21113 40284
rect 20817 40230 20863 40282
rect 20863 40230 20873 40282
rect 20897 40230 20927 40282
rect 20927 40230 20939 40282
rect 20939 40230 20953 40282
rect 20977 40230 20991 40282
rect 20991 40230 21003 40282
rect 21003 40230 21033 40282
rect 21057 40230 21067 40282
rect 21067 40230 21113 40282
rect 20817 40228 20873 40230
rect 20897 40228 20953 40230
rect 20977 40228 21033 40230
rect 21057 40228 21113 40230
rect 20817 39194 20873 39196
rect 20897 39194 20953 39196
rect 20977 39194 21033 39196
rect 21057 39194 21113 39196
rect 20817 39142 20863 39194
rect 20863 39142 20873 39194
rect 20897 39142 20927 39194
rect 20927 39142 20939 39194
rect 20939 39142 20953 39194
rect 20977 39142 20991 39194
rect 20991 39142 21003 39194
rect 21003 39142 21033 39194
rect 21057 39142 21067 39194
rect 21067 39142 21113 39194
rect 20817 39140 20873 39142
rect 20897 39140 20953 39142
rect 20977 39140 21033 39142
rect 21057 39140 21113 39142
rect 20817 38106 20873 38108
rect 20897 38106 20953 38108
rect 20977 38106 21033 38108
rect 21057 38106 21113 38108
rect 20817 38054 20863 38106
rect 20863 38054 20873 38106
rect 20897 38054 20927 38106
rect 20927 38054 20939 38106
rect 20939 38054 20953 38106
rect 20977 38054 20991 38106
rect 20991 38054 21003 38106
rect 21003 38054 21033 38106
rect 21057 38054 21067 38106
rect 21067 38054 21113 38106
rect 20817 38052 20873 38054
rect 20897 38052 20953 38054
rect 20977 38052 21033 38054
rect 21057 38052 21113 38054
rect 18050 25220 18106 25256
rect 18050 25200 18052 25220
rect 18052 25200 18104 25220
rect 18104 25200 18106 25220
rect 17866 15020 17922 15056
rect 17866 15000 17868 15020
rect 17868 15000 17920 15020
rect 17920 15000 17922 15020
rect 16302 8880 16358 8936
rect 16210 6704 16266 6760
rect 15852 6010 15908 6012
rect 15932 6010 15988 6012
rect 16012 6010 16068 6012
rect 16092 6010 16148 6012
rect 15852 5958 15898 6010
rect 15898 5958 15908 6010
rect 15932 5958 15962 6010
rect 15962 5958 15974 6010
rect 15974 5958 15988 6010
rect 16012 5958 16026 6010
rect 16026 5958 16038 6010
rect 16038 5958 16068 6010
rect 16092 5958 16102 6010
rect 16102 5958 16148 6010
rect 15852 5956 15908 5958
rect 15932 5956 15988 5958
rect 16012 5956 16068 5958
rect 16092 5956 16148 5958
rect 15852 4922 15908 4924
rect 15932 4922 15988 4924
rect 16012 4922 16068 4924
rect 16092 4922 16148 4924
rect 15852 4870 15898 4922
rect 15898 4870 15908 4922
rect 15932 4870 15962 4922
rect 15962 4870 15974 4922
rect 15974 4870 15988 4922
rect 16012 4870 16026 4922
rect 16026 4870 16038 4922
rect 16038 4870 16068 4922
rect 16092 4870 16102 4922
rect 16102 4870 16148 4922
rect 15852 4868 15908 4870
rect 15932 4868 15988 4870
rect 16012 4868 16068 4870
rect 16092 4868 16148 4870
rect 15852 3834 15908 3836
rect 15932 3834 15988 3836
rect 16012 3834 16068 3836
rect 16092 3834 16148 3836
rect 15852 3782 15898 3834
rect 15898 3782 15908 3834
rect 15932 3782 15962 3834
rect 15962 3782 15974 3834
rect 15974 3782 15988 3834
rect 16012 3782 16026 3834
rect 16026 3782 16038 3834
rect 16038 3782 16068 3834
rect 16092 3782 16102 3834
rect 16102 3782 16148 3834
rect 15852 3780 15908 3782
rect 15932 3780 15988 3782
rect 16012 3780 16068 3782
rect 16092 3780 16148 3782
rect 15852 2746 15908 2748
rect 15932 2746 15988 2748
rect 16012 2746 16068 2748
rect 16092 2746 16148 2748
rect 15852 2694 15898 2746
rect 15898 2694 15908 2746
rect 15932 2694 15962 2746
rect 15962 2694 15974 2746
rect 15974 2694 15988 2746
rect 16012 2694 16026 2746
rect 16026 2694 16038 2746
rect 16038 2694 16068 2746
rect 16092 2694 16102 2746
rect 16102 2694 16148 2746
rect 15852 2692 15908 2694
rect 15932 2692 15988 2694
rect 16012 2692 16068 2694
rect 16092 2692 16148 2694
rect 17774 9016 17830 9072
rect 18326 15272 18382 15328
rect 18602 13912 18658 13968
rect 19062 27412 19064 27432
rect 19064 27412 19116 27432
rect 19116 27412 19118 27432
rect 19062 27376 19118 27412
rect 19154 27240 19210 27296
rect 20817 37018 20873 37020
rect 20897 37018 20953 37020
rect 20977 37018 21033 37020
rect 21057 37018 21113 37020
rect 20817 36966 20863 37018
rect 20863 36966 20873 37018
rect 20897 36966 20927 37018
rect 20927 36966 20939 37018
rect 20939 36966 20953 37018
rect 20977 36966 20991 37018
rect 20991 36966 21003 37018
rect 21003 36966 21033 37018
rect 21057 36966 21067 37018
rect 21067 36966 21113 37018
rect 20817 36964 20873 36966
rect 20897 36964 20953 36966
rect 20977 36964 21033 36966
rect 21057 36964 21113 36966
rect 20817 35930 20873 35932
rect 20897 35930 20953 35932
rect 20977 35930 21033 35932
rect 21057 35930 21113 35932
rect 20817 35878 20863 35930
rect 20863 35878 20873 35930
rect 20897 35878 20927 35930
rect 20927 35878 20939 35930
rect 20939 35878 20953 35930
rect 20977 35878 20991 35930
rect 20991 35878 21003 35930
rect 21003 35878 21033 35930
rect 21057 35878 21067 35930
rect 21067 35878 21113 35930
rect 20817 35876 20873 35878
rect 20897 35876 20953 35878
rect 20977 35876 21033 35878
rect 21057 35876 21113 35878
rect 20817 34842 20873 34844
rect 20897 34842 20953 34844
rect 20977 34842 21033 34844
rect 21057 34842 21113 34844
rect 20817 34790 20863 34842
rect 20863 34790 20873 34842
rect 20897 34790 20927 34842
rect 20927 34790 20939 34842
rect 20939 34790 20953 34842
rect 20977 34790 20991 34842
rect 20991 34790 21003 34842
rect 21003 34790 21033 34842
rect 21057 34790 21067 34842
rect 21067 34790 21113 34842
rect 20817 34788 20873 34790
rect 20897 34788 20953 34790
rect 20977 34788 21033 34790
rect 21057 34788 21113 34790
rect 20817 33754 20873 33756
rect 20897 33754 20953 33756
rect 20977 33754 21033 33756
rect 21057 33754 21113 33756
rect 20817 33702 20863 33754
rect 20863 33702 20873 33754
rect 20897 33702 20927 33754
rect 20927 33702 20939 33754
rect 20939 33702 20953 33754
rect 20977 33702 20991 33754
rect 20991 33702 21003 33754
rect 21003 33702 21033 33754
rect 21057 33702 21067 33754
rect 21067 33702 21113 33754
rect 20817 33700 20873 33702
rect 20897 33700 20953 33702
rect 20977 33700 21033 33702
rect 21057 33700 21113 33702
rect 20817 32666 20873 32668
rect 20897 32666 20953 32668
rect 20977 32666 21033 32668
rect 21057 32666 21113 32668
rect 20817 32614 20863 32666
rect 20863 32614 20873 32666
rect 20897 32614 20927 32666
rect 20927 32614 20939 32666
rect 20939 32614 20953 32666
rect 20977 32614 20991 32666
rect 20991 32614 21003 32666
rect 21003 32614 21033 32666
rect 21057 32614 21067 32666
rect 21067 32614 21113 32666
rect 20817 32612 20873 32614
rect 20897 32612 20953 32614
rect 20977 32612 21033 32614
rect 21057 32612 21113 32614
rect 20817 31578 20873 31580
rect 20897 31578 20953 31580
rect 20977 31578 21033 31580
rect 21057 31578 21113 31580
rect 20817 31526 20863 31578
rect 20863 31526 20873 31578
rect 20897 31526 20927 31578
rect 20927 31526 20939 31578
rect 20939 31526 20953 31578
rect 20977 31526 20991 31578
rect 20991 31526 21003 31578
rect 21003 31526 21033 31578
rect 21057 31526 21067 31578
rect 21067 31526 21113 31578
rect 20817 31524 20873 31526
rect 20897 31524 20953 31526
rect 20977 31524 21033 31526
rect 21057 31524 21113 31526
rect 20817 30490 20873 30492
rect 20897 30490 20953 30492
rect 20977 30490 21033 30492
rect 21057 30490 21113 30492
rect 20817 30438 20863 30490
rect 20863 30438 20873 30490
rect 20897 30438 20927 30490
rect 20927 30438 20939 30490
rect 20939 30438 20953 30490
rect 20977 30438 20991 30490
rect 20991 30438 21003 30490
rect 21003 30438 21033 30490
rect 21057 30438 21067 30490
rect 21067 30438 21113 30490
rect 20817 30436 20873 30438
rect 20897 30436 20953 30438
rect 20977 30436 21033 30438
rect 21057 30436 21113 30438
rect 19338 17212 19340 17232
rect 19340 17212 19392 17232
rect 19392 17212 19394 17232
rect 19338 17176 19394 17212
rect 20817 29402 20873 29404
rect 20897 29402 20953 29404
rect 20977 29402 21033 29404
rect 21057 29402 21113 29404
rect 20817 29350 20863 29402
rect 20863 29350 20873 29402
rect 20897 29350 20927 29402
rect 20927 29350 20939 29402
rect 20939 29350 20953 29402
rect 20977 29350 20991 29402
rect 20991 29350 21003 29402
rect 21003 29350 21033 29402
rect 21057 29350 21067 29402
rect 21067 29350 21113 29402
rect 20817 29348 20873 29350
rect 20897 29348 20953 29350
rect 20977 29348 21033 29350
rect 21057 29348 21113 29350
rect 20817 28314 20873 28316
rect 20897 28314 20953 28316
rect 20977 28314 21033 28316
rect 21057 28314 21113 28316
rect 20817 28262 20863 28314
rect 20863 28262 20873 28314
rect 20897 28262 20927 28314
rect 20927 28262 20939 28314
rect 20939 28262 20953 28314
rect 20977 28262 20991 28314
rect 20991 28262 21003 28314
rect 21003 28262 21033 28314
rect 21057 28262 21067 28314
rect 21067 28262 21113 28314
rect 20817 28260 20873 28262
rect 20897 28260 20953 28262
rect 20977 28260 21033 28262
rect 21057 28260 21113 28262
rect 20817 27226 20873 27228
rect 20897 27226 20953 27228
rect 20977 27226 21033 27228
rect 21057 27226 21113 27228
rect 20817 27174 20863 27226
rect 20863 27174 20873 27226
rect 20897 27174 20927 27226
rect 20927 27174 20939 27226
rect 20939 27174 20953 27226
rect 20977 27174 20991 27226
rect 20991 27174 21003 27226
rect 21003 27174 21033 27226
rect 21057 27174 21067 27226
rect 21067 27174 21113 27226
rect 20817 27172 20873 27174
rect 20897 27172 20953 27174
rect 20977 27172 21033 27174
rect 21057 27172 21113 27174
rect 18234 9052 18236 9072
rect 18236 9052 18288 9072
rect 18288 9052 18290 9072
rect 18234 9016 18290 9052
rect 20817 26138 20873 26140
rect 20897 26138 20953 26140
rect 20977 26138 21033 26140
rect 21057 26138 21113 26140
rect 20817 26086 20863 26138
rect 20863 26086 20873 26138
rect 20897 26086 20927 26138
rect 20927 26086 20939 26138
rect 20939 26086 20953 26138
rect 20977 26086 20991 26138
rect 20991 26086 21003 26138
rect 21003 26086 21033 26138
rect 21057 26086 21067 26138
rect 21067 26086 21113 26138
rect 20817 26084 20873 26086
rect 20897 26084 20953 26086
rect 20977 26084 21033 26086
rect 21057 26084 21113 26086
rect 20817 25050 20873 25052
rect 20897 25050 20953 25052
rect 20977 25050 21033 25052
rect 21057 25050 21113 25052
rect 20817 24998 20863 25050
rect 20863 24998 20873 25050
rect 20897 24998 20927 25050
rect 20927 24998 20939 25050
rect 20939 24998 20953 25050
rect 20977 24998 20991 25050
rect 20991 24998 21003 25050
rect 21003 24998 21033 25050
rect 21057 24998 21067 25050
rect 21067 24998 21113 25050
rect 20817 24996 20873 24998
rect 20897 24996 20953 24998
rect 20977 24996 21033 24998
rect 21057 24996 21113 24998
rect 20817 23962 20873 23964
rect 20897 23962 20953 23964
rect 20977 23962 21033 23964
rect 21057 23962 21113 23964
rect 20817 23910 20863 23962
rect 20863 23910 20873 23962
rect 20897 23910 20927 23962
rect 20927 23910 20939 23962
rect 20939 23910 20953 23962
rect 20977 23910 20991 23962
rect 20991 23910 21003 23962
rect 21003 23910 21033 23962
rect 21057 23910 21067 23962
rect 21067 23910 21113 23962
rect 20817 23908 20873 23910
rect 20897 23908 20953 23910
rect 20977 23908 21033 23910
rect 21057 23908 21113 23910
rect 20817 22874 20873 22876
rect 20897 22874 20953 22876
rect 20977 22874 21033 22876
rect 21057 22874 21113 22876
rect 20817 22822 20863 22874
rect 20863 22822 20873 22874
rect 20897 22822 20927 22874
rect 20927 22822 20939 22874
rect 20939 22822 20953 22874
rect 20977 22822 20991 22874
rect 20991 22822 21003 22874
rect 21003 22822 21033 22874
rect 21057 22822 21067 22874
rect 21067 22822 21113 22874
rect 20817 22820 20873 22822
rect 20897 22820 20953 22822
rect 20977 22820 21033 22822
rect 21057 22820 21113 22822
rect 20817 21786 20873 21788
rect 20897 21786 20953 21788
rect 20977 21786 21033 21788
rect 21057 21786 21113 21788
rect 20817 21734 20863 21786
rect 20863 21734 20873 21786
rect 20897 21734 20927 21786
rect 20927 21734 20939 21786
rect 20939 21734 20953 21786
rect 20977 21734 20991 21786
rect 20991 21734 21003 21786
rect 21003 21734 21033 21786
rect 21057 21734 21067 21786
rect 21067 21734 21113 21786
rect 20817 21732 20873 21734
rect 20897 21732 20953 21734
rect 20977 21732 21033 21734
rect 21057 21732 21113 21734
rect 25782 41914 25838 41916
rect 25862 41914 25918 41916
rect 25942 41914 25998 41916
rect 26022 41914 26078 41916
rect 25782 41862 25828 41914
rect 25828 41862 25838 41914
rect 25862 41862 25892 41914
rect 25892 41862 25904 41914
rect 25904 41862 25918 41914
rect 25942 41862 25956 41914
rect 25956 41862 25968 41914
rect 25968 41862 25998 41914
rect 26022 41862 26032 41914
rect 26032 41862 26078 41914
rect 25782 41860 25838 41862
rect 25862 41860 25918 41862
rect 25942 41860 25998 41862
rect 26022 41860 26078 41862
rect 30102 40976 30158 41032
rect 25782 40826 25838 40828
rect 25862 40826 25918 40828
rect 25942 40826 25998 40828
rect 26022 40826 26078 40828
rect 25782 40774 25828 40826
rect 25828 40774 25838 40826
rect 25862 40774 25892 40826
rect 25892 40774 25904 40826
rect 25904 40774 25918 40826
rect 25942 40774 25956 40826
rect 25956 40774 25968 40826
rect 25968 40774 25998 40826
rect 26022 40774 26032 40826
rect 26032 40774 26078 40826
rect 25782 40772 25838 40774
rect 25862 40772 25918 40774
rect 25942 40772 25998 40774
rect 26022 40772 26078 40774
rect 25782 39738 25838 39740
rect 25862 39738 25918 39740
rect 25942 39738 25998 39740
rect 26022 39738 26078 39740
rect 25782 39686 25828 39738
rect 25828 39686 25838 39738
rect 25862 39686 25892 39738
rect 25892 39686 25904 39738
rect 25904 39686 25918 39738
rect 25942 39686 25956 39738
rect 25956 39686 25968 39738
rect 25968 39686 25998 39738
rect 26022 39686 26032 39738
rect 26032 39686 26078 39738
rect 25782 39684 25838 39686
rect 25862 39684 25918 39686
rect 25942 39684 25998 39686
rect 26022 39684 26078 39686
rect 30102 38936 30158 38992
rect 25782 38650 25838 38652
rect 25862 38650 25918 38652
rect 25942 38650 25998 38652
rect 26022 38650 26078 38652
rect 25782 38598 25828 38650
rect 25828 38598 25838 38650
rect 25862 38598 25892 38650
rect 25892 38598 25904 38650
rect 25904 38598 25918 38650
rect 25942 38598 25956 38650
rect 25956 38598 25968 38650
rect 25968 38598 25998 38650
rect 26022 38598 26032 38650
rect 26032 38598 26078 38650
rect 25782 38596 25838 38598
rect 25862 38596 25918 38598
rect 25942 38596 25998 38598
rect 26022 38596 26078 38598
rect 25782 37562 25838 37564
rect 25862 37562 25918 37564
rect 25942 37562 25998 37564
rect 26022 37562 26078 37564
rect 25782 37510 25828 37562
rect 25828 37510 25838 37562
rect 25862 37510 25892 37562
rect 25892 37510 25904 37562
rect 25904 37510 25918 37562
rect 25942 37510 25956 37562
rect 25956 37510 25968 37562
rect 25968 37510 25998 37562
rect 26022 37510 26032 37562
rect 26032 37510 26078 37562
rect 25782 37508 25838 37510
rect 25862 37508 25918 37510
rect 25942 37508 25998 37510
rect 26022 37508 26078 37510
rect 30102 36896 30158 36952
rect 25782 36474 25838 36476
rect 25862 36474 25918 36476
rect 25942 36474 25998 36476
rect 26022 36474 26078 36476
rect 25782 36422 25828 36474
rect 25828 36422 25838 36474
rect 25862 36422 25892 36474
rect 25892 36422 25904 36474
rect 25904 36422 25918 36474
rect 25942 36422 25956 36474
rect 25956 36422 25968 36474
rect 25968 36422 25998 36474
rect 26022 36422 26032 36474
rect 26032 36422 26078 36474
rect 25782 36420 25838 36422
rect 25862 36420 25918 36422
rect 25942 36420 25998 36422
rect 26022 36420 26078 36422
rect 25782 35386 25838 35388
rect 25862 35386 25918 35388
rect 25942 35386 25998 35388
rect 26022 35386 26078 35388
rect 25782 35334 25828 35386
rect 25828 35334 25838 35386
rect 25862 35334 25892 35386
rect 25892 35334 25904 35386
rect 25904 35334 25918 35386
rect 25942 35334 25956 35386
rect 25956 35334 25968 35386
rect 25968 35334 25998 35386
rect 26022 35334 26032 35386
rect 26032 35334 26078 35386
rect 25782 35332 25838 35334
rect 25862 35332 25918 35334
rect 25942 35332 25998 35334
rect 26022 35332 26078 35334
rect 30102 35028 30104 35048
rect 30104 35028 30156 35048
rect 30156 35028 30158 35048
rect 30102 34992 30158 35028
rect 25782 34298 25838 34300
rect 25862 34298 25918 34300
rect 25942 34298 25998 34300
rect 26022 34298 26078 34300
rect 25782 34246 25828 34298
rect 25828 34246 25838 34298
rect 25862 34246 25892 34298
rect 25892 34246 25904 34298
rect 25904 34246 25918 34298
rect 25942 34246 25956 34298
rect 25956 34246 25968 34298
rect 25968 34246 25998 34298
rect 26022 34246 26032 34298
rect 26032 34246 26078 34298
rect 25782 34244 25838 34246
rect 25862 34244 25918 34246
rect 25942 34244 25998 34246
rect 26022 34244 26078 34246
rect 20817 20698 20873 20700
rect 20897 20698 20953 20700
rect 20977 20698 21033 20700
rect 21057 20698 21113 20700
rect 20817 20646 20863 20698
rect 20863 20646 20873 20698
rect 20897 20646 20927 20698
rect 20927 20646 20939 20698
rect 20939 20646 20953 20698
rect 20977 20646 20991 20698
rect 20991 20646 21003 20698
rect 21003 20646 21033 20698
rect 21057 20646 21067 20698
rect 21067 20646 21113 20698
rect 20817 20644 20873 20646
rect 20897 20644 20953 20646
rect 20977 20644 21033 20646
rect 21057 20644 21113 20646
rect 20817 19610 20873 19612
rect 20897 19610 20953 19612
rect 20977 19610 21033 19612
rect 21057 19610 21113 19612
rect 20817 19558 20863 19610
rect 20863 19558 20873 19610
rect 20897 19558 20927 19610
rect 20927 19558 20939 19610
rect 20939 19558 20953 19610
rect 20977 19558 20991 19610
rect 20991 19558 21003 19610
rect 21003 19558 21033 19610
rect 21057 19558 21067 19610
rect 21067 19558 21113 19610
rect 20817 19556 20873 19558
rect 20897 19556 20953 19558
rect 20977 19556 21033 19558
rect 21057 19556 21113 19558
rect 20817 18522 20873 18524
rect 20897 18522 20953 18524
rect 20977 18522 21033 18524
rect 21057 18522 21113 18524
rect 20817 18470 20863 18522
rect 20863 18470 20873 18522
rect 20897 18470 20927 18522
rect 20927 18470 20939 18522
rect 20939 18470 20953 18522
rect 20977 18470 20991 18522
rect 20991 18470 21003 18522
rect 21003 18470 21033 18522
rect 21057 18470 21067 18522
rect 21067 18470 21113 18522
rect 20817 18468 20873 18470
rect 20897 18468 20953 18470
rect 20977 18468 21033 18470
rect 21057 18468 21113 18470
rect 20817 17434 20873 17436
rect 20897 17434 20953 17436
rect 20977 17434 21033 17436
rect 21057 17434 21113 17436
rect 20817 17382 20863 17434
rect 20863 17382 20873 17434
rect 20897 17382 20927 17434
rect 20927 17382 20939 17434
rect 20939 17382 20953 17434
rect 20977 17382 20991 17434
rect 20991 17382 21003 17434
rect 21003 17382 21033 17434
rect 21057 17382 21067 17434
rect 21067 17382 21113 17434
rect 20817 17380 20873 17382
rect 20897 17380 20953 17382
rect 20977 17380 21033 17382
rect 21057 17380 21113 17382
rect 20626 17176 20682 17232
rect 20817 16346 20873 16348
rect 20897 16346 20953 16348
rect 20977 16346 21033 16348
rect 21057 16346 21113 16348
rect 20817 16294 20863 16346
rect 20863 16294 20873 16346
rect 20897 16294 20927 16346
rect 20927 16294 20939 16346
rect 20939 16294 20953 16346
rect 20977 16294 20991 16346
rect 20991 16294 21003 16346
rect 21003 16294 21033 16346
rect 21057 16294 21067 16346
rect 21067 16294 21113 16346
rect 20817 16292 20873 16294
rect 20897 16292 20953 16294
rect 20977 16292 21033 16294
rect 21057 16292 21113 16294
rect 20817 15258 20873 15260
rect 20897 15258 20953 15260
rect 20977 15258 21033 15260
rect 21057 15258 21113 15260
rect 20817 15206 20863 15258
rect 20863 15206 20873 15258
rect 20897 15206 20927 15258
rect 20927 15206 20939 15258
rect 20939 15206 20953 15258
rect 20977 15206 20991 15258
rect 20991 15206 21003 15258
rect 21003 15206 21033 15258
rect 21057 15206 21067 15258
rect 21067 15206 21113 15258
rect 20817 15204 20873 15206
rect 20897 15204 20953 15206
rect 20977 15204 21033 15206
rect 21057 15204 21113 15206
rect 25782 33210 25838 33212
rect 25862 33210 25918 33212
rect 25942 33210 25998 33212
rect 26022 33210 26078 33212
rect 25782 33158 25828 33210
rect 25828 33158 25838 33210
rect 25862 33158 25892 33210
rect 25892 33158 25904 33210
rect 25904 33158 25918 33210
rect 25942 33158 25956 33210
rect 25956 33158 25968 33210
rect 25968 33158 25998 33210
rect 26022 33158 26032 33210
rect 26032 33158 26078 33210
rect 25782 33156 25838 33158
rect 25862 33156 25918 33158
rect 25942 33156 25998 33158
rect 26022 33156 26078 33158
rect 30102 32952 30158 33008
rect 25782 32122 25838 32124
rect 25862 32122 25918 32124
rect 25942 32122 25998 32124
rect 26022 32122 26078 32124
rect 25782 32070 25828 32122
rect 25828 32070 25838 32122
rect 25862 32070 25892 32122
rect 25892 32070 25904 32122
rect 25904 32070 25918 32122
rect 25942 32070 25956 32122
rect 25956 32070 25968 32122
rect 25968 32070 25998 32122
rect 26022 32070 26032 32122
rect 26032 32070 26078 32122
rect 25782 32068 25838 32070
rect 25862 32068 25918 32070
rect 25942 32068 25998 32070
rect 26022 32068 26078 32070
rect 25782 31034 25838 31036
rect 25862 31034 25918 31036
rect 25942 31034 25998 31036
rect 26022 31034 26078 31036
rect 25782 30982 25828 31034
rect 25828 30982 25838 31034
rect 25862 30982 25892 31034
rect 25892 30982 25904 31034
rect 25904 30982 25918 31034
rect 25942 30982 25956 31034
rect 25956 30982 25968 31034
rect 25968 30982 25998 31034
rect 26022 30982 26032 31034
rect 26032 30982 26078 31034
rect 25782 30980 25838 30982
rect 25862 30980 25918 30982
rect 25942 30980 25998 30982
rect 26022 30980 26078 30982
rect 30102 30912 30158 30968
rect 25782 29946 25838 29948
rect 25862 29946 25918 29948
rect 25942 29946 25998 29948
rect 26022 29946 26078 29948
rect 25782 29894 25828 29946
rect 25828 29894 25838 29946
rect 25862 29894 25892 29946
rect 25892 29894 25904 29946
rect 25904 29894 25918 29946
rect 25942 29894 25956 29946
rect 25956 29894 25968 29946
rect 25968 29894 25998 29946
rect 26022 29894 26032 29946
rect 26032 29894 26078 29946
rect 25782 29892 25838 29894
rect 25862 29892 25918 29894
rect 25942 29892 25998 29894
rect 26022 29892 26078 29894
rect 25782 28858 25838 28860
rect 25862 28858 25918 28860
rect 25942 28858 25998 28860
rect 26022 28858 26078 28860
rect 25782 28806 25828 28858
rect 25828 28806 25838 28858
rect 25862 28806 25892 28858
rect 25892 28806 25904 28858
rect 25904 28806 25918 28858
rect 25942 28806 25956 28858
rect 25956 28806 25968 28858
rect 25968 28806 25998 28858
rect 26022 28806 26032 28858
rect 26032 28806 26078 28858
rect 25782 28804 25838 28806
rect 25862 28804 25918 28806
rect 25942 28804 25998 28806
rect 26022 28804 26078 28806
rect 25782 27770 25838 27772
rect 25862 27770 25918 27772
rect 25942 27770 25998 27772
rect 26022 27770 26078 27772
rect 25782 27718 25828 27770
rect 25828 27718 25838 27770
rect 25862 27718 25892 27770
rect 25892 27718 25904 27770
rect 25904 27718 25918 27770
rect 25942 27718 25956 27770
rect 25956 27718 25968 27770
rect 25968 27718 25998 27770
rect 26022 27718 26032 27770
rect 26032 27718 26078 27770
rect 25782 27716 25838 27718
rect 25862 27716 25918 27718
rect 25942 27716 25998 27718
rect 26022 27716 26078 27718
rect 25782 26682 25838 26684
rect 25862 26682 25918 26684
rect 25942 26682 25998 26684
rect 26022 26682 26078 26684
rect 25782 26630 25828 26682
rect 25828 26630 25838 26682
rect 25862 26630 25892 26682
rect 25892 26630 25904 26682
rect 25904 26630 25918 26682
rect 25942 26630 25956 26682
rect 25956 26630 25968 26682
rect 25968 26630 25998 26682
rect 26022 26630 26032 26682
rect 26032 26630 26078 26682
rect 25782 26628 25838 26630
rect 25862 26628 25918 26630
rect 25942 26628 25998 26630
rect 26022 26628 26078 26630
rect 25782 25594 25838 25596
rect 25862 25594 25918 25596
rect 25942 25594 25998 25596
rect 26022 25594 26078 25596
rect 25782 25542 25828 25594
rect 25828 25542 25838 25594
rect 25862 25542 25892 25594
rect 25892 25542 25904 25594
rect 25904 25542 25918 25594
rect 25942 25542 25956 25594
rect 25956 25542 25968 25594
rect 25968 25542 25998 25594
rect 26022 25542 26032 25594
rect 26032 25542 26078 25594
rect 25782 25540 25838 25542
rect 25862 25540 25918 25542
rect 25942 25540 25998 25542
rect 26022 25540 26078 25542
rect 25782 24506 25838 24508
rect 25862 24506 25918 24508
rect 25942 24506 25998 24508
rect 26022 24506 26078 24508
rect 25782 24454 25828 24506
rect 25828 24454 25838 24506
rect 25862 24454 25892 24506
rect 25892 24454 25904 24506
rect 25904 24454 25918 24506
rect 25942 24454 25956 24506
rect 25956 24454 25968 24506
rect 25968 24454 25998 24506
rect 26022 24454 26032 24506
rect 26032 24454 26078 24506
rect 25782 24452 25838 24454
rect 25862 24452 25918 24454
rect 25942 24452 25998 24454
rect 26022 24452 26078 24454
rect 25782 23418 25838 23420
rect 25862 23418 25918 23420
rect 25942 23418 25998 23420
rect 26022 23418 26078 23420
rect 25782 23366 25828 23418
rect 25828 23366 25838 23418
rect 25862 23366 25892 23418
rect 25892 23366 25904 23418
rect 25904 23366 25918 23418
rect 25942 23366 25956 23418
rect 25956 23366 25968 23418
rect 25968 23366 25998 23418
rect 26022 23366 26032 23418
rect 26032 23366 26078 23418
rect 25782 23364 25838 23366
rect 25862 23364 25918 23366
rect 25942 23364 25998 23366
rect 26022 23364 26078 23366
rect 25782 22330 25838 22332
rect 25862 22330 25918 22332
rect 25942 22330 25998 22332
rect 26022 22330 26078 22332
rect 25782 22278 25828 22330
rect 25828 22278 25838 22330
rect 25862 22278 25892 22330
rect 25892 22278 25904 22330
rect 25904 22278 25918 22330
rect 25942 22278 25956 22330
rect 25956 22278 25968 22330
rect 25968 22278 25998 22330
rect 26022 22278 26032 22330
rect 26032 22278 26078 22330
rect 25782 22276 25838 22278
rect 25862 22276 25918 22278
rect 25942 22276 25998 22278
rect 26022 22276 26078 22278
rect 25782 21242 25838 21244
rect 25862 21242 25918 21244
rect 25942 21242 25998 21244
rect 26022 21242 26078 21244
rect 25782 21190 25828 21242
rect 25828 21190 25838 21242
rect 25862 21190 25892 21242
rect 25892 21190 25904 21242
rect 25904 21190 25918 21242
rect 25942 21190 25956 21242
rect 25956 21190 25968 21242
rect 25968 21190 25998 21242
rect 26022 21190 26032 21242
rect 26032 21190 26078 21242
rect 25782 21188 25838 21190
rect 25862 21188 25918 21190
rect 25942 21188 25998 21190
rect 26022 21188 26078 21190
rect 25782 20154 25838 20156
rect 25862 20154 25918 20156
rect 25942 20154 25998 20156
rect 26022 20154 26078 20156
rect 25782 20102 25828 20154
rect 25828 20102 25838 20154
rect 25862 20102 25892 20154
rect 25892 20102 25904 20154
rect 25904 20102 25918 20154
rect 25942 20102 25956 20154
rect 25956 20102 25968 20154
rect 25968 20102 25998 20154
rect 26022 20102 26032 20154
rect 26032 20102 26078 20154
rect 25782 20100 25838 20102
rect 25862 20100 25918 20102
rect 25942 20100 25998 20102
rect 26022 20100 26078 20102
rect 25782 19066 25838 19068
rect 25862 19066 25918 19068
rect 25942 19066 25998 19068
rect 26022 19066 26078 19068
rect 25782 19014 25828 19066
rect 25828 19014 25838 19066
rect 25862 19014 25892 19066
rect 25892 19014 25904 19066
rect 25904 19014 25918 19066
rect 25942 19014 25956 19066
rect 25956 19014 25968 19066
rect 25968 19014 25998 19066
rect 26022 19014 26032 19066
rect 26032 19014 26078 19066
rect 25782 19012 25838 19014
rect 25862 19012 25918 19014
rect 25942 19012 25998 19014
rect 26022 19012 26078 19014
rect 25782 17978 25838 17980
rect 25862 17978 25918 17980
rect 25942 17978 25998 17980
rect 26022 17978 26078 17980
rect 25782 17926 25828 17978
rect 25828 17926 25838 17978
rect 25862 17926 25892 17978
rect 25892 17926 25904 17978
rect 25904 17926 25918 17978
rect 25942 17926 25956 17978
rect 25956 17926 25968 17978
rect 25968 17926 25998 17978
rect 26022 17926 26032 17978
rect 26032 17926 26078 17978
rect 25782 17924 25838 17926
rect 25862 17924 25918 17926
rect 25942 17924 25998 17926
rect 26022 17924 26078 17926
rect 25782 16890 25838 16892
rect 25862 16890 25918 16892
rect 25942 16890 25998 16892
rect 26022 16890 26078 16892
rect 25782 16838 25828 16890
rect 25828 16838 25838 16890
rect 25862 16838 25892 16890
rect 25892 16838 25904 16890
rect 25904 16838 25918 16890
rect 25942 16838 25956 16890
rect 25956 16838 25968 16890
rect 25968 16838 25998 16890
rect 26022 16838 26032 16890
rect 26032 16838 26078 16890
rect 25782 16836 25838 16838
rect 25862 16836 25918 16838
rect 25942 16836 25998 16838
rect 26022 16836 26078 16838
rect 25782 15802 25838 15804
rect 25862 15802 25918 15804
rect 25942 15802 25998 15804
rect 26022 15802 26078 15804
rect 25782 15750 25828 15802
rect 25828 15750 25838 15802
rect 25862 15750 25892 15802
rect 25892 15750 25904 15802
rect 25904 15750 25918 15802
rect 25942 15750 25956 15802
rect 25956 15750 25968 15802
rect 25968 15750 25998 15802
rect 26022 15750 26032 15802
rect 26032 15750 26078 15802
rect 25782 15748 25838 15750
rect 25862 15748 25918 15750
rect 25942 15748 25998 15750
rect 26022 15748 26078 15750
rect 20817 14170 20873 14172
rect 20897 14170 20953 14172
rect 20977 14170 21033 14172
rect 21057 14170 21113 14172
rect 20817 14118 20863 14170
rect 20863 14118 20873 14170
rect 20897 14118 20927 14170
rect 20927 14118 20939 14170
rect 20939 14118 20953 14170
rect 20977 14118 20991 14170
rect 20991 14118 21003 14170
rect 21003 14118 21033 14170
rect 21057 14118 21067 14170
rect 21067 14118 21113 14170
rect 20817 14116 20873 14118
rect 20897 14116 20953 14118
rect 20977 14116 21033 14118
rect 21057 14116 21113 14118
rect 20817 13082 20873 13084
rect 20897 13082 20953 13084
rect 20977 13082 21033 13084
rect 21057 13082 21113 13084
rect 20817 13030 20863 13082
rect 20863 13030 20873 13082
rect 20897 13030 20927 13082
rect 20927 13030 20939 13082
rect 20939 13030 20953 13082
rect 20977 13030 20991 13082
rect 20991 13030 21003 13082
rect 21003 13030 21033 13082
rect 21057 13030 21067 13082
rect 21067 13030 21113 13082
rect 20817 13028 20873 13030
rect 20897 13028 20953 13030
rect 20977 13028 21033 13030
rect 21057 13028 21113 13030
rect 25782 14714 25838 14716
rect 25862 14714 25918 14716
rect 25942 14714 25998 14716
rect 26022 14714 26078 14716
rect 25782 14662 25828 14714
rect 25828 14662 25838 14714
rect 25862 14662 25892 14714
rect 25892 14662 25904 14714
rect 25904 14662 25918 14714
rect 25942 14662 25956 14714
rect 25956 14662 25968 14714
rect 25968 14662 25998 14714
rect 26022 14662 26032 14714
rect 26032 14662 26078 14714
rect 25782 14660 25838 14662
rect 25862 14660 25918 14662
rect 25942 14660 25998 14662
rect 26022 14660 26078 14662
rect 25782 13626 25838 13628
rect 25862 13626 25918 13628
rect 25942 13626 25998 13628
rect 26022 13626 26078 13628
rect 25782 13574 25828 13626
rect 25828 13574 25838 13626
rect 25862 13574 25892 13626
rect 25892 13574 25904 13626
rect 25904 13574 25918 13626
rect 25942 13574 25956 13626
rect 25956 13574 25968 13626
rect 25968 13574 25998 13626
rect 26022 13574 26032 13626
rect 26032 13574 26078 13626
rect 25782 13572 25838 13574
rect 25862 13572 25918 13574
rect 25942 13572 25998 13574
rect 26022 13572 26078 13574
rect 25782 12538 25838 12540
rect 25862 12538 25918 12540
rect 25942 12538 25998 12540
rect 26022 12538 26078 12540
rect 25782 12486 25828 12538
rect 25828 12486 25838 12538
rect 25862 12486 25892 12538
rect 25892 12486 25904 12538
rect 25904 12486 25918 12538
rect 25942 12486 25956 12538
rect 25956 12486 25968 12538
rect 25968 12486 25998 12538
rect 26022 12486 26032 12538
rect 26032 12486 26078 12538
rect 25782 12484 25838 12486
rect 25862 12484 25918 12486
rect 25942 12484 25998 12486
rect 26022 12484 26078 12486
rect 20817 11994 20873 11996
rect 20897 11994 20953 11996
rect 20977 11994 21033 11996
rect 21057 11994 21113 11996
rect 20817 11942 20863 11994
rect 20863 11942 20873 11994
rect 20897 11942 20927 11994
rect 20927 11942 20939 11994
rect 20939 11942 20953 11994
rect 20977 11942 20991 11994
rect 20991 11942 21003 11994
rect 21003 11942 21033 11994
rect 21057 11942 21067 11994
rect 21067 11942 21113 11994
rect 20817 11940 20873 11942
rect 20897 11940 20953 11942
rect 20977 11940 21033 11942
rect 21057 11940 21113 11942
rect 20817 10906 20873 10908
rect 20897 10906 20953 10908
rect 20977 10906 21033 10908
rect 21057 10906 21113 10908
rect 20817 10854 20863 10906
rect 20863 10854 20873 10906
rect 20897 10854 20927 10906
rect 20927 10854 20939 10906
rect 20939 10854 20953 10906
rect 20977 10854 20991 10906
rect 20991 10854 21003 10906
rect 21003 10854 21033 10906
rect 21057 10854 21067 10906
rect 21067 10854 21113 10906
rect 20817 10852 20873 10854
rect 20897 10852 20953 10854
rect 20977 10852 21033 10854
rect 21057 10852 21113 10854
rect 20817 9818 20873 9820
rect 20897 9818 20953 9820
rect 20977 9818 21033 9820
rect 21057 9818 21113 9820
rect 20817 9766 20863 9818
rect 20863 9766 20873 9818
rect 20897 9766 20927 9818
rect 20927 9766 20939 9818
rect 20939 9766 20953 9818
rect 20977 9766 20991 9818
rect 20991 9766 21003 9818
rect 21003 9766 21033 9818
rect 21057 9766 21067 9818
rect 21067 9766 21113 9818
rect 20817 9764 20873 9766
rect 20897 9764 20953 9766
rect 20977 9764 21033 9766
rect 21057 9764 21113 9766
rect 20534 8336 20590 8392
rect 20817 8730 20873 8732
rect 20897 8730 20953 8732
rect 20977 8730 21033 8732
rect 21057 8730 21113 8732
rect 20817 8678 20863 8730
rect 20863 8678 20873 8730
rect 20897 8678 20927 8730
rect 20927 8678 20939 8730
rect 20939 8678 20953 8730
rect 20977 8678 20991 8730
rect 20991 8678 21003 8730
rect 21003 8678 21033 8730
rect 21057 8678 21067 8730
rect 21067 8678 21113 8730
rect 20817 8676 20873 8678
rect 20897 8676 20953 8678
rect 20977 8676 21033 8678
rect 21057 8676 21113 8678
rect 20817 7642 20873 7644
rect 20897 7642 20953 7644
rect 20977 7642 21033 7644
rect 21057 7642 21113 7644
rect 20817 7590 20863 7642
rect 20863 7590 20873 7642
rect 20897 7590 20927 7642
rect 20927 7590 20939 7642
rect 20939 7590 20953 7642
rect 20977 7590 20991 7642
rect 20991 7590 21003 7642
rect 21003 7590 21033 7642
rect 21057 7590 21067 7642
rect 21067 7590 21113 7642
rect 20817 7588 20873 7590
rect 20897 7588 20953 7590
rect 20977 7588 21033 7590
rect 21057 7588 21113 7590
rect 20817 6554 20873 6556
rect 20897 6554 20953 6556
rect 20977 6554 21033 6556
rect 21057 6554 21113 6556
rect 20817 6502 20863 6554
rect 20863 6502 20873 6554
rect 20897 6502 20927 6554
rect 20927 6502 20939 6554
rect 20939 6502 20953 6554
rect 20977 6502 20991 6554
rect 20991 6502 21003 6554
rect 21003 6502 21033 6554
rect 21057 6502 21067 6554
rect 21067 6502 21113 6554
rect 20817 6500 20873 6502
rect 20897 6500 20953 6502
rect 20977 6500 21033 6502
rect 21057 6500 21113 6502
rect 20817 5466 20873 5468
rect 20897 5466 20953 5468
rect 20977 5466 21033 5468
rect 21057 5466 21113 5468
rect 20817 5414 20863 5466
rect 20863 5414 20873 5466
rect 20897 5414 20927 5466
rect 20927 5414 20939 5466
rect 20939 5414 20953 5466
rect 20977 5414 20991 5466
rect 20991 5414 21003 5466
rect 21003 5414 21033 5466
rect 21057 5414 21067 5466
rect 21067 5414 21113 5466
rect 20817 5412 20873 5414
rect 20897 5412 20953 5414
rect 20977 5412 21033 5414
rect 21057 5412 21113 5414
rect 20817 4378 20873 4380
rect 20897 4378 20953 4380
rect 20977 4378 21033 4380
rect 21057 4378 21113 4380
rect 20817 4326 20863 4378
rect 20863 4326 20873 4378
rect 20897 4326 20927 4378
rect 20927 4326 20939 4378
rect 20939 4326 20953 4378
rect 20977 4326 20991 4378
rect 20991 4326 21003 4378
rect 21003 4326 21033 4378
rect 21057 4326 21067 4378
rect 21067 4326 21113 4378
rect 20817 4324 20873 4326
rect 20897 4324 20953 4326
rect 20977 4324 21033 4326
rect 21057 4324 21113 4326
rect 25782 11450 25838 11452
rect 25862 11450 25918 11452
rect 25942 11450 25998 11452
rect 26022 11450 26078 11452
rect 25782 11398 25828 11450
rect 25828 11398 25838 11450
rect 25862 11398 25892 11450
rect 25892 11398 25904 11450
rect 25904 11398 25918 11450
rect 25942 11398 25956 11450
rect 25956 11398 25968 11450
rect 25968 11398 25998 11450
rect 26022 11398 26032 11450
rect 26032 11398 26078 11450
rect 25782 11396 25838 11398
rect 25862 11396 25918 11398
rect 25942 11396 25998 11398
rect 26022 11396 26078 11398
rect 25782 10362 25838 10364
rect 25862 10362 25918 10364
rect 25942 10362 25998 10364
rect 26022 10362 26078 10364
rect 25782 10310 25828 10362
rect 25828 10310 25838 10362
rect 25862 10310 25892 10362
rect 25892 10310 25904 10362
rect 25904 10310 25918 10362
rect 25942 10310 25956 10362
rect 25956 10310 25968 10362
rect 25968 10310 25998 10362
rect 26022 10310 26032 10362
rect 26032 10310 26078 10362
rect 25782 10308 25838 10310
rect 25862 10308 25918 10310
rect 25942 10308 25998 10310
rect 26022 10308 26078 10310
rect 25782 9274 25838 9276
rect 25862 9274 25918 9276
rect 25942 9274 25998 9276
rect 26022 9274 26078 9276
rect 25782 9222 25828 9274
rect 25828 9222 25838 9274
rect 25862 9222 25892 9274
rect 25892 9222 25904 9274
rect 25904 9222 25918 9274
rect 25942 9222 25956 9274
rect 25956 9222 25968 9274
rect 25968 9222 25998 9274
rect 26022 9222 26032 9274
rect 26032 9222 26078 9274
rect 25782 9220 25838 9222
rect 25862 9220 25918 9222
rect 25942 9220 25998 9222
rect 26022 9220 26078 9222
rect 22282 8336 22338 8392
rect 20817 3290 20873 3292
rect 20897 3290 20953 3292
rect 20977 3290 21033 3292
rect 21057 3290 21113 3292
rect 20817 3238 20863 3290
rect 20863 3238 20873 3290
rect 20897 3238 20927 3290
rect 20927 3238 20939 3290
rect 20939 3238 20953 3290
rect 20977 3238 20991 3290
rect 20991 3238 21003 3290
rect 21003 3238 21033 3290
rect 21057 3238 21067 3290
rect 21067 3238 21113 3290
rect 20817 3236 20873 3238
rect 20897 3236 20953 3238
rect 20977 3236 21033 3238
rect 21057 3236 21113 3238
rect 20817 2202 20873 2204
rect 20897 2202 20953 2204
rect 20977 2202 21033 2204
rect 21057 2202 21113 2204
rect 20817 2150 20863 2202
rect 20863 2150 20873 2202
rect 20897 2150 20927 2202
rect 20927 2150 20939 2202
rect 20939 2150 20953 2202
rect 20977 2150 20991 2202
rect 20991 2150 21003 2202
rect 21003 2150 21033 2202
rect 21057 2150 21067 2202
rect 21067 2150 21113 2202
rect 20817 2148 20873 2150
rect 20897 2148 20953 2150
rect 20977 2148 21033 2150
rect 21057 2148 21113 2150
rect 2962 312 3018 368
rect 25782 8186 25838 8188
rect 25862 8186 25918 8188
rect 25942 8186 25998 8188
rect 26022 8186 26078 8188
rect 25782 8134 25828 8186
rect 25828 8134 25838 8186
rect 25862 8134 25892 8186
rect 25892 8134 25904 8186
rect 25904 8134 25918 8186
rect 25942 8134 25956 8186
rect 25956 8134 25968 8186
rect 25968 8134 25998 8186
rect 26022 8134 26032 8186
rect 26032 8134 26078 8186
rect 25782 8132 25838 8134
rect 25862 8132 25918 8134
rect 25942 8132 25998 8134
rect 26022 8132 26078 8134
rect 25782 7098 25838 7100
rect 25862 7098 25918 7100
rect 25942 7098 25998 7100
rect 26022 7098 26078 7100
rect 25782 7046 25828 7098
rect 25828 7046 25838 7098
rect 25862 7046 25892 7098
rect 25892 7046 25904 7098
rect 25904 7046 25918 7098
rect 25942 7046 25956 7098
rect 25956 7046 25968 7098
rect 25968 7046 25998 7098
rect 26022 7046 26032 7098
rect 26032 7046 26078 7098
rect 25782 7044 25838 7046
rect 25862 7044 25918 7046
rect 25942 7044 25998 7046
rect 26022 7044 26078 7046
rect 25782 6010 25838 6012
rect 25862 6010 25918 6012
rect 25942 6010 25998 6012
rect 26022 6010 26078 6012
rect 25782 5958 25828 6010
rect 25828 5958 25838 6010
rect 25862 5958 25892 6010
rect 25892 5958 25904 6010
rect 25904 5958 25918 6010
rect 25942 5958 25956 6010
rect 25956 5958 25968 6010
rect 25968 5958 25998 6010
rect 26022 5958 26032 6010
rect 26032 5958 26078 6010
rect 25782 5956 25838 5958
rect 25862 5956 25918 5958
rect 25942 5956 25998 5958
rect 26022 5956 26078 5958
rect 25782 4922 25838 4924
rect 25862 4922 25918 4924
rect 25942 4922 25998 4924
rect 26022 4922 26078 4924
rect 25782 4870 25828 4922
rect 25828 4870 25838 4922
rect 25862 4870 25892 4922
rect 25892 4870 25904 4922
rect 25904 4870 25918 4922
rect 25942 4870 25956 4922
rect 25956 4870 25968 4922
rect 25968 4870 25998 4922
rect 26022 4870 26032 4922
rect 26032 4870 26078 4922
rect 25782 4868 25838 4870
rect 25862 4868 25918 4870
rect 25942 4868 25998 4870
rect 26022 4868 26078 4870
rect 25782 3834 25838 3836
rect 25862 3834 25918 3836
rect 25942 3834 25998 3836
rect 26022 3834 26078 3836
rect 25782 3782 25828 3834
rect 25828 3782 25838 3834
rect 25862 3782 25892 3834
rect 25892 3782 25904 3834
rect 25904 3782 25918 3834
rect 25942 3782 25956 3834
rect 25956 3782 25968 3834
rect 25968 3782 25998 3834
rect 26022 3782 26032 3834
rect 26032 3782 26078 3834
rect 25782 3780 25838 3782
rect 25862 3780 25918 3782
rect 25942 3780 25998 3782
rect 26022 3780 26078 3782
rect 25782 2746 25838 2748
rect 25862 2746 25918 2748
rect 25942 2746 25998 2748
rect 26022 2746 26078 2748
rect 25782 2694 25828 2746
rect 25828 2694 25838 2746
rect 25862 2694 25892 2746
rect 25892 2694 25904 2746
rect 25904 2694 25918 2746
rect 25942 2694 25956 2746
rect 25956 2694 25968 2746
rect 25968 2694 25998 2746
rect 26022 2694 26032 2746
rect 26032 2694 26078 2746
rect 25782 2692 25838 2694
rect 25862 2692 25918 2694
rect 25942 2692 25998 2694
rect 26022 2692 26078 2694
rect 30010 28872 30066 28928
rect 30010 26968 30066 27024
rect 30010 24928 30066 24984
rect 30010 22924 30012 22944
rect 30012 22924 30064 22944
rect 30064 22924 30066 22944
rect 30010 22888 30066 22924
rect 30010 20984 30066 21040
rect 30010 18944 30066 19000
rect 30010 16940 30012 16960
rect 30012 16940 30064 16960
rect 30064 16940 30066 16960
rect 30010 16904 30066 16940
rect 30010 14884 30066 14920
rect 30010 14864 30012 14884
rect 30012 14864 30064 14884
rect 30064 14864 30066 14884
rect 30010 12960 30066 13016
rect 30010 10956 30012 10976
rect 30012 10956 30064 10976
rect 30064 10956 30066 10976
rect 30010 10920 30066 10956
rect 30010 8880 30066 8936
rect 30010 6976 30066 7032
rect 30010 4972 30012 4992
rect 30012 4972 30064 4992
rect 30064 4972 30066 4992
rect 30010 4936 30066 4972
rect 28906 992 28962 1048
rect 30010 2896 30066 2952
<< metal3 >>
rect 0 47562 800 47592
rect 2773 47562 2839 47565
rect 0 47560 2839 47562
rect 0 47504 2778 47560
rect 2834 47504 2839 47560
rect 0 47502 2839 47504
rect 0 47472 800 47502
rect 2773 47499 2839 47502
rect 30005 47018 30071 47021
rect 31200 47018 32000 47048
rect 30005 47016 32000 47018
rect 30005 46960 30010 47016
rect 30066 46960 32000 47016
rect 30005 46958 32000 46960
rect 30005 46955 30071 46958
rect 31200 46928 32000 46958
rect 0 46882 800 46912
rect 2865 46882 2931 46885
rect 0 46880 2931 46882
rect 0 46824 2870 46880
rect 2926 46824 2931 46880
rect 0 46822 2931 46824
rect 0 46792 800 46822
rect 2865 46819 2931 46822
rect 0 46066 800 46096
rect 2957 46066 3023 46069
rect 0 46064 3023 46066
rect 0 46008 2962 46064
rect 3018 46008 3023 46064
rect 0 46006 3023 46008
rect 0 45976 800 46006
rect 2957 46003 3023 46006
rect 10874 45728 11194 45729
rect 10874 45664 10882 45728
rect 10946 45664 10962 45728
rect 11026 45664 11042 45728
rect 11106 45664 11122 45728
rect 11186 45664 11194 45728
rect 10874 45663 11194 45664
rect 20805 45728 21125 45729
rect 20805 45664 20813 45728
rect 20877 45664 20893 45728
rect 20957 45664 20973 45728
rect 21037 45664 21053 45728
rect 21117 45664 21125 45728
rect 20805 45663 21125 45664
rect 0 45386 800 45416
rect 2221 45386 2287 45389
rect 0 45384 2287 45386
rect 0 45328 2226 45384
rect 2282 45328 2287 45384
rect 0 45326 2287 45328
rect 0 45296 800 45326
rect 2221 45323 2287 45326
rect 5909 45184 6229 45185
rect 5909 45120 5917 45184
rect 5981 45120 5997 45184
rect 6061 45120 6077 45184
rect 6141 45120 6157 45184
rect 6221 45120 6229 45184
rect 5909 45119 6229 45120
rect 15840 45184 16160 45185
rect 15840 45120 15848 45184
rect 15912 45120 15928 45184
rect 15992 45120 16008 45184
rect 16072 45120 16088 45184
rect 16152 45120 16160 45184
rect 15840 45119 16160 45120
rect 25770 45184 26090 45185
rect 25770 45120 25778 45184
rect 25842 45120 25858 45184
rect 25922 45120 25938 45184
rect 26002 45120 26018 45184
rect 26082 45120 26090 45184
rect 25770 45119 26090 45120
rect 30097 44978 30163 44981
rect 31200 44978 32000 45008
rect 30097 44976 32000 44978
rect 30097 44920 30102 44976
rect 30158 44920 32000 44976
rect 30097 44918 32000 44920
rect 30097 44915 30163 44918
rect 31200 44888 32000 44918
rect 2405 44842 2471 44845
rect 8017 44842 8083 44845
rect 2405 44840 8083 44842
rect 2405 44784 2410 44840
rect 2466 44784 8022 44840
rect 8078 44784 8083 44840
rect 2405 44782 8083 44784
rect 2405 44779 2471 44782
rect 8017 44779 8083 44782
rect 10874 44640 11194 44641
rect 0 44570 800 44600
rect 10874 44576 10882 44640
rect 10946 44576 10962 44640
rect 11026 44576 11042 44640
rect 11106 44576 11122 44640
rect 11186 44576 11194 44640
rect 10874 44575 11194 44576
rect 20805 44640 21125 44641
rect 20805 44576 20813 44640
rect 20877 44576 20893 44640
rect 20957 44576 20973 44640
rect 21037 44576 21053 44640
rect 21117 44576 21125 44640
rect 20805 44575 21125 44576
rect 1485 44570 1551 44573
rect 0 44568 1551 44570
rect 0 44512 1490 44568
rect 1546 44512 1551 44568
rect 0 44510 1551 44512
rect 0 44480 800 44510
rect 1485 44507 1551 44510
rect 4429 44570 4495 44573
rect 8201 44570 8267 44573
rect 4429 44568 8267 44570
rect 4429 44512 4434 44568
rect 4490 44512 8206 44568
rect 8262 44512 8267 44568
rect 4429 44510 8267 44512
rect 4429 44507 4495 44510
rect 8201 44507 8267 44510
rect 5909 44096 6229 44097
rect 5909 44032 5917 44096
rect 5981 44032 5997 44096
rect 6061 44032 6077 44096
rect 6141 44032 6157 44096
rect 6221 44032 6229 44096
rect 5909 44031 6229 44032
rect 15840 44096 16160 44097
rect 15840 44032 15848 44096
rect 15912 44032 15928 44096
rect 15992 44032 16008 44096
rect 16072 44032 16088 44096
rect 16152 44032 16160 44096
rect 15840 44031 16160 44032
rect 25770 44096 26090 44097
rect 25770 44032 25778 44096
rect 25842 44032 25858 44096
rect 25922 44032 25938 44096
rect 26002 44032 26018 44096
rect 26082 44032 26090 44096
rect 25770 44031 26090 44032
rect 0 43890 800 43920
rect 1485 43890 1551 43893
rect 0 43888 1551 43890
rect 0 43832 1490 43888
rect 1546 43832 1551 43888
rect 0 43830 1551 43832
rect 0 43800 800 43830
rect 1485 43827 1551 43830
rect 10874 43552 11194 43553
rect 10874 43488 10882 43552
rect 10946 43488 10962 43552
rect 11026 43488 11042 43552
rect 11106 43488 11122 43552
rect 11186 43488 11194 43552
rect 10874 43487 11194 43488
rect 20805 43552 21125 43553
rect 20805 43488 20813 43552
rect 20877 43488 20893 43552
rect 20957 43488 20973 43552
rect 21037 43488 21053 43552
rect 21117 43488 21125 43552
rect 20805 43487 21125 43488
rect 0 43074 800 43104
rect 1485 43074 1551 43077
rect 0 43072 1551 43074
rect 0 43016 1490 43072
rect 1546 43016 1551 43072
rect 0 43014 1551 43016
rect 0 42984 800 43014
rect 1485 43011 1551 43014
rect 5909 43008 6229 43009
rect 5909 42944 5917 43008
rect 5981 42944 5997 43008
rect 6061 42944 6077 43008
rect 6141 42944 6157 43008
rect 6221 42944 6229 43008
rect 5909 42943 6229 42944
rect 15840 43008 16160 43009
rect 15840 42944 15848 43008
rect 15912 42944 15928 43008
rect 15992 42944 16008 43008
rect 16072 42944 16088 43008
rect 16152 42944 16160 43008
rect 15840 42943 16160 42944
rect 25770 43008 26090 43009
rect 25770 42944 25778 43008
rect 25842 42944 25858 43008
rect 25922 42944 25938 43008
rect 26002 42944 26018 43008
rect 26082 42944 26090 43008
rect 25770 42943 26090 42944
rect 30097 42938 30163 42941
rect 31200 42938 32000 42968
rect 30097 42936 32000 42938
rect 30097 42880 30102 42936
rect 30158 42880 32000 42936
rect 30097 42878 32000 42880
rect 30097 42875 30163 42878
rect 31200 42848 32000 42878
rect 10874 42464 11194 42465
rect 0 42394 800 42424
rect 10874 42400 10882 42464
rect 10946 42400 10962 42464
rect 11026 42400 11042 42464
rect 11106 42400 11122 42464
rect 11186 42400 11194 42464
rect 10874 42399 11194 42400
rect 20805 42464 21125 42465
rect 20805 42400 20813 42464
rect 20877 42400 20893 42464
rect 20957 42400 20973 42464
rect 21037 42400 21053 42464
rect 21117 42400 21125 42464
rect 20805 42399 21125 42400
rect 1393 42394 1459 42397
rect 0 42392 1459 42394
rect 0 42336 1398 42392
rect 1454 42336 1459 42392
rect 0 42334 1459 42336
rect 0 42304 800 42334
rect 1393 42331 1459 42334
rect 5909 41920 6229 41921
rect 5909 41856 5917 41920
rect 5981 41856 5997 41920
rect 6061 41856 6077 41920
rect 6141 41856 6157 41920
rect 6221 41856 6229 41920
rect 5909 41855 6229 41856
rect 15840 41920 16160 41921
rect 15840 41856 15848 41920
rect 15912 41856 15928 41920
rect 15992 41856 16008 41920
rect 16072 41856 16088 41920
rect 16152 41856 16160 41920
rect 15840 41855 16160 41856
rect 25770 41920 26090 41921
rect 25770 41856 25778 41920
rect 25842 41856 25858 41920
rect 25922 41856 25938 41920
rect 26002 41856 26018 41920
rect 26082 41856 26090 41920
rect 25770 41855 26090 41856
rect 0 41714 800 41744
rect 1485 41714 1551 41717
rect 0 41712 1551 41714
rect 0 41656 1490 41712
rect 1546 41656 1551 41712
rect 0 41654 1551 41656
rect 0 41624 800 41654
rect 1485 41651 1551 41654
rect 10874 41376 11194 41377
rect 10874 41312 10882 41376
rect 10946 41312 10962 41376
rect 11026 41312 11042 41376
rect 11106 41312 11122 41376
rect 11186 41312 11194 41376
rect 10874 41311 11194 41312
rect 20805 41376 21125 41377
rect 20805 41312 20813 41376
rect 20877 41312 20893 41376
rect 20957 41312 20973 41376
rect 21037 41312 21053 41376
rect 21117 41312 21125 41376
rect 20805 41311 21125 41312
rect 30097 41034 30163 41037
rect 31200 41034 32000 41064
rect 30097 41032 32000 41034
rect 30097 40976 30102 41032
rect 30158 40976 32000 41032
rect 30097 40974 32000 40976
rect 30097 40971 30163 40974
rect 31200 40944 32000 40974
rect 0 40898 800 40928
rect 1393 40898 1459 40901
rect 0 40896 1459 40898
rect 0 40840 1398 40896
rect 1454 40840 1459 40896
rect 0 40838 1459 40840
rect 0 40808 800 40838
rect 1393 40835 1459 40838
rect 5909 40832 6229 40833
rect 5909 40768 5917 40832
rect 5981 40768 5997 40832
rect 6061 40768 6077 40832
rect 6141 40768 6157 40832
rect 6221 40768 6229 40832
rect 5909 40767 6229 40768
rect 15840 40832 16160 40833
rect 15840 40768 15848 40832
rect 15912 40768 15928 40832
rect 15992 40768 16008 40832
rect 16072 40768 16088 40832
rect 16152 40768 16160 40832
rect 15840 40767 16160 40768
rect 25770 40832 26090 40833
rect 25770 40768 25778 40832
rect 25842 40768 25858 40832
rect 25922 40768 25938 40832
rect 26002 40768 26018 40832
rect 26082 40768 26090 40832
rect 25770 40767 26090 40768
rect 3509 40626 3575 40629
rect 4245 40626 4311 40629
rect 4797 40626 4863 40629
rect 3509 40624 4863 40626
rect 3509 40568 3514 40624
rect 3570 40568 4250 40624
rect 4306 40568 4802 40624
rect 4858 40568 4863 40624
rect 3509 40566 4863 40568
rect 3509 40563 3575 40566
rect 4245 40563 4311 40566
rect 4797 40563 4863 40566
rect 10874 40288 11194 40289
rect 0 40218 800 40248
rect 10874 40224 10882 40288
rect 10946 40224 10962 40288
rect 11026 40224 11042 40288
rect 11106 40224 11122 40288
rect 11186 40224 11194 40288
rect 10874 40223 11194 40224
rect 20805 40288 21125 40289
rect 20805 40224 20813 40288
rect 20877 40224 20893 40288
rect 20957 40224 20973 40288
rect 21037 40224 21053 40288
rect 21117 40224 21125 40288
rect 20805 40223 21125 40224
rect 1301 40218 1367 40221
rect 0 40216 1367 40218
rect 0 40160 1306 40216
rect 1362 40160 1367 40216
rect 0 40158 1367 40160
rect 0 40128 800 40158
rect 1301 40155 1367 40158
rect 5909 39744 6229 39745
rect 5909 39680 5917 39744
rect 5981 39680 5997 39744
rect 6061 39680 6077 39744
rect 6141 39680 6157 39744
rect 6221 39680 6229 39744
rect 5909 39679 6229 39680
rect 15840 39744 16160 39745
rect 15840 39680 15848 39744
rect 15912 39680 15928 39744
rect 15992 39680 16008 39744
rect 16072 39680 16088 39744
rect 16152 39680 16160 39744
rect 15840 39679 16160 39680
rect 25770 39744 26090 39745
rect 25770 39680 25778 39744
rect 25842 39680 25858 39744
rect 25922 39680 25938 39744
rect 26002 39680 26018 39744
rect 26082 39680 26090 39744
rect 25770 39679 26090 39680
rect 0 39402 800 39432
rect 1485 39402 1551 39405
rect 0 39400 1551 39402
rect 0 39344 1490 39400
rect 1546 39344 1551 39400
rect 0 39342 1551 39344
rect 0 39312 800 39342
rect 1485 39339 1551 39342
rect 10874 39200 11194 39201
rect 10874 39136 10882 39200
rect 10946 39136 10962 39200
rect 11026 39136 11042 39200
rect 11106 39136 11122 39200
rect 11186 39136 11194 39200
rect 10874 39135 11194 39136
rect 20805 39200 21125 39201
rect 20805 39136 20813 39200
rect 20877 39136 20893 39200
rect 20957 39136 20973 39200
rect 21037 39136 21053 39200
rect 21117 39136 21125 39200
rect 20805 39135 21125 39136
rect 30097 38994 30163 38997
rect 31200 38994 32000 39024
rect 30097 38992 32000 38994
rect 30097 38936 30102 38992
rect 30158 38936 32000 38992
rect 30097 38934 32000 38936
rect 30097 38931 30163 38934
rect 31200 38904 32000 38934
rect 0 38722 800 38752
rect 1393 38722 1459 38725
rect 0 38720 1459 38722
rect 0 38664 1398 38720
rect 1454 38664 1459 38720
rect 0 38662 1459 38664
rect 0 38632 800 38662
rect 1393 38659 1459 38662
rect 5909 38656 6229 38657
rect 5909 38592 5917 38656
rect 5981 38592 5997 38656
rect 6061 38592 6077 38656
rect 6141 38592 6157 38656
rect 6221 38592 6229 38656
rect 5909 38591 6229 38592
rect 15840 38656 16160 38657
rect 15840 38592 15848 38656
rect 15912 38592 15928 38656
rect 15992 38592 16008 38656
rect 16072 38592 16088 38656
rect 16152 38592 16160 38656
rect 15840 38591 16160 38592
rect 25770 38656 26090 38657
rect 25770 38592 25778 38656
rect 25842 38592 25858 38656
rect 25922 38592 25938 38656
rect 26002 38592 26018 38656
rect 26082 38592 26090 38656
rect 25770 38591 26090 38592
rect 10874 38112 11194 38113
rect 10874 38048 10882 38112
rect 10946 38048 10962 38112
rect 11026 38048 11042 38112
rect 11106 38048 11122 38112
rect 11186 38048 11194 38112
rect 10874 38047 11194 38048
rect 20805 38112 21125 38113
rect 20805 38048 20813 38112
rect 20877 38048 20893 38112
rect 20957 38048 20973 38112
rect 21037 38048 21053 38112
rect 21117 38048 21125 38112
rect 20805 38047 21125 38048
rect 0 37906 800 37936
rect 3141 37906 3207 37909
rect 0 37904 3207 37906
rect 0 37848 3146 37904
rect 3202 37848 3207 37904
rect 0 37846 3207 37848
rect 0 37816 800 37846
rect 3141 37843 3207 37846
rect 5909 37568 6229 37569
rect 5909 37504 5917 37568
rect 5981 37504 5997 37568
rect 6061 37504 6077 37568
rect 6141 37504 6157 37568
rect 6221 37504 6229 37568
rect 5909 37503 6229 37504
rect 15840 37568 16160 37569
rect 15840 37504 15848 37568
rect 15912 37504 15928 37568
rect 15992 37504 16008 37568
rect 16072 37504 16088 37568
rect 16152 37504 16160 37568
rect 15840 37503 16160 37504
rect 25770 37568 26090 37569
rect 25770 37504 25778 37568
rect 25842 37504 25858 37568
rect 25922 37504 25938 37568
rect 26002 37504 26018 37568
rect 26082 37504 26090 37568
rect 25770 37503 26090 37504
rect 0 37226 800 37256
rect 3141 37226 3207 37229
rect 0 37224 3207 37226
rect 0 37168 3146 37224
rect 3202 37168 3207 37224
rect 0 37166 3207 37168
rect 0 37136 800 37166
rect 3141 37163 3207 37166
rect 10874 37024 11194 37025
rect 10874 36960 10882 37024
rect 10946 36960 10962 37024
rect 11026 36960 11042 37024
rect 11106 36960 11122 37024
rect 11186 36960 11194 37024
rect 10874 36959 11194 36960
rect 20805 37024 21125 37025
rect 20805 36960 20813 37024
rect 20877 36960 20893 37024
rect 20957 36960 20973 37024
rect 21037 36960 21053 37024
rect 21117 36960 21125 37024
rect 20805 36959 21125 36960
rect 30097 36954 30163 36957
rect 31200 36954 32000 36984
rect 30097 36952 32000 36954
rect 30097 36896 30102 36952
rect 30158 36896 32000 36952
rect 30097 36894 32000 36896
rect 30097 36891 30163 36894
rect 31200 36864 32000 36894
rect 0 36546 800 36576
rect 1485 36546 1551 36549
rect 0 36544 1551 36546
rect 0 36488 1490 36544
rect 1546 36488 1551 36544
rect 0 36486 1551 36488
rect 0 36456 800 36486
rect 1485 36483 1551 36486
rect 5909 36480 6229 36481
rect 5909 36416 5917 36480
rect 5981 36416 5997 36480
rect 6061 36416 6077 36480
rect 6141 36416 6157 36480
rect 6221 36416 6229 36480
rect 5909 36415 6229 36416
rect 15840 36480 16160 36481
rect 15840 36416 15848 36480
rect 15912 36416 15928 36480
rect 15992 36416 16008 36480
rect 16072 36416 16088 36480
rect 16152 36416 16160 36480
rect 15840 36415 16160 36416
rect 25770 36480 26090 36481
rect 25770 36416 25778 36480
rect 25842 36416 25858 36480
rect 25922 36416 25938 36480
rect 26002 36416 26018 36480
rect 26082 36416 26090 36480
rect 25770 36415 26090 36416
rect 10874 35936 11194 35937
rect 10874 35872 10882 35936
rect 10946 35872 10962 35936
rect 11026 35872 11042 35936
rect 11106 35872 11122 35936
rect 11186 35872 11194 35936
rect 10874 35871 11194 35872
rect 20805 35936 21125 35937
rect 20805 35872 20813 35936
rect 20877 35872 20893 35936
rect 20957 35872 20973 35936
rect 21037 35872 21053 35936
rect 21117 35872 21125 35936
rect 20805 35871 21125 35872
rect 0 35730 800 35760
rect 2221 35730 2287 35733
rect 0 35728 2287 35730
rect 0 35672 2226 35728
rect 2282 35672 2287 35728
rect 0 35670 2287 35672
rect 0 35640 800 35670
rect 2221 35667 2287 35670
rect 5909 35392 6229 35393
rect 5909 35328 5917 35392
rect 5981 35328 5997 35392
rect 6061 35328 6077 35392
rect 6141 35328 6157 35392
rect 6221 35328 6229 35392
rect 5909 35327 6229 35328
rect 15840 35392 16160 35393
rect 15840 35328 15848 35392
rect 15912 35328 15928 35392
rect 15992 35328 16008 35392
rect 16072 35328 16088 35392
rect 16152 35328 16160 35392
rect 15840 35327 16160 35328
rect 25770 35392 26090 35393
rect 25770 35328 25778 35392
rect 25842 35328 25858 35392
rect 25922 35328 25938 35392
rect 26002 35328 26018 35392
rect 26082 35328 26090 35392
rect 25770 35327 26090 35328
rect 0 35050 800 35080
rect 1485 35050 1551 35053
rect 0 35048 1551 35050
rect 0 34992 1490 35048
rect 1546 34992 1551 35048
rect 0 34990 1551 34992
rect 0 34960 800 34990
rect 1485 34987 1551 34990
rect 30097 35050 30163 35053
rect 31200 35050 32000 35080
rect 30097 35048 32000 35050
rect 30097 34992 30102 35048
rect 30158 34992 32000 35048
rect 30097 34990 32000 34992
rect 30097 34987 30163 34990
rect 31200 34960 32000 34990
rect 10874 34848 11194 34849
rect 10874 34784 10882 34848
rect 10946 34784 10962 34848
rect 11026 34784 11042 34848
rect 11106 34784 11122 34848
rect 11186 34784 11194 34848
rect 10874 34783 11194 34784
rect 20805 34848 21125 34849
rect 20805 34784 20813 34848
rect 20877 34784 20893 34848
rect 20957 34784 20973 34848
rect 21037 34784 21053 34848
rect 21117 34784 21125 34848
rect 20805 34783 21125 34784
rect 6637 34642 6703 34645
rect 8937 34642 9003 34645
rect 6637 34640 9003 34642
rect 6637 34584 6642 34640
rect 6698 34584 8942 34640
rect 8998 34584 9003 34640
rect 6637 34582 9003 34584
rect 6637 34579 6703 34582
rect 8937 34579 9003 34582
rect 5909 34304 6229 34305
rect 0 34234 800 34264
rect 5909 34240 5917 34304
rect 5981 34240 5997 34304
rect 6061 34240 6077 34304
rect 6141 34240 6157 34304
rect 6221 34240 6229 34304
rect 5909 34239 6229 34240
rect 15840 34304 16160 34305
rect 15840 34240 15848 34304
rect 15912 34240 15928 34304
rect 15992 34240 16008 34304
rect 16072 34240 16088 34304
rect 16152 34240 16160 34304
rect 15840 34239 16160 34240
rect 25770 34304 26090 34305
rect 25770 34240 25778 34304
rect 25842 34240 25858 34304
rect 25922 34240 25938 34304
rect 26002 34240 26018 34304
rect 26082 34240 26090 34304
rect 25770 34239 26090 34240
rect 3049 34234 3115 34237
rect 0 34232 3115 34234
rect 0 34176 3054 34232
rect 3110 34176 3115 34232
rect 0 34174 3115 34176
rect 0 34144 800 34174
rect 3049 34171 3115 34174
rect 6177 34098 6243 34101
rect 8293 34098 8359 34101
rect 6177 34096 8359 34098
rect 6177 34040 6182 34096
rect 6238 34040 8298 34096
rect 8354 34040 8359 34096
rect 6177 34038 8359 34040
rect 6177 34035 6243 34038
rect 8293 34035 8359 34038
rect 10874 33760 11194 33761
rect 10874 33696 10882 33760
rect 10946 33696 10962 33760
rect 11026 33696 11042 33760
rect 11106 33696 11122 33760
rect 11186 33696 11194 33760
rect 10874 33695 11194 33696
rect 20805 33760 21125 33761
rect 20805 33696 20813 33760
rect 20877 33696 20893 33760
rect 20957 33696 20973 33760
rect 21037 33696 21053 33760
rect 21117 33696 21125 33760
rect 20805 33695 21125 33696
rect 0 33554 800 33584
rect 2957 33554 3023 33557
rect 0 33552 3023 33554
rect 0 33496 2962 33552
rect 3018 33496 3023 33552
rect 0 33494 3023 33496
rect 0 33464 800 33494
rect 2957 33491 3023 33494
rect 10041 33418 10107 33421
rect 16941 33418 17007 33421
rect 10041 33416 17007 33418
rect 10041 33360 10046 33416
rect 10102 33360 16946 33416
rect 17002 33360 17007 33416
rect 10041 33358 17007 33360
rect 10041 33355 10107 33358
rect 16941 33355 17007 33358
rect 5909 33216 6229 33217
rect 5909 33152 5917 33216
rect 5981 33152 5997 33216
rect 6061 33152 6077 33216
rect 6141 33152 6157 33216
rect 6221 33152 6229 33216
rect 5909 33151 6229 33152
rect 15840 33216 16160 33217
rect 15840 33152 15848 33216
rect 15912 33152 15928 33216
rect 15992 33152 16008 33216
rect 16072 33152 16088 33216
rect 16152 33152 16160 33216
rect 15840 33151 16160 33152
rect 25770 33216 26090 33217
rect 25770 33152 25778 33216
rect 25842 33152 25858 33216
rect 25922 33152 25938 33216
rect 26002 33152 26018 33216
rect 26082 33152 26090 33216
rect 25770 33151 26090 33152
rect 30097 33010 30163 33013
rect 31200 33010 32000 33040
rect 30097 33008 32000 33010
rect 30097 32952 30102 33008
rect 30158 32952 32000 33008
rect 30097 32950 32000 32952
rect 30097 32947 30163 32950
rect 31200 32920 32000 32950
rect 0 32738 800 32768
rect 1485 32738 1551 32741
rect 0 32736 1551 32738
rect 0 32680 1490 32736
rect 1546 32680 1551 32736
rect 0 32678 1551 32680
rect 0 32648 800 32678
rect 1485 32675 1551 32678
rect 10874 32672 11194 32673
rect 10874 32608 10882 32672
rect 10946 32608 10962 32672
rect 11026 32608 11042 32672
rect 11106 32608 11122 32672
rect 11186 32608 11194 32672
rect 10874 32607 11194 32608
rect 20805 32672 21125 32673
rect 20805 32608 20813 32672
rect 20877 32608 20893 32672
rect 20957 32608 20973 32672
rect 21037 32608 21053 32672
rect 21117 32608 21125 32672
rect 20805 32607 21125 32608
rect 5909 32128 6229 32129
rect 0 32058 800 32088
rect 5909 32064 5917 32128
rect 5981 32064 5997 32128
rect 6061 32064 6077 32128
rect 6141 32064 6157 32128
rect 6221 32064 6229 32128
rect 5909 32063 6229 32064
rect 15840 32128 16160 32129
rect 15840 32064 15848 32128
rect 15912 32064 15928 32128
rect 15992 32064 16008 32128
rect 16072 32064 16088 32128
rect 16152 32064 16160 32128
rect 15840 32063 16160 32064
rect 25770 32128 26090 32129
rect 25770 32064 25778 32128
rect 25842 32064 25858 32128
rect 25922 32064 25938 32128
rect 26002 32064 26018 32128
rect 26082 32064 26090 32128
rect 25770 32063 26090 32064
rect 1577 32058 1643 32061
rect 0 32056 1643 32058
rect 0 32000 1582 32056
rect 1638 32000 1643 32056
rect 0 31998 1643 32000
rect 0 31968 800 31998
rect 1577 31995 1643 31998
rect 11278 31724 11284 31788
rect 11348 31786 11354 31788
rect 11513 31786 11579 31789
rect 11348 31784 11579 31786
rect 11348 31728 11518 31784
rect 11574 31728 11579 31784
rect 11348 31726 11579 31728
rect 11348 31724 11354 31726
rect 11513 31723 11579 31726
rect 10874 31584 11194 31585
rect 10874 31520 10882 31584
rect 10946 31520 10962 31584
rect 11026 31520 11042 31584
rect 11106 31520 11122 31584
rect 11186 31520 11194 31584
rect 10874 31519 11194 31520
rect 20805 31584 21125 31585
rect 20805 31520 20813 31584
rect 20877 31520 20893 31584
rect 20957 31520 20973 31584
rect 21037 31520 21053 31584
rect 21117 31520 21125 31584
rect 20805 31519 21125 31520
rect 0 31378 800 31408
rect 1485 31378 1551 31381
rect 0 31376 1551 31378
rect 0 31320 1490 31376
rect 1546 31320 1551 31376
rect 0 31318 1551 31320
rect 0 31288 800 31318
rect 1485 31315 1551 31318
rect 5909 31040 6229 31041
rect 5909 30976 5917 31040
rect 5981 30976 5997 31040
rect 6061 30976 6077 31040
rect 6141 30976 6157 31040
rect 6221 30976 6229 31040
rect 5909 30975 6229 30976
rect 15840 31040 16160 31041
rect 15840 30976 15848 31040
rect 15912 30976 15928 31040
rect 15992 30976 16008 31040
rect 16072 30976 16088 31040
rect 16152 30976 16160 31040
rect 15840 30975 16160 30976
rect 25770 31040 26090 31041
rect 25770 30976 25778 31040
rect 25842 30976 25858 31040
rect 25922 30976 25938 31040
rect 26002 30976 26018 31040
rect 26082 30976 26090 31040
rect 25770 30975 26090 30976
rect 30097 30970 30163 30973
rect 31200 30970 32000 31000
rect 30097 30968 32000 30970
rect 30097 30912 30102 30968
rect 30158 30912 32000 30968
rect 30097 30910 32000 30912
rect 30097 30907 30163 30910
rect 31200 30880 32000 30910
rect 0 30562 800 30592
rect 3969 30562 4035 30565
rect 0 30560 4035 30562
rect 0 30504 3974 30560
rect 4030 30504 4035 30560
rect 0 30502 4035 30504
rect 0 30472 800 30502
rect 3969 30499 4035 30502
rect 10874 30496 11194 30497
rect 10874 30432 10882 30496
rect 10946 30432 10962 30496
rect 11026 30432 11042 30496
rect 11106 30432 11122 30496
rect 11186 30432 11194 30496
rect 10874 30431 11194 30432
rect 20805 30496 21125 30497
rect 20805 30432 20813 30496
rect 20877 30432 20893 30496
rect 20957 30432 20973 30496
rect 21037 30432 21053 30496
rect 21117 30432 21125 30496
rect 20805 30431 21125 30432
rect 5909 29952 6229 29953
rect 0 29882 800 29912
rect 5909 29888 5917 29952
rect 5981 29888 5997 29952
rect 6061 29888 6077 29952
rect 6141 29888 6157 29952
rect 6221 29888 6229 29952
rect 5909 29887 6229 29888
rect 15840 29952 16160 29953
rect 15840 29888 15848 29952
rect 15912 29888 15928 29952
rect 15992 29888 16008 29952
rect 16072 29888 16088 29952
rect 16152 29888 16160 29952
rect 15840 29887 16160 29888
rect 25770 29952 26090 29953
rect 25770 29888 25778 29952
rect 25842 29888 25858 29952
rect 25922 29888 25938 29952
rect 26002 29888 26018 29952
rect 26082 29888 26090 29952
rect 25770 29887 26090 29888
rect 2773 29882 2839 29885
rect 0 29880 2839 29882
rect 0 29824 2778 29880
rect 2834 29824 2839 29880
rect 0 29822 2839 29824
rect 0 29792 800 29822
rect 2773 29819 2839 29822
rect 10874 29408 11194 29409
rect 10874 29344 10882 29408
rect 10946 29344 10962 29408
rect 11026 29344 11042 29408
rect 11106 29344 11122 29408
rect 11186 29344 11194 29408
rect 10874 29343 11194 29344
rect 20805 29408 21125 29409
rect 20805 29344 20813 29408
rect 20877 29344 20893 29408
rect 20957 29344 20973 29408
rect 21037 29344 21053 29408
rect 21117 29344 21125 29408
rect 20805 29343 21125 29344
rect 0 29066 800 29096
rect 1485 29066 1551 29069
rect 0 29064 1551 29066
rect 0 29008 1490 29064
rect 1546 29008 1551 29064
rect 0 29006 1551 29008
rect 0 28976 800 29006
rect 1485 29003 1551 29006
rect 30005 28930 30071 28933
rect 31200 28930 32000 28960
rect 30005 28928 32000 28930
rect 30005 28872 30010 28928
rect 30066 28872 32000 28928
rect 30005 28870 32000 28872
rect 30005 28867 30071 28870
rect 5909 28864 6229 28865
rect 5909 28800 5917 28864
rect 5981 28800 5997 28864
rect 6061 28800 6077 28864
rect 6141 28800 6157 28864
rect 6221 28800 6229 28864
rect 5909 28799 6229 28800
rect 15840 28864 16160 28865
rect 15840 28800 15848 28864
rect 15912 28800 15928 28864
rect 15992 28800 16008 28864
rect 16072 28800 16088 28864
rect 16152 28800 16160 28864
rect 15840 28799 16160 28800
rect 25770 28864 26090 28865
rect 25770 28800 25778 28864
rect 25842 28800 25858 28864
rect 25922 28800 25938 28864
rect 26002 28800 26018 28864
rect 26082 28800 26090 28864
rect 31200 28840 32000 28870
rect 25770 28799 26090 28800
rect 0 28386 800 28416
rect 1485 28386 1551 28389
rect 0 28384 1551 28386
rect 0 28328 1490 28384
rect 1546 28328 1551 28384
rect 0 28326 1551 28328
rect 0 28296 800 28326
rect 1485 28323 1551 28326
rect 10874 28320 11194 28321
rect 10874 28256 10882 28320
rect 10946 28256 10962 28320
rect 11026 28256 11042 28320
rect 11106 28256 11122 28320
rect 11186 28256 11194 28320
rect 10874 28255 11194 28256
rect 20805 28320 21125 28321
rect 20805 28256 20813 28320
rect 20877 28256 20893 28320
rect 20957 28256 20973 28320
rect 21037 28256 21053 28320
rect 21117 28256 21125 28320
rect 20805 28255 21125 28256
rect 5909 27776 6229 27777
rect 5909 27712 5917 27776
rect 5981 27712 5997 27776
rect 6061 27712 6077 27776
rect 6141 27712 6157 27776
rect 6221 27712 6229 27776
rect 5909 27711 6229 27712
rect 15840 27776 16160 27777
rect 15840 27712 15848 27776
rect 15912 27712 15928 27776
rect 15992 27712 16008 27776
rect 16072 27712 16088 27776
rect 16152 27712 16160 27776
rect 15840 27711 16160 27712
rect 25770 27776 26090 27777
rect 25770 27712 25778 27776
rect 25842 27712 25858 27776
rect 25922 27712 25938 27776
rect 26002 27712 26018 27776
rect 26082 27712 26090 27776
rect 25770 27711 26090 27712
rect 7925 27706 7991 27709
rect 9489 27706 9555 27709
rect 7925 27704 9555 27706
rect 7925 27648 7930 27704
rect 7986 27648 9494 27704
rect 9550 27648 9555 27704
rect 7925 27646 9555 27648
rect 7925 27643 7991 27646
rect 9489 27643 9555 27646
rect 0 27570 800 27600
rect 1485 27570 1551 27573
rect 0 27568 1551 27570
rect 0 27512 1490 27568
rect 1546 27512 1551 27568
rect 0 27510 1551 27512
rect 0 27480 800 27510
rect 1485 27507 1551 27510
rect 8661 27570 8727 27573
rect 10685 27570 10751 27573
rect 8661 27568 10751 27570
rect 8661 27512 8666 27568
rect 8722 27512 10690 27568
rect 10746 27512 10751 27568
rect 8661 27510 10751 27512
rect 8661 27507 8727 27510
rect 10685 27507 10751 27510
rect 17534 27372 17540 27436
rect 17604 27434 17610 27436
rect 17677 27434 17743 27437
rect 19057 27434 19123 27437
rect 17604 27432 19123 27434
rect 17604 27376 17682 27432
rect 17738 27376 19062 27432
rect 19118 27376 19123 27432
rect 17604 27374 19123 27376
rect 17604 27372 17610 27374
rect 17677 27371 17743 27374
rect 19057 27371 19123 27374
rect 15561 27298 15627 27301
rect 19149 27298 19215 27301
rect 15561 27296 19215 27298
rect 15561 27240 15566 27296
rect 15622 27240 19154 27296
rect 19210 27240 19215 27296
rect 15561 27238 19215 27240
rect 15561 27235 15627 27238
rect 19149 27235 19215 27238
rect 10874 27232 11194 27233
rect 10874 27168 10882 27232
rect 10946 27168 10962 27232
rect 11026 27168 11042 27232
rect 11106 27168 11122 27232
rect 11186 27168 11194 27232
rect 10874 27167 11194 27168
rect 20805 27232 21125 27233
rect 20805 27168 20813 27232
rect 20877 27168 20893 27232
rect 20957 27168 20973 27232
rect 21037 27168 21053 27232
rect 21117 27168 21125 27232
rect 20805 27167 21125 27168
rect 30005 27026 30071 27029
rect 31200 27026 32000 27056
rect 30005 27024 32000 27026
rect 30005 26968 30010 27024
rect 30066 26968 32000 27024
rect 30005 26966 32000 26968
rect 30005 26963 30071 26966
rect 31200 26936 32000 26966
rect 0 26890 800 26920
rect 1485 26890 1551 26893
rect 0 26888 1551 26890
rect 0 26832 1490 26888
rect 1546 26832 1551 26888
rect 0 26830 1551 26832
rect 0 26800 800 26830
rect 1485 26827 1551 26830
rect 5909 26688 6229 26689
rect 5909 26624 5917 26688
rect 5981 26624 5997 26688
rect 6061 26624 6077 26688
rect 6141 26624 6157 26688
rect 6221 26624 6229 26688
rect 5909 26623 6229 26624
rect 15840 26688 16160 26689
rect 15840 26624 15848 26688
rect 15912 26624 15928 26688
rect 15992 26624 16008 26688
rect 16072 26624 16088 26688
rect 16152 26624 16160 26688
rect 15840 26623 16160 26624
rect 25770 26688 26090 26689
rect 25770 26624 25778 26688
rect 25842 26624 25858 26688
rect 25922 26624 25938 26688
rect 26002 26624 26018 26688
rect 26082 26624 26090 26688
rect 25770 26623 26090 26624
rect 8937 26482 9003 26485
rect 13445 26482 13511 26485
rect 8937 26480 13511 26482
rect 8937 26424 8942 26480
rect 8998 26424 13450 26480
rect 13506 26424 13511 26480
rect 8937 26422 13511 26424
rect 8937 26419 9003 26422
rect 13445 26419 13511 26422
rect 4245 26346 4311 26349
rect 4521 26346 4587 26349
rect 7966 26346 7972 26348
rect 4245 26344 7972 26346
rect 4245 26288 4250 26344
rect 4306 26288 4526 26344
rect 4582 26288 7972 26344
rect 4245 26286 7972 26288
rect 4245 26283 4311 26286
rect 4521 26283 4587 26286
rect 7966 26284 7972 26286
rect 8036 26346 8042 26348
rect 8661 26346 8727 26349
rect 8036 26344 8727 26346
rect 8036 26288 8666 26344
rect 8722 26288 8727 26344
rect 8036 26286 8727 26288
rect 8036 26284 8042 26286
rect 8661 26283 8727 26286
rect 0 26210 800 26240
rect 1485 26210 1551 26213
rect 0 26208 1551 26210
rect 0 26152 1490 26208
rect 1546 26152 1551 26208
rect 0 26150 1551 26152
rect 0 26120 800 26150
rect 1485 26147 1551 26150
rect 10874 26144 11194 26145
rect 10874 26080 10882 26144
rect 10946 26080 10962 26144
rect 11026 26080 11042 26144
rect 11106 26080 11122 26144
rect 11186 26080 11194 26144
rect 10874 26079 11194 26080
rect 20805 26144 21125 26145
rect 20805 26080 20813 26144
rect 20877 26080 20893 26144
rect 20957 26080 20973 26144
rect 21037 26080 21053 26144
rect 21117 26080 21125 26144
rect 20805 26079 21125 26080
rect 5909 25600 6229 25601
rect 5909 25536 5917 25600
rect 5981 25536 5997 25600
rect 6061 25536 6077 25600
rect 6141 25536 6157 25600
rect 6221 25536 6229 25600
rect 5909 25535 6229 25536
rect 15840 25600 16160 25601
rect 15840 25536 15848 25600
rect 15912 25536 15928 25600
rect 15992 25536 16008 25600
rect 16072 25536 16088 25600
rect 16152 25536 16160 25600
rect 15840 25535 16160 25536
rect 25770 25600 26090 25601
rect 25770 25536 25778 25600
rect 25842 25536 25858 25600
rect 25922 25536 25938 25600
rect 26002 25536 26018 25600
rect 26082 25536 26090 25600
rect 25770 25535 26090 25536
rect 0 25394 800 25424
rect 1485 25394 1551 25397
rect 0 25392 1551 25394
rect 0 25336 1490 25392
rect 1546 25336 1551 25392
rect 0 25334 1551 25336
rect 0 25304 800 25334
rect 1485 25331 1551 25334
rect 13353 25258 13419 25261
rect 18045 25258 18111 25261
rect 13353 25256 18111 25258
rect 13353 25200 13358 25256
rect 13414 25200 18050 25256
rect 18106 25200 18111 25256
rect 13353 25198 18111 25200
rect 13353 25195 13419 25198
rect 18045 25195 18111 25198
rect 10874 25056 11194 25057
rect 10874 24992 10882 25056
rect 10946 24992 10962 25056
rect 11026 24992 11042 25056
rect 11106 24992 11122 25056
rect 11186 24992 11194 25056
rect 10874 24991 11194 24992
rect 20805 25056 21125 25057
rect 20805 24992 20813 25056
rect 20877 24992 20893 25056
rect 20957 24992 20973 25056
rect 21037 24992 21053 25056
rect 21117 24992 21125 25056
rect 20805 24991 21125 24992
rect 30005 24986 30071 24989
rect 31200 24986 32000 25016
rect 30005 24984 32000 24986
rect 30005 24928 30010 24984
rect 30066 24928 32000 24984
rect 30005 24926 32000 24928
rect 30005 24923 30071 24926
rect 31200 24896 32000 24926
rect 0 24714 800 24744
rect 1485 24714 1551 24717
rect 0 24712 1551 24714
rect 0 24656 1490 24712
rect 1546 24656 1551 24712
rect 0 24654 1551 24656
rect 0 24624 800 24654
rect 1485 24651 1551 24654
rect 5909 24512 6229 24513
rect 5909 24448 5917 24512
rect 5981 24448 5997 24512
rect 6061 24448 6077 24512
rect 6141 24448 6157 24512
rect 6221 24448 6229 24512
rect 5909 24447 6229 24448
rect 15840 24512 16160 24513
rect 15840 24448 15848 24512
rect 15912 24448 15928 24512
rect 15992 24448 16008 24512
rect 16072 24448 16088 24512
rect 16152 24448 16160 24512
rect 15840 24447 16160 24448
rect 25770 24512 26090 24513
rect 25770 24448 25778 24512
rect 25842 24448 25858 24512
rect 25922 24448 25938 24512
rect 26002 24448 26018 24512
rect 26082 24448 26090 24512
rect 25770 24447 26090 24448
rect 4153 24170 4219 24173
rect 4521 24170 4587 24173
rect 5533 24170 5599 24173
rect 4153 24168 5599 24170
rect 4153 24112 4158 24168
rect 4214 24112 4526 24168
rect 4582 24112 5538 24168
rect 5594 24112 5599 24168
rect 4153 24110 5599 24112
rect 4153 24107 4219 24110
rect 4521 24107 4587 24110
rect 5533 24107 5599 24110
rect 10874 23968 11194 23969
rect 0 23898 800 23928
rect 10874 23904 10882 23968
rect 10946 23904 10962 23968
rect 11026 23904 11042 23968
rect 11106 23904 11122 23968
rect 11186 23904 11194 23968
rect 10874 23903 11194 23904
rect 20805 23968 21125 23969
rect 20805 23904 20813 23968
rect 20877 23904 20893 23968
rect 20957 23904 20973 23968
rect 21037 23904 21053 23968
rect 21117 23904 21125 23968
rect 20805 23903 21125 23904
rect 1485 23898 1551 23901
rect 0 23896 1551 23898
rect 0 23840 1490 23896
rect 1546 23840 1551 23896
rect 0 23838 1551 23840
rect 0 23808 800 23838
rect 1485 23835 1551 23838
rect 5909 23424 6229 23425
rect 5909 23360 5917 23424
rect 5981 23360 5997 23424
rect 6061 23360 6077 23424
rect 6141 23360 6157 23424
rect 6221 23360 6229 23424
rect 5909 23359 6229 23360
rect 15840 23424 16160 23425
rect 15840 23360 15848 23424
rect 15912 23360 15928 23424
rect 15992 23360 16008 23424
rect 16072 23360 16088 23424
rect 16152 23360 16160 23424
rect 15840 23359 16160 23360
rect 25770 23424 26090 23425
rect 25770 23360 25778 23424
rect 25842 23360 25858 23424
rect 25922 23360 25938 23424
rect 26002 23360 26018 23424
rect 26082 23360 26090 23424
rect 25770 23359 26090 23360
rect 0 23218 800 23248
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 800 23158
rect 1393 23155 1459 23158
rect 16665 23218 16731 23221
rect 17534 23218 17540 23220
rect 16665 23216 17540 23218
rect 16665 23160 16670 23216
rect 16726 23160 17540 23216
rect 16665 23158 17540 23160
rect 16665 23155 16731 23158
rect 17534 23156 17540 23158
rect 17604 23156 17610 23220
rect 30005 22946 30071 22949
rect 31200 22946 32000 22976
rect 30005 22944 32000 22946
rect 30005 22888 30010 22944
rect 30066 22888 32000 22944
rect 30005 22886 32000 22888
rect 30005 22883 30071 22886
rect 10874 22880 11194 22881
rect 10874 22816 10882 22880
rect 10946 22816 10962 22880
rect 11026 22816 11042 22880
rect 11106 22816 11122 22880
rect 11186 22816 11194 22880
rect 10874 22815 11194 22816
rect 20805 22880 21125 22881
rect 20805 22816 20813 22880
rect 20877 22816 20893 22880
rect 20957 22816 20973 22880
rect 21037 22816 21053 22880
rect 21117 22816 21125 22880
rect 31200 22856 32000 22886
rect 20805 22815 21125 22816
rect 9397 22676 9463 22677
rect 9397 22674 9444 22676
rect 9352 22672 9444 22674
rect 9352 22616 9402 22672
rect 9352 22614 9444 22616
rect 9397 22612 9444 22614
rect 9508 22612 9514 22676
rect 9397 22611 9463 22612
rect 0 22402 800 22432
rect 2037 22402 2103 22405
rect 0 22400 2103 22402
rect 0 22344 2042 22400
rect 2098 22344 2103 22400
rect 0 22342 2103 22344
rect 0 22312 800 22342
rect 2037 22339 2103 22342
rect 16941 22402 17007 22405
rect 16941 22400 17050 22402
rect 16941 22344 16946 22400
rect 17002 22344 17050 22400
rect 16941 22339 17050 22344
rect 5909 22336 6229 22337
rect 5909 22272 5917 22336
rect 5981 22272 5997 22336
rect 6061 22272 6077 22336
rect 6141 22272 6157 22336
rect 6221 22272 6229 22336
rect 5909 22271 6229 22272
rect 15840 22336 16160 22337
rect 15840 22272 15848 22336
rect 15912 22272 15928 22336
rect 15992 22272 16008 22336
rect 16072 22272 16088 22336
rect 16152 22272 16160 22336
rect 15840 22271 16160 22272
rect 8109 22266 8175 22269
rect 7974 22264 8175 22266
rect 7974 22208 8114 22264
rect 8170 22208 8175 22264
rect 7974 22206 8175 22208
rect 7974 21997 8034 22206
rect 8109 22203 8175 22206
rect 8569 22130 8635 22133
rect 9029 22130 9095 22133
rect 8569 22128 9095 22130
rect 8569 22072 8574 22128
rect 8630 22072 9034 22128
rect 9090 22072 9095 22128
rect 8569 22070 9095 22072
rect 8569 22067 8635 22070
rect 9029 22067 9095 22070
rect 7925 21992 8034 21997
rect 7925 21936 7930 21992
rect 7986 21936 8034 21992
rect 7925 21934 8034 21936
rect 16990 21994 17050 22339
rect 25770 22336 26090 22337
rect 25770 22272 25778 22336
rect 25842 22272 25858 22336
rect 25922 22272 25938 22336
rect 26002 22272 26018 22336
rect 26082 22272 26090 22336
rect 25770 22271 26090 22272
rect 17585 21994 17651 21997
rect 16990 21992 17651 21994
rect 16990 21936 17590 21992
rect 17646 21936 17651 21992
rect 16990 21934 17651 21936
rect 7925 21931 7991 21934
rect 17585 21931 17651 21934
rect 7833 21858 7899 21861
rect 9397 21858 9463 21861
rect 7833 21856 9463 21858
rect 7833 21800 7838 21856
rect 7894 21800 9402 21856
rect 9458 21800 9463 21856
rect 7833 21798 9463 21800
rect 7833 21795 7899 21798
rect 9397 21795 9463 21798
rect 10874 21792 11194 21793
rect 0 21722 800 21752
rect 10874 21728 10882 21792
rect 10946 21728 10962 21792
rect 11026 21728 11042 21792
rect 11106 21728 11122 21792
rect 11186 21728 11194 21792
rect 10874 21727 11194 21728
rect 20805 21792 21125 21793
rect 20805 21728 20813 21792
rect 20877 21728 20893 21792
rect 20957 21728 20973 21792
rect 21037 21728 21053 21792
rect 21117 21728 21125 21792
rect 20805 21727 21125 21728
rect 2957 21722 3023 21725
rect 0 21720 3023 21722
rect 0 21664 2962 21720
rect 3018 21664 3023 21720
rect 0 21662 3023 21664
rect 0 21632 800 21662
rect 2957 21659 3023 21662
rect 7833 21722 7899 21725
rect 7966 21722 7972 21724
rect 7833 21720 7972 21722
rect 7833 21664 7838 21720
rect 7894 21664 7972 21720
rect 7833 21662 7972 21664
rect 7833 21659 7899 21662
rect 7966 21660 7972 21662
rect 8036 21660 8042 21724
rect 8201 21722 8267 21725
rect 9581 21722 9647 21725
rect 8201 21720 9506 21722
rect 8201 21664 8206 21720
rect 8262 21664 9506 21720
rect 8201 21662 9506 21664
rect 8201 21659 8267 21662
rect 9446 21589 9506 21662
rect 9581 21720 9690 21722
rect 9581 21664 9586 21720
rect 9642 21664 9690 21720
rect 9581 21659 9690 21664
rect 9446 21584 9555 21589
rect 9446 21528 9494 21584
rect 9550 21528 9555 21584
rect 9446 21526 9555 21528
rect 9489 21523 9555 21526
rect 9630 21453 9690 21659
rect 9581 21448 9690 21453
rect 9581 21392 9586 21448
rect 9642 21392 9690 21448
rect 9581 21390 9690 21392
rect 9581 21387 9647 21390
rect 5909 21248 6229 21249
rect 5909 21184 5917 21248
rect 5981 21184 5997 21248
rect 6061 21184 6077 21248
rect 6141 21184 6157 21248
rect 6221 21184 6229 21248
rect 5909 21183 6229 21184
rect 15840 21248 16160 21249
rect 15840 21184 15848 21248
rect 15912 21184 15928 21248
rect 15992 21184 16008 21248
rect 16072 21184 16088 21248
rect 16152 21184 16160 21248
rect 15840 21183 16160 21184
rect 25770 21248 26090 21249
rect 25770 21184 25778 21248
rect 25842 21184 25858 21248
rect 25922 21184 25938 21248
rect 26002 21184 26018 21248
rect 26082 21184 26090 21248
rect 25770 21183 26090 21184
rect 9397 21180 9463 21181
rect 9397 21176 9444 21180
rect 9508 21178 9514 21180
rect 9397 21120 9402 21176
rect 9397 21116 9444 21120
rect 9508 21118 9554 21178
rect 9508 21116 9514 21118
rect 9397 21115 9463 21116
rect 0 21042 800 21072
rect 1853 21042 1919 21045
rect 0 21040 1919 21042
rect 0 20984 1858 21040
rect 1914 20984 1919 21040
rect 0 20982 1919 20984
rect 0 20952 800 20982
rect 1853 20979 1919 20982
rect 30005 21042 30071 21045
rect 31200 21042 32000 21072
rect 30005 21040 32000 21042
rect 30005 20984 30010 21040
rect 30066 20984 32000 21040
rect 30005 20982 32000 20984
rect 30005 20979 30071 20982
rect 31200 20952 32000 20982
rect 10874 20704 11194 20705
rect 10874 20640 10882 20704
rect 10946 20640 10962 20704
rect 11026 20640 11042 20704
rect 11106 20640 11122 20704
rect 11186 20640 11194 20704
rect 10874 20639 11194 20640
rect 20805 20704 21125 20705
rect 20805 20640 20813 20704
rect 20877 20640 20893 20704
rect 20957 20640 20973 20704
rect 21037 20640 21053 20704
rect 21117 20640 21125 20704
rect 20805 20639 21125 20640
rect 0 20226 800 20256
rect 2773 20226 2839 20229
rect 0 20224 2839 20226
rect 0 20168 2778 20224
rect 2834 20168 2839 20224
rect 0 20166 2839 20168
rect 0 20136 800 20166
rect 2773 20163 2839 20166
rect 5909 20160 6229 20161
rect 5909 20096 5917 20160
rect 5981 20096 5997 20160
rect 6061 20096 6077 20160
rect 6141 20096 6157 20160
rect 6221 20096 6229 20160
rect 5909 20095 6229 20096
rect 15840 20160 16160 20161
rect 15840 20096 15848 20160
rect 15912 20096 15928 20160
rect 15992 20096 16008 20160
rect 16072 20096 16088 20160
rect 16152 20096 16160 20160
rect 15840 20095 16160 20096
rect 25770 20160 26090 20161
rect 25770 20096 25778 20160
rect 25842 20096 25858 20160
rect 25922 20096 25938 20160
rect 26002 20096 26018 20160
rect 26082 20096 26090 20160
rect 25770 20095 26090 20096
rect 15469 19954 15535 19957
rect 15837 19954 15903 19957
rect 15469 19952 15903 19954
rect 15469 19896 15474 19952
rect 15530 19896 15842 19952
rect 15898 19896 15903 19952
rect 15469 19894 15903 19896
rect 15469 19891 15535 19894
rect 15837 19891 15903 19894
rect 10874 19616 11194 19617
rect 0 19546 800 19576
rect 10874 19552 10882 19616
rect 10946 19552 10962 19616
rect 11026 19552 11042 19616
rect 11106 19552 11122 19616
rect 11186 19552 11194 19616
rect 10874 19551 11194 19552
rect 20805 19616 21125 19617
rect 20805 19552 20813 19616
rect 20877 19552 20893 19616
rect 20957 19552 20973 19616
rect 21037 19552 21053 19616
rect 21117 19552 21125 19616
rect 20805 19551 21125 19552
rect 3141 19546 3207 19549
rect 0 19544 3207 19546
rect 0 19488 3146 19544
rect 3202 19488 3207 19544
rect 0 19486 3207 19488
rect 0 19456 800 19486
rect 3141 19483 3207 19486
rect 11053 19138 11119 19141
rect 11278 19138 11284 19140
rect 11053 19136 11284 19138
rect 11053 19080 11058 19136
rect 11114 19080 11284 19136
rect 11053 19078 11284 19080
rect 11053 19075 11119 19078
rect 11278 19076 11284 19078
rect 11348 19076 11354 19140
rect 5909 19072 6229 19073
rect 5909 19008 5917 19072
rect 5981 19008 5997 19072
rect 6061 19008 6077 19072
rect 6141 19008 6157 19072
rect 6221 19008 6229 19072
rect 5909 19007 6229 19008
rect 15840 19072 16160 19073
rect 15840 19008 15848 19072
rect 15912 19008 15928 19072
rect 15992 19008 16008 19072
rect 16072 19008 16088 19072
rect 16152 19008 16160 19072
rect 15840 19007 16160 19008
rect 25770 19072 26090 19073
rect 25770 19008 25778 19072
rect 25842 19008 25858 19072
rect 25922 19008 25938 19072
rect 26002 19008 26018 19072
rect 26082 19008 26090 19072
rect 25770 19007 26090 19008
rect 30005 19002 30071 19005
rect 31200 19002 32000 19032
rect 30005 19000 32000 19002
rect 30005 18944 30010 19000
rect 30066 18944 32000 19000
rect 30005 18942 32000 18944
rect 30005 18939 30071 18942
rect 31200 18912 32000 18942
rect 0 18730 800 18760
rect 2957 18730 3023 18733
rect 0 18728 3023 18730
rect 0 18672 2962 18728
rect 3018 18672 3023 18728
rect 0 18670 3023 18672
rect 0 18640 800 18670
rect 2957 18667 3023 18670
rect 10874 18528 11194 18529
rect 10874 18464 10882 18528
rect 10946 18464 10962 18528
rect 11026 18464 11042 18528
rect 11106 18464 11122 18528
rect 11186 18464 11194 18528
rect 10874 18463 11194 18464
rect 20805 18528 21125 18529
rect 20805 18464 20813 18528
rect 20877 18464 20893 18528
rect 20957 18464 20973 18528
rect 21037 18464 21053 18528
rect 21117 18464 21125 18528
rect 20805 18463 21125 18464
rect 0 18050 800 18080
rect 3877 18050 3943 18053
rect 0 18048 3943 18050
rect 0 17992 3882 18048
rect 3938 17992 3943 18048
rect 0 17990 3943 17992
rect 0 17960 800 17990
rect 3877 17987 3943 17990
rect 5909 17984 6229 17985
rect 5909 17920 5917 17984
rect 5981 17920 5997 17984
rect 6061 17920 6077 17984
rect 6141 17920 6157 17984
rect 6221 17920 6229 17984
rect 5909 17919 6229 17920
rect 15840 17984 16160 17985
rect 15840 17920 15848 17984
rect 15912 17920 15928 17984
rect 15992 17920 16008 17984
rect 16072 17920 16088 17984
rect 16152 17920 16160 17984
rect 15840 17919 16160 17920
rect 25770 17984 26090 17985
rect 25770 17920 25778 17984
rect 25842 17920 25858 17984
rect 25922 17920 25938 17984
rect 26002 17920 26018 17984
rect 26082 17920 26090 17984
rect 25770 17919 26090 17920
rect 10874 17440 11194 17441
rect 10874 17376 10882 17440
rect 10946 17376 10962 17440
rect 11026 17376 11042 17440
rect 11106 17376 11122 17440
rect 11186 17376 11194 17440
rect 10874 17375 11194 17376
rect 20805 17440 21125 17441
rect 20805 17376 20813 17440
rect 20877 17376 20893 17440
rect 20957 17376 20973 17440
rect 21037 17376 21053 17440
rect 21117 17376 21125 17440
rect 20805 17375 21125 17376
rect 10133 17372 10199 17373
rect 10133 17370 10180 17372
rect 10088 17368 10180 17370
rect 10088 17312 10138 17368
rect 10088 17310 10180 17312
rect 10133 17308 10180 17310
rect 10244 17308 10250 17372
rect 10133 17307 10199 17308
rect 0 17234 800 17264
rect 3969 17234 4035 17237
rect 0 17232 4035 17234
rect 0 17176 3974 17232
rect 4030 17176 4035 17232
rect 0 17174 4035 17176
rect 0 17144 800 17174
rect 3969 17171 4035 17174
rect 19333 17234 19399 17237
rect 20621 17234 20687 17237
rect 19333 17232 20687 17234
rect 19333 17176 19338 17232
rect 19394 17176 20626 17232
rect 20682 17176 20687 17232
rect 19333 17174 20687 17176
rect 19333 17171 19399 17174
rect 20621 17171 20687 17174
rect 30005 16962 30071 16965
rect 31200 16962 32000 16992
rect 30005 16960 32000 16962
rect 30005 16904 30010 16960
rect 30066 16904 32000 16960
rect 30005 16902 32000 16904
rect 30005 16899 30071 16902
rect 5909 16896 6229 16897
rect 5909 16832 5917 16896
rect 5981 16832 5997 16896
rect 6061 16832 6077 16896
rect 6141 16832 6157 16896
rect 6221 16832 6229 16896
rect 5909 16831 6229 16832
rect 15840 16896 16160 16897
rect 15840 16832 15848 16896
rect 15912 16832 15928 16896
rect 15992 16832 16008 16896
rect 16072 16832 16088 16896
rect 16152 16832 16160 16896
rect 15840 16831 16160 16832
rect 25770 16896 26090 16897
rect 25770 16832 25778 16896
rect 25842 16832 25858 16896
rect 25922 16832 25938 16896
rect 26002 16832 26018 16896
rect 26082 16832 26090 16896
rect 31200 16872 32000 16902
rect 25770 16831 26090 16832
rect 0 16554 800 16584
rect 2773 16554 2839 16557
rect 0 16552 2839 16554
rect 0 16496 2778 16552
rect 2834 16496 2839 16552
rect 0 16494 2839 16496
rect 0 16464 800 16494
rect 2773 16491 2839 16494
rect 10874 16352 11194 16353
rect 10874 16288 10882 16352
rect 10946 16288 10962 16352
rect 11026 16288 11042 16352
rect 11106 16288 11122 16352
rect 11186 16288 11194 16352
rect 10874 16287 11194 16288
rect 20805 16352 21125 16353
rect 20805 16288 20813 16352
rect 20877 16288 20893 16352
rect 20957 16288 20973 16352
rect 21037 16288 21053 16352
rect 21117 16288 21125 16352
rect 20805 16287 21125 16288
rect 3233 16282 3299 16285
rect 7189 16282 7255 16285
rect 3233 16280 7255 16282
rect 3233 16224 3238 16280
rect 3294 16224 7194 16280
rect 7250 16224 7255 16280
rect 3233 16222 7255 16224
rect 3233 16219 3299 16222
rect 7189 16219 7255 16222
rect 0 15874 800 15904
rect 1393 15874 1459 15877
rect 0 15872 1459 15874
rect 0 15816 1398 15872
rect 1454 15816 1459 15872
rect 0 15814 1459 15816
rect 0 15784 800 15814
rect 1393 15811 1459 15814
rect 5909 15808 6229 15809
rect 5909 15744 5917 15808
rect 5981 15744 5997 15808
rect 6061 15744 6077 15808
rect 6141 15744 6157 15808
rect 6221 15744 6229 15808
rect 5909 15743 6229 15744
rect 15840 15808 16160 15809
rect 15840 15744 15848 15808
rect 15912 15744 15928 15808
rect 15992 15744 16008 15808
rect 16072 15744 16088 15808
rect 16152 15744 16160 15808
rect 15840 15743 16160 15744
rect 25770 15808 26090 15809
rect 25770 15744 25778 15808
rect 25842 15744 25858 15808
rect 25922 15744 25938 15808
rect 26002 15744 26018 15808
rect 26082 15744 26090 15808
rect 25770 15743 26090 15744
rect 5073 15602 5139 15605
rect 6177 15602 6243 15605
rect 5073 15600 6243 15602
rect 5073 15544 5078 15600
rect 5134 15544 6182 15600
rect 6238 15544 6243 15600
rect 5073 15542 6243 15544
rect 5073 15539 5139 15542
rect 6177 15539 6243 15542
rect 9121 15468 9187 15469
rect 9070 15404 9076 15468
rect 9140 15466 9187 15468
rect 16389 15466 16455 15469
rect 17401 15466 17467 15469
rect 9140 15464 9232 15466
rect 9182 15408 9232 15464
rect 9140 15406 9232 15408
rect 16389 15464 17467 15466
rect 16389 15408 16394 15464
rect 16450 15408 17406 15464
rect 17462 15408 17467 15464
rect 16389 15406 17467 15408
rect 9140 15404 9187 15406
rect 9121 15403 9187 15404
rect 16389 15403 16455 15406
rect 17401 15403 17467 15406
rect 17125 15330 17191 15333
rect 17401 15330 17467 15333
rect 18321 15330 18387 15333
rect 17125 15328 18387 15330
rect 17125 15272 17130 15328
rect 17186 15272 17406 15328
rect 17462 15272 18326 15328
rect 18382 15272 18387 15328
rect 17125 15270 18387 15272
rect 17125 15267 17191 15270
rect 17401 15267 17467 15270
rect 18321 15267 18387 15270
rect 10874 15264 11194 15265
rect 10874 15200 10882 15264
rect 10946 15200 10962 15264
rect 11026 15200 11042 15264
rect 11106 15200 11122 15264
rect 11186 15200 11194 15264
rect 10874 15199 11194 15200
rect 20805 15264 21125 15265
rect 20805 15200 20813 15264
rect 20877 15200 20893 15264
rect 20957 15200 20973 15264
rect 21037 15200 21053 15264
rect 21117 15200 21125 15264
rect 20805 15199 21125 15200
rect 12065 15194 12131 15197
rect 17217 15194 17283 15197
rect 12065 15192 17283 15194
rect 12065 15136 12070 15192
rect 12126 15136 17222 15192
rect 17278 15136 17283 15192
rect 12065 15134 17283 15136
rect 12065 15131 12131 15134
rect 17217 15131 17283 15134
rect 0 15058 800 15088
rect 3141 15058 3207 15061
rect 0 15056 3207 15058
rect 0 15000 3146 15056
rect 3202 15000 3207 15056
rect 0 14998 3207 15000
rect 0 14968 800 14998
rect 3141 14995 3207 14998
rect 17033 15058 17099 15061
rect 17861 15058 17927 15061
rect 17033 15056 17927 15058
rect 17033 15000 17038 15056
rect 17094 15000 17866 15056
rect 17922 15000 17927 15056
rect 17033 14998 17927 15000
rect 17033 14995 17099 14998
rect 17861 14995 17927 14998
rect 30005 14922 30071 14925
rect 31200 14922 32000 14952
rect 30005 14920 32000 14922
rect 30005 14864 30010 14920
rect 30066 14864 32000 14920
rect 30005 14862 32000 14864
rect 30005 14859 30071 14862
rect 31200 14832 32000 14862
rect 5909 14720 6229 14721
rect 5909 14656 5917 14720
rect 5981 14656 5997 14720
rect 6061 14656 6077 14720
rect 6141 14656 6157 14720
rect 6221 14656 6229 14720
rect 5909 14655 6229 14656
rect 15840 14720 16160 14721
rect 15840 14656 15848 14720
rect 15912 14656 15928 14720
rect 15992 14656 16008 14720
rect 16072 14656 16088 14720
rect 16152 14656 16160 14720
rect 15840 14655 16160 14656
rect 25770 14720 26090 14721
rect 25770 14656 25778 14720
rect 25842 14656 25858 14720
rect 25922 14656 25938 14720
rect 26002 14656 26018 14720
rect 26082 14656 26090 14720
rect 25770 14655 26090 14656
rect 6913 14514 6979 14517
rect 9581 14514 9647 14517
rect 6913 14512 9647 14514
rect 6913 14456 6918 14512
rect 6974 14456 9586 14512
rect 9642 14456 9647 14512
rect 6913 14454 9647 14456
rect 6913 14451 6979 14454
rect 9581 14451 9647 14454
rect 0 14378 800 14408
rect 1209 14378 1275 14381
rect 0 14376 1275 14378
rect 0 14320 1214 14376
rect 1270 14320 1275 14376
rect 0 14318 1275 14320
rect 0 14288 800 14318
rect 1209 14315 1275 14318
rect 5901 14378 5967 14381
rect 7097 14378 7163 14381
rect 5901 14376 7163 14378
rect 5901 14320 5906 14376
rect 5962 14320 7102 14376
rect 7158 14320 7163 14376
rect 5901 14318 7163 14320
rect 5901 14315 5967 14318
rect 7097 14315 7163 14318
rect 10874 14176 11194 14177
rect 10874 14112 10882 14176
rect 10946 14112 10962 14176
rect 11026 14112 11042 14176
rect 11106 14112 11122 14176
rect 11186 14112 11194 14176
rect 10874 14111 11194 14112
rect 20805 14176 21125 14177
rect 20805 14112 20813 14176
rect 20877 14112 20893 14176
rect 20957 14112 20973 14176
rect 21037 14112 21053 14176
rect 21117 14112 21125 14176
rect 20805 14111 21125 14112
rect 4981 13970 5047 13973
rect 6821 13970 6887 13973
rect 4981 13968 6887 13970
rect 4981 13912 4986 13968
rect 5042 13912 6826 13968
rect 6882 13912 6887 13968
rect 4981 13910 6887 13912
rect 4981 13907 5047 13910
rect 6821 13907 6887 13910
rect 11421 13970 11487 13973
rect 18597 13970 18663 13973
rect 11421 13968 18663 13970
rect 11421 13912 11426 13968
rect 11482 13912 18602 13968
rect 18658 13912 18663 13968
rect 11421 13910 18663 13912
rect 11421 13907 11487 13910
rect 18597 13907 18663 13910
rect 5909 13632 6229 13633
rect 0 13562 800 13592
rect 5909 13568 5917 13632
rect 5981 13568 5997 13632
rect 6061 13568 6077 13632
rect 6141 13568 6157 13632
rect 6221 13568 6229 13632
rect 5909 13567 6229 13568
rect 15840 13632 16160 13633
rect 15840 13568 15848 13632
rect 15912 13568 15928 13632
rect 15992 13568 16008 13632
rect 16072 13568 16088 13632
rect 16152 13568 16160 13632
rect 15840 13567 16160 13568
rect 25770 13632 26090 13633
rect 25770 13568 25778 13632
rect 25842 13568 25858 13632
rect 25922 13568 25938 13632
rect 26002 13568 26018 13632
rect 26082 13568 26090 13632
rect 25770 13567 26090 13568
rect 1393 13562 1459 13565
rect 0 13560 1459 13562
rect 0 13504 1398 13560
rect 1454 13504 1459 13560
rect 0 13502 1459 13504
rect 0 13472 800 13502
rect 1393 13499 1459 13502
rect 10874 13088 11194 13089
rect 10874 13024 10882 13088
rect 10946 13024 10962 13088
rect 11026 13024 11042 13088
rect 11106 13024 11122 13088
rect 11186 13024 11194 13088
rect 10874 13023 11194 13024
rect 20805 13088 21125 13089
rect 20805 13024 20813 13088
rect 20877 13024 20893 13088
rect 20957 13024 20973 13088
rect 21037 13024 21053 13088
rect 21117 13024 21125 13088
rect 20805 13023 21125 13024
rect 30005 13018 30071 13021
rect 31200 13018 32000 13048
rect 30005 13016 32000 13018
rect 30005 12960 30010 13016
rect 30066 12960 32000 13016
rect 30005 12958 32000 12960
rect 30005 12955 30071 12958
rect 31200 12928 32000 12958
rect 0 12882 800 12912
rect 1393 12882 1459 12885
rect 0 12880 1459 12882
rect 0 12824 1398 12880
rect 1454 12824 1459 12880
rect 0 12822 1459 12824
rect 0 12792 800 12822
rect 1393 12819 1459 12822
rect 9213 12882 9279 12885
rect 9213 12880 9322 12882
rect 9213 12824 9218 12880
rect 9274 12824 9322 12880
rect 9213 12819 9322 12824
rect 9262 12746 9322 12819
rect 9581 12746 9647 12749
rect 9262 12744 9647 12746
rect 9262 12688 9586 12744
rect 9642 12688 9647 12744
rect 9262 12686 9647 12688
rect 9581 12683 9647 12686
rect 5909 12544 6229 12545
rect 5909 12480 5917 12544
rect 5981 12480 5997 12544
rect 6061 12480 6077 12544
rect 6141 12480 6157 12544
rect 6221 12480 6229 12544
rect 5909 12479 6229 12480
rect 15840 12544 16160 12545
rect 15840 12480 15848 12544
rect 15912 12480 15928 12544
rect 15992 12480 16008 12544
rect 16072 12480 16088 12544
rect 16152 12480 16160 12544
rect 15840 12479 16160 12480
rect 25770 12544 26090 12545
rect 25770 12480 25778 12544
rect 25842 12480 25858 12544
rect 25922 12480 25938 12544
rect 26002 12480 26018 12544
rect 26082 12480 26090 12544
rect 25770 12479 26090 12480
rect 9581 12448 9647 12453
rect 9581 12392 9586 12448
rect 9642 12392 9647 12448
rect 9581 12387 9647 12392
rect 0 12066 800 12096
rect 1393 12066 1459 12069
rect 0 12064 1459 12066
rect 0 12008 1398 12064
rect 1454 12008 1459 12064
rect 0 12006 1459 12008
rect 0 11976 800 12006
rect 1393 12003 1459 12006
rect 9121 11794 9187 11797
rect 9078 11792 9187 11794
rect 9078 11736 9126 11792
rect 9182 11736 9187 11792
rect 9078 11731 9187 11736
rect 5909 11456 6229 11457
rect 0 11386 800 11416
rect 5909 11392 5917 11456
rect 5981 11392 5997 11456
rect 6061 11392 6077 11456
rect 6141 11392 6157 11456
rect 6221 11392 6229 11456
rect 5909 11391 6229 11392
rect 9078 11389 9138 11731
rect 9213 11658 9279 11661
rect 9584 11658 9644 12387
rect 10501 12338 10567 12341
rect 11237 12338 11303 12341
rect 10501 12336 11303 12338
rect 10501 12280 10506 12336
rect 10562 12280 11242 12336
rect 11298 12280 11303 12336
rect 10501 12278 11303 12280
rect 10501 12275 10567 12278
rect 11237 12275 11303 12278
rect 10174 12004 10180 12068
rect 10244 12066 10250 12068
rect 10317 12066 10383 12069
rect 10244 12064 10383 12066
rect 10244 12008 10322 12064
rect 10378 12008 10383 12064
rect 10244 12006 10383 12008
rect 10244 12004 10250 12006
rect 10317 12003 10383 12006
rect 10874 12000 11194 12001
rect 10874 11936 10882 12000
rect 10946 11936 10962 12000
rect 11026 11936 11042 12000
rect 11106 11936 11122 12000
rect 11186 11936 11194 12000
rect 10874 11935 11194 11936
rect 20805 12000 21125 12001
rect 20805 11936 20813 12000
rect 20877 11936 20893 12000
rect 20957 11936 20973 12000
rect 21037 11936 21053 12000
rect 21117 11936 21125 12000
rect 20805 11935 21125 11936
rect 9213 11656 9644 11658
rect 9213 11600 9218 11656
rect 9274 11600 9644 11656
rect 9213 11598 9644 11600
rect 9213 11595 9279 11598
rect 9857 11522 9923 11525
rect 10593 11522 10659 11525
rect 9857 11520 10659 11522
rect 9857 11464 9862 11520
rect 9918 11464 10598 11520
rect 10654 11464 10659 11520
rect 9857 11462 10659 11464
rect 9857 11459 9923 11462
rect 10593 11459 10659 11462
rect 15840 11456 16160 11457
rect 15840 11392 15848 11456
rect 15912 11392 15928 11456
rect 15992 11392 16008 11456
rect 16072 11392 16088 11456
rect 16152 11392 16160 11456
rect 15840 11391 16160 11392
rect 25770 11456 26090 11457
rect 25770 11392 25778 11456
rect 25842 11392 25858 11456
rect 25922 11392 25938 11456
rect 26002 11392 26018 11456
rect 26082 11392 26090 11456
rect 25770 11391 26090 11392
rect 1209 11386 1275 11389
rect 0 11384 1275 11386
rect 0 11328 1214 11384
rect 1270 11328 1275 11384
rect 0 11326 1275 11328
rect 9078 11384 9187 11389
rect 9078 11328 9126 11384
rect 9182 11328 9187 11384
rect 9078 11326 9187 11328
rect 0 11296 800 11326
rect 1209 11323 1275 11326
rect 9121 11323 9187 11326
rect 9029 11252 9095 11253
rect 9029 11248 9076 11252
rect 9140 11250 9146 11252
rect 9029 11192 9034 11248
rect 9029 11188 9076 11192
rect 9140 11190 9186 11250
rect 9140 11188 9146 11190
rect 9029 11187 9095 11188
rect 30005 10978 30071 10981
rect 31200 10978 32000 11008
rect 30005 10976 32000 10978
rect 30005 10920 30010 10976
rect 30066 10920 32000 10976
rect 30005 10918 32000 10920
rect 30005 10915 30071 10918
rect 10874 10912 11194 10913
rect 10874 10848 10882 10912
rect 10946 10848 10962 10912
rect 11026 10848 11042 10912
rect 11106 10848 11122 10912
rect 11186 10848 11194 10912
rect 10874 10847 11194 10848
rect 20805 10912 21125 10913
rect 20805 10848 20813 10912
rect 20877 10848 20893 10912
rect 20957 10848 20973 10912
rect 21037 10848 21053 10912
rect 21117 10848 21125 10912
rect 31200 10888 32000 10918
rect 20805 10847 21125 10848
rect 0 10706 800 10736
rect 1393 10706 1459 10709
rect 0 10704 1459 10706
rect 0 10648 1398 10704
rect 1454 10648 1459 10704
rect 0 10646 1459 10648
rect 0 10616 800 10646
rect 1393 10643 1459 10646
rect 5909 10368 6229 10369
rect 5909 10304 5917 10368
rect 5981 10304 5997 10368
rect 6061 10304 6077 10368
rect 6141 10304 6157 10368
rect 6221 10304 6229 10368
rect 5909 10303 6229 10304
rect 15840 10368 16160 10369
rect 15840 10304 15848 10368
rect 15912 10304 15928 10368
rect 15992 10304 16008 10368
rect 16072 10304 16088 10368
rect 16152 10304 16160 10368
rect 15840 10303 16160 10304
rect 25770 10368 26090 10369
rect 25770 10304 25778 10368
rect 25842 10304 25858 10368
rect 25922 10304 25938 10368
rect 26002 10304 26018 10368
rect 26082 10304 26090 10368
rect 25770 10303 26090 10304
rect 0 9890 800 9920
rect 3049 9890 3115 9893
rect 0 9888 3115 9890
rect 0 9832 3054 9888
rect 3110 9832 3115 9888
rect 0 9830 3115 9832
rect 0 9800 800 9830
rect 3049 9827 3115 9830
rect 10874 9824 11194 9825
rect 10874 9760 10882 9824
rect 10946 9760 10962 9824
rect 11026 9760 11042 9824
rect 11106 9760 11122 9824
rect 11186 9760 11194 9824
rect 10874 9759 11194 9760
rect 20805 9824 21125 9825
rect 20805 9760 20813 9824
rect 20877 9760 20893 9824
rect 20957 9760 20973 9824
rect 21037 9760 21053 9824
rect 21117 9760 21125 9824
rect 20805 9759 21125 9760
rect 5441 9618 5507 9621
rect 5901 9618 5967 9621
rect 5441 9616 5967 9618
rect 5441 9560 5446 9616
rect 5502 9560 5906 9616
rect 5962 9560 5967 9616
rect 5441 9558 5967 9560
rect 5441 9555 5507 9558
rect 5901 9555 5967 9558
rect 13721 9618 13787 9621
rect 15101 9618 15167 9621
rect 13721 9616 15167 9618
rect 13721 9560 13726 9616
rect 13782 9560 15106 9616
rect 15162 9560 15167 9616
rect 13721 9558 15167 9560
rect 13721 9555 13787 9558
rect 15101 9555 15167 9558
rect 2313 9482 2379 9485
rect 6177 9482 6243 9485
rect 2313 9480 6243 9482
rect 2313 9424 2318 9480
rect 2374 9424 6182 9480
rect 6238 9424 6243 9480
rect 2313 9422 6243 9424
rect 2313 9419 2379 9422
rect 6177 9419 6243 9422
rect 5909 9280 6229 9281
rect 0 9210 800 9240
rect 5909 9216 5917 9280
rect 5981 9216 5997 9280
rect 6061 9216 6077 9280
rect 6141 9216 6157 9280
rect 6221 9216 6229 9280
rect 5909 9215 6229 9216
rect 15840 9280 16160 9281
rect 15840 9216 15848 9280
rect 15912 9216 15928 9280
rect 15992 9216 16008 9280
rect 16072 9216 16088 9280
rect 16152 9216 16160 9280
rect 15840 9215 16160 9216
rect 25770 9280 26090 9281
rect 25770 9216 25778 9280
rect 25842 9216 25858 9280
rect 25922 9216 25938 9280
rect 26002 9216 26018 9280
rect 26082 9216 26090 9280
rect 25770 9215 26090 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 17769 9074 17835 9077
rect 18229 9074 18295 9077
rect 17769 9072 18295 9074
rect 17769 9016 17774 9072
rect 17830 9016 18234 9072
rect 18290 9016 18295 9072
rect 17769 9014 18295 9016
rect 17769 9011 17835 9014
rect 18229 9011 18295 9014
rect 14089 8938 14155 8941
rect 16297 8938 16363 8941
rect 14089 8936 16363 8938
rect 14089 8880 14094 8936
rect 14150 8880 16302 8936
rect 16358 8880 16363 8936
rect 14089 8878 16363 8880
rect 14089 8875 14155 8878
rect 16297 8875 16363 8878
rect 30005 8938 30071 8941
rect 31200 8938 32000 8968
rect 30005 8936 32000 8938
rect 30005 8880 30010 8936
rect 30066 8880 32000 8936
rect 30005 8878 32000 8880
rect 30005 8875 30071 8878
rect 31200 8848 32000 8878
rect 10874 8736 11194 8737
rect 10874 8672 10882 8736
rect 10946 8672 10962 8736
rect 11026 8672 11042 8736
rect 11106 8672 11122 8736
rect 11186 8672 11194 8736
rect 10874 8671 11194 8672
rect 20805 8736 21125 8737
rect 20805 8672 20813 8736
rect 20877 8672 20893 8736
rect 20957 8672 20973 8736
rect 21037 8672 21053 8736
rect 21117 8672 21125 8736
rect 20805 8671 21125 8672
rect 0 8394 800 8424
rect 1393 8394 1459 8397
rect 0 8392 1459 8394
rect 0 8336 1398 8392
rect 1454 8336 1459 8392
rect 0 8334 1459 8336
rect 0 8304 800 8334
rect 1393 8331 1459 8334
rect 20529 8394 20595 8397
rect 22277 8394 22343 8397
rect 20529 8392 22343 8394
rect 20529 8336 20534 8392
rect 20590 8336 22282 8392
rect 22338 8336 22343 8392
rect 20529 8334 22343 8336
rect 20529 8331 20595 8334
rect 22277 8331 22343 8334
rect 5909 8192 6229 8193
rect 5909 8128 5917 8192
rect 5981 8128 5997 8192
rect 6061 8128 6077 8192
rect 6141 8128 6157 8192
rect 6221 8128 6229 8192
rect 5909 8127 6229 8128
rect 15840 8192 16160 8193
rect 15840 8128 15848 8192
rect 15912 8128 15928 8192
rect 15992 8128 16008 8192
rect 16072 8128 16088 8192
rect 16152 8128 16160 8192
rect 15840 8127 16160 8128
rect 25770 8192 26090 8193
rect 25770 8128 25778 8192
rect 25842 8128 25858 8192
rect 25922 8128 25938 8192
rect 26002 8128 26018 8192
rect 26082 8128 26090 8192
rect 25770 8127 26090 8128
rect 10041 7986 10107 7989
rect 10317 7986 10383 7989
rect 10041 7984 10383 7986
rect 10041 7928 10046 7984
rect 10102 7928 10322 7984
rect 10378 7928 10383 7984
rect 10041 7926 10383 7928
rect 10041 7923 10107 7926
rect 10317 7923 10383 7926
rect 0 7714 800 7744
rect 1393 7714 1459 7717
rect 0 7712 1459 7714
rect 0 7656 1398 7712
rect 1454 7656 1459 7712
rect 0 7654 1459 7656
rect 0 7624 800 7654
rect 1393 7651 1459 7654
rect 10874 7648 11194 7649
rect 10874 7584 10882 7648
rect 10946 7584 10962 7648
rect 11026 7584 11042 7648
rect 11106 7584 11122 7648
rect 11186 7584 11194 7648
rect 10874 7583 11194 7584
rect 20805 7648 21125 7649
rect 20805 7584 20813 7648
rect 20877 7584 20893 7648
rect 20957 7584 20973 7648
rect 21037 7584 21053 7648
rect 21117 7584 21125 7648
rect 20805 7583 21125 7584
rect 5909 7104 6229 7105
rect 5909 7040 5917 7104
rect 5981 7040 5997 7104
rect 6061 7040 6077 7104
rect 6141 7040 6157 7104
rect 6221 7040 6229 7104
rect 5909 7039 6229 7040
rect 15840 7104 16160 7105
rect 15840 7040 15848 7104
rect 15912 7040 15928 7104
rect 15992 7040 16008 7104
rect 16072 7040 16088 7104
rect 16152 7040 16160 7104
rect 15840 7039 16160 7040
rect 25770 7104 26090 7105
rect 25770 7040 25778 7104
rect 25842 7040 25858 7104
rect 25922 7040 25938 7104
rect 26002 7040 26018 7104
rect 26082 7040 26090 7104
rect 25770 7039 26090 7040
rect 30005 7034 30071 7037
rect 31200 7034 32000 7064
rect 30005 7032 32000 7034
rect 30005 6976 30010 7032
rect 30066 6976 32000 7032
rect 30005 6974 32000 6976
rect 30005 6971 30071 6974
rect 31200 6944 32000 6974
rect 0 6898 800 6928
rect 2037 6898 2103 6901
rect 0 6896 2103 6898
rect 0 6840 2042 6896
rect 2098 6840 2103 6896
rect 0 6838 2103 6840
rect 0 6808 800 6838
rect 2037 6835 2103 6838
rect 10593 6762 10659 6765
rect 16205 6762 16271 6765
rect 10593 6760 16271 6762
rect 10593 6704 10598 6760
rect 10654 6704 16210 6760
rect 16266 6704 16271 6760
rect 10593 6702 16271 6704
rect 10593 6699 10659 6702
rect 16205 6699 16271 6702
rect 10874 6560 11194 6561
rect 10874 6496 10882 6560
rect 10946 6496 10962 6560
rect 11026 6496 11042 6560
rect 11106 6496 11122 6560
rect 11186 6496 11194 6560
rect 10874 6495 11194 6496
rect 20805 6560 21125 6561
rect 20805 6496 20813 6560
rect 20877 6496 20893 6560
rect 20957 6496 20973 6560
rect 21037 6496 21053 6560
rect 21117 6496 21125 6560
rect 20805 6495 21125 6496
rect 6085 6354 6151 6357
rect 6913 6354 6979 6357
rect 6085 6352 6979 6354
rect 6085 6296 6090 6352
rect 6146 6296 6918 6352
rect 6974 6296 6979 6352
rect 6085 6294 6979 6296
rect 6085 6291 6151 6294
rect 6913 6291 6979 6294
rect 0 6218 800 6248
rect 2773 6218 2839 6221
rect 0 6216 2839 6218
rect 0 6160 2778 6216
rect 2834 6160 2839 6216
rect 0 6158 2839 6160
rect 0 6128 800 6158
rect 2773 6155 2839 6158
rect 5909 6016 6229 6017
rect 5909 5952 5917 6016
rect 5981 5952 5997 6016
rect 6061 5952 6077 6016
rect 6141 5952 6157 6016
rect 6221 5952 6229 6016
rect 5909 5951 6229 5952
rect 15840 6016 16160 6017
rect 15840 5952 15848 6016
rect 15912 5952 15928 6016
rect 15992 5952 16008 6016
rect 16072 5952 16088 6016
rect 16152 5952 16160 6016
rect 15840 5951 16160 5952
rect 25770 6016 26090 6017
rect 25770 5952 25778 6016
rect 25842 5952 25858 6016
rect 25922 5952 25938 6016
rect 26002 5952 26018 6016
rect 26082 5952 26090 6016
rect 25770 5951 26090 5952
rect 0 5538 800 5568
rect 1209 5538 1275 5541
rect 0 5536 1275 5538
rect 0 5480 1214 5536
rect 1270 5480 1275 5536
rect 0 5478 1275 5480
rect 0 5448 800 5478
rect 1209 5475 1275 5478
rect 10874 5472 11194 5473
rect 10874 5408 10882 5472
rect 10946 5408 10962 5472
rect 11026 5408 11042 5472
rect 11106 5408 11122 5472
rect 11186 5408 11194 5472
rect 10874 5407 11194 5408
rect 20805 5472 21125 5473
rect 20805 5408 20813 5472
rect 20877 5408 20893 5472
rect 20957 5408 20973 5472
rect 21037 5408 21053 5472
rect 21117 5408 21125 5472
rect 20805 5407 21125 5408
rect 30005 4994 30071 4997
rect 31200 4994 32000 5024
rect 30005 4992 32000 4994
rect 30005 4936 30010 4992
rect 30066 4936 32000 4992
rect 30005 4934 32000 4936
rect 30005 4931 30071 4934
rect 5909 4928 6229 4929
rect 5909 4864 5917 4928
rect 5981 4864 5997 4928
rect 6061 4864 6077 4928
rect 6141 4864 6157 4928
rect 6221 4864 6229 4928
rect 5909 4863 6229 4864
rect 15840 4928 16160 4929
rect 15840 4864 15848 4928
rect 15912 4864 15928 4928
rect 15992 4864 16008 4928
rect 16072 4864 16088 4928
rect 16152 4864 16160 4928
rect 15840 4863 16160 4864
rect 25770 4928 26090 4929
rect 25770 4864 25778 4928
rect 25842 4864 25858 4928
rect 25922 4864 25938 4928
rect 26002 4864 26018 4928
rect 26082 4864 26090 4928
rect 31200 4904 32000 4934
rect 25770 4863 26090 4864
rect 0 4722 800 4752
rect 1393 4722 1459 4725
rect 0 4720 1459 4722
rect 0 4664 1398 4720
rect 1454 4664 1459 4720
rect 0 4662 1459 4664
rect 0 4632 800 4662
rect 1393 4659 1459 4662
rect 10874 4384 11194 4385
rect 10874 4320 10882 4384
rect 10946 4320 10962 4384
rect 11026 4320 11042 4384
rect 11106 4320 11122 4384
rect 11186 4320 11194 4384
rect 10874 4319 11194 4320
rect 20805 4384 21125 4385
rect 20805 4320 20813 4384
rect 20877 4320 20893 4384
rect 20957 4320 20973 4384
rect 21037 4320 21053 4384
rect 21117 4320 21125 4384
rect 20805 4319 21125 4320
rect 0 4042 800 4072
rect 1393 4042 1459 4045
rect 0 4040 1459 4042
rect 0 3984 1398 4040
rect 1454 3984 1459 4040
rect 0 3982 1459 3984
rect 0 3952 800 3982
rect 1393 3979 1459 3982
rect 3049 4042 3115 4045
rect 5809 4042 5875 4045
rect 3049 4040 5875 4042
rect 3049 3984 3054 4040
rect 3110 3984 5814 4040
rect 5870 3984 5875 4040
rect 3049 3982 5875 3984
rect 3049 3979 3115 3982
rect 5809 3979 5875 3982
rect 5909 3840 6229 3841
rect 5909 3776 5917 3840
rect 5981 3776 5997 3840
rect 6061 3776 6077 3840
rect 6141 3776 6157 3840
rect 6221 3776 6229 3840
rect 5909 3775 6229 3776
rect 15840 3840 16160 3841
rect 15840 3776 15848 3840
rect 15912 3776 15928 3840
rect 15992 3776 16008 3840
rect 16072 3776 16088 3840
rect 16152 3776 16160 3840
rect 15840 3775 16160 3776
rect 25770 3840 26090 3841
rect 25770 3776 25778 3840
rect 25842 3776 25858 3840
rect 25922 3776 25938 3840
rect 26002 3776 26018 3840
rect 26082 3776 26090 3840
rect 25770 3775 26090 3776
rect 10874 3296 11194 3297
rect 0 3226 800 3256
rect 10874 3232 10882 3296
rect 10946 3232 10962 3296
rect 11026 3232 11042 3296
rect 11106 3232 11122 3296
rect 11186 3232 11194 3296
rect 10874 3231 11194 3232
rect 20805 3296 21125 3297
rect 20805 3232 20813 3296
rect 20877 3232 20893 3296
rect 20957 3232 20973 3296
rect 21037 3232 21053 3296
rect 21117 3232 21125 3296
rect 20805 3231 21125 3232
rect 2773 3226 2839 3229
rect 0 3224 2839 3226
rect 0 3168 2778 3224
rect 2834 3168 2839 3224
rect 0 3166 2839 3168
rect 0 3136 800 3166
rect 2773 3163 2839 3166
rect 30005 2954 30071 2957
rect 31200 2954 32000 2984
rect 30005 2952 32000 2954
rect 30005 2896 30010 2952
rect 30066 2896 32000 2952
rect 30005 2894 32000 2896
rect 30005 2891 30071 2894
rect 31200 2864 32000 2894
rect 5909 2752 6229 2753
rect 5909 2688 5917 2752
rect 5981 2688 5997 2752
rect 6061 2688 6077 2752
rect 6141 2688 6157 2752
rect 6221 2688 6229 2752
rect 5909 2687 6229 2688
rect 15840 2752 16160 2753
rect 15840 2688 15848 2752
rect 15912 2688 15928 2752
rect 15992 2688 16008 2752
rect 16072 2688 16088 2752
rect 16152 2688 16160 2752
rect 15840 2687 16160 2688
rect 25770 2752 26090 2753
rect 25770 2688 25778 2752
rect 25842 2688 25858 2752
rect 25922 2688 25938 2752
rect 26002 2688 26018 2752
rect 26082 2688 26090 2752
rect 25770 2687 26090 2688
rect 0 2546 800 2576
rect 1853 2546 1919 2549
rect 0 2544 1919 2546
rect 0 2488 1858 2544
rect 1914 2488 1919 2544
rect 0 2486 1919 2488
rect 0 2456 800 2486
rect 1853 2483 1919 2486
rect 10874 2208 11194 2209
rect 10874 2144 10882 2208
rect 10946 2144 10962 2208
rect 11026 2144 11042 2208
rect 11106 2144 11122 2208
rect 11186 2144 11194 2208
rect 10874 2143 11194 2144
rect 20805 2208 21125 2209
rect 20805 2144 20813 2208
rect 20877 2144 20893 2208
rect 20957 2144 20973 2208
rect 21037 2144 21053 2208
rect 21117 2144 21125 2208
rect 20805 2143 21125 2144
rect 0 1730 800 1760
rect 2773 1730 2839 1733
rect 0 1728 2839 1730
rect 0 1672 2778 1728
rect 2834 1672 2839 1728
rect 0 1670 2839 1672
rect 0 1640 800 1670
rect 2773 1667 2839 1670
rect 0 1050 800 1080
rect 2865 1050 2931 1053
rect 0 1048 2931 1050
rect 0 992 2870 1048
rect 2926 992 2931 1048
rect 0 990 2931 992
rect 0 960 800 990
rect 2865 987 2931 990
rect 28901 1050 28967 1053
rect 31200 1050 32000 1080
rect 28901 1048 32000 1050
rect 28901 992 28906 1048
rect 28962 992 32000 1048
rect 28901 990 32000 992
rect 28901 987 28967 990
rect 31200 960 32000 990
rect 0 370 800 400
rect 2957 370 3023 373
rect 0 368 3023 370
rect 0 312 2962 368
rect 3018 312 3023 368
rect 0 310 3023 312
rect 0 280 800 310
rect 2957 307 3023 310
<< via3 >>
rect 10882 45724 10946 45728
rect 10882 45668 10886 45724
rect 10886 45668 10942 45724
rect 10942 45668 10946 45724
rect 10882 45664 10946 45668
rect 10962 45724 11026 45728
rect 10962 45668 10966 45724
rect 10966 45668 11022 45724
rect 11022 45668 11026 45724
rect 10962 45664 11026 45668
rect 11042 45724 11106 45728
rect 11042 45668 11046 45724
rect 11046 45668 11102 45724
rect 11102 45668 11106 45724
rect 11042 45664 11106 45668
rect 11122 45724 11186 45728
rect 11122 45668 11126 45724
rect 11126 45668 11182 45724
rect 11182 45668 11186 45724
rect 11122 45664 11186 45668
rect 20813 45724 20877 45728
rect 20813 45668 20817 45724
rect 20817 45668 20873 45724
rect 20873 45668 20877 45724
rect 20813 45664 20877 45668
rect 20893 45724 20957 45728
rect 20893 45668 20897 45724
rect 20897 45668 20953 45724
rect 20953 45668 20957 45724
rect 20893 45664 20957 45668
rect 20973 45724 21037 45728
rect 20973 45668 20977 45724
rect 20977 45668 21033 45724
rect 21033 45668 21037 45724
rect 20973 45664 21037 45668
rect 21053 45724 21117 45728
rect 21053 45668 21057 45724
rect 21057 45668 21113 45724
rect 21113 45668 21117 45724
rect 21053 45664 21117 45668
rect 5917 45180 5981 45184
rect 5917 45124 5921 45180
rect 5921 45124 5977 45180
rect 5977 45124 5981 45180
rect 5917 45120 5981 45124
rect 5997 45180 6061 45184
rect 5997 45124 6001 45180
rect 6001 45124 6057 45180
rect 6057 45124 6061 45180
rect 5997 45120 6061 45124
rect 6077 45180 6141 45184
rect 6077 45124 6081 45180
rect 6081 45124 6137 45180
rect 6137 45124 6141 45180
rect 6077 45120 6141 45124
rect 6157 45180 6221 45184
rect 6157 45124 6161 45180
rect 6161 45124 6217 45180
rect 6217 45124 6221 45180
rect 6157 45120 6221 45124
rect 15848 45180 15912 45184
rect 15848 45124 15852 45180
rect 15852 45124 15908 45180
rect 15908 45124 15912 45180
rect 15848 45120 15912 45124
rect 15928 45180 15992 45184
rect 15928 45124 15932 45180
rect 15932 45124 15988 45180
rect 15988 45124 15992 45180
rect 15928 45120 15992 45124
rect 16008 45180 16072 45184
rect 16008 45124 16012 45180
rect 16012 45124 16068 45180
rect 16068 45124 16072 45180
rect 16008 45120 16072 45124
rect 16088 45180 16152 45184
rect 16088 45124 16092 45180
rect 16092 45124 16148 45180
rect 16148 45124 16152 45180
rect 16088 45120 16152 45124
rect 25778 45180 25842 45184
rect 25778 45124 25782 45180
rect 25782 45124 25838 45180
rect 25838 45124 25842 45180
rect 25778 45120 25842 45124
rect 25858 45180 25922 45184
rect 25858 45124 25862 45180
rect 25862 45124 25918 45180
rect 25918 45124 25922 45180
rect 25858 45120 25922 45124
rect 25938 45180 26002 45184
rect 25938 45124 25942 45180
rect 25942 45124 25998 45180
rect 25998 45124 26002 45180
rect 25938 45120 26002 45124
rect 26018 45180 26082 45184
rect 26018 45124 26022 45180
rect 26022 45124 26078 45180
rect 26078 45124 26082 45180
rect 26018 45120 26082 45124
rect 10882 44636 10946 44640
rect 10882 44580 10886 44636
rect 10886 44580 10942 44636
rect 10942 44580 10946 44636
rect 10882 44576 10946 44580
rect 10962 44636 11026 44640
rect 10962 44580 10966 44636
rect 10966 44580 11022 44636
rect 11022 44580 11026 44636
rect 10962 44576 11026 44580
rect 11042 44636 11106 44640
rect 11042 44580 11046 44636
rect 11046 44580 11102 44636
rect 11102 44580 11106 44636
rect 11042 44576 11106 44580
rect 11122 44636 11186 44640
rect 11122 44580 11126 44636
rect 11126 44580 11182 44636
rect 11182 44580 11186 44636
rect 11122 44576 11186 44580
rect 20813 44636 20877 44640
rect 20813 44580 20817 44636
rect 20817 44580 20873 44636
rect 20873 44580 20877 44636
rect 20813 44576 20877 44580
rect 20893 44636 20957 44640
rect 20893 44580 20897 44636
rect 20897 44580 20953 44636
rect 20953 44580 20957 44636
rect 20893 44576 20957 44580
rect 20973 44636 21037 44640
rect 20973 44580 20977 44636
rect 20977 44580 21033 44636
rect 21033 44580 21037 44636
rect 20973 44576 21037 44580
rect 21053 44636 21117 44640
rect 21053 44580 21057 44636
rect 21057 44580 21113 44636
rect 21113 44580 21117 44636
rect 21053 44576 21117 44580
rect 5917 44092 5981 44096
rect 5917 44036 5921 44092
rect 5921 44036 5977 44092
rect 5977 44036 5981 44092
rect 5917 44032 5981 44036
rect 5997 44092 6061 44096
rect 5997 44036 6001 44092
rect 6001 44036 6057 44092
rect 6057 44036 6061 44092
rect 5997 44032 6061 44036
rect 6077 44092 6141 44096
rect 6077 44036 6081 44092
rect 6081 44036 6137 44092
rect 6137 44036 6141 44092
rect 6077 44032 6141 44036
rect 6157 44092 6221 44096
rect 6157 44036 6161 44092
rect 6161 44036 6217 44092
rect 6217 44036 6221 44092
rect 6157 44032 6221 44036
rect 15848 44092 15912 44096
rect 15848 44036 15852 44092
rect 15852 44036 15908 44092
rect 15908 44036 15912 44092
rect 15848 44032 15912 44036
rect 15928 44092 15992 44096
rect 15928 44036 15932 44092
rect 15932 44036 15988 44092
rect 15988 44036 15992 44092
rect 15928 44032 15992 44036
rect 16008 44092 16072 44096
rect 16008 44036 16012 44092
rect 16012 44036 16068 44092
rect 16068 44036 16072 44092
rect 16008 44032 16072 44036
rect 16088 44092 16152 44096
rect 16088 44036 16092 44092
rect 16092 44036 16148 44092
rect 16148 44036 16152 44092
rect 16088 44032 16152 44036
rect 25778 44092 25842 44096
rect 25778 44036 25782 44092
rect 25782 44036 25838 44092
rect 25838 44036 25842 44092
rect 25778 44032 25842 44036
rect 25858 44092 25922 44096
rect 25858 44036 25862 44092
rect 25862 44036 25918 44092
rect 25918 44036 25922 44092
rect 25858 44032 25922 44036
rect 25938 44092 26002 44096
rect 25938 44036 25942 44092
rect 25942 44036 25998 44092
rect 25998 44036 26002 44092
rect 25938 44032 26002 44036
rect 26018 44092 26082 44096
rect 26018 44036 26022 44092
rect 26022 44036 26078 44092
rect 26078 44036 26082 44092
rect 26018 44032 26082 44036
rect 10882 43548 10946 43552
rect 10882 43492 10886 43548
rect 10886 43492 10942 43548
rect 10942 43492 10946 43548
rect 10882 43488 10946 43492
rect 10962 43548 11026 43552
rect 10962 43492 10966 43548
rect 10966 43492 11022 43548
rect 11022 43492 11026 43548
rect 10962 43488 11026 43492
rect 11042 43548 11106 43552
rect 11042 43492 11046 43548
rect 11046 43492 11102 43548
rect 11102 43492 11106 43548
rect 11042 43488 11106 43492
rect 11122 43548 11186 43552
rect 11122 43492 11126 43548
rect 11126 43492 11182 43548
rect 11182 43492 11186 43548
rect 11122 43488 11186 43492
rect 20813 43548 20877 43552
rect 20813 43492 20817 43548
rect 20817 43492 20873 43548
rect 20873 43492 20877 43548
rect 20813 43488 20877 43492
rect 20893 43548 20957 43552
rect 20893 43492 20897 43548
rect 20897 43492 20953 43548
rect 20953 43492 20957 43548
rect 20893 43488 20957 43492
rect 20973 43548 21037 43552
rect 20973 43492 20977 43548
rect 20977 43492 21033 43548
rect 21033 43492 21037 43548
rect 20973 43488 21037 43492
rect 21053 43548 21117 43552
rect 21053 43492 21057 43548
rect 21057 43492 21113 43548
rect 21113 43492 21117 43548
rect 21053 43488 21117 43492
rect 5917 43004 5981 43008
rect 5917 42948 5921 43004
rect 5921 42948 5977 43004
rect 5977 42948 5981 43004
rect 5917 42944 5981 42948
rect 5997 43004 6061 43008
rect 5997 42948 6001 43004
rect 6001 42948 6057 43004
rect 6057 42948 6061 43004
rect 5997 42944 6061 42948
rect 6077 43004 6141 43008
rect 6077 42948 6081 43004
rect 6081 42948 6137 43004
rect 6137 42948 6141 43004
rect 6077 42944 6141 42948
rect 6157 43004 6221 43008
rect 6157 42948 6161 43004
rect 6161 42948 6217 43004
rect 6217 42948 6221 43004
rect 6157 42944 6221 42948
rect 15848 43004 15912 43008
rect 15848 42948 15852 43004
rect 15852 42948 15908 43004
rect 15908 42948 15912 43004
rect 15848 42944 15912 42948
rect 15928 43004 15992 43008
rect 15928 42948 15932 43004
rect 15932 42948 15988 43004
rect 15988 42948 15992 43004
rect 15928 42944 15992 42948
rect 16008 43004 16072 43008
rect 16008 42948 16012 43004
rect 16012 42948 16068 43004
rect 16068 42948 16072 43004
rect 16008 42944 16072 42948
rect 16088 43004 16152 43008
rect 16088 42948 16092 43004
rect 16092 42948 16148 43004
rect 16148 42948 16152 43004
rect 16088 42944 16152 42948
rect 25778 43004 25842 43008
rect 25778 42948 25782 43004
rect 25782 42948 25838 43004
rect 25838 42948 25842 43004
rect 25778 42944 25842 42948
rect 25858 43004 25922 43008
rect 25858 42948 25862 43004
rect 25862 42948 25918 43004
rect 25918 42948 25922 43004
rect 25858 42944 25922 42948
rect 25938 43004 26002 43008
rect 25938 42948 25942 43004
rect 25942 42948 25998 43004
rect 25998 42948 26002 43004
rect 25938 42944 26002 42948
rect 26018 43004 26082 43008
rect 26018 42948 26022 43004
rect 26022 42948 26078 43004
rect 26078 42948 26082 43004
rect 26018 42944 26082 42948
rect 10882 42460 10946 42464
rect 10882 42404 10886 42460
rect 10886 42404 10942 42460
rect 10942 42404 10946 42460
rect 10882 42400 10946 42404
rect 10962 42460 11026 42464
rect 10962 42404 10966 42460
rect 10966 42404 11022 42460
rect 11022 42404 11026 42460
rect 10962 42400 11026 42404
rect 11042 42460 11106 42464
rect 11042 42404 11046 42460
rect 11046 42404 11102 42460
rect 11102 42404 11106 42460
rect 11042 42400 11106 42404
rect 11122 42460 11186 42464
rect 11122 42404 11126 42460
rect 11126 42404 11182 42460
rect 11182 42404 11186 42460
rect 11122 42400 11186 42404
rect 20813 42460 20877 42464
rect 20813 42404 20817 42460
rect 20817 42404 20873 42460
rect 20873 42404 20877 42460
rect 20813 42400 20877 42404
rect 20893 42460 20957 42464
rect 20893 42404 20897 42460
rect 20897 42404 20953 42460
rect 20953 42404 20957 42460
rect 20893 42400 20957 42404
rect 20973 42460 21037 42464
rect 20973 42404 20977 42460
rect 20977 42404 21033 42460
rect 21033 42404 21037 42460
rect 20973 42400 21037 42404
rect 21053 42460 21117 42464
rect 21053 42404 21057 42460
rect 21057 42404 21113 42460
rect 21113 42404 21117 42460
rect 21053 42400 21117 42404
rect 5917 41916 5981 41920
rect 5917 41860 5921 41916
rect 5921 41860 5977 41916
rect 5977 41860 5981 41916
rect 5917 41856 5981 41860
rect 5997 41916 6061 41920
rect 5997 41860 6001 41916
rect 6001 41860 6057 41916
rect 6057 41860 6061 41916
rect 5997 41856 6061 41860
rect 6077 41916 6141 41920
rect 6077 41860 6081 41916
rect 6081 41860 6137 41916
rect 6137 41860 6141 41916
rect 6077 41856 6141 41860
rect 6157 41916 6221 41920
rect 6157 41860 6161 41916
rect 6161 41860 6217 41916
rect 6217 41860 6221 41916
rect 6157 41856 6221 41860
rect 15848 41916 15912 41920
rect 15848 41860 15852 41916
rect 15852 41860 15908 41916
rect 15908 41860 15912 41916
rect 15848 41856 15912 41860
rect 15928 41916 15992 41920
rect 15928 41860 15932 41916
rect 15932 41860 15988 41916
rect 15988 41860 15992 41916
rect 15928 41856 15992 41860
rect 16008 41916 16072 41920
rect 16008 41860 16012 41916
rect 16012 41860 16068 41916
rect 16068 41860 16072 41916
rect 16008 41856 16072 41860
rect 16088 41916 16152 41920
rect 16088 41860 16092 41916
rect 16092 41860 16148 41916
rect 16148 41860 16152 41916
rect 16088 41856 16152 41860
rect 25778 41916 25842 41920
rect 25778 41860 25782 41916
rect 25782 41860 25838 41916
rect 25838 41860 25842 41916
rect 25778 41856 25842 41860
rect 25858 41916 25922 41920
rect 25858 41860 25862 41916
rect 25862 41860 25918 41916
rect 25918 41860 25922 41916
rect 25858 41856 25922 41860
rect 25938 41916 26002 41920
rect 25938 41860 25942 41916
rect 25942 41860 25998 41916
rect 25998 41860 26002 41916
rect 25938 41856 26002 41860
rect 26018 41916 26082 41920
rect 26018 41860 26022 41916
rect 26022 41860 26078 41916
rect 26078 41860 26082 41916
rect 26018 41856 26082 41860
rect 10882 41372 10946 41376
rect 10882 41316 10886 41372
rect 10886 41316 10942 41372
rect 10942 41316 10946 41372
rect 10882 41312 10946 41316
rect 10962 41372 11026 41376
rect 10962 41316 10966 41372
rect 10966 41316 11022 41372
rect 11022 41316 11026 41372
rect 10962 41312 11026 41316
rect 11042 41372 11106 41376
rect 11042 41316 11046 41372
rect 11046 41316 11102 41372
rect 11102 41316 11106 41372
rect 11042 41312 11106 41316
rect 11122 41372 11186 41376
rect 11122 41316 11126 41372
rect 11126 41316 11182 41372
rect 11182 41316 11186 41372
rect 11122 41312 11186 41316
rect 20813 41372 20877 41376
rect 20813 41316 20817 41372
rect 20817 41316 20873 41372
rect 20873 41316 20877 41372
rect 20813 41312 20877 41316
rect 20893 41372 20957 41376
rect 20893 41316 20897 41372
rect 20897 41316 20953 41372
rect 20953 41316 20957 41372
rect 20893 41312 20957 41316
rect 20973 41372 21037 41376
rect 20973 41316 20977 41372
rect 20977 41316 21033 41372
rect 21033 41316 21037 41372
rect 20973 41312 21037 41316
rect 21053 41372 21117 41376
rect 21053 41316 21057 41372
rect 21057 41316 21113 41372
rect 21113 41316 21117 41372
rect 21053 41312 21117 41316
rect 5917 40828 5981 40832
rect 5917 40772 5921 40828
rect 5921 40772 5977 40828
rect 5977 40772 5981 40828
rect 5917 40768 5981 40772
rect 5997 40828 6061 40832
rect 5997 40772 6001 40828
rect 6001 40772 6057 40828
rect 6057 40772 6061 40828
rect 5997 40768 6061 40772
rect 6077 40828 6141 40832
rect 6077 40772 6081 40828
rect 6081 40772 6137 40828
rect 6137 40772 6141 40828
rect 6077 40768 6141 40772
rect 6157 40828 6221 40832
rect 6157 40772 6161 40828
rect 6161 40772 6217 40828
rect 6217 40772 6221 40828
rect 6157 40768 6221 40772
rect 15848 40828 15912 40832
rect 15848 40772 15852 40828
rect 15852 40772 15908 40828
rect 15908 40772 15912 40828
rect 15848 40768 15912 40772
rect 15928 40828 15992 40832
rect 15928 40772 15932 40828
rect 15932 40772 15988 40828
rect 15988 40772 15992 40828
rect 15928 40768 15992 40772
rect 16008 40828 16072 40832
rect 16008 40772 16012 40828
rect 16012 40772 16068 40828
rect 16068 40772 16072 40828
rect 16008 40768 16072 40772
rect 16088 40828 16152 40832
rect 16088 40772 16092 40828
rect 16092 40772 16148 40828
rect 16148 40772 16152 40828
rect 16088 40768 16152 40772
rect 25778 40828 25842 40832
rect 25778 40772 25782 40828
rect 25782 40772 25838 40828
rect 25838 40772 25842 40828
rect 25778 40768 25842 40772
rect 25858 40828 25922 40832
rect 25858 40772 25862 40828
rect 25862 40772 25918 40828
rect 25918 40772 25922 40828
rect 25858 40768 25922 40772
rect 25938 40828 26002 40832
rect 25938 40772 25942 40828
rect 25942 40772 25998 40828
rect 25998 40772 26002 40828
rect 25938 40768 26002 40772
rect 26018 40828 26082 40832
rect 26018 40772 26022 40828
rect 26022 40772 26078 40828
rect 26078 40772 26082 40828
rect 26018 40768 26082 40772
rect 10882 40284 10946 40288
rect 10882 40228 10886 40284
rect 10886 40228 10942 40284
rect 10942 40228 10946 40284
rect 10882 40224 10946 40228
rect 10962 40284 11026 40288
rect 10962 40228 10966 40284
rect 10966 40228 11022 40284
rect 11022 40228 11026 40284
rect 10962 40224 11026 40228
rect 11042 40284 11106 40288
rect 11042 40228 11046 40284
rect 11046 40228 11102 40284
rect 11102 40228 11106 40284
rect 11042 40224 11106 40228
rect 11122 40284 11186 40288
rect 11122 40228 11126 40284
rect 11126 40228 11182 40284
rect 11182 40228 11186 40284
rect 11122 40224 11186 40228
rect 20813 40284 20877 40288
rect 20813 40228 20817 40284
rect 20817 40228 20873 40284
rect 20873 40228 20877 40284
rect 20813 40224 20877 40228
rect 20893 40284 20957 40288
rect 20893 40228 20897 40284
rect 20897 40228 20953 40284
rect 20953 40228 20957 40284
rect 20893 40224 20957 40228
rect 20973 40284 21037 40288
rect 20973 40228 20977 40284
rect 20977 40228 21033 40284
rect 21033 40228 21037 40284
rect 20973 40224 21037 40228
rect 21053 40284 21117 40288
rect 21053 40228 21057 40284
rect 21057 40228 21113 40284
rect 21113 40228 21117 40284
rect 21053 40224 21117 40228
rect 5917 39740 5981 39744
rect 5917 39684 5921 39740
rect 5921 39684 5977 39740
rect 5977 39684 5981 39740
rect 5917 39680 5981 39684
rect 5997 39740 6061 39744
rect 5997 39684 6001 39740
rect 6001 39684 6057 39740
rect 6057 39684 6061 39740
rect 5997 39680 6061 39684
rect 6077 39740 6141 39744
rect 6077 39684 6081 39740
rect 6081 39684 6137 39740
rect 6137 39684 6141 39740
rect 6077 39680 6141 39684
rect 6157 39740 6221 39744
rect 6157 39684 6161 39740
rect 6161 39684 6217 39740
rect 6217 39684 6221 39740
rect 6157 39680 6221 39684
rect 15848 39740 15912 39744
rect 15848 39684 15852 39740
rect 15852 39684 15908 39740
rect 15908 39684 15912 39740
rect 15848 39680 15912 39684
rect 15928 39740 15992 39744
rect 15928 39684 15932 39740
rect 15932 39684 15988 39740
rect 15988 39684 15992 39740
rect 15928 39680 15992 39684
rect 16008 39740 16072 39744
rect 16008 39684 16012 39740
rect 16012 39684 16068 39740
rect 16068 39684 16072 39740
rect 16008 39680 16072 39684
rect 16088 39740 16152 39744
rect 16088 39684 16092 39740
rect 16092 39684 16148 39740
rect 16148 39684 16152 39740
rect 16088 39680 16152 39684
rect 25778 39740 25842 39744
rect 25778 39684 25782 39740
rect 25782 39684 25838 39740
rect 25838 39684 25842 39740
rect 25778 39680 25842 39684
rect 25858 39740 25922 39744
rect 25858 39684 25862 39740
rect 25862 39684 25918 39740
rect 25918 39684 25922 39740
rect 25858 39680 25922 39684
rect 25938 39740 26002 39744
rect 25938 39684 25942 39740
rect 25942 39684 25998 39740
rect 25998 39684 26002 39740
rect 25938 39680 26002 39684
rect 26018 39740 26082 39744
rect 26018 39684 26022 39740
rect 26022 39684 26078 39740
rect 26078 39684 26082 39740
rect 26018 39680 26082 39684
rect 10882 39196 10946 39200
rect 10882 39140 10886 39196
rect 10886 39140 10942 39196
rect 10942 39140 10946 39196
rect 10882 39136 10946 39140
rect 10962 39196 11026 39200
rect 10962 39140 10966 39196
rect 10966 39140 11022 39196
rect 11022 39140 11026 39196
rect 10962 39136 11026 39140
rect 11042 39196 11106 39200
rect 11042 39140 11046 39196
rect 11046 39140 11102 39196
rect 11102 39140 11106 39196
rect 11042 39136 11106 39140
rect 11122 39196 11186 39200
rect 11122 39140 11126 39196
rect 11126 39140 11182 39196
rect 11182 39140 11186 39196
rect 11122 39136 11186 39140
rect 20813 39196 20877 39200
rect 20813 39140 20817 39196
rect 20817 39140 20873 39196
rect 20873 39140 20877 39196
rect 20813 39136 20877 39140
rect 20893 39196 20957 39200
rect 20893 39140 20897 39196
rect 20897 39140 20953 39196
rect 20953 39140 20957 39196
rect 20893 39136 20957 39140
rect 20973 39196 21037 39200
rect 20973 39140 20977 39196
rect 20977 39140 21033 39196
rect 21033 39140 21037 39196
rect 20973 39136 21037 39140
rect 21053 39196 21117 39200
rect 21053 39140 21057 39196
rect 21057 39140 21113 39196
rect 21113 39140 21117 39196
rect 21053 39136 21117 39140
rect 5917 38652 5981 38656
rect 5917 38596 5921 38652
rect 5921 38596 5977 38652
rect 5977 38596 5981 38652
rect 5917 38592 5981 38596
rect 5997 38652 6061 38656
rect 5997 38596 6001 38652
rect 6001 38596 6057 38652
rect 6057 38596 6061 38652
rect 5997 38592 6061 38596
rect 6077 38652 6141 38656
rect 6077 38596 6081 38652
rect 6081 38596 6137 38652
rect 6137 38596 6141 38652
rect 6077 38592 6141 38596
rect 6157 38652 6221 38656
rect 6157 38596 6161 38652
rect 6161 38596 6217 38652
rect 6217 38596 6221 38652
rect 6157 38592 6221 38596
rect 15848 38652 15912 38656
rect 15848 38596 15852 38652
rect 15852 38596 15908 38652
rect 15908 38596 15912 38652
rect 15848 38592 15912 38596
rect 15928 38652 15992 38656
rect 15928 38596 15932 38652
rect 15932 38596 15988 38652
rect 15988 38596 15992 38652
rect 15928 38592 15992 38596
rect 16008 38652 16072 38656
rect 16008 38596 16012 38652
rect 16012 38596 16068 38652
rect 16068 38596 16072 38652
rect 16008 38592 16072 38596
rect 16088 38652 16152 38656
rect 16088 38596 16092 38652
rect 16092 38596 16148 38652
rect 16148 38596 16152 38652
rect 16088 38592 16152 38596
rect 25778 38652 25842 38656
rect 25778 38596 25782 38652
rect 25782 38596 25838 38652
rect 25838 38596 25842 38652
rect 25778 38592 25842 38596
rect 25858 38652 25922 38656
rect 25858 38596 25862 38652
rect 25862 38596 25918 38652
rect 25918 38596 25922 38652
rect 25858 38592 25922 38596
rect 25938 38652 26002 38656
rect 25938 38596 25942 38652
rect 25942 38596 25998 38652
rect 25998 38596 26002 38652
rect 25938 38592 26002 38596
rect 26018 38652 26082 38656
rect 26018 38596 26022 38652
rect 26022 38596 26078 38652
rect 26078 38596 26082 38652
rect 26018 38592 26082 38596
rect 10882 38108 10946 38112
rect 10882 38052 10886 38108
rect 10886 38052 10942 38108
rect 10942 38052 10946 38108
rect 10882 38048 10946 38052
rect 10962 38108 11026 38112
rect 10962 38052 10966 38108
rect 10966 38052 11022 38108
rect 11022 38052 11026 38108
rect 10962 38048 11026 38052
rect 11042 38108 11106 38112
rect 11042 38052 11046 38108
rect 11046 38052 11102 38108
rect 11102 38052 11106 38108
rect 11042 38048 11106 38052
rect 11122 38108 11186 38112
rect 11122 38052 11126 38108
rect 11126 38052 11182 38108
rect 11182 38052 11186 38108
rect 11122 38048 11186 38052
rect 20813 38108 20877 38112
rect 20813 38052 20817 38108
rect 20817 38052 20873 38108
rect 20873 38052 20877 38108
rect 20813 38048 20877 38052
rect 20893 38108 20957 38112
rect 20893 38052 20897 38108
rect 20897 38052 20953 38108
rect 20953 38052 20957 38108
rect 20893 38048 20957 38052
rect 20973 38108 21037 38112
rect 20973 38052 20977 38108
rect 20977 38052 21033 38108
rect 21033 38052 21037 38108
rect 20973 38048 21037 38052
rect 21053 38108 21117 38112
rect 21053 38052 21057 38108
rect 21057 38052 21113 38108
rect 21113 38052 21117 38108
rect 21053 38048 21117 38052
rect 5917 37564 5981 37568
rect 5917 37508 5921 37564
rect 5921 37508 5977 37564
rect 5977 37508 5981 37564
rect 5917 37504 5981 37508
rect 5997 37564 6061 37568
rect 5997 37508 6001 37564
rect 6001 37508 6057 37564
rect 6057 37508 6061 37564
rect 5997 37504 6061 37508
rect 6077 37564 6141 37568
rect 6077 37508 6081 37564
rect 6081 37508 6137 37564
rect 6137 37508 6141 37564
rect 6077 37504 6141 37508
rect 6157 37564 6221 37568
rect 6157 37508 6161 37564
rect 6161 37508 6217 37564
rect 6217 37508 6221 37564
rect 6157 37504 6221 37508
rect 15848 37564 15912 37568
rect 15848 37508 15852 37564
rect 15852 37508 15908 37564
rect 15908 37508 15912 37564
rect 15848 37504 15912 37508
rect 15928 37564 15992 37568
rect 15928 37508 15932 37564
rect 15932 37508 15988 37564
rect 15988 37508 15992 37564
rect 15928 37504 15992 37508
rect 16008 37564 16072 37568
rect 16008 37508 16012 37564
rect 16012 37508 16068 37564
rect 16068 37508 16072 37564
rect 16008 37504 16072 37508
rect 16088 37564 16152 37568
rect 16088 37508 16092 37564
rect 16092 37508 16148 37564
rect 16148 37508 16152 37564
rect 16088 37504 16152 37508
rect 25778 37564 25842 37568
rect 25778 37508 25782 37564
rect 25782 37508 25838 37564
rect 25838 37508 25842 37564
rect 25778 37504 25842 37508
rect 25858 37564 25922 37568
rect 25858 37508 25862 37564
rect 25862 37508 25918 37564
rect 25918 37508 25922 37564
rect 25858 37504 25922 37508
rect 25938 37564 26002 37568
rect 25938 37508 25942 37564
rect 25942 37508 25998 37564
rect 25998 37508 26002 37564
rect 25938 37504 26002 37508
rect 26018 37564 26082 37568
rect 26018 37508 26022 37564
rect 26022 37508 26078 37564
rect 26078 37508 26082 37564
rect 26018 37504 26082 37508
rect 10882 37020 10946 37024
rect 10882 36964 10886 37020
rect 10886 36964 10942 37020
rect 10942 36964 10946 37020
rect 10882 36960 10946 36964
rect 10962 37020 11026 37024
rect 10962 36964 10966 37020
rect 10966 36964 11022 37020
rect 11022 36964 11026 37020
rect 10962 36960 11026 36964
rect 11042 37020 11106 37024
rect 11042 36964 11046 37020
rect 11046 36964 11102 37020
rect 11102 36964 11106 37020
rect 11042 36960 11106 36964
rect 11122 37020 11186 37024
rect 11122 36964 11126 37020
rect 11126 36964 11182 37020
rect 11182 36964 11186 37020
rect 11122 36960 11186 36964
rect 20813 37020 20877 37024
rect 20813 36964 20817 37020
rect 20817 36964 20873 37020
rect 20873 36964 20877 37020
rect 20813 36960 20877 36964
rect 20893 37020 20957 37024
rect 20893 36964 20897 37020
rect 20897 36964 20953 37020
rect 20953 36964 20957 37020
rect 20893 36960 20957 36964
rect 20973 37020 21037 37024
rect 20973 36964 20977 37020
rect 20977 36964 21033 37020
rect 21033 36964 21037 37020
rect 20973 36960 21037 36964
rect 21053 37020 21117 37024
rect 21053 36964 21057 37020
rect 21057 36964 21113 37020
rect 21113 36964 21117 37020
rect 21053 36960 21117 36964
rect 5917 36476 5981 36480
rect 5917 36420 5921 36476
rect 5921 36420 5977 36476
rect 5977 36420 5981 36476
rect 5917 36416 5981 36420
rect 5997 36476 6061 36480
rect 5997 36420 6001 36476
rect 6001 36420 6057 36476
rect 6057 36420 6061 36476
rect 5997 36416 6061 36420
rect 6077 36476 6141 36480
rect 6077 36420 6081 36476
rect 6081 36420 6137 36476
rect 6137 36420 6141 36476
rect 6077 36416 6141 36420
rect 6157 36476 6221 36480
rect 6157 36420 6161 36476
rect 6161 36420 6217 36476
rect 6217 36420 6221 36476
rect 6157 36416 6221 36420
rect 15848 36476 15912 36480
rect 15848 36420 15852 36476
rect 15852 36420 15908 36476
rect 15908 36420 15912 36476
rect 15848 36416 15912 36420
rect 15928 36476 15992 36480
rect 15928 36420 15932 36476
rect 15932 36420 15988 36476
rect 15988 36420 15992 36476
rect 15928 36416 15992 36420
rect 16008 36476 16072 36480
rect 16008 36420 16012 36476
rect 16012 36420 16068 36476
rect 16068 36420 16072 36476
rect 16008 36416 16072 36420
rect 16088 36476 16152 36480
rect 16088 36420 16092 36476
rect 16092 36420 16148 36476
rect 16148 36420 16152 36476
rect 16088 36416 16152 36420
rect 25778 36476 25842 36480
rect 25778 36420 25782 36476
rect 25782 36420 25838 36476
rect 25838 36420 25842 36476
rect 25778 36416 25842 36420
rect 25858 36476 25922 36480
rect 25858 36420 25862 36476
rect 25862 36420 25918 36476
rect 25918 36420 25922 36476
rect 25858 36416 25922 36420
rect 25938 36476 26002 36480
rect 25938 36420 25942 36476
rect 25942 36420 25998 36476
rect 25998 36420 26002 36476
rect 25938 36416 26002 36420
rect 26018 36476 26082 36480
rect 26018 36420 26022 36476
rect 26022 36420 26078 36476
rect 26078 36420 26082 36476
rect 26018 36416 26082 36420
rect 10882 35932 10946 35936
rect 10882 35876 10886 35932
rect 10886 35876 10942 35932
rect 10942 35876 10946 35932
rect 10882 35872 10946 35876
rect 10962 35932 11026 35936
rect 10962 35876 10966 35932
rect 10966 35876 11022 35932
rect 11022 35876 11026 35932
rect 10962 35872 11026 35876
rect 11042 35932 11106 35936
rect 11042 35876 11046 35932
rect 11046 35876 11102 35932
rect 11102 35876 11106 35932
rect 11042 35872 11106 35876
rect 11122 35932 11186 35936
rect 11122 35876 11126 35932
rect 11126 35876 11182 35932
rect 11182 35876 11186 35932
rect 11122 35872 11186 35876
rect 20813 35932 20877 35936
rect 20813 35876 20817 35932
rect 20817 35876 20873 35932
rect 20873 35876 20877 35932
rect 20813 35872 20877 35876
rect 20893 35932 20957 35936
rect 20893 35876 20897 35932
rect 20897 35876 20953 35932
rect 20953 35876 20957 35932
rect 20893 35872 20957 35876
rect 20973 35932 21037 35936
rect 20973 35876 20977 35932
rect 20977 35876 21033 35932
rect 21033 35876 21037 35932
rect 20973 35872 21037 35876
rect 21053 35932 21117 35936
rect 21053 35876 21057 35932
rect 21057 35876 21113 35932
rect 21113 35876 21117 35932
rect 21053 35872 21117 35876
rect 5917 35388 5981 35392
rect 5917 35332 5921 35388
rect 5921 35332 5977 35388
rect 5977 35332 5981 35388
rect 5917 35328 5981 35332
rect 5997 35388 6061 35392
rect 5997 35332 6001 35388
rect 6001 35332 6057 35388
rect 6057 35332 6061 35388
rect 5997 35328 6061 35332
rect 6077 35388 6141 35392
rect 6077 35332 6081 35388
rect 6081 35332 6137 35388
rect 6137 35332 6141 35388
rect 6077 35328 6141 35332
rect 6157 35388 6221 35392
rect 6157 35332 6161 35388
rect 6161 35332 6217 35388
rect 6217 35332 6221 35388
rect 6157 35328 6221 35332
rect 15848 35388 15912 35392
rect 15848 35332 15852 35388
rect 15852 35332 15908 35388
rect 15908 35332 15912 35388
rect 15848 35328 15912 35332
rect 15928 35388 15992 35392
rect 15928 35332 15932 35388
rect 15932 35332 15988 35388
rect 15988 35332 15992 35388
rect 15928 35328 15992 35332
rect 16008 35388 16072 35392
rect 16008 35332 16012 35388
rect 16012 35332 16068 35388
rect 16068 35332 16072 35388
rect 16008 35328 16072 35332
rect 16088 35388 16152 35392
rect 16088 35332 16092 35388
rect 16092 35332 16148 35388
rect 16148 35332 16152 35388
rect 16088 35328 16152 35332
rect 25778 35388 25842 35392
rect 25778 35332 25782 35388
rect 25782 35332 25838 35388
rect 25838 35332 25842 35388
rect 25778 35328 25842 35332
rect 25858 35388 25922 35392
rect 25858 35332 25862 35388
rect 25862 35332 25918 35388
rect 25918 35332 25922 35388
rect 25858 35328 25922 35332
rect 25938 35388 26002 35392
rect 25938 35332 25942 35388
rect 25942 35332 25998 35388
rect 25998 35332 26002 35388
rect 25938 35328 26002 35332
rect 26018 35388 26082 35392
rect 26018 35332 26022 35388
rect 26022 35332 26078 35388
rect 26078 35332 26082 35388
rect 26018 35328 26082 35332
rect 10882 34844 10946 34848
rect 10882 34788 10886 34844
rect 10886 34788 10942 34844
rect 10942 34788 10946 34844
rect 10882 34784 10946 34788
rect 10962 34844 11026 34848
rect 10962 34788 10966 34844
rect 10966 34788 11022 34844
rect 11022 34788 11026 34844
rect 10962 34784 11026 34788
rect 11042 34844 11106 34848
rect 11042 34788 11046 34844
rect 11046 34788 11102 34844
rect 11102 34788 11106 34844
rect 11042 34784 11106 34788
rect 11122 34844 11186 34848
rect 11122 34788 11126 34844
rect 11126 34788 11182 34844
rect 11182 34788 11186 34844
rect 11122 34784 11186 34788
rect 20813 34844 20877 34848
rect 20813 34788 20817 34844
rect 20817 34788 20873 34844
rect 20873 34788 20877 34844
rect 20813 34784 20877 34788
rect 20893 34844 20957 34848
rect 20893 34788 20897 34844
rect 20897 34788 20953 34844
rect 20953 34788 20957 34844
rect 20893 34784 20957 34788
rect 20973 34844 21037 34848
rect 20973 34788 20977 34844
rect 20977 34788 21033 34844
rect 21033 34788 21037 34844
rect 20973 34784 21037 34788
rect 21053 34844 21117 34848
rect 21053 34788 21057 34844
rect 21057 34788 21113 34844
rect 21113 34788 21117 34844
rect 21053 34784 21117 34788
rect 5917 34300 5981 34304
rect 5917 34244 5921 34300
rect 5921 34244 5977 34300
rect 5977 34244 5981 34300
rect 5917 34240 5981 34244
rect 5997 34300 6061 34304
rect 5997 34244 6001 34300
rect 6001 34244 6057 34300
rect 6057 34244 6061 34300
rect 5997 34240 6061 34244
rect 6077 34300 6141 34304
rect 6077 34244 6081 34300
rect 6081 34244 6137 34300
rect 6137 34244 6141 34300
rect 6077 34240 6141 34244
rect 6157 34300 6221 34304
rect 6157 34244 6161 34300
rect 6161 34244 6217 34300
rect 6217 34244 6221 34300
rect 6157 34240 6221 34244
rect 15848 34300 15912 34304
rect 15848 34244 15852 34300
rect 15852 34244 15908 34300
rect 15908 34244 15912 34300
rect 15848 34240 15912 34244
rect 15928 34300 15992 34304
rect 15928 34244 15932 34300
rect 15932 34244 15988 34300
rect 15988 34244 15992 34300
rect 15928 34240 15992 34244
rect 16008 34300 16072 34304
rect 16008 34244 16012 34300
rect 16012 34244 16068 34300
rect 16068 34244 16072 34300
rect 16008 34240 16072 34244
rect 16088 34300 16152 34304
rect 16088 34244 16092 34300
rect 16092 34244 16148 34300
rect 16148 34244 16152 34300
rect 16088 34240 16152 34244
rect 25778 34300 25842 34304
rect 25778 34244 25782 34300
rect 25782 34244 25838 34300
rect 25838 34244 25842 34300
rect 25778 34240 25842 34244
rect 25858 34300 25922 34304
rect 25858 34244 25862 34300
rect 25862 34244 25918 34300
rect 25918 34244 25922 34300
rect 25858 34240 25922 34244
rect 25938 34300 26002 34304
rect 25938 34244 25942 34300
rect 25942 34244 25998 34300
rect 25998 34244 26002 34300
rect 25938 34240 26002 34244
rect 26018 34300 26082 34304
rect 26018 34244 26022 34300
rect 26022 34244 26078 34300
rect 26078 34244 26082 34300
rect 26018 34240 26082 34244
rect 10882 33756 10946 33760
rect 10882 33700 10886 33756
rect 10886 33700 10942 33756
rect 10942 33700 10946 33756
rect 10882 33696 10946 33700
rect 10962 33756 11026 33760
rect 10962 33700 10966 33756
rect 10966 33700 11022 33756
rect 11022 33700 11026 33756
rect 10962 33696 11026 33700
rect 11042 33756 11106 33760
rect 11042 33700 11046 33756
rect 11046 33700 11102 33756
rect 11102 33700 11106 33756
rect 11042 33696 11106 33700
rect 11122 33756 11186 33760
rect 11122 33700 11126 33756
rect 11126 33700 11182 33756
rect 11182 33700 11186 33756
rect 11122 33696 11186 33700
rect 20813 33756 20877 33760
rect 20813 33700 20817 33756
rect 20817 33700 20873 33756
rect 20873 33700 20877 33756
rect 20813 33696 20877 33700
rect 20893 33756 20957 33760
rect 20893 33700 20897 33756
rect 20897 33700 20953 33756
rect 20953 33700 20957 33756
rect 20893 33696 20957 33700
rect 20973 33756 21037 33760
rect 20973 33700 20977 33756
rect 20977 33700 21033 33756
rect 21033 33700 21037 33756
rect 20973 33696 21037 33700
rect 21053 33756 21117 33760
rect 21053 33700 21057 33756
rect 21057 33700 21113 33756
rect 21113 33700 21117 33756
rect 21053 33696 21117 33700
rect 5917 33212 5981 33216
rect 5917 33156 5921 33212
rect 5921 33156 5977 33212
rect 5977 33156 5981 33212
rect 5917 33152 5981 33156
rect 5997 33212 6061 33216
rect 5997 33156 6001 33212
rect 6001 33156 6057 33212
rect 6057 33156 6061 33212
rect 5997 33152 6061 33156
rect 6077 33212 6141 33216
rect 6077 33156 6081 33212
rect 6081 33156 6137 33212
rect 6137 33156 6141 33212
rect 6077 33152 6141 33156
rect 6157 33212 6221 33216
rect 6157 33156 6161 33212
rect 6161 33156 6217 33212
rect 6217 33156 6221 33212
rect 6157 33152 6221 33156
rect 15848 33212 15912 33216
rect 15848 33156 15852 33212
rect 15852 33156 15908 33212
rect 15908 33156 15912 33212
rect 15848 33152 15912 33156
rect 15928 33212 15992 33216
rect 15928 33156 15932 33212
rect 15932 33156 15988 33212
rect 15988 33156 15992 33212
rect 15928 33152 15992 33156
rect 16008 33212 16072 33216
rect 16008 33156 16012 33212
rect 16012 33156 16068 33212
rect 16068 33156 16072 33212
rect 16008 33152 16072 33156
rect 16088 33212 16152 33216
rect 16088 33156 16092 33212
rect 16092 33156 16148 33212
rect 16148 33156 16152 33212
rect 16088 33152 16152 33156
rect 25778 33212 25842 33216
rect 25778 33156 25782 33212
rect 25782 33156 25838 33212
rect 25838 33156 25842 33212
rect 25778 33152 25842 33156
rect 25858 33212 25922 33216
rect 25858 33156 25862 33212
rect 25862 33156 25918 33212
rect 25918 33156 25922 33212
rect 25858 33152 25922 33156
rect 25938 33212 26002 33216
rect 25938 33156 25942 33212
rect 25942 33156 25998 33212
rect 25998 33156 26002 33212
rect 25938 33152 26002 33156
rect 26018 33212 26082 33216
rect 26018 33156 26022 33212
rect 26022 33156 26078 33212
rect 26078 33156 26082 33212
rect 26018 33152 26082 33156
rect 10882 32668 10946 32672
rect 10882 32612 10886 32668
rect 10886 32612 10942 32668
rect 10942 32612 10946 32668
rect 10882 32608 10946 32612
rect 10962 32668 11026 32672
rect 10962 32612 10966 32668
rect 10966 32612 11022 32668
rect 11022 32612 11026 32668
rect 10962 32608 11026 32612
rect 11042 32668 11106 32672
rect 11042 32612 11046 32668
rect 11046 32612 11102 32668
rect 11102 32612 11106 32668
rect 11042 32608 11106 32612
rect 11122 32668 11186 32672
rect 11122 32612 11126 32668
rect 11126 32612 11182 32668
rect 11182 32612 11186 32668
rect 11122 32608 11186 32612
rect 20813 32668 20877 32672
rect 20813 32612 20817 32668
rect 20817 32612 20873 32668
rect 20873 32612 20877 32668
rect 20813 32608 20877 32612
rect 20893 32668 20957 32672
rect 20893 32612 20897 32668
rect 20897 32612 20953 32668
rect 20953 32612 20957 32668
rect 20893 32608 20957 32612
rect 20973 32668 21037 32672
rect 20973 32612 20977 32668
rect 20977 32612 21033 32668
rect 21033 32612 21037 32668
rect 20973 32608 21037 32612
rect 21053 32668 21117 32672
rect 21053 32612 21057 32668
rect 21057 32612 21113 32668
rect 21113 32612 21117 32668
rect 21053 32608 21117 32612
rect 5917 32124 5981 32128
rect 5917 32068 5921 32124
rect 5921 32068 5977 32124
rect 5977 32068 5981 32124
rect 5917 32064 5981 32068
rect 5997 32124 6061 32128
rect 5997 32068 6001 32124
rect 6001 32068 6057 32124
rect 6057 32068 6061 32124
rect 5997 32064 6061 32068
rect 6077 32124 6141 32128
rect 6077 32068 6081 32124
rect 6081 32068 6137 32124
rect 6137 32068 6141 32124
rect 6077 32064 6141 32068
rect 6157 32124 6221 32128
rect 6157 32068 6161 32124
rect 6161 32068 6217 32124
rect 6217 32068 6221 32124
rect 6157 32064 6221 32068
rect 15848 32124 15912 32128
rect 15848 32068 15852 32124
rect 15852 32068 15908 32124
rect 15908 32068 15912 32124
rect 15848 32064 15912 32068
rect 15928 32124 15992 32128
rect 15928 32068 15932 32124
rect 15932 32068 15988 32124
rect 15988 32068 15992 32124
rect 15928 32064 15992 32068
rect 16008 32124 16072 32128
rect 16008 32068 16012 32124
rect 16012 32068 16068 32124
rect 16068 32068 16072 32124
rect 16008 32064 16072 32068
rect 16088 32124 16152 32128
rect 16088 32068 16092 32124
rect 16092 32068 16148 32124
rect 16148 32068 16152 32124
rect 16088 32064 16152 32068
rect 25778 32124 25842 32128
rect 25778 32068 25782 32124
rect 25782 32068 25838 32124
rect 25838 32068 25842 32124
rect 25778 32064 25842 32068
rect 25858 32124 25922 32128
rect 25858 32068 25862 32124
rect 25862 32068 25918 32124
rect 25918 32068 25922 32124
rect 25858 32064 25922 32068
rect 25938 32124 26002 32128
rect 25938 32068 25942 32124
rect 25942 32068 25998 32124
rect 25998 32068 26002 32124
rect 25938 32064 26002 32068
rect 26018 32124 26082 32128
rect 26018 32068 26022 32124
rect 26022 32068 26078 32124
rect 26078 32068 26082 32124
rect 26018 32064 26082 32068
rect 11284 31724 11348 31788
rect 10882 31580 10946 31584
rect 10882 31524 10886 31580
rect 10886 31524 10942 31580
rect 10942 31524 10946 31580
rect 10882 31520 10946 31524
rect 10962 31580 11026 31584
rect 10962 31524 10966 31580
rect 10966 31524 11022 31580
rect 11022 31524 11026 31580
rect 10962 31520 11026 31524
rect 11042 31580 11106 31584
rect 11042 31524 11046 31580
rect 11046 31524 11102 31580
rect 11102 31524 11106 31580
rect 11042 31520 11106 31524
rect 11122 31580 11186 31584
rect 11122 31524 11126 31580
rect 11126 31524 11182 31580
rect 11182 31524 11186 31580
rect 11122 31520 11186 31524
rect 20813 31580 20877 31584
rect 20813 31524 20817 31580
rect 20817 31524 20873 31580
rect 20873 31524 20877 31580
rect 20813 31520 20877 31524
rect 20893 31580 20957 31584
rect 20893 31524 20897 31580
rect 20897 31524 20953 31580
rect 20953 31524 20957 31580
rect 20893 31520 20957 31524
rect 20973 31580 21037 31584
rect 20973 31524 20977 31580
rect 20977 31524 21033 31580
rect 21033 31524 21037 31580
rect 20973 31520 21037 31524
rect 21053 31580 21117 31584
rect 21053 31524 21057 31580
rect 21057 31524 21113 31580
rect 21113 31524 21117 31580
rect 21053 31520 21117 31524
rect 5917 31036 5981 31040
rect 5917 30980 5921 31036
rect 5921 30980 5977 31036
rect 5977 30980 5981 31036
rect 5917 30976 5981 30980
rect 5997 31036 6061 31040
rect 5997 30980 6001 31036
rect 6001 30980 6057 31036
rect 6057 30980 6061 31036
rect 5997 30976 6061 30980
rect 6077 31036 6141 31040
rect 6077 30980 6081 31036
rect 6081 30980 6137 31036
rect 6137 30980 6141 31036
rect 6077 30976 6141 30980
rect 6157 31036 6221 31040
rect 6157 30980 6161 31036
rect 6161 30980 6217 31036
rect 6217 30980 6221 31036
rect 6157 30976 6221 30980
rect 15848 31036 15912 31040
rect 15848 30980 15852 31036
rect 15852 30980 15908 31036
rect 15908 30980 15912 31036
rect 15848 30976 15912 30980
rect 15928 31036 15992 31040
rect 15928 30980 15932 31036
rect 15932 30980 15988 31036
rect 15988 30980 15992 31036
rect 15928 30976 15992 30980
rect 16008 31036 16072 31040
rect 16008 30980 16012 31036
rect 16012 30980 16068 31036
rect 16068 30980 16072 31036
rect 16008 30976 16072 30980
rect 16088 31036 16152 31040
rect 16088 30980 16092 31036
rect 16092 30980 16148 31036
rect 16148 30980 16152 31036
rect 16088 30976 16152 30980
rect 25778 31036 25842 31040
rect 25778 30980 25782 31036
rect 25782 30980 25838 31036
rect 25838 30980 25842 31036
rect 25778 30976 25842 30980
rect 25858 31036 25922 31040
rect 25858 30980 25862 31036
rect 25862 30980 25918 31036
rect 25918 30980 25922 31036
rect 25858 30976 25922 30980
rect 25938 31036 26002 31040
rect 25938 30980 25942 31036
rect 25942 30980 25998 31036
rect 25998 30980 26002 31036
rect 25938 30976 26002 30980
rect 26018 31036 26082 31040
rect 26018 30980 26022 31036
rect 26022 30980 26078 31036
rect 26078 30980 26082 31036
rect 26018 30976 26082 30980
rect 10882 30492 10946 30496
rect 10882 30436 10886 30492
rect 10886 30436 10942 30492
rect 10942 30436 10946 30492
rect 10882 30432 10946 30436
rect 10962 30492 11026 30496
rect 10962 30436 10966 30492
rect 10966 30436 11022 30492
rect 11022 30436 11026 30492
rect 10962 30432 11026 30436
rect 11042 30492 11106 30496
rect 11042 30436 11046 30492
rect 11046 30436 11102 30492
rect 11102 30436 11106 30492
rect 11042 30432 11106 30436
rect 11122 30492 11186 30496
rect 11122 30436 11126 30492
rect 11126 30436 11182 30492
rect 11182 30436 11186 30492
rect 11122 30432 11186 30436
rect 20813 30492 20877 30496
rect 20813 30436 20817 30492
rect 20817 30436 20873 30492
rect 20873 30436 20877 30492
rect 20813 30432 20877 30436
rect 20893 30492 20957 30496
rect 20893 30436 20897 30492
rect 20897 30436 20953 30492
rect 20953 30436 20957 30492
rect 20893 30432 20957 30436
rect 20973 30492 21037 30496
rect 20973 30436 20977 30492
rect 20977 30436 21033 30492
rect 21033 30436 21037 30492
rect 20973 30432 21037 30436
rect 21053 30492 21117 30496
rect 21053 30436 21057 30492
rect 21057 30436 21113 30492
rect 21113 30436 21117 30492
rect 21053 30432 21117 30436
rect 5917 29948 5981 29952
rect 5917 29892 5921 29948
rect 5921 29892 5977 29948
rect 5977 29892 5981 29948
rect 5917 29888 5981 29892
rect 5997 29948 6061 29952
rect 5997 29892 6001 29948
rect 6001 29892 6057 29948
rect 6057 29892 6061 29948
rect 5997 29888 6061 29892
rect 6077 29948 6141 29952
rect 6077 29892 6081 29948
rect 6081 29892 6137 29948
rect 6137 29892 6141 29948
rect 6077 29888 6141 29892
rect 6157 29948 6221 29952
rect 6157 29892 6161 29948
rect 6161 29892 6217 29948
rect 6217 29892 6221 29948
rect 6157 29888 6221 29892
rect 15848 29948 15912 29952
rect 15848 29892 15852 29948
rect 15852 29892 15908 29948
rect 15908 29892 15912 29948
rect 15848 29888 15912 29892
rect 15928 29948 15992 29952
rect 15928 29892 15932 29948
rect 15932 29892 15988 29948
rect 15988 29892 15992 29948
rect 15928 29888 15992 29892
rect 16008 29948 16072 29952
rect 16008 29892 16012 29948
rect 16012 29892 16068 29948
rect 16068 29892 16072 29948
rect 16008 29888 16072 29892
rect 16088 29948 16152 29952
rect 16088 29892 16092 29948
rect 16092 29892 16148 29948
rect 16148 29892 16152 29948
rect 16088 29888 16152 29892
rect 25778 29948 25842 29952
rect 25778 29892 25782 29948
rect 25782 29892 25838 29948
rect 25838 29892 25842 29948
rect 25778 29888 25842 29892
rect 25858 29948 25922 29952
rect 25858 29892 25862 29948
rect 25862 29892 25918 29948
rect 25918 29892 25922 29948
rect 25858 29888 25922 29892
rect 25938 29948 26002 29952
rect 25938 29892 25942 29948
rect 25942 29892 25998 29948
rect 25998 29892 26002 29948
rect 25938 29888 26002 29892
rect 26018 29948 26082 29952
rect 26018 29892 26022 29948
rect 26022 29892 26078 29948
rect 26078 29892 26082 29948
rect 26018 29888 26082 29892
rect 10882 29404 10946 29408
rect 10882 29348 10886 29404
rect 10886 29348 10942 29404
rect 10942 29348 10946 29404
rect 10882 29344 10946 29348
rect 10962 29404 11026 29408
rect 10962 29348 10966 29404
rect 10966 29348 11022 29404
rect 11022 29348 11026 29404
rect 10962 29344 11026 29348
rect 11042 29404 11106 29408
rect 11042 29348 11046 29404
rect 11046 29348 11102 29404
rect 11102 29348 11106 29404
rect 11042 29344 11106 29348
rect 11122 29404 11186 29408
rect 11122 29348 11126 29404
rect 11126 29348 11182 29404
rect 11182 29348 11186 29404
rect 11122 29344 11186 29348
rect 20813 29404 20877 29408
rect 20813 29348 20817 29404
rect 20817 29348 20873 29404
rect 20873 29348 20877 29404
rect 20813 29344 20877 29348
rect 20893 29404 20957 29408
rect 20893 29348 20897 29404
rect 20897 29348 20953 29404
rect 20953 29348 20957 29404
rect 20893 29344 20957 29348
rect 20973 29404 21037 29408
rect 20973 29348 20977 29404
rect 20977 29348 21033 29404
rect 21033 29348 21037 29404
rect 20973 29344 21037 29348
rect 21053 29404 21117 29408
rect 21053 29348 21057 29404
rect 21057 29348 21113 29404
rect 21113 29348 21117 29404
rect 21053 29344 21117 29348
rect 5917 28860 5981 28864
rect 5917 28804 5921 28860
rect 5921 28804 5977 28860
rect 5977 28804 5981 28860
rect 5917 28800 5981 28804
rect 5997 28860 6061 28864
rect 5997 28804 6001 28860
rect 6001 28804 6057 28860
rect 6057 28804 6061 28860
rect 5997 28800 6061 28804
rect 6077 28860 6141 28864
rect 6077 28804 6081 28860
rect 6081 28804 6137 28860
rect 6137 28804 6141 28860
rect 6077 28800 6141 28804
rect 6157 28860 6221 28864
rect 6157 28804 6161 28860
rect 6161 28804 6217 28860
rect 6217 28804 6221 28860
rect 6157 28800 6221 28804
rect 15848 28860 15912 28864
rect 15848 28804 15852 28860
rect 15852 28804 15908 28860
rect 15908 28804 15912 28860
rect 15848 28800 15912 28804
rect 15928 28860 15992 28864
rect 15928 28804 15932 28860
rect 15932 28804 15988 28860
rect 15988 28804 15992 28860
rect 15928 28800 15992 28804
rect 16008 28860 16072 28864
rect 16008 28804 16012 28860
rect 16012 28804 16068 28860
rect 16068 28804 16072 28860
rect 16008 28800 16072 28804
rect 16088 28860 16152 28864
rect 16088 28804 16092 28860
rect 16092 28804 16148 28860
rect 16148 28804 16152 28860
rect 16088 28800 16152 28804
rect 25778 28860 25842 28864
rect 25778 28804 25782 28860
rect 25782 28804 25838 28860
rect 25838 28804 25842 28860
rect 25778 28800 25842 28804
rect 25858 28860 25922 28864
rect 25858 28804 25862 28860
rect 25862 28804 25918 28860
rect 25918 28804 25922 28860
rect 25858 28800 25922 28804
rect 25938 28860 26002 28864
rect 25938 28804 25942 28860
rect 25942 28804 25998 28860
rect 25998 28804 26002 28860
rect 25938 28800 26002 28804
rect 26018 28860 26082 28864
rect 26018 28804 26022 28860
rect 26022 28804 26078 28860
rect 26078 28804 26082 28860
rect 26018 28800 26082 28804
rect 10882 28316 10946 28320
rect 10882 28260 10886 28316
rect 10886 28260 10942 28316
rect 10942 28260 10946 28316
rect 10882 28256 10946 28260
rect 10962 28316 11026 28320
rect 10962 28260 10966 28316
rect 10966 28260 11022 28316
rect 11022 28260 11026 28316
rect 10962 28256 11026 28260
rect 11042 28316 11106 28320
rect 11042 28260 11046 28316
rect 11046 28260 11102 28316
rect 11102 28260 11106 28316
rect 11042 28256 11106 28260
rect 11122 28316 11186 28320
rect 11122 28260 11126 28316
rect 11126 28260 11182 28316
rect 11182 28260 11186 28316
rect 11122 28256 11186 28260
rect 20813 28316 20877 28320
rect 20813 28260 20817 28316
rect 20817 28260 20873 28316
rect 20873 28260 20877 28316
rect 20813 28256 20877 28260
rect 20893 28316 20957 28320
rect 20893 28260 20897 28316
rect 20897 28260 20953 28316
rect 20953 28260 20957 28316
rect 20893 28256 20957 28260
rect 20973 28316 21037 28320
rect 20973 28260 20977 28316
rect 20977 28260 21033 28316
rect 21033 28260 21037 28316
rect 20973 28256 21037 28260
rect 21053 28316 21117 28320
rect 21053 28260 21057 28316
rect 21057 28260 21113 28316
rect 21113 28260 21117 28316
rect 21053 28256 21117 28260
rect 5917 27772 5981 27776
rect 5917 27716 5921 27772
rect 5921 27716 5977 27772
rect 5977 27716 5981 27772
rect 5917 27712 5981 27716
rect 5997 27772 6061 27776
rect 5997 27716 6001 27772
rect 6001 27716 6057 27772
rect 6057 27716 6061 27772
rect 5997 27712 6061 27716
rect 6077 27772 6141 27776
rect 6077 27716 6081 27772
rect 6081 27716 6137 27772
rect 6137 27716 6141 27772
rect 6077 27712 6141 27716
rect 6157 27772 6221 27776
rect 6157 27716 6161 27772
rect 6161 27716 6217 27772
rect 6217 27716 6221 27772
rect 6157 27712 6221 27716
rect 15848 27772 15912 27776
rect 15848 27716 15852 27772
rect 15852 27716 15908 27772
rect 15908 27716 15912 27772
rect 15848 27712 15912 27716
rect 15928 27772 15992 27776
rect 15928 27716 15932 27772
rect 15932 27716 15988 27772
rect 15988 27716 15992 27772
rect 15928 27712 15992 27716
rect 16008 27772 16072 27776
rect 16008 27716 16012 27772
rect 16012 27716 16068 27772
rect 16068 27716 16072 27772
rect 16008 27712 16072 27716
rect 16088 27772 16152 27776
rect 16088 27716 16092 27772
rect 16092 27716 16148 27772
rect 16148 27716 16152 27772
rect 16088 27712 16152 27716
rect 25778 27772 25842 27776
rect 25778 27716 25782 27772
rect 25782 27716 25838 27772
rect 25838 27716 25842 27772
rect 25778 27712 25842 27716
rect 25858 27772 25922 27776
rect 25858 27716 25862 27772
rect 25862 27716 25918 27772
rect 25918 27716 25922 27772
rect 25858 27712 25922 27716
rect 25938 27772 26002 27776
rect 25938 27716 25942 27772
rect 25942 27716 25998 27772
rect 25998 27716 26002 27772
rect 25938 27712 26002 27716
rect 26018 27772 26082 27776
rect 26018 27716 26022 27772
rect 26022 27716 26078 27772
rect 26078 27716 26082 27772
rect 26018 27712 26082 27716
rect 17540 27372 17604 27436
rect 10882 27228 10946 27232
rect 10882 27172 10886 27228
rect 10886 27172 10942 27228
rect 10942 27172 10946 27228
rect 10882 27168 10946 27172
rect 10962 27228 11026 27232
rect 10962 27172 10966 27228
rect 10966 27172 11022 27228
rect 11022 27172 11026 27228
rect 10962 27168 11026 27172
rect 11042 27228 11106 27232
rect 11042 27172 11046 27228
rect 11046 27172 11102 27228
rect 11102 27172 11106 27228
rect 11042 27168 11106 27172
rect 11122 27228 11186 27232
rect 11122 27172 11126 27228
rect 11126 27172 11182 27228
rect 11182 27172 11186 27228
rect 11122 27168 11186 27172
rect 20813 27228 20877 27232
rect 20813 27172 20817 27228
rect 20817 27172 20873 27228
rect 20873 27172 20877 27228
rect 20813 27168 20877 27172
rect 20893 27228 20957 27232
rect 20893 27172 20897 27228
rect 20897 27172 20953 27228
rect 20953 27172 20957 27228
rect 20893 27168 20957 27172
rect 20973 27228 21037 27232
rect 20973 27172 20977 27228
rect 20977 27172 21033 27228
rect 21033 27172 21037 27228
rect 20973 27168 21037 27172
rect 21053 27228 21117 27232
rect 21053 27172 21057 27228
rect 21057 27172 21113 27228
rect 21113 27172 21117 27228
rect 21053 27168 21117 27172
rect 5917 26684 5981 26688
rect 5917 26628 5921 26684
rect 5921 26628 5977 26684
rect 5977 26628 5981 26684
rect 5917 26624 5981 26628
rect 5997 26684 6061 26688
rect 5997 26628 6001 26684
rect 6001 26628 6057 26684
rect 6057 26628 6061 26684
rect 5997 26624 6061 26628
rect 6077 26684 6141 26688
rect 6077 26628 6081 26684
rect 6081 26628 6137 26684
rect 6137 26628 6141 26684
rect 6077 26624 6141 26628
rect 6157 26684 6221 26688
rect 6157 26628 6161 26684
rect 6161 26628 6217 26684
rect 6217 26628 6221 26684
rect 6157 26624 6221 26628
rect 15848 26684 15912 26688
rect 15848 26628 15852 26684
rect 15852 26628 15908 26684
rect 15908 26628 15912 26684
rect 15848 26624 15912 26628
rect 15928 26684 15992 26688
rect 15928 26628 15932 26684
rect 15932 26628 15988 26684
rect 15988 26628 15992 26684
rect 15928 26624 15992 26628
rect 16008 26684 16072 26688
rect 16008 26628 16012 26684
rect 16012 26628 16068 26684
rect 16068 26628 16072 26684
rect 16008 26624 16072 26628
rect 16088 26684 16152 26688
rect 16088 26628 16092 26684
rect 16092 26628 16148 26684
rect 16148 26628 16152 26684
rect 16088 26624 16152 26628
rect 25778 26684 25842 26688
rect 25778 26628 25782 26684
rect 25782 26628 25838 26684
rect 25838 26628 25842 26684
rect 25778 26624 25842 26628
rect 25858 26684 25922 26688
rect 25858 26628 25862 26684
rect 25862 26628 25918 26684
rect 25918 26628 25922 26684
rect 25858 26624 25922 26628
rect 25938 26684 26002 26688
rect 25938 26628 25942 26684
rect 25942 26628 25998 26684
rect 25998 26628 26002 26684
rect 25938 26624 26002 26628
rect 26018 26684 26082 26688
rect 26018 26628 26022 26684
rect 26022 26628 26078 26684
rect 26078 26628 26082 26684
rect 26018 26624 26082 26628
rect 7972 26284 8036 26348
rect 10882 26140 10946 26144
rect 10882 26084 10886 26140
rect 10886 26084 10942 26140
rect 10942 26084 10946 26140
rect 10882 26080 10946 26084
rect 10962 26140 11026 26144
rect 10962 26084 10966 26140
rect 10966 26084 11022 26140
rect 11022 26084 11026 26140
rect 10962 26080 11026 26084
rect 11042 26140 11106 26144
rect 11042 26084 11046 26140
rect 11046 26084 11102 26140
rect 11102 26084 11106 26140
rect 11042 26080 11106 26084
rect 11122 26140 11186 26144
rect 11122 26084 11126 26140
rect 11126 26084 11182 26140
rect 11182 26084 11186 26140
rect 11122 26080 11186 26084
rect 20813 26140 20877 26144
rect 20813 26084 20817 26140
rect 20817 26084 20873 26140
rect 20873 26084 20877 26140
rect 20813 26080 20877 26084
rect 20893 26140 20957 26144
rect 20893 26084 20897 26140
rect 20897 26084 20953 26140
rect 20953 26084 20957 26140
rect 20893 26080 20957 26084
rect 20973 26140 21037 26144
rect 20973 26084 20977 26140
rect 20977 26084 21033 26140
rect 21033 26084 21037 26140
rect 20973 26080 21037 26084
rect 21053 26140 21117 26144
rect 21053 26084 21057 26140
rect 21057 26084 21113 26140
rect 21113 26084 21117 26140
rect 21053 26080 21117 26084
rect 5917 25596 5981 25600
rect 5917 25540 5921 25596
rect 5921 25540 5977 25596
rect 5977 25540 5981 25596
rect 5917 25536 5981 25540
rect 5997 25596 6061 25600
rect 5997 25540 6001 25596
rect 6001 25540 6057 25596
rect 6057 25540 6061 25596
rect 5997 25536 6061 25540
rect 6077 25596 6141 25600
rect 6077 25540 6081 25596
rect 6081 25540 6137 25596
rect 6137 25540 6141 25596
rect 6077 25536 6141 25540
rect 6157 25596 6221 25600
rect 6157 25540 6161 25596
rect 6161 25540 6217 25596
rect 6217 25540 6221 25596
rect 6157 25536 6221 25540
rect 15848 25596 15912 25600
rect 15848 25540 15852 25596
rect 15852 25540 15908 25596
rect 15908 25540 15912 25596
rect 15848 25536 15912 25540
rect 15928 25596 15992 25600
rect 15928 25540 15932 25596
rect 15932 25540 15988 25596
rect 15988 25540 15992 25596
rect 15928 25536 15992 25540
rect 16008 25596 16072 25600
rect 16008 25540 16012 25596
rect 16012 25540 16068 25596
rect 16068 25540 16072 25596
rect 16008 25536 16072 25540
rect 16088 25596 16152 25600
rect 16088 25540 16092 25596
rect 16092 25540 16148 25596
rect 16148 25540 16152 25596
rect 16088 25536 16152 25540
rect 25778 25596 25842 25600
rect 25778 25540 25782 25596
rect 25782 25540 25838 25596
rect 25838 25540 25842 25596
rect 25778 25536 25842 25540
rect 25858 25596 25922 25600
rect 25858 25540 25862 25596
rect 25862 25540 25918 25596
rect 25918 25540 25922 25596
rect 25858 25536 25922 25540
rect 25938 25596 26002 25600
rect 25938 25540 25942 25596
rect 25942 25540 25998 25596
rect 25998 25540 26002 25596
rect 25938 25536 26002 25540
rect 26018 25596 26082 25600
rect 26018 25540 26022 25596
rect 26022 25540 26078 25596
rect 26078 25540 26082 25596
rect 26018 25536 26082 25540
rect 10882 25052 10946 25056
rect 10882 24996 10886 25052
rect 10886 24996 10942 25052
rect 10942 24996 10946 25052
rect 10882 24992 10946 24996
rect 10962 25052 11026 25056
rect 10962 24996 10966 25052
rect 10966 24996 11022 25052
rect 11022 24996 11026 25052
rect 10962 24992 11026 24996
rect 11042 25052 11106 25056
rect 11042 24996 11046 25052
rect 11046 24996 11102 25052
rect 11102 24996 11106 25052
rect 11042 24992 11106 24996
rect 11122 25052 11186 25056
rect 11122 24996 11126 25052
rect 11126 24996 11182 25052
rect 11182 24996 11186 25052
rect 11122 24992 11186 24996
rect 20813 25052 20877 25056
rect 20813 24996 20817 25052
rect 20817 24996 20873 25052
rect 20873 24996 20877 25052
rect 20813 24992 20877 24996
rect 20893 25052 20957 25056
rect 20893 24996 20897 25052
rect 20897 24996 20953 25052
rect 20953 24996 20957 25052
rect 20893 24992 20957 24996
rect 20973 25052 21037 25056
rect 20973 24996 20977 25052
rect 20977 24996 21033 25052
rect 21033 24996 21037 25052
rect 20973 24992 21037 24996
rect 21053 25052 21117 25056
rect 21053 24996 21057 25052
rect 21057 24996 21113 25052
rect 21113 24996 21117 25052
rect 21053 24992 21117 24996
rect 5917 24508 5981 24512
rect 5917 24452 5921 24508
rect 5921 24452 5977 24508
rect 5977 24452 5981 24508
rect 5917 24448 5981 24452
rect 5997 24508 6061 24512
rect 5997 24452 6001 24508
rect 6001 24452 6057 24508
rect 6057 24452 6061 24508
rect 5997 24448 6061 24452
rect 6077 24508 6141 24512
rect 6077 24452 6081 24508
rect 6081 24452 6137 24508
rect 6137 24452 6141 24508
rect 6077 24448 6141 24452
rect 6157 24508 6221 24512
rect 6157 24452 6161 24508
rect 6161 24452 6217 24508
rect 6217 24452 6221 24508
rect 6157 24448 6221 24452
rect 15848 24508 15912 24512
rect 15848 24452 15852 24508
rect 15852 24452 15908 24508
rect 15908 24452 15912 24508
rect 15848 24448 15912 24452
rect 15928 24508 15992 24512
rect 15928 24452 15932 24508
rect 15932 24452 15988 24508
rect 15988 24452 15992 24508
rect 15928 24448 15992 24452
rect 16008 24508 16072 24512
rect 16008 24452 16012 24508
rect 16012 24452 16068 24508
rect 16068 24452 16072 24508
rect 16008 24448 16072 24452
rect 16088 24508 16152 24512
rect 16088 24452 16092 24508
rect 16092 24452 16148 24508
rect 16148 24452 16152 24508
rect 16088 24448 16152 24452
rect 25778 24508 25842 24512
rect 25778 24452 25782 24508
rect 25782 24452 25838 24508
rect 25838 24452 25842 24508
rect 25778 24448 25842 24452
rect 25858 24508 25922 24512
rect 25858 24452 25862 24508
rect 25862 24452 25918 24508
rect 25918 24452 25922 24508
rect 25858 24448 25922 24452
rect 25938 24508 26002 24512
rect 25938 24452 25942 24508
rect 25942 24452 25998 24508
rect 25998 24452 26002 24508
rect 25938 24448 26002 24452
rect 26018 24508 26082 24512
rect 26018 24452 26022 24508
rect 26022 24452 26078 24508
rect 26078 24452 26082 24508
rect 26018 24448 26082 24452
rect 10882 23964 10946 23968
rect 10882 23908 10886 23964
rect 10886 23908 10942 23964
rect 10942 23908 10946 23964
rect 10882 23904 10946 23908
rect 10962 23964 11026 23968
rect 10962 23908 10966 23964
rect 10966 23908 11022 23964
rect 11022 23908 11026 23964
rect 10962 23904 11026 23908
rect 11042 23964 11106 23968
rect 11042 23908 11046 23964
rect 11046 23908 11102 23964
rect 11102 23908 11106 23964
rect 11042 23904 11106 23908
rect 11122 23964 11186 23968
rect 11122 23908 11126 23964
rect 11126 23908 11182 23964
rect 11182 23908 11186 23964
rect 11122 23904 11186 23908
rect 20813 23964 20877 23968
rect 20813 23908 20817 23964
rect 20817 23908 20873 23964
rect 20873 23908 20877 23964
rect 20813 23904 20877 23908
rect 20893 23964 20957 23968
rect 20893 23908 20897 23964
rect 20897 23908 20953 23964
rect 20953 23908 20957 23964
rect 20893 23904 20957 23908
rect 20973 23964 21037 23968
rect 20973 23908 20977 23964
rect 20977 23908 21033 23964
rect 21033 23908 21037 23964
rect 20973 23904 21037 23908
rect 21053 23964 21117 23968
rect 21053 23908 21057 23964
rect 21057 23908 21113 23964
rect 21113 23908 21117 23964
rect 21053 23904 21117 23908
rect 5917 23420 5981 23424
rect 5917 23364 5921 23420
rect 5921 23364 5977 23420
rect 5977 23364 5981 23420
rect 5917 23360 5981 23364
rect 5997 23420 6061 23424
rect 5997 23364 6001 23420
rect 6001 23364 6057 23420
rect 6057 23364 6061 23420
rect 5997 23360 6061 23364
rect 6077 23420 6141 23424
rect 6077 23364 6081 23420
rect 6081 23364 6137 23420
rect 6137 23364 6141 23420
rect 6077 23360 6141 23364
rect 6157 23420 6221 23424
rect 6157 23364 6161 23420
rect 6161 23364 6217 23420
rect 6217 23364 6221 23420
rect 6157 23360 6221 23364
rect 15848 23420 15912 23424
rect 15848 23364 15852 23420
rect 15852 23364 15908 23420
rect 15908 23364 15912 23420
rect 15848 23360 15912 23364
rect 15928 23420 15992 23424
rect 15928 23364 15932 23420
rect 15932 23364 15988 23420
rect 15988 23364 15992 23420
rect 15928 23360 15992 23364
rect 16008 23420 16072 23424
rect 16008 23364 16012 23420
rect 16012 23364 16068 23420
rect 16068 23364 16072 23420
rect 16008 23360 16072 23364
rect 16088 23420 16152 23424
rect 16088 23364 16092 23420
rect 16092 23364 16148 23420
rect 16148 23364 16152 23420
rect 16088 23360 16152 23364
rect 25778 23420 25842 23424
rect 25778 23364 25782 23420
rect 25782 23364 25838 23420
rect 25838 23364 25842 23420
rect 25778 23360 25842 23364
rect 25858 23420 25922 23424
rect 25858 23364 25862 23420
rect 25862 23364 25918 23420
rect 25918 23364 25922 23420
rect 25858 23360 25922 23364
rect 25938 23420 26002 23424
rect 25938 23364 25942 23420
rect 25942 23364 25998 23420
rect 25998 23364 26002 23420
rect 25938 23360 26002 23364
rect 26018 23420 26082 23424
rect 26018 23364 26022 23420
rect 26022 23364 26078 23420
rect 26078 23364 26082 23420
rect 26018 23360 26082 23364
rect 17540 23156 17604 23220
rect 10882 22876 10946 22880
rect 10882 22820 10886 22876
rect 10886 22820 10942 22876
rect 10942 22820 10946 22876
rect 10882 22816 10946 22820
rect 10962 22876 11026 22880
rect 10962 22820 10966 22876
rect 10966 22820 11022 22876
rect 11022 22820 11026 22876
rect 10962 22816 11026 22820
rect 11042 22876 11106 22880
rect 11042 22820 11046 22876
rect 11046 22820 11102 22876
rect 11102 22820 11106 22876
rect 11042 22816 11106 22820
rect 11122 22876 11186 22880
rect 11122 22820 11126 22876
rect 11126 22820 11182 22876
rect 11182 22820 11186 22876
rect 11122 22816 11186 22820
rect 20813 22876 20877 22880
rect 20813 22820 20817 22876
rect 20817 22820 20873 22876
rect 20873 22820 20877 22876
rect 20813 22816 20877 22820
rect 20893 22876 20957 22880
rect 20893 22820 20897 22876
rect 20897 22820 20953 22876
rect 20953 22820 20957 22876
rect 20893 22816 20957 22820
rect 20973 22876 21037 22880
rect 20973 22820 20977 22876
rect 20977 22820 21033 22876
rect 21033 22820 21037 22876
rect 20973 22816 21037 22820
rect 21053 22876 21117 22880
rect 21053 22820 21057 22876
rect 21057 22820 21113 22876
rect 21113 22820 21117 22876
rect 21053 22816 21117 22820
rect 9444 22672 9508 22676
rect 9444 22616 9458 22672
rect 9458 22616 9508 22672
rect 9444 22612 9508 22616
rect 5917 22332 5981 22336
rect 5917 22276 5921 22332
rect 5921 22276 5977 22332
rect 5977 22276 5981 22332
rect 5917 22272 5981 22276
rect 5997 22332 6061 22336
rect 5997 22276 6001 22332
rect 6001 22276 6057 22332
rect 6057 22276 6061 22332
rect 5997 22272 6061 22276
rect 6077 22332 6141 22336
rect 6077 22276 6081 22332
rect 6081 22276 6137 22332
rect 6137 22276 6141 22332
rect 6077 22272 6141 22276
rect 6157 22332 6221 22336
rect 6157 22276 6161 22332
rect 6161 22276 6217 22332
rect 6217 22276 6221 22332
rect 6157 22272 6221 22276
rect 15848 22332 15912 22336
rect 15848 22276 15852 22332
rect 15852 22276 15908 22332
rect 15908 22276 15912 22332
rect 15848 22272 15912 22276
rect 15928 22332 15992 22336
rect 15928 22276 15932 22332
rect 15932 22276 15988 22332
rect 15988 22276 15992 22332
rect 15928 22272 15992 22276
rect 16008 22332 16072 22336
rect 16008 22276 16012 22332
rect 16012 22276 16068 22332
rect 16068 22276 16072 22332
rect 16008 22272 16072 22276
rect 16088 22332 16152 22336
rect 16088 22276 16092 22332
rect 16092 22276 16148 22332
rect 16148 22276 16152 22332
rect 16088 22272 16152 22276
rect 25778 22332 25842 22336
rect 25778 22276 25782 22332
rect 25782 22276 25838 22332
rect 25838 22276 25842 22332
rect 25778 22272 25842 22276
rect 25858 22332 25922 22336
rect 25858 22276 25862 22332
rect 25862 22276 25918 22332
rect 25918 22276 25922 22332
rect 25858 22272 25922 22276
rect 25938 22332 26002 22336
rect 25938 22276 25942 22332
rect 25942 22276 25998 22332
rect 25998 22276 26002 22332
rect 25938 22272 26002 22276
rect 26018 22332 26082 22336
rect 26018 22276 26022 22332
rect 26022 22276 26078 22332
rect 26078 22276 26082 22332
rect 26018 22272 26082 22276
rect 10882 21788 10946 21792
rect 10882 21732 10886 21788
rect 10886 21732 10942 21788
rect 10942 21732 10946 21788
rect 10882 21728 10946 21732
rect 10962 21788 11026 21792
rect 10962 21732 10966 21788
rect 10966 21732 11022 21788
rect 11022 21732 11026 21788
rect 10962 21728 11026 21732
rect 11042 21788 11106 21792
rect 11042 21732 11046 21788
rect 11046 21732 11102 21788
rect 11102 21732 11106 21788
rect 11042 21728 11106 21732
rect 11122 21788 11186 21792
rect 11122 21732 11126 21788
rect 11126 21732 11182 21788
rect 11182 21732 11186 21788
rect 11122 21728 11186 21732
rect 20813 21788 20877 21792
rect 20813 21732 20817 21788
rect 20817 21732 20873 21788
rect 20873 21732 20877 21788
rect 20813 21728 20877 21732
rect 20893 21788 20957 21792
rect 20893 21732 20897 21788
rect 20897 21732 20953 21788
rect 20953 21732 20957 21788
rect 20893 21728 20957 21732
rect 20973 21788 21037 21792
rect 20973 21732 20977 21788
rect 20977 21732 21033 21788
rect 21033 21732 21037 21788
rect 20973 21728 21037 21732
rect 21053 21788 21117 21792
rect 21053 21732 21057 21788
rect 21057 21732 21113 21788
rect 21113 21732 21117 21788
rect 21053 21728 21117 21732
rect 7972 21660 8036 21724
rect 5917 21244 5981 21248
rect 5917 21188 5921 21244
rect 5921 21188 5977 21244
rect 5977 21188 5981 21244
rect 5917 21184 5981 21188
rect 5997 21244 6061 21248
rect 5997 21188 6001 21244
rect 6001 21188 6057 21244
rect 6057 21188 6061 21244
rect 5997 21184 6061 21188
rect 6077 21244 6141 21248
rect 6077 21188 6081 21244
rect 6081 21188 6137 21244
rect 6137 21188 6141 21244
rect 6077 21184 6141 21188
rect 6157 21244 6221 21248
rect 6157 21188 6161 21244
rect 6161 21188 6217 21244
rect 6217 21188 6221 21244
rect 6157 21184 6221 21188
rect 15848 21244 15912 21248
rect 15848 21188 15852 21244
rect 15852 21188 15908 21244
rect 15908 21188 15912 21244
rect 15848 21184 15912 21188
rect 15928 21244 15992 21248
rect 15928 21188 15932 21244
rect 15932 21188 15988 21244
rect 15988 21188 15992 21244
rect 15928 21184 15992 21188
rect 16008 21244 16072 21248
rect 16008 21188 16012 21244
rect 16012 21188 16068 21244
rect 16068 21188 16072 21244
rect 16008 21184 16072 21188
rect 16088 21244 16152 21248
rect 16088 21188 16092 21244
rect 16092 21188 16148 21244
rect 16148 21188 16152 21244
rect 16088 21184 16152 21188
rect 25778 21244 25842 21248
rect 25778 21188 25782 21244
rect 25782 21188 25838 21244
rect 25838 21188 25842 21244
rect 25778 21184 25842 21188
rect 25858 21244 25922 21248
rect 25858 21188 25862 21244
rect 25862 21188 25918 21244
rect 25918 21188 25922 21244
rect 25858 21184 25922 21188
rect 25938 21244 26002 21248
rect 25938 21188 25942 21244
rect 25942 21188 25998 21244
rect 25998 21188 26002 21244
rect 25938 21184 26002 21188
rect 26018 21244 26082 21248
rect 26018 21188 26022 21244
rect 26022 21188 26078 21244
rect 26078 21188 26082 21244
rect 26018 21184 26082 21188
rect 9444 21176 9508 21180
rect 9444 21120 9458 21176
rect 9458 21120 9508 21176
rect 9444 21116 9508 21120
rect 10882 20700 10946 20704
rect 10882 20644 10886 20700
rect 10886 20644 10942 20700
rect 10942 20644 10946 20700
rect 10882 20640 10946 20644
rect 10962 20700 11026 20704
rect 10962 20644 10966 20700
rect 10966 20644 11022 20700
rect 11022 20644 11026 20700
rect 10962 20640 11026 20644
rect 11042 20700 11106 20704
rect 11042 20644 11046 20700
rect 11046 20644 11102 20700
rect 11102 20644 11106 20700
rect 11042 20640 11106 20644
rect 11122 20700 11186 20704
rect 11122 20644 11126 20700
rect 11126 20644 11182 20700
rect 11182 20644 11186 20700
rect 11122 20640 11186 20644
rect 20813 20700 20877 20704
rect 20813 20644 20817 20700
rect 20817 20644 20873 20700
rect 20873 20644 20877 20700
rect 20813 20640 20877 20644
rect 20893 20700 20957 20704
rect 20893 20644 20897 20700
rect 20897 20644 20953 20700
rect 20953 20644 20957 20700
rect 20893 20640 20957 20644
rect 20973 20700 21037 20704
rect 20973 20644 20977 20700
rect 20977 20644 21033 20700
rect 21033 20644 21037 20700
rect 20973 20640 21037 20644
rect 21053 20700 21117 20704
rect 21053 20644 21057 20700
rect 21057 20644 21113 20700
rect 21113 20644 21117 20700
rect 21053 20640 21117 20644
rect 5917 20156 5981 20160
rect 5917 20100 5921 20156
rect 5921 20100 5977 20156
rect 5977 20100 5981 20156
rect 5917 20096 5981 20100
rect 5997 20156 6061 20160
rect 5997 20100 6001 20156
rect 6001 20100 6057 20156
rect 6057 20100 6061 20156
rect 5997 20096 6061 20100
rect 6077 20156 6141 20160
rect 6077 20100 6081 20156
rect 6081 20100 6137 20156
rect 6137 20100 6141 20156
rect 6077 20096 6141 20100
rect 6157 20156 6221 20160
rect 6157 20100 6161 20156
rect 6161 20100 6217 20156
rect 6217 20100 6221 20156
rect 6157 20096 6221 20100
rect 15848 20156 15912 20160
rect 15848 20100 15852 20156
rect 15852 20100 15908 20156
rect 15908 20100 15912 20156
rect 15848 20096 15912 20100
rect 15928 20156 15992 20160
rect 15928 20100 15932 20156
rect 15932 20100 15988 20156
rect 15988 20100 15992 20156
rect 15928 20096 15992 20100
rect 16008 20156 16072 20160
rect 16008 20100 16012 20156
rect 16012 20100 16068 20156
rect 16068 20100 16072 20156
rect 16008 20096 16072 20100
rect 16088 20156 16152 20160
rect 16088 20100 16092 20156
rect 16092 20100 16148 20156
rect 16148 20100 16152 20156
rect 16088 20096 16152 20100
rect 25778 20156 25842 20160
rect 25778 20100 25782 20156
rect 25782 20100 25838 20156
rect 25838 20100 25842 20156
rect 25778 20096 25842 20100
rect 25858 20156 25922 20160
rect 25858 20100 25862 20156
rect 25862 20100 25918 20156
rect 25918 20100 25922 20156
rect 25858 20096 25922 20100
rect 25938 20156 26002 20160
rect 25938 20100 25942 20156
rect 25942 20100 25998 20156
rect 25998 20100 26002 20156
rect 25938 20096 26002 20100
rect 26018 20156 26082 20160
rect 26018 20100 26022 20156
rect 26022 20100 26078 20156
rect 26078 20100 26082 20156
rect 26018 20096 26082 20100
rect 10882 19612 10946 19616
rect 10882 19556 10886 19612
rect 10886 19556 10942 19612
rect 10942 19556 10946 19612
rect 10882 19552 10946 19556
rect 10962 19612 11026 19616
rect 10962 19556 10966 19612
rect 10966 19556 11022 19612
rect 11022 19556 11026 19612
rect 10962 19552 11026 19556
rect 11042 19612 11106 19616
rect 11042 19556 11046 19612
rect 11046 19556 11102 19612
rect 11102 19556 11106 19612
rect 11042 19552 11106 19556
rect 11122 19612 11186 19616
rect 11122 19556 11126 19612
rect 11126 19556 11182 19612
rect 11182 19556 11186 19612
rect 11122 19552 11186 19556
rect 20813 19612 20877 19616
rect 20813 19556 20817 19612
rect 20817 19556 20873 19612
rect 20873 19556 20877 19612
rect 20813 19552 20877 19556
rect 20893 19612 20957 19616
rect 20893 19556 20897 19612
rect 20897 19556 20953 19612
rect 20953 19556 20957 19612
rect 20893 19552 20957 19556
rect 20973 19612 21037 19616
rect 20973 19556 20977 19612
rect 20977 19556 21033 19612
rect 21033 19556 21037 19612
rect 20973 19552 21037 19556
rect 21053 19612 21117 19616
rect 21053 19556 21057 19612
rect 21057 19556 21113 19612
rect 21113 19556 21117 19612
rect 21053 19552 21117 19556
rect 11284 19076 11348 19140
rect 5917 19068 5981 19072
rect 5917 19012 5921 19068
rect 5921 19012 5977 19068
rect 5977 19012 5981 19068
rect 5917 19008 5981 19012
rect 5997 19068 6061 19072
rect 5997 19012 6001 19068
rect 6001 19012 6057 19068
rect 6057 19012 6061 19068
rect 5997 19008 6061 19012
rect 6077 19068 6141 19072
rect 6077 19012 6081 19068
rect 6081 19012 6137 19068
rect 6137 19012 6141 19068
rect 6077 19008 6141 19012
rect 6157 19068 6221 19072
rect 6157 19012 6161 19068
rect 6161 19012 6217 19068
rect 6217 19012 6221 19068
rect 6157 19008 6221 19012
rect 15848 19068 15912 19072
rect 15848 19012 15852 19068
rect 15852 19012 15908 19068
rect 15908 19012 15912 19068
rect 15848 19008 15912 19012
rect 15928 19068 15992 19072
rect 15928 19012 15932 19068
rect 15932 19012 15988 19068
rect 15988 19012 15992 19068
rect 15928 19008 15992 19012
rect 16008 19068 16072 19072
rect 16008 19012 16012 19068
rect 16012 19012 16068 19068
rect 16068 19012 16072 19068
rect 16008 19008 16072 19012
rect 16088 19068 16152 19072
rect 16088 19012 16092 19068
rect 16092 19012 16148 19068
rect 16148 19012 16152 19068
rect 16088 19008 16152 19012
rect 25778 19068 25842 19072
rect 25778 19012 25782 19068
rect 25782 19012 25838 19068
rect 25838 19012 25842 19068
rect 25778 19008 25842 19012
rect 25858 19068 25922 19072
rect 25858 19012 25862 19068
rect 25862 19012 25918 19068
rect 25918 19012 25922 19068
rect 25858 19008 25922 19012
rect 25938 19068 26002 19072
rect 25938 19012 25942 19068
rect 25942 19012 25998 19068
rect 25998 19012 26002 19068
rect 25938 19008 26002 19012
rect 26018 19068 26082 19072
rect 26018 19012 26022 19068
rect 26022 19012 26078 19068
rect 26078 19012 26082 19068
rect 26018 19008 26082 19012
rect 10882 18524 10946 18528
rect 10882 18468 10886 18524
rect 10886 18468 10942 18524
rect 10942 18468 10946 18524
rect 10882 18464 10946 18468
rect 10962 18524 11026 18528
rect 10962 18468 10966 18524
rect 10966 18468 11022 18524
rect 11022 18468 11026 18524
rect 10962 18464 11026 18468
rect 11042 18524 11106 18528
rect 11042 18468 11046 18524
rect 11046 18468 11102 18524
rect 11102 18468 11106 18524
rect 11042 18464 11106 18468
rect 11122 18524 11186 18528
rect 11122 18468 11126 18524
rect 11126 18468 11182 18524
rect 11182 18468 11186 18524
rect 11122 18464 11186 18468
rect 20813 18524 20877 18528
rect 20813 18468 20817 18524
rect 20817 18468 20873 18524
rect 20873 18468 20877 18524
rect 20813 18464 20877 18468
rect 20893 18524 20957 18528
rect 20893 18468 20897 18524
rect 20897 18468 20953 18524
rect 20953 18468 20957 18524
rect 20893 18464 20957 18468
rect 20973 18524 21037 18528
rect 20973 18468 20977 18524
rect 20977 18468 21033 18524
rect 21033 18468 21037 18524
rect 20973 18464 21037 18468
rect 21053 18524 21117 18528
rect 21053 18468 21057 18524
rect 21057 18468 21113 18524
rect 21113 18468 21117 18524
rect 21053 18464 21117 18468
rect 5917 17980 5981 17984
rect 5917 17924 5921 17980
rect 5921 17924 5977 17980
rect 5977 17924 5981 17980
rect 5917 17920 5981 17924
rect 5997 17980 6061 17984
rect 5997 17924 6001 17980
rect 6001 17924 6057 17980
rect 6057 17924 6061 17980
rect 5997 17920 6061 17924
rect 6077 17980 6141 17984
rect 6077 17924 6081 17980
rect 6081 17924 6137 17980
rect 6137 17924 6141 17980
rect 6077 17920 6141 17924
rect 6157 17980 6221 17984
rect 6157 17924 6161 17980
rect 6161 17924 6217 17980
rect 6217 17924 6221 17980
rect 6157 17920 6221 17924
rect 15848 17980 15912 17984
rect 15848 17924 15852 17980
rect 15852 17924 15908 17980
rect 15908 17924 15912 17980
rect 15848 17920 15912 17924
rect 15928 17980 15992 17984
rect 15928 17924 15932 17980
rect 15932 17924 15988 17980
rect 15988 17924 15992 17980
rect 15928 17920 15992 17924
rect 16008 17980 16072 17984
rect 16008 17924 16012 17980
rect 16012 17924 16068 17980
rect 16068 17924 16072 17980
rect 16008 17920 16072 17924
rect 16088 17980 16152 17984
rect 16088 17924 16092 17980
rect 16092 17924 16148 17980
rect 16148 17924 16152 17980
rect 16088 17920 16152 17924
rect 25778 17980 25842 17984
rect 25778 17924 25782 17980
rect 25782 17924 25838 17980
rect 25838 17924 25842 17980
rect 25778 17920 25842 17924
rect 25858 17980 25922 17984
rect 25858 17924 25862 17980
rect 25862 17924 25918 17980
rect 25918 17924 25922 17980
rect 25858 17920 25922 17924
rect 25938 17980 26002 17984
rect 25938 17924 25942 17980
rect 25942 17924 25998 17980
rect 25998 17924 26002 17980
rect 25938 17920 26002 17924
rect 26018 17980 26082 17984
rect 26018 17924 26022 17980
rect 26022 17924 26078 17980
rect 26078 17924 26082 17980
rect 26018 17920 26082 17924
rect 10882 17436 10946 17440
rect 10882 17380 10886 17436
rect 10886 17380 10942 17436
rect 10942 17380 10946 17436
rect 10882 17376 10946 17380
rect 10962 17436 11026 17440
rect 10962 17380 10966 17436
rect 10966 17380 11022 17436
rect 11022 17380 11026 17436
rect 10962 17376 11026 17380
rect 11042 17436 11106 17440
rect 11042 17380 11046 17436
rect 11046 17380 11102 17436
rect 11102 17380 11106 17436
rect 11042 17376 11106 17380
rect 11122 17436 11186 17440
rect 11122 17380 11126 17436
rect 11126 17380 11182 17436
rect 11182 17380 11186 17436
rect 11122 17376 11186 17380
rect 20813 17436 20877 17440
rect 20813 17380 20817 17436
rect 20817 17380 20873 17436
rect 20873 17380 20877 17436
rect 20813 17376 20877 17380
rect 20893 17436 20957 17440
rect 20893 17380 20897 17436
rect 20897 17380 20953 17436
rect 20953 17380 20957 17436
rect 20893 17376 20957 17380
rect 20973 17436 21037 17440
rect 20973 17380 20977 17436
rect 20977 17380 21033 17436
rect 21033 17380 21037 17436
rect 20973 17376 21037 17380
rect 21053 17436 21117 17440
rect 21053 17380 21057 17436
rect 21057 17380 21113 17436
rect 21113 17380 21117 17436
rect 21053 17376 21117 17380
rect 10180 17368 10244 17372
rect 10180 17312 10194 17368
rect 10194 17312 10244 17368
rect 10180 17308 10244 17312
rect 5917 16892 5981 16896
rect 5917 16836 5921 16892
rect 5921 16836 5977 16892
rect 5977 16836 5981 16892
rect 5917 16832 5981 16836
rect 5997 16892 6061 16896
rect 5997 16836 6001 16892
rect 6001 16836 6057 16892
rect 6057 16836 6061 16892
rect 5997 16832 6061 16836
rect 6077 16892 6141 16896
rect 6077 16836 6081 16892
rect 6081 16836 6137 16892
rect 6137 16836 6141 16892
rect 6077 16832 6141 16836
rect 6157 16892 6221 16896
rect 6157 16836 6161 16892
rect 6161 16836 6217 16892
rect 6217 16836 6221 16892
rect 6157 16832 6221 16836
rect 15848 16892 15912 16896
rect 15848 16836 15852 16892
rect 15852 16836 15908 16892
rect 15908 16836 15912 16892
rect 15848 16832 15912 16836
rect 15928 16892 15992 16896
rect 15928 16836 15932 16892
rect 15932 16836 15988 16892
rect 15988 16836 15992 16892
rect 15928 16832 15992 16836
rect 16008 16892 16072 16896
rect 16008 16836 16012 16892
rect 16012 16836 16068 16892
rect 16068 16836 16072 16892
rect 16008 16832 16072 16836
rect 16088 16892 16152 16896
rect 16088 16836 16092 16892
rect 16092 16836 16148 16892
rect 16148 16836 16152 16892
rect 16088 16832 16152 16836
rect 25778 16892 25842 16896
rect 25778 16836 25782 16892
rect 25782 16836 25838 16892
rect 25838 16836 25842 16892
rect 25778 16832 25842 16836
rect 25858 16892 25922 16896
rect 25858 16836 25862 16892
rect 25862 16836 25918 16892
rect 25918 16836 25922 16892
rect 25858 16832 25922 16836
rect 25938 16892 26002 16896
rect 25938 16836 25942 16892
rect 25942 16836 25998 16892
rect 25998 16836 26002 16892
rect 25938 16832 26002 16836
rect 26018 16892 26082 16896
rect 26018 16836 26022 16892
rect 26022 16836 26078 16892
rect 26078 16836 26082 16892
rect 26018 16832 26082 16836
rect 10882 16348 10946 16352
rect 10882 16292 10886 16348
rect 10886 16292 10942 16348
rect 10942 16292 10946 16348
rect 10882 16288 10946 16292
rect 10962 16348 11026 16352
rect 10962 16292 10966 16348
rect 10966 16292 11022 16348
rect 11022 16292 11026 16348
rect 10962 16288 11026 16292
rect 11042 16348 11106 16352
rect 11042 16292 11046 16348
rect 11046 16292 11102 16348
rect 11102 16292 11106 16348
rect 11042 16288 11106 16292
rect 11122 16348 11186 16352
rect 11122 16292 11126 16348
rect 11126 16292 11182 16348
rect 11182 16292 11186 16348
rect 11122 16288 11186 16292
rect 20813 16348 20877 16352
rect 20813 16292 20817 16348
rect 20817 16292 20873 16348
rect 20873 16292 20877 16348
rect 20813 16288 20877 16292
rect 20893 16348 20957 16352
rect 20893 16292 20897 16348
rect 20897 16292 20953 16348
rect 20953 16292 20957 16348
rect 20893 16288 20957 16292
rect 20973 16348 21037 16352
rect 20973 16292 20977 16348
rect 20977 16292 21033 16348
rect 21033 16292 21037 16348
rect 20973 16288 21037 16292
rect 21053 16348 21117 16352
rect 21053 16292 21057 16348
rect 21057 16292 21113 16348
rect 21113 16292 21117 16348
rect 21053 16288 21117 16292
rect 5917 15804 5981 15808
rect 5917 15748 5921 15804
rect 5921 15748 5977 15804
rect 5977 15748 5981 15804
rect 5917 15744 5981 15748
rect 5997 15804 6061 15808
rect 5997 15748 6001 15804
rect 6001 15748 6057 15804
rect 6057 15748 6061 15804
rect 5997 15744 6061 15748
rect 6077 15804 6141 15808
rect 6077 15748 6081 15804
rect 6081 15748 6137 15804
rect 6137 15748 6141 15804
rect 6077 15744 6141 15748
rect 6157 15804 6221 15808
rect 6157 15748 6161 15804
rect 6161 15748 6217 15804
rect 6217 15748 6221 15804
rect 6157 15744 6221 15748
rect 15848 15804 15912 15808
rect 15848 15748 15852 15804
rect 15852 15748 15908 15804
rect 15908 15748 15912 15804
rect 15848 15744 15912 15748
rect 15928 15804 15992 15808
rect 15928 15748 15932 15804
rect 15932 15748 15988 15804
rect 15988 15748 15992 15804
rect 15928 15744 15992 15748
rect 16008 15804 16072 15808
rect 16008 15748 16012 15804
rect 16012 15748 16068 15804
rect 16068 15748 16072 15804
rect 16008 15744 16072 15748
rect 16088 15804 16152 15808
rect 16088 15748 16092 15804
rect 16092 15748 16148 15804
rect 16148 15748 16152 15804
rect 16088 15744 16152 15748
rect 25778 15804 25842 15808
rect 25778 15748 25782 15804
rect 25782 15748 25838 15804
rect 25838 15748 25842 15804
rect 25778 15744 25842 15748
rect 25858 15804 25922 15808
rect 25858 15748 25862 15804
rect 25862 15748 25918 15804
rect 25918 15748 25922 15804
rect 25858 15744 25922 15748
rect 25938 15804 26002 15808
rect 25938 15748 25942 15804
rect 25942 15748 25998 15804
rect 25998 15748 26002 15804
rect 25938 15744 26002 15748
rect 26018 15804 26082 15808
rect 26018 15748 26022 15804
rect 26022 15748 26078 15804
rect 26078 15748 26082 15804
rect 26018 15744 26082 15748
rect 9076 15464 9140 15468
rect 9076 15408 9126 15464
rect 9126 15408 9140 15464
rect 9076 15404 9140 15408
rect 10882 15260 10946 15264
rect 10882 15204 10886 15260
rect 10886 15204 10942 15260
rect 10942 15204 10946 15260
rect 10882 15200 10946 15204
rect 10962 15260 11026 15264
rect 10962 15204 10966 15260
rect 10966 15204 11022 15260
rect 11022 15204 11026 15260
rect 10962 15200 11026 15204
rect 11042 15260 11106 15264
rect 11042 15204 11046 15260
rect 11046 15204 11102 15260
rect 11102 15204 11106 15260
rect 11042 15200 11106 15204
rect 11122 15260 11186 15264
rect 11122 15204 11126 15260
rect 11126 15204 11182 15260
rect 11182 15204 11186 15260
rect 11122 15200 11186 15204
rect 20813 15260 20877 15264
rect 20813 15204 20817 15260
rect 20817 15204 20873 15260
rect 20873 15204 20877 15260
rect 20813 15200 20877 15204
rect 20893 15260 20957 15264
rect 20893 15204 20897 15260
rect 20897 15204 20953 15260
rect 20953 15204 20957 15260
rect 20893 15200 20957 15204
rect 20973 15260 21037 15264
rect 20973 15204 20977 15260
rect 20977 15204 21033 15260
rect 21033 15204 21037 15260
rect 20973 15200 21037 15204
rect 21053 15260 21117 15264
rect 21053 15204 21057 15260
rect 21057 15204 21113 15260
rect 21113 15204 21117 15260
rect 21053 15200 21117 15204
rect 5917 14716 5981 14720
rect 5917 14660 5921 14716
rect 5921 14660 5977 14716
rect 5977 14660 5981 14716
rect 5917 14656 5981 14660
rect 5997 14716 6061 14720
rect 5997 14660 6001 14716
rect 6001 14660 6057 14716
rect 6057 14660 6061 14716
rect 5997 14656 6061 14660
rect 6077 14716 6141 14720
rect 6077 14660 6081 14716
rect 6081 14660 6137 14716
rect 6137 14660 6141 14716
rect 6077 14656 6141 14660
rect 6157 14716 6221 14720
rect 6157 14660 6161 14716
rect 6161 14660 6217 14716
rect 6217 14660 6221 14716
rect 6157 14656 6221 14660
rect 15848 14716 15912 14720
rect 15848 14660 15852 14716
rect 15852 14660 15908 14716
rect 15908 14660 15912 14716
rect 15848 14656 15912 14660
rect 15928 14716 15992 14720
rect 15928 14660 15932 14716
rect 15932 14660 15988 14716
rect 15988 14660 15992 14716
rect 15928 14656 15992 14660
rect 16008 14716 16072 14720
rect 16008 14660 16012 14716
rect 16012 14660 16068 14716
rect 16068 14660 16072 14716
rect 16008 14656 16072 14660
rect 16088 14716 16152 14720
rect 16088 14660 16092 14716
rect 16092 14660 16148 14716
rect 16148 14660 16152 14716
rect 16088 14656 16152 14660
rect 25778 14716 25842 14720
rect 25778 14660 25782 14716
rect 25782 14660 25838 14716
rect 25838 14660 25842 14716
rect 25778 14656 25842 14660
rect 25858 14716 25922 14720
rect 25858 14660 25862 14716
rect 25862 14660 25918 14716
rect 25918 14660 25922 14716
rect 25858 14656 25922 14660
rect 25938 14716 26002 14720
rect 25938 14660 25942 14716
rect 25942 14660 25998 14716
rect 25998 14660 26002 14716
rect 25938 14656 26002 14660
rect 26018 14716 26082 14720
rect 26018 14660 26022 14716
rect 26022 14660 26078 14716
rect 26078 14660 26082 14716
rect 26018 14656 26082 14660
rect 10882 14172 10946 14176
rect 10882 14116 10886 14172
rect 10886 14116 10942 14172
rect 10942 14116 10946 14172
rect 10882 14112 10946 14116
rect 10962 14172 11026 14176
rect 10962 14116 10966 14172
rect 10966 14116 11022 14172
rect 11022 14116 11026 14172
rect 10962 14112 11026 14116
rect 11042 14172 11106 14176
rect 11042 14116 11046 14172
rect 11046 14116 11102 14172
rect 11102 14116 11106 14172
rect 11042 14112 11106 14116
rect 11122 14172 11186 14176
rect 11122 14116 11126 14172
rect 11126 14116 11182 14172
rect 11182 14116 11186 14172
rect 11122 14112 11186 14116
rect 20813 14172 20877 14176
rect 20813 14116 20817 14172
rect 20817 14116 20873 14172
rect 20873 14116 20877 14172
rect 20813 14112 20877 14116
rect 20893 14172 20957 14176
rect 20893 14116 20897 14172
rect 20897 14116 20953 14172
rect 20953 14116 20957 14172
rect 20893 14112 20957 14116
rect 20973 14172 21037 14176
rect 20973 14116 20977 14172
rect 20977 14116 21033 14172
rect 21033 14116 21037 14172
rect 20973 14112 21037 14116
rect 21053 14172 21117 14176
rect 21053 14116 21057 14172
rect 21057 14116 21113 14172
rect 21113 14116 21117 14172
rect 21053 14112 21117 14116
rect 5917 13628 5981 13632
rect 5917 13572 5921 13628
rect 5921 13572 5977 13628
rect 5977 13572 5981 13628
rect 5917 13568 5981 13572
rect 5997 13628 6061 13632
rect 5997 13572 6001 13628
rect 6001 13572 6057 13628
rect 6057 13572 6061 13628
rect 5997 13568 6061 13572
rect 6077 13628 6141 13632
rect 6077 13572 6081 13628
rect 6081 13572 6137 13628
rect 6137 13572 6141 13628
rect 6077 13568 6141 13572
rect 6157 13628 6221 13632
rect 6157 13572 6161 13628
rect 6161 13572 6217 13628
rect 6217 13572 6221 13628
rect 6157 13568 6221 13572
rect 15848 13628 15912 13632
rect 15848 13572 15852 13628
rect 15852 13572 15908 13628
rect 15908 13572 15912 13628
rect 15848 13568 15912 13572
rect 15928 13628 15992 13632
rect 15928 13572 15932 13628
rect 15932 13572 15988 13628
rect 15988 13572 15992 13628
rect 15928 13568 15992 13572
rect 16008 13628 16072 13632
rect 16008 13572 16012 13628
rect 16012 13572 16068 13628
rect 16068 13572 16072 13628
rect 16008 13568 16072 13572
rect 16088 13628 16152 13632
rect 16088 13572 16092 13628
rect 16092 13572 16148 13628
rect 16148 13572 16152 13628
rect 16088 13568 16152 13572
rect 25778 13628 25842 13632
rect 25778 13572 25782 13628
rect 25782 13572 25838 13628
rect 25838 13572 25842 13628
rect 25778 13568 25842 13572
rect 25858 13628 25922 13632
rect 25858 13572 25862 13628
rect 25862 13572 25918 13628
rect 25918 13572 25922 13628
rect 25858 13568 25922 13572
rect 25938 13628 26002 13632
rect 25938 13572 25942 13628
rect 25942 13572 25998 13628
rect 25998 13572 26002 13628
rect 25938 13568 26002 13572
rect 26018 13628 26082 13632
rect 26018 13572 26022 13628
rect 26022 13572 26078 13628
rect 26078 13572 26082 13628
rect 26018 13568 26082 13572
rect 10882 13084 10946 13088
rect 10882 13028 10886 13084
rect 10886 13028 10942 13084
rect 10942 13028 10946 13084
rect 10882 13024 10946 13028
rect 10962 13084 11026 13088
rect 10962 13028 10966 13084
rect 10966 13028 11022 13084
rect 11022 13028 11026 13084
rect 10962 13024 11026 13028
rect 11042 13084 11106 13088
rect 11042 13028 11046 13084
rect 11046 13028 11102 13084
rect 11102 13028 11106 13084
rect 11042 13024 11106 13028
rect 11122 13084 11186 13088
rect 11122 13028 11126 13084
rect 11126 13028 11182 13084
rect 11182 13028 11186 13084
rect 11122 13024 11186 13028
rect 20813 13084 20877 13088
rect 20813 13028 20817 13084
rect 20817 13028 20873 13084
rect 20873 13028 20877 13084
rect 20813 13024 20877 13028
rect 20893 13084 20957 13088
rect 20893 13028 20897 13084
rect 20897 13028 20953 13084
rect 20953 13028 20957 13084
rect 20893 13024 20957 13028
rect 20973 13084 21037 13088
rect 20973 13028 20977 13084
rect 20977 13028 21033 13084
rect 21033 13028 21037 13084
rect 20973 13024 21037 13028
rect 21053 13084 21117 13088
rect 21053 13028 21057 13084
rect 21057 13028 21113 13084
rect 21113 13028 21117 13084
rect 21053 13024 21117 13028
rect 5917 12540 5981 12544
rect 5917 12484 5921 12540
rect 5921 12484 5977 12540
rect 5977 12484 5981 12540
rect 5917 12480 5981 12484
rect 5997 12540 6061 12544
rect 5997 12484 6001 12540
rect 6001 12484 6057 12540
rect 6057 12484 6061 12540
rect 5997 12480 6061 12484
rect 6077 12540 6141 12544
rect 6077 12484 6081 12540
rect 6081 12484 6137 12540
rect 6137 12484 6141 12540
rect 6077 12480 6141 12484
rect 6157 12540 6221 12544
rect 6157 12484 6161 12540
rect 6161 12484 6217 12540
rect 6217 12484 6221 12540
rect 6157 12480 6221 12484
rect 15848 12540 15912 12544
rect 15848 12484 15852 12540
rect 15852 12484 15908 12540
rect 15908 12484 15912 12540
rect 15848 12480 15912 12484
rect 15928 12540 15992 12544
rect 15928 12484 15932 12540
rect 15932 12484 15988 12540
rect 15988 12484 15992 12540
rect 15928 12480 15992 12484
rect 16008 12540 16072 12544
rect 16008 12484 16012 12540
rect 16012 12484 16068 12540
rect 16068 12484 16072 12540
rect 16008 12480 16072 12484
rect 16088 12540 16152 12544
rect 16088 12484 16092 12540
rect 16092 12484 16148 12540
rect 16148 12484 16152 12540
rect 16088 12480 16152 12484
rect 25778 12540 25842 12544
rect 25778 12484 25782 12540
rect 25782 12484 25838 12540
rect 25838 12484 25842 12540
rect 25778 12480 25842 12484
rect 25858 12540 25922 12544
rect 25858 12484 25862 12540
rect 25862 12484 25918 12540
rect 25918 12484 25922 12540
rect 25858 12480 25922 12484
rect 25938 12540 26002 12544
rect 25938 12484 25942 12540
rect 25942 12484 25998 12540
rect 25998 12484 26002 12540
rect 25938 12480 26002 12484
rect 26018 12540 26082 12544
rect 26018 12484 26022 12540
rect 26022 12484 26078 12540
rect 26078 12484 26082 12540
rect 26018 12480 26082 12484
rect 5917 11452 5981 11456
rect 5917 11396 5921 11452
rect 5921 11396 5977 11452
rect 5977 11396 5981 11452
rect 5917 11392 5981 11396
rect 5997 11452 6061 11456
rect 5997 11396 6001 11452
rect 6001 11396 6057 11452
rect 6057 11396 6061 11452
rect 5997 11392 6061 11396
rect 6077 11452 6141 11456
rect 6077 11396 6081 11452
rect 6081 11396 6137 11452
rect 6137 11396 6141 11452
rect 6077 11392 6141 11396
rect 6157 11452 6221 11456
rect 6157 11396 6161 11452
rect 6161 11396 6217 11452
rect 6217 11396 6221 11452
rect 6157 11392 6221 11396
rect 10180 12004 10244 12068
rect 10882 11996 10946 12000
rect 10882 11940 10886 11996
rect 10886 11940 10942 11996
rect 10942 11940 10946 11996
rect 10882 11936 10946 11940
rect 10962 11996 11026 12000
rect 10962 11940 10966 11996
rect 10966 11940 11022 11996
rect 11022 11940 11026 11996
rect 10962 11936 11026 11940
rect 11042 11996 11106 12000
rect 11042 11940 11046 11996
rect 11046 11940 11102 11996
rect 11102 11940 11106 11996
rect 11042 11936 11106 11940
rect 11122 11996 11186 12000
rect 11122 11940 11126 11996
rect 11126 11940 11182 11996
rect 11182 11940 11186 11996
rect 11122 11936 11186 11940
rect 20813 11996 20877 12000
rect 20813 11940 20817 11996
rect 20817 11940 20873 11996
rect 20873 11940 20877 11996
rect 20813 11936 20877 11940
rect 20893 11996 20957 12000
rect 20893 11940 20897 11996
rect 20897 11940 20953 11996
rect 20953 11940 20957 11996
rect 20893 11936 20957 11940
rect 20973 11996 21037 12000
rect 20973 11940 20977 11996
rect 20977 11940 21033 11996
rect 21033 11940 21037 11996
rect 20973 11936 21037 11940
rect 21053 11996 21117 12000
rect 21053 11940 21057 11996
rect 21057 11940 21113 11996
rect 21113 11940 21117 11996
rect 21053 11936 21117 11940
rect 15848 11452 15912 11456
rect 15848 11396 15852 11452
rect 15852 11396 15908 11452
rect 15908 11396 15912 11452
rect 15848 11392 15912 11396
rect 15928 11452 15992 11456
rect 15928 11396 15932 11452
rect 15932 11396 15988 11452
rect 15988 11396 15992 11452
rect 15928 11392 15992 11396
rect 16008 11452 16072 11456
rect 16008 11396 16012 11452
rect 16012 11396 16068 11452
rect 16068 11396 16072 11452
rect 16008 11392 16072 11396
rect 16088 11452 16152 11456
rect 16088 11396 16092 11452
rect 16092 11396 16148 11452
rect 16148 11396 16152 11452
rect 16088 11392 16152 11396
rect 25778 11452 25842 11456
rect 25778 11396 25782 11452
rect 25782 11396 25838 11452
rect 25838 11396 25842 11452
rect 25778 11392 25842 11396
rect 25858 11452 25922 11456
rect 25858 11396 25862 11452
rect 25862 11396 25918 11452
rect 25918 11396 25922 11452
rect 25858 11392 25922 11396
rect 25938 11452 26002 11456
rect 25938 11396 25942 11452
rect 25942 11396 25998 11452
rect 25998 11396 26002 11452
rect 25938 11392 26002 11396
rect 26018 11452 26082 11456
rect 26018 11396 26022 11452
rect 26022 11396 26078 11452
rect 26078 11396 26082 11452
rect 26018 11392 26082 11396
rect 9076 11248 9140 11252
rect 9076 11192 9090 11248
rect 9090 11192 9140 11248
rect 9076 11188 9140 11192
rect 10882 10908 10946 10912
rect 10882 10852 10886 10908
rect 10886 10852 10942 10908
rect 10942 10852 10946 10908
rect 10882 10848 10946 10852
rect 10962 10908 11026 10912
rect 10962 10852 10966 10908
rect 10966 10852 11022 10908
rect 11022 10852 11026 10908
rect 10962 10848 11026 10852
rect 11042 10908 11106 10912
rect 11042 10852 11046 10908
rect 11046 10852 11102 10908
rect 11102 10852 11106 10908
rect 11042 10848 11106 10852
rect 11122 10908 11186 10912
rect 11122 10852 11126 10908
rect 11126 10852 11182 10908
rect 11182 10852 11186 10908
rect 11122 10848 11186 10852
rect 20813 10908 20877 10912
rect 20813 10852 20817 10908
rect 20817 10852 20873 10908
rect 20873 10852 20877 10908
rect 20813 10848 20877 10852
rect 20893 10908 20957 10912
rect 20893 10852 20897 10908
rect 20897 10852 20953 10908
rect 20953 10852 20957 10908
rect 20893 10848 20957 10852
rect 20973 10908 21037 10912
rect 20973 10852 20977 10908
rect 20977 10852 21033 10908
rect 21033 10852 21037 10908
rect 20973 10848 21037 10852
rect 21053 10908 21117 10912
rect 21053 10852 21057 10908
rect 21057 10852 21113 10908
rect 21113 10852 21117 10908
rect 21053 10848 21117 10852
rect 5917 10364 5981 10368
rect 5917 10308 5921 10364
rect 5921 10308 5977 10364
rect 5977 10308 5981 10364
rect 5917 10304 5981 10308
rect 5997 10364 6061 10368
rect 5997 10308 6001 10364
rect 6001 10308 6057 10364
rect 6057 10308 6061 10364
rect 5997 10304 6061 10308
rect 6077 10364 6141 10368
rect 6077 10308 6081 10364
rect 6081 10308 6137 10364
rect 6137 10308 6141 10364
rect 6077 10304 6141 10308
rect 6157 10364 6221 10368
rect 6157 10308 6161 10364
rect 6161 10308 6217 10364
rect 6217 10308 6221 10364
rect 6157 10304 6221 10308
rect 15848 10364 15912 10368
rect 15848 10308 15852 10364
rect 15852 10308 15908 10364
rect 15908 10308 15912 10364
rect 15848 10304 15912 10308
rect 15928 10364 15992 10368
rect 15928 10308 15932 10364
rect 15932 10308 15988 10364
rect 15988 10308 15992 10364
rect 15928 10304 15992 10308
rect 16008 10364 16072 10368
rect 16008 10308 16012 10364
rect 16012 10308 16068 10364
rect 16068 10308 16072 10364
rect 16008 10304 16072 10308
rect 16088 10364 16152 10368
rect 16088 10308 16092 10364
rect 16092 10308 16148 10364
rect 16148 10308 16152 10364
rect 16088 10304 16152 10308
rect 25778 10364 25842 10368
rect 25778 10308 25782 10364
rect 25782 10308 25838 10364
rect 25838 10308 25842 10364
rect 25778 10304 25842 10308
rect 25858 10364 25922 10368
rect 25858 10308 25862 10364
rect 25862 10308 25918 10364
rect 25918 10308 25922 10364
rect 25858 10304 25922 10308
rect 25938 10364 26002 10368
rect 25938 10308 25942 10364
rect 25942 10308 25998 10364
rect 25998 10308 26002 10364
rect 25938 10304 26002 10308
rect 26018 10364 26082 10368
rect 26018 10308 26022 10364
rect 26022 10308 26078 10364
rect 26078 10308 26082 10364
rect 26018 10304 26082 10308
rect 10882 9820 10946 9824
rect 10882 9764 10886 9820
rect 10886 9764 10942 9820
rect 10942 9764 10946 9820
rect 10882 9760 10946 9764
rect 10962 9820 11026 9824
rect 10962 9764 10966 9820
rect 10966 9764 11022 9820
rect 11022 9764 11026 9820
rect 10962 9760 11026 9764
rect 11042 9820 11106 9824
rect 11042 9764 11046 9820
rect 11046 9764 11102 9820
rect 11102 9764 11106 9820
rect 11042 9760 11106 9764
rect 11122 9820 11186 9824
rect 11122 9764 11126 9820
rect 11126 9764 11182 9820
rect 11182 9764 11186 9820
rect 11122 9760 11186 9764
rect 20813 9820 20877 9824
rect 20813 9764 20817 9820
rect 20817 9764 20873 9820
rect 20873 9764 20877 9820
rect 20813 9760 20877 9764
rect 20893 9820 20957 9824
rect 20893 9764 20897 9820
rect 20897 9764 20953 9820
rect 20953 9764 20957 9820
rect 20893 9760 20957 9764
rect 20973 9820 21037 9824
rect 20973 9764 20977 9820
rect 20977 9764 21033 9820
rect 21033 9764 21037 9820
rect 20973 9760 21037 9764
rect 21053 9820 21117 9824
rect 21053 9764 21057 9820
rect 21057 9764 21113 9820
rect 21113 9764 21117 9820
rect 21053 9760 21117 9764
rect 5917 9276 5981 9280
rect 5917 9220 5921 9276
rect 5921 9220 5977 9276
rect 5977 9220 5981 9276
rect 5917 9216 5981 9220
rect 5997 9276 6061 9280
rect 5997 9220 6001 9276
rect 6001 9220 6057 9276
rect 6057 9220 6061 9276
rect 5997 9216 6061 9220
rect 6077 9276 6141 9280
rect 6077 9220 6081 9276
rect 6081 9220 6137 9276
rect 6137 9220 6141 9276
rect 6077 9216 6141 9220
rect 6157 9276 6221 9280
rect 6157 9220 6161 9276
rect 6161 9220 6217 9276
rect 6217 9220 6221 9276
rect 6157 9216 6221 9220
rect 15848 9276 15912 9280
rect 15848 9220 15852 9276
rect 15852 9220 15908 9276
rect 15908 9220 15912 9276
rect 15848 9216 15912 9220
rect 15928 9276 15992 9280
rect 15928 9220 15932 9276
rect 15932 9220 15988 9276
rect 15988 9220 15992 9276
rect 15928 9216 15992 9220
rect 16008 9276 16072 9280
rect 16008 9220 16012 9276
rect 16012 9220 16068 9276
rect 16068 9220 16072 9276
rect 16008 9216 16072 9220
rect 16088 9276 16152 9280
rect 16088 9220 16092 9276
rect 16092 9220 16148 9276
rect 16148 9220 16152 9276
rect 16088 9216 16152 9220
rect 25778 9276 25842 9280
rect 25778 9220 25782 9276
rect 25782 9220 25838 9276
rect 25838 9220 25842 9276
rect 25778 9216 25842 9220
rect 25858 9276 25922 9280
rect 25858 9220 25862 9276
rect 25862 9220 25918 9276
rect 25918 9220 25922 9276
rect 25858 9216 25922 9220
rect 25938 9276 26002 9280
rect 25938 9220 25942 9276
rect 25942 9220 25998 9276
rect 25998 9220 26002 9276
rect 25938 9216 26002 9220
rect 26018 9276 26082 9280
rect 26018 9220 26022 9276
rect 26022 9220 26078 9276
rect 26078 9220 26082 9276
rect 26018 9216 26082 9220
rect 10882 8732 10946 8736
rect 10882 8676 10886 8732
rect 10886 8676 10942 8732
rect 10942 8676 10946 8732
rect 10882 8672 10946 8676
rect 10962 8732 11026 8736
rect 10962 8676 10966 8732
rect 10966 8676 11022 8732
rect 11022 8676 11026 8732
rect 10962 8672 11026 8676
rect 11042 8732 11106 8736
rect 11042 8676 11046 8732
rect 11046 8676 11102 8732
rect 11102 8676 11106 8732
rect 11042 8672 11106 8676
rect 11122 8732 11186 8736
rect 11122 8676 11126 8732
rect 11126 8676 11182 8732
rect 11182 8676 11186 8732
rect 11122 8672 11186 8676
rect 20813 8732 20877 8736
rect 20813 8676 20817 8732
rect 20817 8676 20873 8732
rect 20873 8676 20877 8732
rect 20813 8672 20877 8676
rect 20893 8732 20957 8736
rect 20893 8676 20897 8732
rect 20897 8676 20953 8732
rect 20953 8676 20957 8732
rect 20893 8672 20957 8676
rect 20973 8732 21037 8736
rect 20973 8676 20977 8732
rect 20977 8676 21033 8732
rect 21033 8676 21037 8732
rect 20973 8672 21037 8676
rect 21053 8732 21117 8736
rect 21053 8676 21057 8732
rect 21057 8676 21113 8732
rect 21113 8676 21117 8732
rect 21053 8672 21117 8676
rect 5917 8188 5981 8192
rect 5917 8132 5921 8188
rect 5921 8132 5977 8188
rect 5977 8132 5981 8188
rect 5917 8128 5981 8132
rect 5997 8188 6061 8192
rect 5997 8132 6001 8188
rect 6001 8132 6057 8188
rect 6057 8132 6061 8188
rect 5997 8128 6061 8132
rect 6077 8188 6141 8192
rect 6077 8132 6081 8188
rect 6081 8132 6137 8188
rect 6137 8132 6141 8188
rect 6077 8128 6141 8132
rect 6157 8188 6221 8192
rect 6157 8132 6161 8188
rect 6161 8132 6217 8188
rect 6217 8132 6221 8188
rect 6157 8128 6221 8132
rect 15848 8188 15912 8192
rect 15848 8132 15852 8188
rect 15852 8132 15908 8188
rect 15908 8132 15912 8188
rect 15848 8128 15912 8132
rect 15928 8188 15992 8192
rect 15928 8132 15932 8188
rect 15932 8132 15988 8188
rect 15988 8132 15992 8188
rect 15928 8128 15992 8132
rect 16008 8188 16072 8192
rect 16008 8132 16012 8188
rect 16012 8132 16068 8188
rect 16068 8132 16072 8188
rect 16008 8128 16072 8132
rect 16088 8188 16152 8192
rect 16088 8132 16092 8188
rect 16092 8132 16148 8188
rect 16148 8132 16152 8188
rect 16088 8128 16152 8132
rect 25778 8188 25842 8192
rect 25778 8132 25782 8188
rect 25782 8132 25838 8188
rect 25838 8132 25842 8188
rect 25778 8128 25842 8132
rect 25858 8188 25922 8192
rect 25858 8132 25862 8188
rect 25862 8132 25918 8188
rect 25918 8132 25922 8188
rect 25858 8128 25922 8132
rect 25938 8188 26002 8192
rect 25938 8132 25942 8188
rect 25942 8132 25998 8188
rect 25998 8132 26002 8188
rect 25938 8128 26002 8132
rect 26018 8188 26082 8192
rect 26018 8132 26022 8188
rect 26022 8132 26078 8188
rect 26078 8132 26082 8188
rect 26018 8128 26082 8132
rect 10882 7644 10946 7648
rect 10882 7588 10886 7644
rect 10886 7588 10942 7644
rect 10942 7588 10946 7644
rect 10882 7584 10946 7588
rect 10962 7644 11026 7648
rect 10962 7588 10966 7644
rect 10966 7588 11022 7644
rect 11022 7588 11026 7644
rect 10962 7584 11026 7588
rect 11042 7644 11106 7648
rect 11042 7588 11046 7644
rect 11046 7588 11102 7644
rect 11102 7588 11106 7644
rect 11042 7584 11106 7588
rect 11122 7644 11186 7648
rect 11122 7588 11126 7644
rect 11126 7588 11182 7644
rect 11182 7588 11186 7644
rect 11122 7584 11186 7588
rect 20813 7644 20877 7648
rect 20813 7588 20817 7644
rect 20817 7588 20873 7644
rect 20873 7588 20877 7644
rect 20813 7584 20877 7588
rect 20893 7644 20957 7648
rect 20893 7588 20897 7644
rect 20897 7588 20953 7644
rect 20953 7588 20957 7644
rect 20893 7584 20957 7588
rect 20973 7644 21037 7648
rect 20973 7588 20977 7644
rect 20977 7588 21033 7644
rect 21033 7588 21037 7644
rect 20973 7584 21037 7588
rect 21053 7644 21117 7648
rect 21053 7588 21057 7644
rect 21057 7588 21113 7644
rect 21113 7588 21117 7644
rect 21053 7584 21117 7588
rect 5917 7100 5981 7104
rect 5917 7044 5921 7100
rect 5921 7044 5977 7100
rect 5977 7044 5981 7100
rect 5917 7040 5981 7044
rect 5997 7100 6061 7104
rect 5997 7044 6001 7100
rect 6001 7044 6057 7100
rect 6057 7044 6061 7100
rect 5997 7040 6061 7044
rect 6077 7100 6141 7104
rect 6077 7044 6081 7100
rect 6081 7044 6137 7100
rect 6137 7044 6141 7100
rect 6077 7040 6141 7044
rect 6157 7100 6221 7104
rect 6157 7044 6161 7100
rect 6161 7044 6217 7100
rect 6217 7044 6221 7100
rect 6157 7040 6221 7044
rect 15848 7100 15912 7104
rect 15848 7044 15852 7100
rect 15852 7044 15908 7100
rect 15908 7044 15912 7100
rect 15848 7040 15912 7044
rect 15928 7100 15992 7104
rect 15928 7044 15932 7100
rect 15932 7044 15988 7100
rect 15988 7044 15992 7100
rect 15928 7040 15992 7044
rect 16008 7100 16072 7104
rect 16008 7044 16012 7100
rect 16012 7044 16068 7100
rect 16068 7044 16072 7100
rect 16008 7040 16072 7044
rect 16088 7100 16152 7104
rect 16088 7044 16092 7100
rect 16092 7044 16148 7100
rect 16148 7044 16152 7100
rect 16088 7040 16152 7044
rect 25778 7100 25842 7104
rect 25778 7044 25782 7100
rect 25782 7044 25838 7100
rect 25838 7044 25842 7100
rect 25778 7040 25842 7044
rect 25858 7100 25922 7104
rect 25858 7044 25862 7100
rect 25862 7044 25918 7100
rect 25918 7044 25922 7100
rect 25858 7040 25922 7044
rect 25938 7100 26002 7104
rect 25938 7044 25942 7100
rect 25942 7044 25998 7100
rect 25998 7044 26002 7100
rect 25938 7040 26002 7044
rect 26018 7100 26082 7104
rect 26018 7044 26022 7100
rect 26022 7044 26078 7100
rect 26078 7044 26082 7100
rect 26018 7040 26082 7044
rect 10882 6556 10946 6560
rect 10882 6500 10886 6556
rect 10886 6500 10942 6556
rect 10942 6500 10946 6556
rect 10882 6496 10946 6500
rect 10962 6556 11026 6560
rect 10962 6500 10966 6556
rect 10966 6500 11022 6556
rect 11022 6500 11026 6556
rect 10962 6496 11026 6500
rect 11042 6556 11106 6560
rect 11042 6500 11046 6556
rect 11046 6500 11102 6556
rect 11102 6500 11106 6556
rect 11042 6496 11106 6500
rect 11122 6556 11186 6560
rect 11122 6500 11126 6556
rect 11126 6500 11182 6556
rect 11182 6500 11186 6556
rect 11122 6496 11186 6500
rect 20813 6556 20877 6560
rect 20813 6500 20817 6556
rect 20817 6500 20873 6556
rect 20873 6500 20877 6556
rect 20813 6496 20877 6500
rect 20893 6556 20957 6560
rect 20893 6500 20897 6556
rect 20897 6500 20953 6556
rect 20953 6500 20957 6556
rect 20893 6496 20957 6500
rect 20973 6556 21037 6560
rect 20973 6500 20977 6556
rect 20977 6500 21033 6556
rect 21033 6500 21037 6556
rect 20973 6496 21037 6500
rect 21053 6556 21117 6560
rect 21053 6500 21057 6556
rect 21057 6500 21113 6556
rect 21113 6500 21117 6556
rect 21053 6496 21117 6500
rect 5917 6012 5981 6016
rect 5917 5956 5921 6012
rect 5921 5956 5977 6012
rect 5977 5956 5981 6012
rect 5917 5952 5981 5956
rect 5997 6012 6061 6016
rect 5997 5956 6001 6012
rect 6001 5956 6057 6012
rect 6057 5956 6061 6012
rect 5997 5952 6061 5956
rect 6077 6012 6141 6016
rect 6077 5956 6081 6012
rect 6081 5956 6137 6012
rect 6137 5956 6141 6012
rect 6077 5952 6141 5956
rect 6157 6012 6221 6016
rect 6157 5956 6161 6012
rect 6161 5956 6217 6012
rect 6217 5956 6221 6012
rect 6157 5952 6221 5956
rect 15848 6012 15912 6016
rect 15848 5956 15852 6012
rect 15852 5956 15908 6012
rect 15908 5956 15912 6012
rect 15848 5952 15912 5956
rect 15928 6012 15992 6016
rect 15928 5956 15932 6012
rect 15932 5956 15988 6012
rect 15988 5956 15992 6012
rect 15928 5952 15992 5956
rect 16008 6012 16072 6016
rect 16008 5956 16012 6012
rect 16012 5956 16068 6012
rect 16068 5956 16072 6012
rect 16008 5952 16072 5956
rect 16088 6012 16152 6016
rect 16088 5956 16092 6012
rect 16092 5956 16148 6012
rect 16148 5956 16152 6012
rect 16088 5952 16152 5956
rect 25778 6012 25842 6016
rect 25778 5956 25782 6012
rect 25782 5956 25838 6012
rect 25838 5956 25842 6012
rect 25778 5952 25842 5956
rect 25858 6012 25922 6016
rect 25858 5956 25862 6012
rect 25862 5956 25918 6012
rect 25918 5956 25922 6012
rect 25858 5952 25922 5956
rect 25938 6012 26002 6016
rect 25938 5956 25942 6012
rect 25942 5956 25998 6012
rect 25998 5956 26002 6012
rect 25938 5952 26002 5956
rect 26018 6012 26082 6016
rect 26018 5956 26022 6012
rect 26022 5956 26078 6012
rect 26078 5956 26082 6012
rect 26018 5952 26082 5956
rect 10882 5468 10946 5472
rect 10882 5412 10886 5468
rect 10886 5412 10942 5468
rect 10942 5412 10946 5468
rect 10882 5408 10946 5412
rect 10962 5468 11026 5472
rect 10962 5412 10966 5468
rect 10966 5412 11022 5468
rect 11022 5412 11026 5468
rect 10962 5408 11026 5412
rect 11042 5468 11106 5472
rect 11042 5412 11046 5468
rect 11046 5412 11102 5468
rect 11102 5412 11106 5468
rect 11042 5408 11106 5412
rect 11122 5468 11186 5472
rect 11122 5412 11126 5468
rect 11126 5412 11182 5468
rect 11182 5412 11186 5468
rect 11122 5408 11186 5412
rect 20813 5468 20877 5472
rect 20813 5412 20817 5468
rect 20817 5412 20873 5468
rect 20873 5412 20877 5468
rect 20813 5408 20877 5412
rect 20893 5468 20957 5472
rect 20893 5412 20897 5468
rect 20897 5412 20953 5468
rect 20953 5412 20957 5468
rect 20893 5408 20957 5412
rect 20973 5468 21037 5472
rect 20973 5412 20977 5468
rect 20977 5412 21033 5468
rect 21033 5412 21037 5468
rect 20973 5408 21037 5412
rect 21053 5468 21117 5472
rect 21053 5412 21057 5468
rect 21057 5412 21113 5468
rect 21113 5412 21117 5468
rect 21053 5408 21117 5412
rect 5917 4924 5981 4928
rect 5917 4868 5921 4924
rect 5921 4868 5977 4924
rect 5977 4868 5981 4924
rect 5917 4864 5981 4868
rect 5997 4924 6061 4928
rect 5997 4868 6001 4924
rect 6001 4868 6057 4924
rect 6057 4868 6061 4924
rect 5997 4864 6061 4868
rect 6077 4924 6141 4928
rect 6077 4868 6081 4924
rect 6081 4868 6137 4924
rect 6137 4868 6141 4924
rect 6077 4864 6141 4868
rect 6157 4924 6221 4928
rect 6157 4868 6161 4924
rect 6161 4868 6217 4924
rect 6217 4868 6221 4924
rect 6157 4864 6221 4868
rect 15848 4924 15912 4928
rect 15848 4868 15852 4924
rect 15852 4868 15908 4924
rect 15908 4868 15912 4924
rect 15848 4864 15912 4868
rect 15928 4924 15992 4928
rect 15928 4868 15932 4924
rect 15932 4868 15988 4924
rect 15988 4868 15992 4924
rect 15928 4864 15992 4868
rect 16008 4924 16072 4928
rect 16008 4868 16012 4924
rect 16012 4868 16068 4924
rect 16068 4868 16072 4924
rect 16008 4864 16072 4868
rect 16088 4924 16152 4928
rect 16088 4868 16092 4924
rect 16092 4868 16148 4924
rect 16148 4868 16152 4924
rect 16088 4864 16152 4868
rect 25778 4924 25842 4928
rect 25778 4868 25782 4924
rect 25782 4868 25838 4924
rect 25838 4868 25842 4924
rect 25778 4864 25842 4868
rect 25858 4924 25922 4928
rect 25858 4868 25862 4924
rect 25862 4868 25918 4924
rect 25918 4868 25922 4924
rect 25858 4864 25922 4868
rect 25938 4924 26002 4928
rect 25938 4868 25942 4924
rect 25942 4868 25998 4924
rect 25998 4868 26002 4924
rect 25938 4864 26002 4868
rect 26018 4924 26082 4928
rect 26018 4868 26022 4924
rect 26022 4868 26078 4924
rect 26078 4868 26082 4924
rect 26018 4864 26082 4868
rect 10882 4380 10946 4384
rect 10882 4324 10886 4380
rect 10886 4324 10942 4380
rect 10942 4324 10946 4380
rect 10882 4320 10946 4324
rect 10962 4380 11026 4384
rect 10962 4324 10966 4380
rect 10966 4324 11022 4380
rect 11022 4324 11026 4380
rect 10962 4320 11026 4324
rect 11042 4380 11106 4384
rect 11042 4324 11046 4380
rect 11046 4324 11102 4380
rect 11102 4324 11106 4380
rect 11042 4320 11106 4324
rect 11122 4380 11186 4384
rect 11122 4324 11126 4380
rect 11126 4324 11182 4380
rect 11182 4324 11186 4380
rect 11122 4320 11186 4324
rect 20813 4380 20877 4384
rect 20813 4324 20817 4380
rect 20817 4324 20873 4380
rect 20873 4324 20877 4380
rect 20813 4320 20877 4324
rect 20893 4380 20957 4384
rect 20893 4324 20897 4380
rect 20897 4324 20953 4380
rect 20953 4324 20957 4380
rect 20893 4320 20957 4324
rect 20973 4380 21037 4384
rect 20973 4324 20977 4380
rect 20977 4324 21033 4380
rect 21033 4324 21037 4380
rect 20973 4320 21037 4324
rect 21053 4380 21117 4384
rect 21053 4324 21057 4380
rect 21057 4324 21113 4380
rect 21113 4324 21117 4380
rect 21053 4320 21117 4324
rect 5917 3836 5981 3840
rect 5917 3780 5921 3836
rect 5921 3780 5977 3836
rect 5977 3780 5981 3836
rect 5917 3776 5981 3780
rect 5997 3836 6061 3840
rect 5997 3780 6001 3836
rect 6001 3780 6057 3836
rect 6057 3780 6061 3836
rect 5997 3776 6061 3780
rect 6077 3836 6141 3840
rect 6077 3780 6081 3836
rect 6081 3780 6137 3836
rect 6137 3780 6141 3836
rect 6077 3776 6141 3780
rect 6157 3836 6221 3840
rect 6157 3780 6161 3836
rect 6161 3780 6217 3836
rect 6217 3780 6221 3836
rect 6157 3776 6221 3780
rect 15848 3836 15912 3840
rect 15848 3780 15852 3836
rect 15852 3780 15908 3836
rect 15908 3780 15912 3836
rect 15848 3776 15912 3780
rect 15928 3836 15992 3840
rect 15928 3780 15932 3836
rect 15932 3780 15988 3836
rect 15988 3780 15992 3836
rect 15928 3776 15992 3780
rect 16008 3836 16072 3840
rect 16008 3780 16012 3836
rect 16012 3780 16068 3836
rect 16068 3780 16072 3836
rect 16008 3776 16072 3780
rect 16088 3836 16152 3840
rect 16088 3780 16092 3836
rect 16092 3780 16148 3836
rect 16148 3780 16152 3836
rect 16088 3776 16152 3780
rect 25778 3836 25842 3840
rect 25778 3780 25782 3836
rect 25782 3780 25838 3836
rect 25838 3780 25842 3836
rect 25778 3776 25842 3780
rect 25858 3836 25922 3840
rect 25858 3780 25862 3836
rect 25862 3780 25918 3836
rect 25918 3780 25922 3836
rect 25858 3776 25922 3780
rect 25938 3836 26002 3840
rect 25938 3780 25942 3836
rect 25942 3780 25998 3836
rect 25998 3780 26002 3836
rect 25938 3776 26002 3780
rect 26018 3836 26082 3840
rect 26018 3780 26022 3836
rect 26022 3780 26078 3836
rect 26078 3780 26082 3836
rect 26018 3776 26082 3780
rect 10882 3292 10946 3296
rect 10882 3236 10886 3292
rect 10886 3236 10942 3292
rect 10942 3236 10946 3292
rect 10882 3232 10946 3236
rect 10962 3292 11026 3296
rect 10962 3236 10966 3292
rect 10966 3236 11022 3292
rect 11022 3236 11026 3292
rect 10962 3232 11026 3236
rect 11042 3292 11106 3296
rect 11042 3236 11046 3292
rect 11046 3236 11102 3292
rect 11102 3236 11106 3292
rect 11042 3232 11106 3236
rect 11122 3292 11186 3296
rect 11122 3236 11126 3292
rect 11126 3236 11182 3292
rect 11182 3236 11186 3292
rect 11122 3232 11186 3236
rect 20813 3292 20877 3296
rect 20813 3236 20817 3292
rect 20817 3236 20873 3292
rect 20873 3236 20877 3292
rect 20813 3232 20877 3236
rect 20893 3292 20957 3296
rect 20893 3236 20897 3292
rect 20897 3236 20953 3292
rect 20953 3236 20957 3292
rect 20893 3232 20957 3236
rect 20973 3292 21037 3296
rect 20973 3236 20977 3292
rect 20977 3236 21033 3292
rect 21033 3236 21037 3292
rect 20973 3232 21037 3236
rect 21053 3292 21117 3296
rect 21053 3236 21057 3292
rect 21057 3236 21113 3292
rect 21113 3236 21117 3292
rect 21053 3232 21117 3236
rect 5917 2748 5981 2752
rect 5917 2692 5921 2748
rect 5921 2692 5977 2748
rect 5977 2692 5981 2748
rect 5917 2688 5981 2692
rect 5997 2748 6061 2752
rect 5997 2692 6001 2748
rect 6001 2692 6057 2748
rect 6057 2692 6061 2748
rect 5997 2688 6061 2692
rect 6077 2748 6141 2752
rect 6077 2692 6081 2748
rect 6081 2692 6137 2748
rect 6137 2692 6141 2748
rect 6077 2688 6141 2692
rect 6157 2748 6221 2752
rect 6157 2692 6161 2748
rect 6161 2692 6217 2748
rect 6217 2692 6221 2748
rect 6157 2688 6221 2692
rect 15848 2748 15912 2752
rect 15848 2692 15852 2748
rect 15852 2692 15908 2748
rect 15908 2692 15912 2748
rect 15848 2688 15912 2692
rect 15928 2748 15992 2752
rect 15928 2692 15932 2748
rect 15932 2692 15988 2748
rect 15988 2692 15992 2748
rect 15928 2688 15992 2692
rect 16008 2748 16072 2752
rect 16008 2692 16012 2748
rect 16012 2692 16068 2748
rect 16068 2692 16072 2748
rect 16008 2688 16072 2692
rect 16088 2748 16152 2752
rect 16088 2692 16092 2748
rect 16092 2692 16148 2748
rect 16148 2692 16152 2748
rect 16088 2688 16152 2692
rect 25778 2748 25842 2752
rect 25778 2692 25782 2748
rect 25782 2692 25838 2748
rect 25838 2692 25842 2748
rect 25778 2688 25842 2692
rect 25858 2748 25922 2752
rect 25858 2692 25862 2748
rect 25862 2692 25918 2748
rect 25918 2692 25922 2748
rect 25858 2688 25922 2692
rect 25938 2748 26002 2752
rect 25938 2692 25942 2748
rect 25942 2692 25998 2748
rect 25998 2692 26002 2748
rect 25938 2688 26002 2692
rect 26018 2748 26082 2752
rect 26018 2692 26022 2748
rect 26022 2692 26078 2748
rect 26078 2692 26082 2748
rect 26018 2688 26082 2692
rect 10882 2204 10946 2208
rect 10882 2148 10886 2204
rect 10886 2148 10942 2204
rect 10942 2148 10946 2204
rect 10882 2144 10946 2148
rect 10962 2204 11026 2208
rect 10962 2148 10966 2204
rect 10966 2148 11022 2204
rect 11022 2148 11026 2204
rect 10962 2144 11026 2148
rect 11042 2204 11106 2208
rect 11042 2148 11046 2204
rect 11046 2148 11102 2204
rect 11102 2148 11106 2204
rect 11042 2144 11106 2148
rect 11122 2204 11186 2208
rect 11122 2148 11126 2204
rect 11126 2148 11182 2204
rect 11182 2148 11186 2204
rect 11122 2144 11186 2148
rect 20813 2204 20877 2208
rect 20813 2148 20817 2204
rect 20817 2148 20873 2204
rect 20873 2148 20877 2204
rect 20813 2144 20877 2148
rect 20893 2204 20957 2208
rect 20893 2148 20897 2204
rect 20897 2148 20953 2204
rect 20953 2148 20957 2204
rect 20893 2144 20957 2148
rect 20973 2204 21037 2208
rect 20973 2148 20977 2204
rect 20977 2148 21033 2204
rect 21033 2148 21037 2204
rect 20973 2144 21037 2148
rect 21053 2204 21117 2208
rect 21053 2148 21057 2204
rect 21057 2148 21113 2204
rect 21113 2148 21117 2204
rect 21053 2144 21117 2148
<< metal4 >>
rect 5909 45184 6229 45744
rect 5909 45120 5917 45184
rect 5981 45120 5997 45184
rect 6061 45120 6077 45184
rect 6141 45120 6157 45184
rect 6221 45120 6229 45184
rect 5909 44096 6229 45120
rect 5909 44032 5917 44096
rect 5981 44032 5997 44096
rect 6061 44032 6077 44096
rect 6141 44032 6157 44096
rect 6221 44032 6229 44096
rect 5909 43008 6229 44032
rect 5909 42944 5917 43008
rect 5981 42944 5997 43008
rect 6061 42944 6077 43008
rect 6141 42944 6157 43008
rect 6221 42944 6229 43008
rect 5909 41920 6229 42944
rect 5909 41856 5917 41920
rect 5981 41856 5997 41920
rect 6061 41856 6077 41920
rect 6141 41856 6157 41920
rect 6221 41856 6229 41920
rect 5909 40832 6229 41856
rect 5909 40768 5917 40832
rect 5981 40768 5997 40832
rect 6061 40768 6077 40832
rect 6141 40768 6157 40832
rect 6221 40768 6229 40832
rect 5909 39744 6229 40768
rect 5909 39680 5917 39744
rect 5981 39680 5997 39744
rect 6061 39680 6077 39744
rect 6141 39680 6157 39744
rect 6221 39680 6229 39744
rect 5909 38656 6229 39680
rect 5909 38592 5917 38656
rect 5981 38592 5997 38656
rect 6061 38592 6077 38656
rect 6141 38592 6157 38656
rect 6221 38592 6229 38656
rect 5909 37568 6229 38592
rect 5909 37504 5917 37568
rect 5981 37504 5997 37568
rect 6061 37504 6077 37568
rect 6141 37504 6157 37568
rect 6221 37504 6229 37568
rect 5909 36480 6229 37504
rect 5909 36416 5917 36480
rect 5981 36416 5997 36480
rect 6061 36416 6077 36480
rect 6141 36416 6157 36480
rect 6221 36416 6229 36480
rect 5909 35392 6229 36416
rect 5909 35328 5917 35392
rect 5981 35328 5997 35392
rect 6061 35328 6077 35392
rect 6141 35328 6157 35392
rect 6221 35328 6229 35392
rect 5909 34304 6229 35328
rect 5909 34240 5917 34304
rect 5981 34240 5997 34304
rect 6061 34240 6077 34304
rect 6141 34240 6157 34304
rect 6221 34240 6229 34304
rect 5909 33216 6229 34240
rect 5909 33152 5917 33216
rect 5981 33152 5997 33216
rect 6061 33152 6077 33216
rect 6141 33152 6157 33216
rect 6221 33152 6229 33216
rect 5909 32128 6229 33152
rect 5909 32064 5917 32128
rect 5981 32064 5997 32128
rect 6061 32064 6077 32128
rect 6141 32064 6157 32128
rect 6221 32064 6229 32128
rect 5909 31040 6229 32064
rect 5909 30976 5917 31040
rect 5981 30976 5997 31040
rect 6061 30976 6077 31040
rect 6141 30976 6157 31040
rect 6221 30976 6229 31040
rect 5909 29952 6229 30976
rect 5909 29888 5917 29952
rect 5981 29888 5997 29952
rect 6061 29888 6077 29952
rect 6141 29888 6157 29952
rect 6221 29888 6229 29952
rect 5909 28864 6229 29888
rect 5909 28800 5917 28864
rect 5981 28800 5997 28864
rect 6061 28800 6077 28864
rect 6141 28800 6157 28864
rect 6221 28800 6229 28864
rect 5909 27776 6229 28800
rect 5909 27712 5917 27776
rect 5981 27712 5997 27776
rect 6061 27712 6077 27776
rect 6141 27712 6157 27776
rect 6221 27712 6229 27776
rect 5909 26688 6229 27712
rect 5909 26624 5917 26688
rect 5981 26624 5997 26688
rect 6061 26624 6077 26688
rect 6141 26624 6157 26688
rect 6221 26624 6229 26688
rect 5909 25600 6229 26624
rect 10874 45728 11194 45744
rect 10874 45664 10882 45728
rect 10946 45664 10962 45728
rect 11026 45664 11042 45728
rect 11106 45664 11122 45728
rect 11186 45664 11194 45728
rect 10874 44640 11194 45664
rect 10874 44576 10882 44640
rect 10946 44576 10962 44640
rect 11026 44576 11042 44640
rect 11106 44576 11122 44640
rect 11186 44576 11194 44640
rect 10874 43552 11194 44576
rect 10874 43488 10882 43552
rect 10946 43488 10962 43552
rect 11026 43488 11042 43552
rect 11106 43488 11122 43552
rect 11186 43488 11194 43552
rect 10874 42464 11194 43488
rect 10874 42400 10882 42464
rect 10946 42400 10962 42464
rect 11026 42400 11042 42464
rect 11106 42400 11122 42464
rect 11186 42400 11194 42464
rect 10874 41376 11194 42400
rect 10874 41312 10882 41376
rect 10946 41312 10962 41376
rect 11026 41312 11042 41376
rect 11106 41312 11122 41376
rect 11186 41312 11194 41376
rect 10874 40288 11194 41312
rect 10874 40224 10882 40288
rect 10946 40224 10962 40288
rect 11026 40224 11042 40288
rect 11106 40224 11122 40288
rect 11186 40224 11194 40288
rect 10874 39200 11194 40224
rect 10874 39136 10882 39200
rect 10946 39136 10962 39200
rect 11026 39136 11042 39200
rect 11106 39136 11122 39200
rect 11186 39136 11194 39200
rect 10874 38112 11194 39136
rect 10874 38048 10882 38112
rect 10946 38048 10962 38112
rect 11026 38048 11042 38112
rect 11106 38048 11122 38112
rect 11186 38048 11194 38112
rect 10874 37024 11194 38048
rect 10874 36960 10882 37024
rect 10946 36960 10962 37024
rect 11026 36960 11042 37024
rect 11106 36960 11122 37024
rect 11186 36960 11194 37024
rect 10874 35936 11194 36960
rect 10874 35872 10882 35936
rect 10946 35872 10962 35936
rect 11026 35872 11042 35936
rect 11106 35872 11122 35936
rect 11186 35872 11194 35936
rect 10874 34848 11194 35872
rect 10874 34784 10882 34848
rect 10946 34784 10962 34848
rect 11026 34784 11042 34848
rect 11106 34784 11122 34848
rect 11186 34784 11194 34848
rect 10874 33760 11194 34784
rect 10874 33696 10882 33760
rect 10946 33696 10962 33760
rect 11026 33696 11042 33760
rect 11106 33696 11122 33760
rect 11186 33696 11194 33760
rect 10874 32672 11194 33696
rect 10874 32608 10882 32672
rect 10946 32608 10962 32672
rect 11026 32608 11042 32672
rect 11106 32608 11122 32672
rect 11186 32608 11194 32672
rect 10874 31584 11194 32608
rect 15839 45184 16160 45744
rect 15839 45120 15848 45184
rect 15912 45120 15928 45184
rect 15992 45120 16008 45184
rect 16072 45120 16088 45184
rect 16152 45120 16160 45184
rect 15839 44096 16160 45120
rect 15839 44032 15848 44096
rect 15912 44032 15928 44096
rect 15992 44032 16008 44096
rect 16072 44032 16088 44096
rect 16152 44032 16160 44096
rect 15839 43008 16160 44032
rect 15839 42944 15848 43008
rect 15912 42944 15928 43008
rect 15992 42944 16008 43008
rect 16072 42944 16088 43008
rect 16152 42944 16160 43008
rect 15839 41920 16160 42944
rect 15839 41856 15848 41920
rect 15912 41856 15928 41920
rect 15992 41856 16008 41920
rect 16072 41856 16088 41920
rect 16152 41856 16160 41920
rect 15839 40832 16160 41856
rect 15839 40768 15848 40832
rect 15912 40768 15928 40832
rect 15992 40768 16008 40832
rect 16072 40768 16088 40832
rect 16152 40768 16160 40832
rect 15839 39744 16160 40768
rect 15839 39680 15848 39744
rect 15912 39680 15928 39744
rect 15992 39680 16008 39744
rect 16072 39680 16088 39744
rect 16152 39680 16160 39744
rect 15839 38656 16160 39680
rect 15839 38592 15848 38656
rect 15912 38592 15928 38656
rect 15992 38592 16008 38656
rect 16072 38592 16088 38656
rect 16152 38592 16160 38656
rect 15839 37568 16160 38592
rect 15839 37504 15848 37568
rect 15912 37504 15928 37568
rect 15992 37504 16008 37568
rect 16072 37504 16088 37568
rect 16152 37504 16160 37568
rect 15839 36480 16160 37504
rect 15839 36416 15848 36480
rect 15912 36416 15928 36480
rect 15992 36416 16008 36480
rect 16072 36416 16088 36480
rect 16152 36416 16160 36480
rect 15839 35392 16160 36416
rect 15839 35328 15848 35392
rect 15912 35328 15928 35392
rect 15992 35328 16008 35392
rect 16072 35328 16088 35392
rect 16152 35328 16160 35392
rect 15839 34304 16160 35328
rect 15839 34240 15848 34304
rect 15912 34240 15928 34304
rect 15992 34240 16008 34304
rect 16072 34240 16088 34304
rect 16152 34240 16160 34304
rect 15839 33216 16160 34240
rect 15839 33152 15848 33216
rect 15912 33152 15928 33216
rect 15992 33152 16008 33216
rect 16072 33152 16088 33216
rect 16152 33152 16160 33216
rect 15839 32128 16160 33152
rect 15839 32064 15848 32128
rect 15912 32064 15928 32128
rect 15992 32064 16008 32128
rect 16072 32064 16088 32128
rect 16152 32064 16160 32128
rect 11283 31788 11349 31789
rect 11283 31724 11284 31788
rect 11348 31724 11349 31788
rect 11283 31723 11349 31724
rect 10874 31520 10882 31584
rect 10946 31520 10962 31584
rect 11026 31520 11042 31584
rect 11106 31520 11122 31584
rect 11186 31520 11194 31584
rect 10874 30496 11194 31520
rect 10874 30432 10882 30496
rect 10946 30432 10962 30496
rect 11026 30432 11042 30496
rect 11106 30432 11122 30496
rect 11186 30432 11194 30496
rect 10874 29408 11194 30432
rect 10874 29344 10882 29408
rect 10946 29344 10962 29408
rect 11026 29344 11042 29408
rect 11106 29344 11122 29408
rect 11186 29344 11194 29408
rect 10874 28320 11194 29344
rect 10874 28256 10882 28320
rect 10946 28256 10962 28320
rect 11026 28256 11042 28320
rect 11106 28256 11122 28320
rect 11186 28256 11194 28320
rect 10874 27232 11194 28256
rect 10874 27168 10882 27232
rect 10946 27168 10962 27232
rect 11026 27168 11042 27232
rect 11106 27168 11122 27232
rect 11186 27168 11194 27232
rect 7971 26348 8037 26349
rect 7971 26284 7972 26348
rect 8036 26284 8037 26348
rect 7971 26283 8037 26284
rect 5909 25536 5917 25600
rect 5981 25536 5997 25600
rect 6061 25536 6077 25600
rect 6141 25536 6157 25600
rect 6221 25536 6229 25600
rect 5909 24512 6229 25536
rect 5909 24448 5917 24512
rect 5981 24448 5997 24512
rect 6061 24448 6077 24512
rect 6141 24448 6157 24512
rect 6221 24448 6229 24512
rect 5909 23424 6229 24448
rect 5909 23360 5917 23424
rect 5981 23360 5997 23424
rect 6061 23360 6077 23424
rect 6141 23360 6157 23424
rect 6221 23360 6229 23424
rect 5909 22336 6229 23360
rect 5909 22272 5917 22336
rect 5981 22272 5997 22336
rect 6061 22272 6077 22336
rect 6141 22272 6157 22336
rect 6221 22272 6229 22336
rect 5909 21248 6229 22272
rect 7974 21725 8034 26283
rect 10874 26144 11194 27168
rect 10874 26080 10882 26144
rect 10946 26080 10962 26144
rect 11026 26080 11042 26144
rect 11106 26080 11122 26144
rect 11186 26080 11194 26144
rect 10874 25056 11194 26080
rect 10874 24992 10882 25056
rect 10946 24992 10962 25056
rect 11026 24992 11042 25056
rect 11106 24992 11122 25056
rect 11186 24992 11194 25056
rect 10874 23968 11194 24992
rect 10874 23904 10882 23968
rect 10946 23904 10962 23968
rect 11026 23904 11042 23968
rect 11106 23904 11122 23968
rect 11186 23904 11194 23968
rect 10874 22880 11194 23904
rect 10874 22816 10882 22880
rect 10946 22816 10962 22880
rect 11026 22816 11042 22880
rect 11106 22816 11122 22880
rect 11186 22816 11194 22880
rect 9443 22676 9509 22677
rect 9443 22612 9444 22676
rect 9508 22612 9509 22676
rect 9443 22611 9509 22612
rect 7971 21724 8037 21725
rect 7971 21660 7972 21724
rect 8036 21660 8037 21724
rect 7971 21659 8037 21660
rect 5909 21184 5917 21248
rect 5981 21184 5997 21248
rect 6061 21184 6077 21248
rect 6141 21184 6157 21248
rect 6221 21184 6229 21248
rect 5909 20160 6229 21184
rect 9446 21181 9506 22611
rect 10874 21792 11194 22816
rect 10874 21728 10882 21792
rect 10946 21728 10962 21792
rect 11026 21728 11042 21792
rect 11106 21728 11122 21792
rect 11186 21728 11194 21792
rect 9443 21180 9509 21181
rect 9443 21116 9444 21180
rect 9508 21116 9509 21180
rect 9443 21115 9509 21116
rect 5909 20096 5917 20160
rect 5981 20096 5997 20160
rect 6061 20096 6077 20160
rect 6141 20096 6157 20160
rect 6221 20096 6229 20160
rect 5909 19072 6229 20096
rect 5909 19008 5917 19072
rect 5981 19008 5997 19072
rect 6061 19008 6077 19072
rect 6141 19008 6157 19072
rect 6221 19008 6229 19072
rect 5909 17984 6229 19008
rect 5909 17920 5917 17984
rect 5981 17920 5997 17984
rect 6061 17920 6077 17984
rect 6141 17920 6157 17984
rect 6221 17920 6229 17984
rect 5909 16896 6229 17920
rect 10874 20704 11194 21728
rect 10874 20640 10882 20704
rect 10946 20640 10962 20704
rect 11026 20640 11042 20704
rect 11106 20640 11122 20704
rect 11186 20640 11194 20704
rect 10874 19616 11194 20640
rect 10874 19552 10882 19616
rect 10946 19552 10962 19616
rect 11026 19552 11042 19616
rect 11106 19552 11122 19616
rect 11186 19552 11194 19616
rect 10874 18528 11194 19552
rect 11286 19141 11346 31723
rect 15839 31040 16160 32064
rect 15839 30976 15848 31040
rect 15912 30976 15928 31040
rect 15992 30976 16008 31040
rect 16072 30976 16088 31040
rect 16152 30976 16160 31040
rect 15839 29952 16160 30976
rect 15839 29888 15848 29952
rect 15912 29888 15928 29952
rect 15992 29888 16008 29952
rect 16072 29888 16088 29952
rect 16152 29888 16160 29952
rect 15839 28864 16160 29888
rect 15839 28800 15848 28864
rect 15912 28800 15928 28864
rect 15992 28800 16008 28864
rect 16072 28800 16088 28864
rect 16152 28800 16160 28864
rect 15839 27776 16160 28800
rect 15839 27712 15848 27776
rect 15912 27712 15928 27776
rect 15992 27712 16008 27776
rect 16072 27712 16088 27776
rect 16152 27712 16160 27776
rect 15839 26688 16160 27712
rect 20805 45728 21125 45744
rect 20805 45664 20813 45728
rect 20877 45664 20893 45728
rect 20957 45664 20973 45728
rect 21037 45664 21053 45728
rect 21117 45664 21125 45728
rect 20805 44640 21125 45664
rect 20805 44576 20813 44640
rect 20877 44576 20893 44640
rect 20957 44576 20973 44640
rect 21037 44576 21053 44640
rect 21117 44576 21125 44640
rect 20805 43552 21125 44576
rect 20805 43488 20813 43552
rect 20877 43488 20893 43552
rect 20957 43488 20973 43552
rect 21037 43488 21053 43552
rect 21117 43488 21125 43552
rect 20805 42464 21125 43488
rect 20805 42400 20813 42464
rect 20877 42400 20893 42464
rect 20957 42400 20973 42464
rect 21037 42400 21053 42464
rect 21117 42400 21125 42464
rect 20805 41376 21125 42400
rect 20805 41312 20813 41376
rect 20877 41312 20893 41376
rect 20957 41312 20973 41376
rect 21037 41312 21053 41376
rect 21117 41312 21125 41376
rect 20805 40288 21125 41312
rect 20805 40224 20813 40288
rect 20877 40224 20893 40288
rect 20957 40224 20973 40288
rect 21037 40224 21053 40288
rect 21117 40224 21125 40288
rect 20805 39200 21125 40224
rect 20805 39136 20813 39200
rect 20877 39136 20893 39200
rect 20957 39136 20973 39200
rect 21037 39136 21053 39200
rect 21117 39136 21125 39200
rect 20805 38112 21125 39136
rect 20805 38048 20813 38112
rect 20877 38048 20893 38112
rect 20957 38048 20973 38112
rect 21037 38048 21053 38112
rect 21117 38048 21125 38112
rect 20805 37024 21125 38048
rect 20805 36960 20813 37024
rect 20877 36960 20893 37024
rect 20957 36960 20973 37024
rect 21037 36960 21053 37024
rect 21117 36960 21125 37024
rect 20805 35936 21125 36960
rect 20805 35872 20813 35936
rect 20877 35872 20893 35936
rect 20957 35872 20973 35936
rect 21037 35872 21053 35936
rect 21117 35872 21125 35936
rect 20805 34848 21125 35872
rect 20805 34784 20813 34848
rect 20877 34784 20893 34848
rect 20957 34784 20973 34848
rect 21037 34784 21053 34848
rect 21117 34784 21125 34848
rect 20805 33760 21125 34784
rect 20805 33696 20813 33760
rect 20877 33696 20893 33760
rect 20957 33696 20973 33760
rect 21037 33696 21053 33760
rect 21117 33696 21125 33760
rect 20805 32672 21125 33696
rect 20805 32608 20813 32672
rect 20877 32608 20893 32672
rect 20957 32608 20973 32672
rect 21037 32608 21053 32672
rect 21117 32608 21125 32672
rect 20805 31584 21125 32608
rect 20805 31520 20813 31584
rect 20877 31520 20893 31584
rect 20957 31520 20973 31584
rect 21037 31520 21053 31584
rect 21117 31520 21125 31584
rect 20805 30496 21125 31520
rect 20805 30432 20813 30496
rect 20877 30432 20893 30496
rect 20957 30432 20973 30496
rect 21037 30432 21053 30496
rect 21117 30432 21125 30496
rect 20805 29408 21125 30432
rect 20805 29344 20813 29408
rect 20877 29344 20893 29408
rect 20957 29344 20973 29408
rect 21037 29344 21053 29408
rect 21117 29344 21125 29408
rect 20805 28320 21125 29344
rect 20805 28256 20813 28320
rect 20877 28256 20893 28320
rect 20957 28256 20973 28320
rect 21037 28256 21053 28320
rect 21117 28256 21125 28320
rect 17539 27436 17605 27437
rect 17539 27372 17540 27436
rect 17604 27372 17605 27436
rect 17539 27371 17605 27372
rect 15839 26624 15848 26688
rect 15912 26624 15928 26688
rect 15992 26624 16008 26688
rect 16072 26624 16088 26688
rect 16152 26624 16160 26688
rect 15839 25600 16160 26624
rect 15839 25536 15848 25600
rect 15912 25536 15928 25600
rect 15992 25536 16008 25600
rect 16072 25536 16088 25600
rect 16152 25536 16160 25600
rect 15839 24512 16160 25536
rect 15839 24448 15848 24512
rect 15912 24448 15928 24512
rect 15992 24448 16008 24512
rect 16072 24448 16088 24512
rect 16152 24448 16160 24512
rect 15839 23424 16160 24448
rect 15839 23360 15848 23424
rect 15912 23360 15928 23424
rect 15992 23360 16008 23424
rect 16072 23360 16088 23424
rect 16152 23360 16160 23424
rect 15839 22336 16160 23360
rect 17542 23221 17602 27371
rect 20805 27232 21125 28256
rect 20805 27168 20813 27232
rect 20877 27168 20893 27232
rect 20957 27168 20973 27232
rect 21037 27168 21053 27232
rect 21117 27168 21125 27232
rect 20805 26144 21125 27168
rect 20805 26080 20813 26144
rect 20877 26080 20893 26144
rect 20957 26080 20973 26144
rect 21037 26080 21053 26144
rect 21117 26080 21125 26144
rect 20805 25056 21125 26080
rect 20805 24992 20813 25056
rect 20877 24992 20893 25056
rect 20957 24992 20973 25056
rect 21037 24992 21053 25056
rect 21117 24992 21125 25056
rect 20805 23968 21125 24992
rect 20805 23904 20813 23968
rect 20877 23904 20893 23968
rect 20957 23904 20973 23968
rect 21037 23904 21053 23968
rect 21117 23904 21125 23968
rect 17539 23220 17605 23221
rect 17539 23156 17540 23220
rect 17604 23156 17605 23220
rect 17539 23155 17605 23156
rect 15839 22272 15848 22336
rect 15912 22272 15928 22336
rect 15992 22272 16008 22336
rect 16072 22272 16088 22336
rect 16152 22272 16160 22336
rect 15839 21248 16160 22272
rect 15839 21184 15848 21248
rect 15912 21184 15928 21248
rect 15992 21184 16008 21248
rect 16072 21184 16088 21248
rect 16152 21184 16160 21248
rect 15839 20160 16160 21184
rect 15839 20096 15848 20160
rect 15912 20096 15928 20160
rect 15992 20096 16008 20160
rect 16072 20096 16088 20160
rect 16152 20096 16160 20160
rect 11283 19140 11349 19141
rect 11283 19076 11284 19140
rect 11348 19076 11349 19140
rect 11283 19075 11349 19076
rect 10874 18464 10882 18528
rect 10946 18464 10962 18528
rect 11026 18464 11042 18528
rect 11106 18464 11122 18528
rect 11186 18464 11194 18528
rect 10874 17440 11194 18464
rect 10874 17376 10882 17440
rect 10946 17376 10962 17440
rect 11026 17376 11042 17440
rect 11106 17376 11122 17440
rect 11186 17376 11194 17440
rect 10179 17372 10245 17373
rect 10179 17308 10180 17372
rect 10244 17308 10245 17372
rect 10179 17307 10245 17308
rect 5909 16832 5917 16896
rect 5981 16832 5997 16896
rect 6061 16832 6077 16896
rect 6141 16832 6157 16896
rect 6221 16832 6229 16896
rect 5909 15808 6229 16832
rect 5909 15744 5917 15808
rect 5981 15744 5997 15808
rect 6061 15744 6077 15808
rect 6141 15744 6157 15808
rect 6221 15744 6229 15808
rect 5909 14720 6229 15744
rect 9075 15468 9141 15469
rect 9075 15404 9076 15468
rect 9140 15404 9141 15468
rect 9075 15403 9141 15404
rect 5909 14656 5917 14720
rect 5981 14656 5997 14720
rect 6061 14656 6077 14720
rect 6141 14656 6157 14720
rect 6221 14656 6229 14720
rect 5909 13632 6229 14656
rect 5909 13568 5917 13632
rect 5981 13568 5997 13632
rect 6061 13568 6077 13632
rect 6141 13568 6157 13632
rect 6221 13568 6229 13632
rect 5909 12544 6229 13568
rect 5909 12480 5917 12544
rect 5981 12480 5997 12544
rect 6061 12480 6077 12544
rect 6141 12480 6157 12544
rect 6221 12480 6229 12544
rect 5909 11456 6229 12480
rect 5909 11392 5917 11456
rect 5981 11392 5997 11456
rect 6061 11392 6077 11456
rect 6141 11392 6157 11456
rect 6221 11392 6229 11456
rect 5909 10368 6229 11392
rect 9078 11253 9138 15403
rect 10182 12069 10242 17307
rect 10874 16352 11194 17376
rect 10874 16288 10882 16352
rect 10946 16288 10962 16352
rect 11026 16288 11042 16352
rect 11106 16288 11122 16352
rect 11186 16288 11194 16352
rect 10874 15264 11194 16288
rect 10874 15200 10882 15264
rect 10946 15200 10962 15264
rect 11026 15200 11042 15264
rect 11106 15200 11122 15264
rect 11186 15200 11194 15264
rect 10874 14176 11194 15200
rect 10874 14112 10882 14176
rect 10946 14112 10962 14176
rect 11026 14112 11042 14176
rect 11106 14112 11122 14176
rect 11186 14112 11194 14176
rect 10874 13088 11194 14112
rect 10874 13024 10882 13088
rect 10946 13024 10962 13088
rect 11026 13024 11042 13088
rect 11106 13024 11122 13088
rect 11186 13024 11194 13088
rect 10179 12068 10245 12069
rect 10179 12004 10180 12068
rect 10244 12004 10245 12068
rect 10179 12003 10245 12004
rect 10874 12000 11194 13024
rect 10874 11936 10882 12000
rect 10946 11936 10962 12000
rect 11026 11936 11042 12000
rect 11106 11936 11122 12000
rect 11186 11936 11194 12000
rect 9075 11252 9141 11253
rect 9075 11188 9076 11252
rect 9140 11188 9141 11252
rect 9075 11187 9141 11188
rect 5909 10304 5917 10368
rect 5981 10304 5997 10368
rect 6061 10304 6077 10368
rect 6141 10304 6157 10368
rect 6221 10304 6229 10368
rect 5909 9280 6229 10304
rect 5909 9216 5917 9280
rect 5981 9216 5997 9280
rect 6061 9216 6077 9280
rect 6141 9216 6157 9280
rect 6221 9216 6229 9280
rect 5909 8192 6229 9216
rect 5909 8128 5917 8192
rect 5981 8128 5997 8192
rect 6061 8128 6077 8192
rect 6141 8128 6157 8192
rect 6221 8128 6229 8192
rect 5909 7104 6229 8128
rect 5909 7040 5917 7104
rect 5981 7040 5997 7104
rect 6061 7040 6077 7104
rect 6141 7040 6157 7104
rect 6221 7040 6229 7104
rect 5909 6016 6229 7040
rect 5909 5952 5917 6016
rect 5981 5952 5997 6016
rect 6061 5952 6077 6016
rect 6141 5952 6157 6016
rect 6221 5952 6229 6016
rect 5909 4928 6229 5952
rect 5909 4864 5917 4928
rect 5981 4864 5997 4928
rect 6061 4864 6077 4928
rect 6141 4864 6157 4928
rect 6221 4864 6229 4928
rect 5909 3840 6229 4864
rect 5909 3776 5917 3840
rect 5981 3776 5997 3840
rect 6061 3776 6077 3840
rect 6141 3776 6157 3840
rect 6221 3776 6229 3840
rect 5909 2752 6229 3776
rect 5909 2688 5917 2752
rect 5981 2688 5997 2752
rect 6061 2688 6077 2752
rect 6141 2688 6157 2752
rect 6221 2688 6229 2752
rect 5909 2128 6229 2688
rect 10874 10912 11194 11936
rect 10874 10848 10882 10912
rect 10946 10848 10962 10912
rect 11026 10848 11042 10912
rect 11106 10848 11122 10912
rect 11186 10848 11194 10912
rect 10874 9824 11194 10848
rect 10874 9760 10882 9824
rect 10946 9760 10962 9824
rect 11026 9760 11042 9824
rect 11106 9760 11122 9824
rect 11186 9760 11194 9824
rect 10874 8736 11194 9760
rect 10874 8672 10882 8736
rect 10946 8672 10962 8736
rect 11026 8672 11042 8736
rect 11106 8672 11122 8736
rect 11186 8672 11194 8736
rect 10874 7648 11194 8672
rect 10874 7584 10882 7648
rect 10946 7584 10962 7648
rect 11026 7584 11042 7648
rect 11106 7584 11122 7648
rect 11186 7584 11194 7648
rect 10874 6560 11194 7584
rect 10874 6496 10882 6560
rect 10946 6496 10962 6560
rect 11026 6496 11042 6560
rect 11106 6496 11122 6560
rect 11186 6496 11194 6560
rect 10874 5472 11194 6496
rect 10874 5408 10882 5472
rect 10946 5408 10962 5472
rect 11026 5408 11042 5472
rect 11106 5408 11122 5472
rect 11186 5408 11194 5472
rect 10874 4384 11194 5408
rect 10874 4320 10882 4384
rect 10946 4320 10962 4384
rect 11026 4320 11042 4384
rect 11106 4320 11122 4384
rect 11186 4320 11194 4384
rect 10874 3296 11194 4320
rect 10874 3232 10882 3296
rect 10946 3232 10962 3296
rect 11026 3232 11042 3296
rect 11106 3232 11122 3296
rect 11186 3232 11194 3296
rect 10874 2208 11194 3232
rect 10874 2144 10882 2208
rect 10946 2144 10962 2208
rect 11026 2144 11042 2208
rect 11106 2144 11122 2208
rect 11186 2144 11194 2208
rect 10874 2128 11194 2144
rect 15839 19072 16160 20096
rect 15839 19008 15848 19072
rect 15912 19008 15928 19072
rect 15992 19008 16008 19072
rect 16072 19008 16088 19072
rect 16152 19008 16160 19072
rect 15839 17984 16160 19008
rect 15839 17920 15848 17984
rect 15912 17920 15928 17984
rect 15992 17920 16008 17984
rect 16072 17920 16088 17984
rect 16152 17920 16160 17984
rect 15839 16896 16160 17920
rect 15839 16832 15848 16896
rect 15912 16832 15928 16896
rect 15992 16832 16008 16896
rect 16072 16832 16088 16896
rect 16152 16832 16160 16896
rect 15839 15808 16160 16832
rect 15839 15744 15848 15808
rect 15912 15744 15928 15808
rect 15992 15744 16008 15808
rect 16072 15744 16088 15808
rect 16152 15744 16160 15808
rect 15839 14720 16160 15744
rect 15839 14656 15848 14720
rect 15912 14656 15928 14720
rect 15992 14656 16008 14720
rect 16072 14656 16088 14720
rect 16152 14656 16160 14720
rect 15839 13632 16160 14656
rect 15839 13568 15848 13632
rect 15912 13568 15928 13632
rect 15992 13568 16008 13632
rect 16072 13568 16088 13632
rect 16152 13568 16160 13632
rect 15839 12544 16160 13568
rect 15839 12480 15848 12544
rect 15912 12480 15928 12544
rect 15992 12480 16008 12544
rect 16072 12480 16088 12544
rect 16152 12480 16160 12544
rect 15839 11456 16160 12480
rect 15839 11392 15848 11456
rect 15912 11392 15928 11456
rect 15992 11392 16008 11456
rect 16072 11392 16088 11456
rect 16152 11392 16160 11456
rect 15839 10368 16160 11392
rect 15839 10304 15848 10368
rect 15912 10304 15928 10368
rect 15992 10304 16008 10368
rect 16072 10304 16088 10368
rect 16152 10304 16160 10368
rect 15839 9280 16160 10304
rect 15839 9216 15848 9280
rect 15912 9216 15928 9280
rect 15992 9216 16008 9280
rect 16072 9216 16088 9280
rect 16152 9216 16160 9280
rect 15839 8192 16160 9216
rect 15839 8128 15848 8192
rect 15912 8128 15928 8192
rect 15992 8128 16008 8192
rect 16072 8128 16088 8192
rect 16152 8128 16160 8192
rect 15839 7104 16160 8128
rect 15839 7040 15848 7104
rect 15912 7040 15928 7104
rect 15992 7040 16008 7104
rect 16072 7040 16088 7104
rect 16152 7040 16160 7104
rect 15839 6016 16160 7040
rect 15839 5952 15848 6016
rect 15912 5952 15928 6016
rect 15992 5952 16008 6016
rect 16072 5952 16088 6016
rect 16152 5952 16160 6016
rect 15839 4928 16160 5952
rect 15839 4864 15848 4928
rect 15912 4864 15928 4928
rect 15992 4864 16008 4928
rect 16072 4864 16088 4928
rect 16152 4864 16160 4928
rect 15839 3840 16160 4864
rect 15839 3776 15848 3840
rect 15912 3776 15928 3840
rect 15992 3776 16008 3840
rect 16072 3776 16088 3840
rect 16152 3776 16160 3840
rect 15839 2752 16160 3776
rect 15839 2688 15848 2752
rect 15912 2688 15928 2752
rect 15992 2688 16008 2752
rect 16072 2688 16088 2752
rect 16152 2688 16160 2752
rect 15839 2128 16160 2688
rect 20805 22880 21125 23904
rect 20805 22816 20813 22880
rect 20877 22816 20893 22880
rect 20957 22816 20973 22880
rect 21037 22816 21053 22880
rect 21117 22816 21125 22880
rect 20805 21792 21125 22816
rect 20805 21728 20813 21792
rect 20877 21728 20893 21792
rect 20957 21728 20973 21792
rect 21037 21728 21053 21792
rect 21117 21728 21125 21792
rect 20805 20704 21125 21728
rect 20805 20640 20813 20704
rect 20877 20640 20893 20704
rect 20957 20640 20973 20704
rect 21037 20640 21053 20704
rect 21117 20640 21125 20704
rect 20805 19616 21125 20640
rect 20805 19552 20813 19616
rect 20877 19552 20893 19616
rect 20957 19552 20973 19616
rect 21037 19552 21053 19616
rect 21117 19552 21125 19616
rect 20805 18528 21125 19552
rect 20805 18464 20813 18528
rect 20877 18464 20893 18528
rect 20957 18464 20973 18528
rect 21037 18464 21053 18528
rect 21117 18464 21125 18528
rect 20805 17440 21125 18464
rect 20805 17376 20813 17440
rect 20877 17376 20893 17440
rect 20957 17376 20973 17440
rect 21037 17376 21053 17440
rect 21117 17376 21125 17440
rect 20805 16352 21125 17376
rect 20805 16288 20813 16352
rect 20877 16288 20893 16352
rect 20957 16288 20973 16352
rect 21037 16288 21053 16352
rect 21117 16288 21125 16352
rect 20805 15264 21125 16288
rect 20805 15200 20813 15264
rect 20877 15200 20893 15264
rect 20957 15200 20973 15264
rect 21037 15200 21053 15264
rect 21117 15200 21125 15264
rect 20805 14176 21125 15200
rect 20805 14112 20813 14176
rect 20877 14112 20893 14176
rect 20957 14112 20973 14176
rect 21037 14112 21053 14176
rect 21117 14112 21125 14176
rect 20805 13088 21125 14112
rect 20805 13024 20813 13088
rect 20877 13024 20893 13088
rect 20957 13024 20973 13088
rect 21037 13024 21053 13088
rect 21117 13024 21125 13088
rect 20805 12000 21125 13024
rect 20805 11936 20813 12000
rect 20877 11936 20893 12000
rect 20957 11936 20973 12000
rect 21037 11936 21053 12000
rect 21117 11936 21125 12000
rect 20805 10912 21125 11936
rect 20805 10848 20813 10912
rect 20877 10848 20893 10912
rect 20957 10848 20973 10912
rect 21037 10848 21053 10912
rect 21117 10848 21125 10912
rect 20805 9824 21125 10848
rect 20805 9760 20813 9824
rect 20877 9760 20893 9824
rect 20957 9760 20973 9824
rect 21037 9760 21053 9824
rect 21117 9760 21125 9824
rect 20805 8736 21125 9760
rect 20805 8672 20813 8736
rect 20877 8672 20893 8736
rect 20957 8672 20973 8736
rect 21037 8672 21053 8736
rect 21117 8672 21125 8736
rect 20805 7648 21125 8672
rect 20805 7584 20813 7648
rect 20877 7584 20893 7648
rect 20957 7584 20973 7648
rect 21037 7584 21053 7648
rect 21117 7584 21125 7648
rect 20805 6560 21125 7584
rect 20805 6496 20813 6560
rect 20877 6496 20893 6560
rect 20957 6496 20973 6560
rect 21037 6496 21053 6560
rect 21117 6496 21125 6560
rect 20805 5472 21125 6496
rect 20805 5408 20813 5472
rect 20877 5408 20893 5472
rect 20957 5408 20973 5472
rect 21037 5408 21053 5472
rect 21117 5408 21125 5472
rect 20805 4384 21125 5408
rect 20805 4320 20813 4384
rect 20877 4320 20893 4384
rect 20957 4320 20973 4384
rect 21037 4320 21053 4384
rect 21117 4320 21125 4384
rect 20805 3296 21125 4320
rect 20805 3232 20813 3296
rect 20877 3232 20893 3296
rect 20957 3232 20973 3296
rect 21037 3232 21053 3296
rect 21117 3232 21125 3296
rect 20805 2208 21125 3232
rect 20805 2144 20813 2208
rect 20877 2144 20893 2208
rect 20957 2144 20973 2208
rect 21037 2144 21053 2208
rect 21117 2144 21125 2208
rect 20805 2128 21125 2144
rect 25770 45184 26090 45744
rect 25770 45120 25778 45184
rect 25842 45120 25858 45184
rect 25922 45120 25938 45184
rect 26002 45120 26018 45184
rect 26082 45120 26090 45184
rect 25770 44096 26090 45120
rect 25770 44032 25778 44096
rect 25842 44032 25858 44096
rect 25922 44032 25938 44096
rect 26002 44032 26018 44096
rect 26082 44032 26090 44096
rect 25770 43008 26090 44032
rect 25770 42944 25778 43008
rect 25842 42944 25858 43008
rect 25922 42944 25938 43008
rect 26002 42944 26018 43008
rect 26082 42944 26090 43008
rect 25770 41920 26090 42944
rect 25770 41856 25778 41920
rect 25842 41856 25858 41920
rect 25922 41856 25938 41920
rect 26002 41856 26018 41920
rect 26082 41856 26090 41920
rect 25770 40832 26090 41856
rect 25770 40768 25778 40832
rect 25842 40768 25858 40832
rect 25922 40768 25938 40832
rect 26002 40768 26018 40832
rect 26082 40768 26090 40832
rect 25770 39744 26090 40768
rect 25770 39680 25778 39744
rect 25842 39680 25858 39744
rect 25922 39680 25938 39744
rect 26002 39680 26018 39744
rect 26082 39680 26090 39744
rect 25770 38656 26090 39680
rect 25770 38592 25778 38656
rect 25842 38592 25858 38656
rect 25922 38592 25938 38656
rect 26002 38592 26018 38656
rect 26082 38592 26090 38656
rect 25770 37568 26090 38592
rect 25770 37504 25778 37568
rect 25842 37504 25858 37568
rect 25922 37504 25938 37568
rect 26002 37504 26018 37568
rect 26082 37504 26090 37568
rect 25770 36480 26090 37504
rect 25770 36416 25778 36480
rect 25842 36416 25858 36480
rect 25922 36416 25938 36480
rect 26002 36416 26018 36480
rect 26082 36416 26090 36480
rect 25770 35392 26090 36416
rect 25770 35328 25778 35392
rect 25842 35328 25858 35392
rect 25922 35328 25938 35392
rect 26002 35328 26018 35392
rect 26082 35328 26090 35392
rect 25770 34304 26090 35328
rect 25770 34240 25778 34304
rect 25842 34240 25858 34304
rect 25922 34240 25938 34304
rect 26002 34240 26018 34304
rect 26082 34240 26090 34304
rect 25770 33216 26090 34240
rect 25770 33152 25778 33216
rect 25842 33152 25858 33216
rect 25922 33152 25938 33216
rect 26002 33152 26018 33216
rect 26082 33152 26090 33216
rect 25770 32128 26090 33152
rect 25770 32064 25778 32128
rect 25842 32064 25858 32128
rect 25922 32064 25938 32128
rect 26002 32064 26018 32128
rect 26082 32064 26090 32128
rect 25770 31040 26090 32064
rect 25770 30976 25778 31040
rect 25842 30976 25858 31040
rect 25922 30976 25938 31040
rect 26002 30976 26018 31040
rect 26082 30976 26090 31040
rect 25770 29952 26090 30976
rect 25770 29888 25778 29952
rect 25842 29888 25858 29952
rect 25922 29888 25938 29952
rect 26002 29888 26018 29952
rect 26082 29888 26090 29952
rect 25770 28864 26090 29888
rect 25770 28800 25778 28864
rect 25842 28800 25858 28864
rect 25922 28800 25938 28864
rect 26002 28800 26018 28864
rect 26082 28800 26090 28864
rect 25770 27776 26090 28800
rect 25770 27712 25778 27776
rect 25842 27712 25858 27776
rect 25922 27712 25938 27776
rect 26002 27712 26018 27776
rect 26082 27712 26090 27776
rect 25770 26688 26090 27712
rect 25770 26624 25778 26688
rect 25842 26624 25858 26688
rect 25922 26624 25938 26688
rect 26002 26624 26018 26688
rect 26082 26624 26090 26688
rect 25770 25600 26090 26624
rect 25770 25536 25778 25600
rect 25842 25536 25858 25600
rect 25922 25536 25938 25600
rect 26002 25536 26018 25600
rect 26082 25536 26090 25600
rect 25770 24512 26090 25536
rect 25770 24448 25778 24512
rect 25842 24448 25858 24512
rect 25922 24448 25938 24512
rect 26002 24448 26018 24512
rect 26082 24448 26090 24512
rect 25770 23424 26090 24448
rect 25770 23360 25778 23424
rect 25842 23360 25858 23424
rect 25922 23360 25938 23424
rect 26002 23360 26018 23424
rect 26082 23360 26090 23424
rect 25770 22336 26090 23360
rect 25770 22272 25778 22336
rect 25842 22272 25858 22336
rect 25922 22272 25938 22336
rect 26002 22272 26018 22336
rect 26082 22272 26090 22336
rect 25770 21248 26090 22272
rect 25770 21184 25778 21248
rect 25842 21184 25858 21248
rect 25922 21184 25938 21248
rect 26002 21184 26018 21248
rect 26082 21184 26090 21248
rect 25770 20160 26090 21184
rect 25770 20096 25778 20160
rect 25842 20096 25858 20160
rect 25922 20096 25938 20160
rect 26002 20096 26018 20160
rect 26082 20096 26090 20160
rect 25770 19072 26090 20096
rect 25770 19008 25778 19072
rect 25842 19008 25858 19072
rect 25922 19008 25938 19072
rect 26002 19008 26018 19072
rect 26082 19008 26090 19072
rect 25770 17984 26090 19008
rect 25770 17920 25778 17984
rect 25842 17920 25858 17984
rect 25922 17920 25938 17984
rect 26002 17920 26018 17984
rect 26082 17920 26090 17984
rect 25770 16896 26090 17920
rect 25770 16832 25778 16896
rect 25842 16832 25858 16896
rect 25922 16832 25938 16896
rect 26002 16832 26018 16896
rect 26082 16832 26090 16896
rect 25770 15808 26090 16832
rect 25770 15744 25778 15808
rect 25842 15744 25858 15808
rect 25922 15744 25938 15808
rect 26002 15744 26018 15808
rect 26082 15744 26090 15808
rect 25770 14720 26090 15744
rect 25770 14656 25778 14720
rect 25842 14656 25858 14720
rect 25922 14656 25938 14720
rect 26002 14656 26018 14720
rect 26082 14656 26090 14720
rect 25770 13632 26090 14656
rect 25770 13568 25778 13632
rect 25842 13568 25858 13632
rect 25922 13568 25938 13632
rect 26002 13568 26018 13632
rect 26082 13568 26090 13632
rect 25770 12544 26090 13568
rect 25770 12480 25778 12544
rect 25842 12480 25858 12544
rect 25922 12480 25938 12544
rect 26002 12480 26018 12544
rect 26082 12480 26090 12544
rect 25770 11456 26090 12480
rect 25770 11392 25778 11456
rect 25842 11392 25858 11456
rect 25922 11392 25938 11456
rect 26002 11392 26018 11456
rect 26082 11392 26090 11456
rect 25770 10368 26090 11392
rect 25770 10304 25778 10368
rect 25842 10304 25858 10368
rect 25922 10304 25938 10368
rect 26002 10304 26018 10368
rect 26082 10304 26090 10368
rect 25770 9280 26090 10304
rect 25770 9216 25778 9280
rect 25842 9216 25858 9280
rect 25922 9216 25938 9280
rect 26002 9216 26018 9280
rect 26082 9216 26090 9280
rect 25770 8192 26090 9216
rect 25770 8128 25778 8192
rect 25842 8128 25858 8192
rect 25922 8128 25938 8192
rect 26002 8128 26018 8192
rect 26082 8128 26090 8192
rect 25770 7104 26090 8128
rect 25770 7040 25778 7104
rect 25842 7040 25858 7104
rect 25922 7040 25938 7104
rect 26002 7040 26018 7104
rect 26082 7040 26090 7104
rect 25770 6016 26090 7040
rect 25770 5952 25778 6016
rect 25842 5952 25858 6016
rect 25922 5952 25938 6016
rect 26002 5952 26018 6016
rect 26082 5952 26090 6016
rect 25770 4928 26090 5952
rect 25770 4864 25778 4928
rect 25842 4864 25858 4928
rect 25922 4864 25938 4928
rect 26002 4864 26018 4928
rect 26082 4864 26090 4928
rect 25770 3840 26090 4864
rect 25770 3776 25778 3840
rect 25842 3776 25858 3840
rect 25922 3776 25938 3840
rect 26002 3776 26018 3840
rect 26082 3776 26090 3840
rect 25770 2752 26090 3776
rect 25770 2688 25778 2752
rect 25842 2688 25858 2752
rect 25922 2688 25938 2752
rect 26002 2688 26018 2752
rect 26082 2688 26090 2752
rect 25770 2128 26090 2688
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1635444444
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1635444444
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1635444444
transform 1 0 2668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1635444444
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input67
timestamp 1635444444
transform 1 0 4048 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1635444444
transform -1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_30
timestamp 1635444444
transform 1 0 3864 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_23
timestamp 1635444444
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp 1635444444
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22
timestamp 1635444444
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 4968 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1635444444
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1893_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 4416 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1635444444
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6624 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1635444444
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1635444444
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1635444444
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1635444444
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1635444444
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1635444444
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1635444444
transform -1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635444444
transform -1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_70
timestamp 1635444444
transform 1 0 7544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68
timestamp 1635444444
transform 1 0 7360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1635444444
transform -1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1635444444
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_77
timestamp 1635444444
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1635444444
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1635444444
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_84
timestamp 1635444444
transform 1 0 8832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1635444444
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102
timestamp 1635444444
transform 1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1635444444
transform 1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_104
timestamp 1635444444
transform 1 0 10672 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1635444444
transform 1 0 9200 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1635444444
transform 1 0 9568 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1635444444
transform 1 0 11500 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 12052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1635444444
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1635444444
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1635444444
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1635444444
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1015_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 13156 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_123
timestamp 1635444444
transform 1 0 12420 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123
timestamp 1635444444
transform 1 0 12420 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_131
timestamp 1635444444
transform 1 0 13156 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1635444444
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1635444444
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_147
timestamp 1635444444
transform 1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_146
timestamp 1635444444
transform 1 0 14536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1635444444
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1087_
timestamp 1635444444
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1258_
timestamp 1635444444
transform -1 0 15456 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1515_
timestamp 1635444444
transform 1 0 14996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1750_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 14536 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1635444444
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_157
timestamp 1635444444
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1635444444
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1635444444
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1635444444
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_160
timestamp 1635444444
transform 1 0 15824 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1635444444
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1518_
timestamp 1635444444
transform -1 0 17204 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1259_
timestamp 1635444444
transform -1 0 17388 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1635444444
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1635444444
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1635444444
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1757_
timestamp 1635444444
transform 1 0 17756 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1519_
timestamp 1635444444
transform 1 0 17572 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_177
timestamp 1635444444
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1635444444
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1635444444
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1520_
timestamp 1635444444
transform -1 0 19504 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_190
timestamp 1635444444
transform 1 0 18584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1635444444
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_185
timestamp 1635444444
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1635444444
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_200
timestamp 1635444444
transform 1 0 19504 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_211
timestamp 1635444444
transform 1 0 20516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_200
timestamp 1635444444
transform 1 0 19504 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_208
timestamp 1635444444
transform 1 0 20240 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1635444444
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1009_
timestamp 1635444444
transform 1 0 20424 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1013_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 21344 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1257_
timestamp 1635444444
transform -1 0 20516 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1635444444
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1014_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 22264 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 22540 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1635444444
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1635444444
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1635444444
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1635444444
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_233
timestamp 1635444444
transform 1 0 22540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1635444444
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1635444444
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1635444444
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1635444444
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244
timestamp 1635444444
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_256
timestamp 1635444444
transform 1 0 24656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_247 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 23828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_259
timestamp 1635444444
transform 1 0 24932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1635444444
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1635444444
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1635444444
transform 1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1635444444
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1635444444
transform 1 0 25024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1635444444
transform 1 0 25668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_270
timestamp 1635444444
transform 1 0 25944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_263
timestamp 1635444444
transform 1 0 25300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1635444444
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_271
timestamp 1635444444
transform 1 0 26036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1635444444
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1635444444
transform -1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1635444444
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1635444444
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1635444444
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1635444444
transform 1 0 27600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 1635444444
transform -1 0 27876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_291
timestamp 1635444444
transform 1 0 27876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_291
timestamp 1635444444
transform 1 0 27876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_284
timestamp 1635444444
transform 1 0 27232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 28704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1012_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 28244 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_1_300
timestamp 1635444444
transform 1 0 28704 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_299
timestamp 1635444444
transform 1 0 28612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1635444444
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_309
timestamp 1635444444
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_316
timestamp 1635444444
transform 1 0 30176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_306
timestamp 1635444444
transform 1 0 29256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_316
timestamp 1635444444
transform 1 0 30176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635444444
transform -1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635444444
transform -1 0 30820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1635444444
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__or4bb_1  _1010_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 30176 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1635444444
transform 1 0 29808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1635444444
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1635444444
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635444444
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0881_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2760 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1635444444
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1635444444
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1635444444
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1635444444
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_40
timestamp 1635444444
transform 1 0 4784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1635444444
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input82
timestamp 1635444444
transform 1 0 4232 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 1635444444
transform 1 0 5152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_61
timestamp 1635444444
transform 1 0 6716 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1635444444
transform 1 0 5244 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp 1635444444
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1635444444
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1635444444
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1635444444
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1635444444
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1635444444
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1635444444
transform 1 0 9384 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1635444444
transform 1 0 11684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1016_
timestamp 1635444444
transform 1 0 11224 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _1372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 12052 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1635444444
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_151
timestamp 1635444444
transform 1 0 14996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1635444444
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1512_
timestamp 1635444444
transform 1 0 14076 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1635444444
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1753_
timestamp 1635444444
transform 1 0 15548 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1755_
timestamp 1635444444
transform 1 0 16744 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1635444444
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1635444444
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1635444444
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1756_
timestamp 1635444444
transform 1 0 17940 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_213
timestamp 1635444444
transform 1 0 20700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1256_
timestamp 1635444444
transform -1 0 21804 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1635444444
transform -1 0 20700 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_225
timestamp 1635444444
transform 1 0 21804 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_232
timestamp 1635444444
transform 1 0 22448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1635444444
transform 1 0 23092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1635444444
transform 1 0 22172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1635444444
transform 1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1635444444
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1635444444
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1635444444
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1635444444
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1635444444
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_289
timestamp 1635444444
transform 1 0 27692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1635444444
transform 1 0 28152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1635444444
transform 1 0 28520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1635444444
transform 1 0 28888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1635444444
transform 1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1635444444
transform 1 0 28612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_312
timestamp 1635444444
transform 1 0 29808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635444444
transform -1 0 30820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1635444444
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1635444444
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1635444444
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1635444444
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635444444
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1635444444
transform 1 0 1748 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1635444444
transform 1 0 2668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_23
timestamp 1635444444
transform 1 0 3220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_30
timestamp 1635444444
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _1174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 5796 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1635444444
transform -1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1635444444
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1635444444
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1635444444
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1176_
timestamp 1635444444
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_66
timestamp 1635444444
transform 1 0 7176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1635444444
transform 1 0 8280 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1635444444
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 1635444444
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1077_
timestamp 1635444444
transform 1 0 10120 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1635444444
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_119
timestamp 1635444444
transform 1 0 12052 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1635444444
transform 1 0 12788 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1635444444
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 12052 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1501_
timestamp 1635444444
transform -1 0 13892 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1635444444
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1513_
timestamp 1635444444
transform 1 0 14260 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1635444444
transform 1 0 15180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1635444444
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1635444444
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1635444444
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1516_
timestamp 1635444444
transform 1 0 15548 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1754_
timestamp 1635444444
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_178
timestamp 1635444444
transform 1 0 17480 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_186
timestamp 1635444444
transform 1 0 18216 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1635444444
transform -1 0 19780 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_203
timestamp 1635444444
transform 1 0 19780 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1635444444
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1101_
timestamp 1635444444
transform 1 0 20148 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_228
timestamp 1635444444
transform 1 0 22080 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_240
timestamp 1635444444
transform 1 0 23184 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1635444444
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1635444444
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_252
timestamp 1635444444
transform 1 0 24288 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_264
timestamp 1635444444
transform 1 0 25392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1635444444
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1635444444
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1635444444
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1635444444
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_305
timestamp 1635444444
transform 1 0 29164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_309
timestamp 1635444444
transform 1 0 29532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_316
timestamp 1635444444
transform 1 0 30176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635444444
transform -1 0 30820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1635444444
transform 1 0 29900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1635444444
transform -1 0 29532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_13
timestamp 1635444444
transform 1 0 2300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635444444
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1635444444
transform 1 0 1380 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1635444444
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1635444444
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1635444444
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1635444444
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_45
timestamp 1635444444
transform 1 0 5244 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_55
timestamp 1635444444
transform 1 0 6164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1177_
timestamp 1635444444
transform -1 0 6164 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1635444444
transform -1 0 8004 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp 1635444444
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1635444444
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1635444444
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1076_
timestamp 1635444444
transform 1 0 8924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_102
timestamp 1635444444
transform 1 0 10488 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_106
timestamp 1635444444
transform 1 0 10856 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_94
timestamp 1635444444
transform 1 0 9752 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1635444444
transform 1 0 10580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_115
timestamp 1635444444
transform 1 0 11684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_125
timestamp 1635444444
transform 1 0 12604 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_131
timestamp 1635444444
transform 1 0 13156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_1  _1086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 12604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1261_
timestamp 1635444444
transform -1 0 11684 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1635444444
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_150
timestamp 1635444444
transform 1 0 14904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1635444444
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1502_
timestamp 1635444444
transform 1 0 13248 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1751_
timestamp 1635444444
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_163
timestamp 1635444444
transform 1 0 16100 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_173
timestamp 1635444444
transform 1 0 17020 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1517_
timestamp 1635444444
transform 1 0 16468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1752_
timestamp 1635444444
transform 1 0 15272 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_181
timestamp 1635444444
transform 1 0 17756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1635444444
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1635444444
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1102_
timestamp 1635444444
transform 1 0 17940 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_200
timestamp 1635444444
transform 1 0 19504 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_213
timestamp 1635444444
transform 1 0 20700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _1100_
timestamp 1635444444
transform 1 0 19872 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1690_
timestamp 1635444444
transform -1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_225
timestamp 1635444444
transform 1 0 21804 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_237
timestamp 1635444444
transform 1 0 22908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1635444444
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1635444444
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1635444444
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1635444444
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1635444444
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1635444444
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1635444444
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1635444444
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp 1635444444
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_316
timestamp 1635444444
transform 1 0 30176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635444444
transform -1 0 30820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1635444444
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1635444444
transform 1 0 29900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_13
timestamp 1635444444
transform 1 0 2300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635444444
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1635444444
transform 1 0 1380 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_5_25
timestamp 1635444444
transform 1 0 3404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_43
timestamp 1635444444
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1635444444
transform 1 0 3588 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1635444444
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1635444444
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_2  _1694_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6348 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_5_67
timestamp 1635444444
transform 1 0 7268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _1078_
timestamp 1635444444
transform 1 0 8372 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_100
timestamp 1635444444
transform 1 0 10304 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_104
timestamp 1635444444
transform 1 0 10672 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1635444444
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_88
timestamp 1635444444
transform 1 0 9200 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1635444444
transform -1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_119
timestamp 1635444444
transform 1 0 12052 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1635444444
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1504_
timestamp 1635444444
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1510_
timestamp 1635444444
transform -1 0 13340 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_133
timestamp 1635444444
transform 1 0 13340 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_140
timestamp 1635444444
transform 1 0 13984 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1635444444
transform 1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1109_
timestamp 1635444444
transform -1 0 15732 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1635444444
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_159
timestamp 1635444444
transform 1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1635444444
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_172
timestamp 1635444444
transform 1 0 16928 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1635444444
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1635444444
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_180
timestamp 1635444444
transform 1 0 17664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_187
timestamp 1635444444
transform 1 0 18308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1521_
timestamp 1635444444
transform -1 0 18308 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_199
timestamp 1635444444
transform 1 0 19412 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_203
timestamp 1635444444
transform 1 0 19780 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1937_
timestamp 1635444444
transform -1 0 21344 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1635444444
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1635444444
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1635444444
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1635444444
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1635444444
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1635444444
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1635444444
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1635444444
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1635444444
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1635444444
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1635444444
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_305
timestamp 1635444444
transform 1 0 29164 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_311
timestamp 1635444444
transform 1 0 29716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_316
timestamp 1635444444
transform 1 0 30176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635444444
transform -1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1635444444
transform 1 0 29808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1635444444
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1635444444
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_20
timestamp 1635444444
transform 1 0 2944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1635444444
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635444444
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635444444
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1635444444
transform 1 0 1840 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1635444444
transform 1 0 1472 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1635444444
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1635444444
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_33
timestamp 1635444444
transform 1 0 4140 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_41
timestamp 1635444444
transform 1 0 4876 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1635444444
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1164_
timestamp 1635444444
transform 1 0 3312 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_2  _1662_
timestamp 1635444444
transform -1 0 5888 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1635444444
transform 1 0 4140 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_49
timestamp 1635444444
transform 1 0 5612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_63
timestamp 1635444444
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1635444444
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1635444444
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1168_
timestamp 1635444444
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_2  _1673_
timestamp 1635444444
transform -1 0 6900 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1635444444
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1635444444
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1635444444
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_66
timestamp 1635444444
transform 1 0 7176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_86
timestamp 1635444444
transform 1 0 9016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1635444444
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1946_
timestamp 1635444444
transform 1 0 7544 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1635444444
transform 1 0 9660 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1635444444
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1079_
timestamp 1635444444
transform -1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1743_
timestamp 1635444444
transform 1 0 10764 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _1821_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 11040 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_6_114
timestamp 1635444444
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 1635444444
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_125
timestamp 1635444444
transform 1 0 12604 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1635444444
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_128
timestamp 1635444444
transform 1 0 12880 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1635444444
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1376_
timestamp 1635444444
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1747_
timestamp 1635444444
transform -1 0 12880 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1748_
timestamp 1635444444
transform -1 0 13524 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1635444444
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1635444444
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_151
timestamp 1635444444
transform 1 0 14996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_138
timestamp 1635444444
transform 1 0 13800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_142
timestamp 1635444444
transform 1 0 14168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1635444444
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1503_
timestamp 1635444444
transform 1 0 14076 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1509_
timestamp 1635444444
transform 1 0 13248 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1635444444
transform 1 0 14260 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_173
timestamp 1635444444
transform 1 0 17020 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_159
timestamp 1635444444
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1635444444
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1635444444
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1635444444
transform 1 0 15548 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1635444444
transform -1 0 18124 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_6_177
timestamp 1635444444
transform 1 0 17388 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_187
timestamp 1635444444
transform 1 0 18308 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1635444444
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_185
timestamp 1635444444
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_193
timestamp 1635444444
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1635444444
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1085_
timestamp 1635444444
transform -1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1104_
timestamp 1635444444
transform 1 0 17480 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_201
timestamp 1635444444
transform 1 0 19596 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_214
timestamp 1635444444
transform 1 0 20792 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_211
timestamp 1635444444
transform 1 0 20516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1091_
timestamp 1635444444
transform 1 0 19596 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1098_
timestamp 1635444444
transform 1 0 19964 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1099_
timestamp 1635444444
transform -1 0 19596 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_226
timestamp 1635444444
transform 1 0 21896 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_238
timestamp 1635444444
transform 1 0 23000 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1635444444
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1635444444
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1635444444
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1635444444
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1635444444
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1635444444
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1635444444
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1635444444
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1635444444
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1635444444
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1635444444
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1635444444
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1635444444
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1635444444
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1635444444
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1635444444
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1635444444
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1635444444
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1635444444
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1635444444
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1635444444
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_317
timestamp 1635444444
transform 1 0 30268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_317
timestamp 1635444444
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635444444
transform -1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635444444
transform -1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1635444444
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1635444444
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1635444444
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635444444
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1161_
timestamp 1635444444
transform 1 0 1380 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1635444444
transform -1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1635444444
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_38
timestamp 1635444444
transform 1 0 4600 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1635444444
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1166_
timestamp 1635444444
transform -1 0 4600 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1167_
timestamp 1635444444
transform -1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_46
timestamp 1635444444
transform 1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1635444444
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_2  _1647_
timestamp 1635444444
transform -1 0 6624 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1635444444
transform -1 0 8464 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1635444444
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1635444444
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1635444444
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_101
timestamp 1635444444
transform 1 0 10396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_109
timestamp 1635444444
transform 1 0 11132 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1073_
timestamp 1635444444
transform -1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1074_
timestamp 1635444444
transform -1 0 10396 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_8_121
timestamp 1635444444
transform 1 0 12236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1508_
timestamp 1635444444
transform 1 0 11684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1749_
timestamp 1635444444
transform 1 0 12788 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1635444444
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1635444444
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1635444444
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1108_
timestamp 1635444444
transform -1 0 15364 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_8_155
timestamp 1635444444
transform 1 0 15364 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_162
timestamp 1635444444
transform 1 0 16008 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_166
timestamp 1635444444
transform 1 0 16376 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1107_
timestamp 1635444444
transform 1 0 16468 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1635444444
transform 1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_176
timestamp 1635444444
transform 1 0 17296 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_180
timestamp 1635444444
transform 1 0 17664 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_185
timestamp 1635444444
transform 1 0 18124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1635444444
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1635444444
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1072_
timestamp 1635444444
transform 1 0 17756 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1635444444
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_202
timestamp 1635444444
transform 1 0 19688 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1713_
timestamp 1635444444
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1938_
timestamp 1635444444
transform 1 0 20056 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_222
timestamp 1635444444
transform 1 0 21528 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_234
timestamp 1635444444
transform 1 0 22632 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1635444444
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1635444444
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1635444444
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1635444444
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1635444444
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1635444444
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1635444444
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1635444444
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_309
timestamp 1635444444
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_317
timestamp 1635444444
transform 1 0 30268 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635444444
transform -1 0 30820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1635444444
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_13
timestamp 1635444444
transform 1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_17
timestamp 1635444444
transform 1 0 2668 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_6
timestamp 1635444444
transform 1 0 1656 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635444444
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1155_
timestamp 1635444444
transform -1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1635444444
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1635444444
transform -1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_22
timestamp 1635444444
transform 1 0 3128 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_38
timestamp 1635444444
transform 1 0 4600 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1159_
timestamp 1635444444
transform -1 0 4600 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_9_46
timestamp 1635444444
transform 1 0 5336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1635444444
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_60
timestamp 1635444444
transform 1 0 6624 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1635444444
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1635444444
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1171_
timestamp 1635444444
transform 1 0 5520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1178_
timestamp 1635444444
transform 1 0 6992 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_73
timestamp 1635444444
transform 1 0 7820 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_79
timestamp 1635444444
transform 1 0 8372 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1080_
timestamp 1635444444
transform 1 0 8464 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1635444444
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_89
timestamp 1635444444
transform 1 0 9292 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_97
timestamp 1635444444
transform 1 0 10028 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1255_
timestamp 1635444444
transform -1 0 10580 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1635444444
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_116
timestamp 1635444444
transform 1 0 11776 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_125
timestamp 1635444444
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1635444444
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _1254_
timestamp 1635444444
transform -1 0 12604 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1506_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1511_
timestamp 1635444444
transform 1 0 12972 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_135
timestamp 1635444444
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_139
timestamp 1635444444
transform 1 0 13892 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_149
timestamp 1635444444
transform 1 0 14812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1114_
timestamp 1635444444
transform 1 0 13984 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1635444444
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1635444444
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1635444444
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1111_
timestamp 1635444444
transform 1 0 15180 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_179
timestamp 1635444444
transform 1 0 17572 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1097_
timestamp 1635444444
transform 1 0 17204 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1635444444
transform -1 0 19412 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_199
timestamp 1635444444
transform 1 0 19412 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_207
timestamp 1635444444
transform 1 0 20148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1094_
timestamp 1635444444
transform 1 0 20516 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1103_
timestamp 1635444444
transform -1 0 20148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1635444444
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1635444444
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1635444444
transform 1 0 21804 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_241
timestamp 1635444444
transform 1 0 23276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_253
timestamp 1635444444
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_265
timestamp 1635444444
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1635444444
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1635444444
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1635444444
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1635444444
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_305
timestamp 1635444444
transform 1 0 29164 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_311
timestamp 1635444444
transform 1 0 29716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_316
timestamp 1635444444
transform 1 0 30176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635444444
transform -1 0 30820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1635444444
transform 1 0 29808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_13
timestamp 1635444444
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1635444444
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635444444
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1162_
timestamp 1635444444
transform 1 0 1472 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1635444444
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_39
timestamp 1635444444
transform 1 0 4692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1635444444
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1163_
timestamp 1635444444
transform 1 0 3772 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1170_
timestamp 1635444444
transform -1 0 5888 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_52
timestamp 1635444444
transform 1 0 5888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_58
timestamp 1635444444
transform 1 0 6440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1175_
timestamp 1635444444
transform 1 0 6532 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1635444444
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1635444444
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1635444444
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1635444444
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1071_
timestamp 1635444444
transform 1 0 7728 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1262_
timestamp 1635444444
transform -1 0 9568 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_10_103
timestamp 1635444444
transform 1 0 10580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_92
timestamp 1635444444
transform 1 0 9568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 10580 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_10_111
timestamp 1635444444
transform 1 0 11316 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1635444444
transform 1 0 12328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_129
timestamp 1635444444
transform 1 0 12972 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1507_
timestamp 1635444444
transform -1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1746_
timestamp 1635444444
transform -1 0 12328 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1635444444
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1635444444
transform 1 0 14352 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_148
timestamp 1635444444
transform 1 0 14720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1635444444
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1110_
timestamp 1635444444
transform 1 0 14812 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1505_
timestamp 1635444444
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1635444444
transform 1 0 15640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1635444444
transform 1 0 16008 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_178
timestamp 1635444444
transform 1 0 17480 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_190
timestamp 1635444444
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1635444444
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1095_
timestamp 1635444444
transform 1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_197
timestamp 1635444444
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_203
timestamp 1635444444
transform 1 0 19780 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1635444444
transform 1 0 19872 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_220
timestamp 1635444444
transform 1 0 21344 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_232
timestamp 1635444444
transform 1 0 22448 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1635444444
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1635444444
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1635444444
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1635444444
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1635444444
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1635444444
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1635444444
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1635444444
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_309
timestamp 1635444444
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_317
timestamp 1635444444
transform 1 0 30268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635444444
transform -1 0 30820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1635444444
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1635444444
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635444444
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1635444444
transform 1 0 1656 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_22
timestamp 1635444444
transform 1 0 3128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1635444444
transform 1 0 3864 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1112_
timestamp 1635444444
transform -1 0 3864 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1635444444
transform 1 0 4232 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_11_50
timestamp 1635444444
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1635444444
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1635444444
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1173_
timestamp 1635444444
transform 1 0 6440 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_11_68
timestamp 1635444444
transform 1 0 7360 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_76
timestamp 1635444444
transform 1 0 8096 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1075_
timestamp 1635444444
transform 1 0 8280 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_11_100
timestamp 1635444444
transform 1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1635444444
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_88
timestamp 1635444444
transform 1 0 9200 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1285_
timestamp 1635444444
transform -1 0 10304 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_wb_clk_i
timestamp 1635444444
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_122
timestamp 1635444444
transform 1 0 12328 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1635444444
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1106_
timestamp 1635444444
transform 1 0 13064 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1745_
timestamp 1635444444
transform 1 0 11500 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_140
timestamp 1635444444
transform 1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1635444444
transform 1 0 14352 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_160
timestamp 1635444444
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1635444444
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_173
timestamp 1635444444
transform 1 0 17020 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1635444444
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1088_
timestamp 1635444444
transform 1 0 17112 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_11_184
timestamp 1635444444
transform 1 0 18032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1944_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 18400 0 -1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1635444444
transform 1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1096_
timestamp 1635444444
transform -1 0 21344 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1635444444
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_234
timestamp 1635444444
transform 1 0 22632 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1635444444
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1092_
timestamp 1635444444
transform -1 0 22632 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_246
timestamp 1635444444
transform 1 0 23736 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_258
timestamp 1635444444
transform 1 0 24840 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_270
timestamp 1635444444
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1635444444
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1635444444
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1635444444
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1635444444
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_305
timestamp 1635444444
transform 1 0 29164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_316
timestamp 1635444444
transform 1 0 30176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635444444
transform -1 0 30820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1729_
timestamp 1635444444
transform 1 0 29900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1635444444
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1635444444
transform 1 0 1656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635444444
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1157_
timestamp 1635444444
transform -1 0 2944 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1635444444
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_39
timestamp 1635444444
transform 1 0 4692 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1635444444
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1165_
timestamp 1635444444
transform 1 0 3772 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1635444444
transform 1 0 5060 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_59
timestamp 1635444444
transform 1 0 6532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1635444444
transform -1 0 8372 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1635444444
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1635444444
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1635444444
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1084_
timestamp 1635444444
transform 1 0 8924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_108
timestamp 1635444444
transform 1 0 11040 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_94
timestamp 1635444444
transform 1 0 9752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_98
timestamp 1635444444
transform 1 0 10120 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1744_
timestamp 1635444444
transform 1 0 10212 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1635444444
transform 1 0 11684 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_119
timestamp 1635444444
transform 1 0 12052 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1253_
timestamp 1635444444
transform -1 0 11684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1635444444
transform -1 0 13616 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1635444444
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1635444444
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1635444444
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1635444444
transform 1 0 14168 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_12_158
timestamp 1635444444
transform 1 0 15640 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_168
timestamp 1635444444
transform 1 0 16560 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_wb_clk_i
timestamp 1635444444
transform -1 0 16560 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_wb_clk_i
timestamp 1635444444
transform 1 0 16928 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_176
timestamp 1635444444
transform 1 0 17296 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_180
timestamp 1635444444
transform 1 0 17664 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_190
timestamp 1635444444
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1635444444
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1089_
timestamp 1635444444
transform 1 0 17756 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1635444444
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_201
timestamp 1635444444
transform 1 0 19596 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_205
timestamp 1635444444
transform 1 0 19964 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1635444444
transform 1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1093_
timestamp 1635444444
transform 1 0 20332 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1723_
timestamp 1635444444
transform 1 0 19688 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_238
timestamp 1635444444
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1635444444
transform 1 0 21528 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1635444444
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1635444444
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1635444444
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1635444444
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1635444444
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1635444444
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1635444444
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1635444444
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_309
timestamp 1635444444
transform 1 0 29532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_316
timestamp 1635444444
transform 1 0 30176 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635444444
transform -1 0 30820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1635444444
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1635444444
transform 1 0 29808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1635444444
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1160_
timestamp 1635444444
transform 1 0 1656 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635444444
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635444444
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1635444444
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_6
timestamp 1635444444
transform 1 0 1656 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_10
timestamp 1635444444
transform 1 0 2024 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1635444444
transform 1 0 2852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1635444444
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1635444444
transform 1 0 2116 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1635444444
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_31
timestamp 1635444444
transform 1 0 3956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_41
timestamp 1635444444
transform 1 0 4876 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1635444444
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1635444444
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1635444444
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1169_
timestamp 1635444444
transform 1 0 4048 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1635444444
transform 1 0 3864 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_wb_clk_i
timestamp 1635444444
transform -1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1172_
timestamp 1635444444
transform -1 0 6532 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_46
timestamp 1635444444
transform 1 0 5336 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1635444444
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _1686_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 7084 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1645_
timestamp 1635444444
transform -1 0 7268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1635444444
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_59
timestamp 1635444444
transform 1 0 6532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1635444444
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1635444444
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_65
timestamp 1635444444
transform 1 0 7084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_73
timestamp 1635444444
transform 1 0 7820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_67
timestamp 1635444444
transform 1 0 7268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1635444444
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1635444444
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 1635444444
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1635444444
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1646_
timestamp 1635444444
transform -1 0 8004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1945_
timestamp 1635444444
transform 1 0 8188 0 -1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1635444444
transform -1 0 7820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1635444444
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_96
timestamp 1635444444
transform 1 0 9936 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_102
timestamp 1635444444
transform 1 0 10488 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1635444444
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1263_
timestamp 1635444444
transform -1 0 9660 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1277_
timestamp 1635444444
transform 1 0 10028 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1635444444
transform -1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_116
timestamp 1635444444
transform 1 0 11776 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_130
timestamp 1635444444
transform 1 0 13064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_126
timestamp 1635444444
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1635444444
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1113_
timestamp 1635444444
transform 1 0 12144 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1252_
timestamp 1635444444
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1635444444
transform 1 0 11224 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1635444444
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_144
timestamp 1635444444
transform 1 0 14352 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1635444444
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_150
timestamp 1635444444
transform 1 0 14904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1635444444
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1115_
timestamp 1635444444
transform 1 0 13432 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1116_
timestamp 1635444444
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1121_
timestamp 1635444444
transform 1 0 14720 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1635444444
transform 1 0 15272 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_158
timestamp 1635444444
transform 1 0 15640 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_157
timestamp 1635444444
transform 1 0 15548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _1667_
timestamp 1635444444
transform 1 0 16284 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1649_
timestamp 1635444444
transform 1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_164
timestamp 1635444444
transform 1 0 16192 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1635444444
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1635444444
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_171
timestamp 1635444444
transform 1 0 16836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1635444444
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1635444444
transform 1 0 17480 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1635444444
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1635444444
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1635444444
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1635444444
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1090_
timestamp 1635444444
transform 1 0 18124 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1665_
timestamp 1635444444
transform 1 0 17204 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _1678_
timestamp 1635444444
transform -1 0 17756 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1635444444
transform 1 0 17848 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_198
timestamp 1635444444
transform 1 0 19320 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1635444444
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1635444444
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1635444444
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_212
timestamp 1635444444
transform 1 0 20608 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_218
timestamp 1635444444
transform 1 0 21160 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1702_
timestamp 1635444444
transform 1 0 19688 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1703_
timestamp 1635444444
transform 1 0 20332 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1635444444
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1635444444
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1635444444
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_235
timestamp 1635444444
transform 1 0 22724 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1635444444
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1635444444
transform 1 0 21252 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1635444444
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1635444444
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_247
timestamp 1635444444
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1635444444
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1635444444
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1635444444
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1635444444
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1635444444
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1635444444
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1635444444
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1635444444
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1635444444
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1635444444
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1635444444
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1635444444
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1635444444
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_317
timestamp 1635444444
transform 1 0 30268 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1635444444
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_309
timestamp 1635444444
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_317
timestamp 1635444444
transform 1 0 30268 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635444444
transform -1 0 30820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635444444
transform -1 0 30820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1635444444
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_12
timestamp 1635444444
transform 1 0 2208 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635444444
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1158_
timestamp 1635444444
transform 1 0 1380 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1635444444
transform 1 0 2760 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_34
timestamp 1635444444
transform 1 0 4232 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1635444444
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_63
timestamp 1635444444
transform 1 0 6900 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1635444444
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_1  _1700_
timestamp 1635444444
transform -1 0 6900 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _1721_
timestamp 1635444444
transform 1 0 5336 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_79
timestamp 1635444444
transform 1 0 8372 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_87
timestamp 1635444444
transform 1 0 9108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1635444444
transform -1 0 8372 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1635444444
transform -1 0 9108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1635444444
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_95
timestamp 1635444444
transform 1 0 9844 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1127_
timestamp 1635444444
transform 1 0 9936 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1635444444
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_122
timestamp 1635444444
transform 1 0 12328 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_128
timestamp 1635444444
transform 1 0 12880 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1635444444
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1120_
timestamp 1635444444
transform 1 0 12972 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1125_
timestamp 1635444444
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_138
timestamp 1635444444
transform 1 0 13800 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1370_
timestamp 1635444444
transform 1 0 14904 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_154
timestamp 1635444444
transform 1 0 15272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1635444444
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1635444444
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_1  _1655_
timestamp 1635444444
transform 1 0 15640 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1668_
timestamp 1635444444
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1635444444
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1635444444
transform 1 0 17848 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_186
timestamp 1635444444
transform 1 0 18216 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_192
timestamp 1635444444
transform 1 0 18768 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1675_
timestamp 1635444444
transform 1 0 17940 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1705_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 18860 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_199
timestamp 1635444444
transform 1 0 19412 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_212
timestamp 1635444444
transform 1 0 20608 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1706_
timestamp 1635444444
transform 1 0 19780 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1714_
timestamp 1635444444
transform -1 0 21252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1635444444
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1635444444
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1635444444
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1635444444
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1635444444
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1635444444
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1635444444
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1635444444
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1635444444
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1635444444
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1635444444
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1635444444
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1635444444
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_317
timestamp 1635444444
transform 1 0 30268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635444444
transform -1 0 30820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1635444444
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635444444
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1635444444
transform 1 0 1380 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1635444444
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_38
timestamp 1635444444
transform 1 0 4600 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1635444444
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1156_
timestamp 1635444444
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_44
timestamp 1635444444
transform 1 0 5152 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_51
timestamp 1635444444
transform 1 0 5796 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_63
timestamp 1635444444
transform 1 0 6900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_1  _1711_
timestamp 1635444444
transform 1 0 5244 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1635444444
transform 1 0 6992 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1635444444
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1635444444
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1635444444
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1360_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 9476 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_91
timestamp 1635444444
transform 1 0 9476 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_97
timestamp 1635444444
transform 1 0 10028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1635444444
transform 1 0 10120 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_114
timestamp 1635444444
transform 1 0 11592 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_126
timestamp 1635444444
transform 1 0 12696 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1119_
timestamp 1635444444
transform 1 0 12788 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1635444444
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1635444444
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1635444444
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_157
timestamp 1635444444
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1635444444
transform 1 0 16744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1656_
timestamp 1635444444
transform 1 0 15916 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1679_
timestamp 1635444444
transform 1 0 17112 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_183
timestamp 1635444444
transform 1 0 17940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_187
timestamp 1635444444
transform 1 0 18308 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1635444444
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1635444444
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1682_
timestamp 1635444444
transform 1 0 18400 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1635444444
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_203
timestamp 1635444444
transform 1 0 19780 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_213
timestamp 1635444444
transform 1 0 20700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1716_
timestamp 1635444444
transform -1 0 20700 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1724_
timestamp 1635444444
transform -1 0 21344 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_220
timestamp 1635444444
transform 1 0 21344 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_232
timestamp 1635444444
transform 1 0 22448 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1635444444
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1635444444
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1635444444
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1635444444
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1635444444
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1635444444
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1635444444
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1635444444
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_309
timestamp 1635444444
transform 1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_316
timestamp 1635444444
transform 1 0 30176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635444444
transform -1 0 30820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1635444444
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1635444444
transform 1 0 29808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_14
timestamp 1635444444
transform 1 0 2392 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_6
timestamp 1635444444
transform 1 0 1656 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635444444
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1154_
timestamp 1635444444
transform 1 0 2576 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1635444444
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1635444444
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_37
timestamp 1635444444
transform 1 0 4508 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_42
timestamp 1635444444
transform 1 0 4968 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1635444444
transform 1 0 4600 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_48
timestamp 1635444444
transform 1 0 5520 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1635444444
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1635444444
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1635444444
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1635444444
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1660_
timestamp 1635444444
transform 1 0 5612 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_75
timestamp 1635444444
transform 1 0 8004 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_81
timestamp 1635444444
transform 1 0 8556 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1129_
timestamp 1635444444
transform 1 0 7176 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_2  _1265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8648 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1635444444
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_90
timestamp 1635444444
transform 1 0 9384 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_98
timestamp 1635444444
transform 1 0 10120 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1128_
timestamp 1635444444
transform 1 0 10212 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1635444444
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1635444444
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1635444444
transform 1 0 12236 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_137
timestamp 1635444444
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1635444444
transform 1 0 14076 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_157
timestamp 1635444444
transform 1 0 15548 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1635444444
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_172
timestamp 1635444444
transform 1 0 16928 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1635444444
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1666_
timestamp 1635444444
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1677_
timestamp 1635444444
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_180
timestamp 1635444444
transform 1 0 17664 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_189
timestamp 1635444444
transform 1 0 18492 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1683_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1715_
timestamp 1635444444
transform 1 0 19044 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_17_200
timestamp 1635444444
transform 1 0 19504 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_213
timestamp 1635444444
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1726_
timestamp 1635444444
transform 1 0 19872 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1635444444
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1635444444
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_239
timestamp 1635444444
transform 1 0 23092 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1635444444
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1375_
timestamp 1635444444
transform 1 0 22172 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_17_251
timestamp 1635444444
transform 1 0 24196 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_263
timestamp 1635444444
transform 1 0 25300 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1635444444
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1635444444
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1635444444
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1635444444
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1635444444
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1635444444
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_317
timestamp 1635444444
transform 1 0 30268 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635444444
transform -1 0 30820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_14
timestamp 1635444444
transform 1 0 2392 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_6
timestamp 1635444444
transform 1 0 1656 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635444444
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1153_
timestamp 1635444444
transform 1 0 2484 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1635444444
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1635444444
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1635444444
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1635444444
transform 1 0 3772 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_45
timestamp 1635444444
transform 1 0 5244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_52
timestamp 1635444444
transform 1 0 5888 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_56
timestamp 1635444444
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_61
timestamp 1635444444
transform 1 0 6716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1638_
timestamp 1635444444
transform 1 0 5612 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1676_
timestamp 1635444444
transform -1 0 6716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1722_
timestamp 1635444444
transform 1 0 7084 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_74
timestamp 1635444444
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1635444444
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1635444444
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1635444444
transform -1 0 10396 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_101
timestamp 1635444444
transform 1 0 10396 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1635444444
transform 1 0 10948 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1635444444
transform 1 0 12420 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 1635444444
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1635444444
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_145
timestamp 1635444444
transform 1 0 14444 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_152
timestamp 1635444444
transform 1 0 15088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1635444444
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1651_
timestamp 1635444444
transform 1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1635444444
transform -1 0 14444 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1635444444
transform 1 0 16376 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1650_
timestamp 1635444444
transform 1 0 15456 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_18_178
timestamp 1635444444
transform 1 0 17480 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1635444444
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1635444444
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _1691_
timestamp 1635444444
transform 1 0 17848 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1635444444
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_204
timestamp 1635444444
transform 1 0 19872 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_217
timestamp 1635444444
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1725_
timestamp 1635444444
transform 1 0 19412 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1727_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 21068 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_18_226
timestamp 1635444444
transform 1 0 21896 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_238
timestamp 1635444444
transform 1 0 23000 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1374_
timestamp 1635444444
transform 1 0 21436 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1635444444
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1635444444
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1635444444
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1635444444
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1635444444
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1635444444
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1635444444
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1635444444
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_309
timestamp 1635444444
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_317
timestamp 1635444444
transform 1 0 30268 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635444444
transform -1 0 30820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1635444444
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_6
timestamp 1635444444
transform 1 0 1656 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_6
timestamp 1635444444
transform 1 0 1656 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635444444
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635444444
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1149_
timestamp 1635444444
transform 1 0 2208 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1151_
timestamp 1635444444
transform -1 0 3128 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1635444444
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1635444444
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1635444444
transform 1 0 4048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1635444444
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_29
timestamp 1635444444
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1635444444
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_26
timestamp 1635444444
transform 1 0 3496 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_22
timestamp 1635444444
transform 1 0 3128 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_wb_clk_i
timestamp 1635444444
transform -1 0 5336 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_41
timestamp 1635444444
transform 1 0 4876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_35
timestamp 1635444444
transform 1 0 4324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_43
timestamp 1635444444
transform 1 0 5060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1635444444
transform 1 0 3588 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_19_47
timestamp 1635444444
transform 1 0 5428 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1635444444
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_46
timestamp 1635444444
transform 1 0 5336 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1635444444
transform 1 0 6532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1635444444
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1642_
timestamp 1635444444
transform 1 0 6900 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1648_
timestamp 1635444444
transform 1 0 5704 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1663_
timestamp 1635444444
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1635444444
transform -1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_66
timestamp 1635444444
transform 1 0 7176 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1635444444
transform 1 0 8832 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_73
timestamp 1635444444
transform 1 0 7820 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1635444444
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1635444444
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1635444444
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1652_
timestamp 1635444444
transform -1 0 8832 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1720_
timestamp 1635444444
transform -1 0 8464 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1635444444
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_88
timestamp 1635444444
transform 1 0 9200 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_94
timestamp 1635444444
transform 1 0 9752 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_96
timestamp 1635444444
transform 1 0 9936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1118_
timestamp 1635444444
transform 1 0 10488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1356_
timestamp 1635444444
transform -1 0 9752 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1358_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9476 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1635444444
transform 1 0 10304 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1635444444
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1635444444
transform 1 0 12696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_116
timestamp 1635444444
transform 1 0 11776 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_124
timestamp 1635444444
transform 1 0 12512 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1635444444
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _1028_
timestamp 1635444444
transform 1 0 12696 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1123_
timestamp 1635444444
transform 1 0 11868 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_wb_clk_i
timestamp 1635444444
transform -1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1635444444
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1635444444
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1635444444
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_wb_clk_i
timestamp 1635444444
transform 1 0 14168 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1575_
timestamp 1635444444
transform 1 0 14996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1574_
timestamp 1635444444
transform -1 0 15364 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_20_146
timestamp 1635444444
transform 1 0 14536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_150
timestamp 1635444444
transform 1 0 14904 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1635444444
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_134
timestamp 1635444444
transform 1 0 13432 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_155
timestamp 1635444444
transform 1 0 15364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1635444444
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_155
timestamp 1635444444
transform 1 0 15364 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_164
timestamp 1635444444
transform 1 0 16192 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1635444444
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1641_
timestamp 1635444444
transform -1 0 16192 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1643_
timestamp 1635444444
transform 1 0 15732 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _1644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 17388 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _1654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 17848 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_19_177
timestamp 1635444444
transform 1 0 17388 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_185
timestamp 1635444444
transform 1 0 18124 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_182
timestamp 1635444444
transform 1 0 17848 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1635444444
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1635444444
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1635444444
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _1704_
timestamp 1635444444
transform 1 0 18216 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 19780 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_19_203
timestamp 1635444444
transform 1 0 19780 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1635444444
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1635444444
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_204
timestamp 1635444444
transform 1 0 19872 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_208
timestamp 1635444444
transform 1 0 20240 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_216
timestamp 1635444444
transform 1 0 20976 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_4  _1044_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 20148 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1635444444
transform -1 0 19872 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1669_
timestamp 1635444444
transform -1 0 20976 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1635444444
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1635444444
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1635444444
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_228
timestamp 1635444444
transform 1 0 22080 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_240
timestamp 1635444444
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1635444444
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1635444444
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1635444444
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1635444444
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1635444444
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1635444444
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1635444444
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1635444444
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1635444444
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1635444444
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1635444444
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1635444444
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_305
timestamp 1635444444
transform 1 0 29164 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1635444444
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1635444444
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_316
timestamp 1635444444
transform 1 0 30176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1635444444
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1635444444
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_316
timestamp 1635444444
transform 1 0 30176 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635444444
transform -1 0 30820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635444444
transform -1 0 30820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1635444444
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1728_
timestamp 1635444444
transform 1 0 29900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1635444444
transform 1 0 29808 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_19
timestamp 1635444444
transform 1 0 2852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635444444
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1635444444
transform 1 0 1380 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_23
timestamp 1635444444
transform 1 0 3220 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_34
timestamp 1635444444
transform 1 0 4232 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_40
timestamp 1635444444
transform 1 0 4784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1146_
timestamp 1635444444
transform 1 0 3312 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1671_
timestamp 1635444444
transform 1 0 4876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_44
timestamp 1635444444
transform 1 0 5152 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1635444444
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1635444444
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1653_
timestamp 1635444444
transform 1 0 5520 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1674_
timestamp 1635444444
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_66
timestamp 1635444444
transform 1 0 7176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_74
timestamp 1635444444
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_80
timestamp 1635444444
transform 1 0 8464 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1357_
timestamp 1635444444
transform 1 0 8832 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1639_
timestamp 1635444444
transform -1 0 8464 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1635444444
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_88
timestamp 1635444444
transform 1 0 9200 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1635444444
transform 1 0 10212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1126_
timestamp 1635444444
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _1384_
timestamp 1635444444
transform -1 0 10212 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1635444444
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1635444444
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_120
timestamp 1635444444
transform 1 0 12144 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_128
timestamp 1635444444
transform 1 0 12880 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1635444444
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1017_
timestamp 1635444444
transform 1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 12144 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_21_132
timestamp 1635444444
transform 1 0 13248 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_136
timestamp 1635444444
transform 1 0 13616 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_148
timestamp 1635444444
transform 1 0 14720 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1635444444
transform -1 0 13616 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _1528_
timestamp 1635444444
transform -1 0 15640 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1635444444
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1635444444
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1635444444
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _1573_
timestamp 1635444444
transform -1 0 17204 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_175
timestamp 1635444444
transform 1 0 17204 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1635444444
transform 1 0 18032 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_191
timestamp 1635444444
transform 1 0 18676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0914_
timestamp 1635444444
transform -1 0 19412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1021_
timestamp 1635444444
transform 1 0 17572 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1560_
timestamp 1635444444
transform -1 0 18676 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_199
timestamp 1635444444
transform 1 0 19412 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_207
timestamp 1635444444
transform 1 0 20148 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1635444444
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1680_
timestamp 1635444444
transform -1 0 20884 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1635444444
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1635444444
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1635444444
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1635444444
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1635444444
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1635444444
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1635444444
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1635444444
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1635444444
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1635444444
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1635444444
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_305
timestamp 1635444444
transform 1 0 29164 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_316
timestamp 1635444444
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635444444
transform -1 0 30820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1670_
timestamp 1635444444
transform 1 0 29900 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_14
timestamp 1635444444
transform 1 0 2392 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_6
timestamp 1635444444
transform 1 0 1656 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635444444
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1150_
timestamp 1635444444
transform 1 0 2484 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1635444444
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1635444444
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1635444444
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1635444444
transform 1 0 3772 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_45
timestamp 1635444444
transform 1 0 5244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_58
timestamp 1635444444
transform 1 0 6440 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1687_
timestamp 1635444444
transform 1 0 6808 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1695_
timestamp 1635444444
transform 1 0 5612 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_71
timestamp 1635444444
transform 1 0 7636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1635444444
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1635444444
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1286_
timestamp 1635444444
transform -1 0 8464 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1295_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_101
timestamp 1635444444
transform 1 0 10396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_108
timestamp 1635444444
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1635444444
transform 1 0 9660 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1359_
timestamp 1635444444
transform 1 0 10764 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_wb_clk_i
timestamp 1635444444
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_112
timestamp 1635444444
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_116
timestamp 1635444444
transform 1 0 11776 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1378_
timestamp 1635444444
transform -1 0 11776 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1635444444
transform 1 0 12144 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1635444444
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1635444444
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1635444444
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0903_
timestamp 1635444444
transform -1 0 15272 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_154
timestamp 1635444444
transform 1 0 15272 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_162
timestamp 1635444444
transform 1 0 16008 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_171
timestamp 1635444444
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1657_
timestamp 1635444444
transform -1 0 16836 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_22_175
timestamp 1635444444
transform 1 0 17204 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_183
timestamp 1635444444
transform 1 0 17940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1635444444
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1635444444
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1539_
timestamp 1635444444
transform 1 0 18308 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1688_
timestamp 1635444444
transform -1 0 17940 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_22_197
timestamp 1635444444
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1635444444
transform 1 0 20424 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1664_
timestamp 1635444444
transform 1 0 20792 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1717_
timestamp 1635444444
transform -1 0 20424 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_22_224
timestamp 1635444444
transform 1 0 21712 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_236
timestamp 1635444444
transform 1 0 22816 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1635444444
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1635444444
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1635444444
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1635444444
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1635444444
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1635444444
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1635444444
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1635444444
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_309
timestamp 1635444444
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_316
timestamp 1635444444
transform 1 0 30176 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635444444
transform -1 0 30820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1635444444
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1658_
timestamp 1635444444
transform 1 0 29900 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_14
timestamp 1635444444
transform 1 0 2392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1635444444
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1635444444
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1147_
timestamp 1635444444
transform 1 0 2760 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1152_
timestamp 1635444444
transform -1 0 2392 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1635444444
transform 1 0 3588 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1635444444
transform 1 0 3956 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1635444444
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1635444444
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1635444444
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1701_
timestamp 1635444444
transform 1 0 6348 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_66
timestamp 1635444444
transform 1 0 7176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_87
timestamp 1635444444
transform 1 0 9108 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1851_
timestamp 1635444444
transform -1 0 9108 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1635444444
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1847_
timestamp 1635444444
transform 1 0 9476 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_23_113
timestamp 1635444444
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_128
timestamp 1635444444
transform 1 0 12880 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1635444444
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _1733_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 12880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_135
timestamp 1635444444
transform 1 0 13524 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_143
timestamp 1635444444
transform 1 0 14260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _1369_
timestamp 1635444444
transform 1 0 13248 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1974_
timestamp 1635444444
transform 1 0 14444 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1635444444
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1635444444
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1635444444
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1635444444
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1696_
timestamp 1635444444
transform -1 0 17756 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_181
timestamp 1635444444
transform 1 0 17756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1635444444
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0902_
timestamp 1635444444
transform 1 0 18124 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_201
timestamp 1635444444
transform 1 0 19596 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_209
timestamp 1635444444
transform 1 0 20332 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1635444444
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0897_
timestamp 1635444444
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1707_
timestamp 1635444444
transform -1 0 21068 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1635444444
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_235
timestamp 1635444444
transform 1 0 22724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1635444444
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1659_
timestamp 1635444444
transform 1 0 21804 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_23_247
timestamp 1635444444
transform 1 0 23828 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_259
timestamp 1635444444
transform 1 0 24932 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_271
timestamp 1635444444
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1635444444
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1635444444
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1635444444
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1635444444
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1708_
timestamp 1635444444
transform 1 0 29164 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_308
timestamp 1635444444
transform 1 0 29440 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_316
timestamp 1635444444
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1635444444
transform -1 0 30820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1635444444
transform 1 0 29808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_16
timestamp 1635444444
transform 1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1635444444
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1635444444
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1145_
timestamp 1635444444
transform -1 0 2576 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1635444444
transform 1 0 2944 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1635444444
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1635444444
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_38
timestamp 1635444444
transform 1 0 4600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_42
timestamp 1635444444
transform 1 0 4968 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1635444444
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1144_
timestamp 1635444444
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1635444444
transform 1 0 5060 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_46
timestamp 1635444444
transform 1 0 5336 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_59
timestamp 1635444444
transform 1 0 6532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1712_
timestamp 1635444444
transform 1 0 5704 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_67
timestamp 1635444444
transform 1 0 7268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_78
timestamp 1635444444
transform 1 0 8280 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1635444444
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1635444444
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1291_
timestamp 1635444444
transform 1 0 7544 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1297_
timestamp 1635444444
transform 1 0 9016 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_102
timestamp 1635444444
transform 1 0 10488 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_95
timestamp 1635444444
transform 1 0 9844 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1635444444
transform 1 0 10212 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_114
timestamp 1635444444
transform 1 0 11592 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_122
timestamp 1635444444
transform 1 0 12328 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_126
timestamp 1635444444
transform 1 0 12696 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1379_
timestamp 1635444444
transform -1 0 13524 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1380_
timestamp 1635444444
transform 1 0 12420 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1635444444
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1635444444
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1635444444
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1635444444
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1635444444
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0905_
timestamp 1635444444
transform -1 0 15364 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_24_155
timestamp 1635444444
transform 1 0 15364 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1635444444
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0899_
timestamp 1635444444
transform 1 0 16652 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1535_
timestamp 1635444444
transform 1 0 15916 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_178
timestamp 1635444444
transform 1 0 17480 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1635444444
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1635444444
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1635444444
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0896_
timestamp 1635444444
transform -1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1635444444
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1635444444
transform 1 0 20884 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1977_
timestamp 1635444444
transform 1 0 19412 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_24_223
timestamp 1635444444
transform 1 0 21620 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_235
timestamp 1635444444
transform 1 0 22724 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1046_
timestamp 1635444444
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1635444444
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1635444444
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1635444444
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1635444444
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1635444444
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1635444444
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1635444444
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1635444444
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1635444444
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_309
timestamp 1635444444
transform 1 0 29532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_316
timestamp 1635444444
transform 1 0 30176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1635444444
transform -1 0 30820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1635444444
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1697_
timestamp 1635444444
transform 1 0 29900 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1635444444
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1635444444
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1635444444
transform 1 0 1656 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_22
timestamp 1635444444
transform 1 0 3128 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_35
timestamp 1635444444
transform 1 0 4324 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_41
timestamp 1635444444
transform 1 0 4876 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1143_
timestamp 1635444444
transform 1 0 3496 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1709_
timestamp 1635444444
transform 1 0 4968 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_45
timestamp 1635444444
transform 1 0 5244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1635444444
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_60
timestamp 1635444444
transform 1 0 6624 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1635444444
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1117_
timestamp 1635444444
transform 1 0 6992 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1685_
timestamp 1635444444
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1698_
timestamp 1635444444
transform 1 0 5612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_68
timestamp 1635444444
transform 1 0 7360 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_76
timestamp 1635444444
transform 1 0 8096 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_87
timestamp 1635444444
transform 1 0 9108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1289_
timestamp 1635444444
transform -1 0 9108 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1635444444
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_91
timestamp 1635444444
transform 1 0 9476 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1635444444
transform 1 0 9568 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1635444444
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_128
timestamp 1635444444
transform 1 0 12880 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1635444444
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1635444444
transform -1 0 12880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_138
timestamp 1635444444
transform 1 0 13800 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_144
timestamp 1635444444
transform 1 0 14352 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1019_
timestamp 1635444444
transform -1 0 13800 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1973_
timestamp 1635444444
transform 1 0 14444 0 -1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1635444444
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_169
timestamp 1635444444
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1635444444
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1976_
timestamp 1635444444
transform 1 0 16928 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_25_189
timestamp 1635444444
transform 1 0 18492 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0898_
timestamp 1635444444
transform 1 0 18860 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_202
timestamp 1635444444
transform 1 0 19688 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_211
timestamp 1635444444
transform 1 0 20516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1020_
timestamp 1635444444
transform -1 0 20516 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1534_
timestamp 1635444444
transform -1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1635444444
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1635444444
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1635444444
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1635444444
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1635444444
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1635444444
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1635444444
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1635444444
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1635444444
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1635444444
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1635444444
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1635444444
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_305
timestamp 1635444444
transform 1 0 29164 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1635444444
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1635444444
transform -1 0 30820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1718_
timestamp 1635444444
transform 1 0 29900 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_6
timestamp 1635444444
transform 1 0 1656 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_20
timestamp 1635444444
transform 1 0 2944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_6
timestamp 1635444444
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1635444444
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1635444444
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1134_
timestamp 1635444444
transform -1 0 2944 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1142_
timestamp 1635444444
transform -1 0 3312 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1635444444
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1635444444
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1635444444
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_29
timestamp 1635444444
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_28
timestamp 1635444444
transform 1 0 3680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1635444444
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1635444444
transform 1 0 3864 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1635444444
transform 1 0 4324 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1635444444
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_46
timestamp 1635444444
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_51
timestamp 1635444444
transform 1 0 5796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1719_
timestamp 1635444444
transform 1 0 6808 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1640_
timestamp 1635444444
transform 1 0 6164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1290_
timestamp 1635444444
transform 1 0 6716 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1635444444
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1635444444
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_58
timestamp 1635444444
transform 1 0 6440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1635444444
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1635444444
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1635444444
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_70
timestamp 1635444444
transform 1 0 7544 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_78
timestamp 1635444444
transform 1 0 8280 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1635444444
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1288_
timestamp 1635444444
transform -1 0 9844 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1294_
timestamp 1635444444
transform 1 0 8372 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_108
timestamp 1635444444
transform 1 0 11040 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_95
timestamp 1635444444
transform 1 0 9844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1635444444
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_88
timestamp 1635444444
transform 1 0 9200 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1296_
timestamp 1635444444
transform 1 0 10212 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1635444444
transform -1 0 11040 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_26_116
timestamp 1635444444
transform 1 0 11776 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_123
timestamp 1635444444
transform 1 0 12420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1635444444
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_131
timestamp 1635444444
transform 1 0 13156 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1635444444
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _0884_
timestamp 1635444444
transform 1 0 11868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 13616 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1950_
timestamp 1635444444
transform 1 0 11684 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__o31a_1  _1060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14076 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1024_
timestamp 1635444444
transform -1 0 14260 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1635444444
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_137
timestamp 1635444444
transform 1 0 13708 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1635444444
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1635444444
transform 1 0 14720 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1026_
timestamp 1635444444
transform -1 0 15456 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_147
timestamp 1635444444
transform 1 0 14628 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_143
timestamp 1635444444
transform 1 0 14260 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1635444444
transform 1 0 14720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_151
timestamp 1635444444
transform 1 0 14996 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_156
timestamp 1635444444
transform 1 0 15456 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_169
timestamp 1635444444
transform 1 0 16652 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1635444444
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1635444444
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_169
timestamp 1635444444
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1635444444
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1022_
timestamp 1635444444
transform 1 0 17020 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1635444444
transform -1 0 16652 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1562_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 17664 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_179
timestamp 1635444444
transform 1 0 17572 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1635444444
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1635444444
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_180
timestamp 1635444444
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_189
timestamp 1635444444
transform 1 0 18492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1635444444
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1561_
timestamp 1635444444
transform 1 0 18032 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_26_200
timestamp 1635444444
transform 1 0 19504 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_208
timestamp 1635444444
transform 1 0 20240 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_206
timestamp 1635444444
transform 1 0 20056 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_214
timestamp 1635444444
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1635444444
transform -1 0 19504 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1730_
timestamp 1635444444
transform 1 0 19228 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1978_
timestamp 1635444444
transform 1 0 20332 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_26_225
timestamp 1635444444
transform 1 0 21804 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_237
timestamp 1635444444
transform 1 0 22908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1635444444
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_228
timestamp 1635444444
transform 1 0 22080 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_240
timestamp 1635444444
transform 1 0 23184 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1635444444
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1623_
timestamp 1635444444
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1635444444
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1635444444
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_252
timestamp 1635444444
transform 1 0 24288 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1635444444
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1635444444
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1635444444
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_264
timestamp 1635444444
transform 1 0 25392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1635444444
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1635444444
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1635444444
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1635444444
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1635444444
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1635444444
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_305
timestamp 1635444444
transform 1 0 29164 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1635444444
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_309
timestamp 1635444444
transform 1 0 29532 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_317
timestamp 1635444444
transform 1 0 30268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_311
timestamp 1635444444
transform 1 0 29716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_316
timestamp 1635444444
transform 1 0 30176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1635444444
transform -1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1635444444
transform -1 0 30820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1635444444
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1635444444
transform 1 0 29808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1635444444
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1635444444
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1635444444
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1635444444
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1635444444
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_39
timestamp 1635444444
transform 1 0 4692 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1635444444
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1140_
timestamp 1635444444
transform 1 0 3772 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1635444444
transform 1 0 5060 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_46
timestamp 1635444444
transform 1 0 5336 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_55
timestamp 1635444444
transform 1 0 6164 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1270_
timestamp 1635444444
transform -1 0 6164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1635444444
transform 1 0 6532 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_28_75
timestamp 1635444444
transform 1 0 8004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1635444444
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1635444444
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1635444444
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_93
timestamp 1635444444
transform 1 0 9660 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1635444444
transform 1 0 9936 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_28_112
timestamp 1635444444
transform 1 0 11408 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_120
timestamp 1635444444
transform 1 0 12144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_126
timestamp 1635444444
transform 1 0 12696 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1068_
timestamp 1635444444
transform 1 0 12420 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1635444444
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1635444444
transform 1 0 14812 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1635444444
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_1  _1066_
timestamp 1635444444
transform 1 0 13248 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 14812 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_153
timestamp 1635444444
transform 1 0 15180 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_158
timestamp 1635444444
transform 1 0 15640 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_171
timestamp 1635444444
transform 1 0 16836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1540_
timestamp 1635444444
transform 1 0 15272 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1802_
timestamp 1635444444
transform -1 0 16836 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1635444444
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1635444444
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1585_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 18768 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_28_204
timestamp 1635444444
transform 1 0 19872 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_213
timestamp 1635444444
transform 1 0 20700 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1584_
timestamp 1635444444
transform 1 0 21068 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1605_
timestamp 1635444444
transform 1 0 19228 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1625_
timestamp 1635444444
transform 1 0 20240 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_28_220
timestamp 1635444444
transform 1 0 21344 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1635444444
transform 1 0 21988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1635444444
transform 1 0 23092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1604_
timestamp 1635444444
transform 1 0 21712 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1635444444
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1635444444
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1635444444
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1635444444
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1635444444
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1635444444
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1635444444
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1635444444
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_309
timestamp 1635444444
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_317
timestamp 1635444444
transform 1 0 30268 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1635444444
transform -1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1635444444
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1635444444
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1635444444
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1635444444
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1139_
timestamp 1635444444
transform 1 0 1656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1141_
timestamp 1635444444
transform -1 0 3680 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_28
timestamp 1635444444
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_36
timestamp 1635444444
transform 1 0 4416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_43
timestamp 1635444444
transform 1 0 5060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1130_
timestamp 1635444444
transform -1 0 4416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1635444444
transform 1 0 4784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_47
timestamp 1635444444
transform 1 0 5428 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1635444444
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_57
timestamp 1635444444
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1635444444
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1271_
timestamp 1635444444
transform 1 0 5520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1635444444
transform 1 0 6900 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_79
timestamp 1635444444
transform 1 0 8372 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_83
timestamp 1635444444
transform 1 0 8740 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1635444444
transform -1 0 10304 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_100
timestamp 1635444444
transform 1 0 10304 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1635444444
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1148_
timestamp 1635444444
transform -1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1635444444
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_121
timestamp 1635444444
transform 1 0 12236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_125
timestamp 1635444444
transform 1 0 12604 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_129
timestamp 1635444444
transform 1 0 12972 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1635444444
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1635444444
transform -1 0 12972 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1189_
timestamp 1635444444
transform 1 0 11868 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_141
timestamp 1635444444
transform 1 0 14076 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_149
timestamp 1635444444
transform 1 0 14812 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1768_
timestamp 1635444444
transform 1 0 14904 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1635444444
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1635444444
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1635444444
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_12  _1371_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 16652 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_185
timestamp 1635444444
transform 1 0 18124 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_193
timestamp 1635444444
transform 1 0 18860 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1782_
timestamp 1635444444
transform 1 0 18952 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_203
timestamp 1635444444
transform 1 0 19780 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1732_
timestamp 1635444444
transform 1 0 20516 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1635444444
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_228
timestamp 1635444444
transform 1 0 22080 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_240
timestamp 1635444444
transform 1 0 23184 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1635444444
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1626_
timestamp 1635444444
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_252
timestamp 1635444444
transform 1 0 24288 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_264
timestamp 1635444444
transform 1 0 25392 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1635444444
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1635444444
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1635444444
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1635444444
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_305
timestamp 1635444444
transform 1 0 29164 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_316
timestamp 1635444444
transform 1 0 30176 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1635444444
transform -1 0 30820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1681_
timestamp 1635444444
transform 1 0 29900 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_13
timestamp 1635444444
transform 1 0 2300 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_19
timestamp 1635444444
transform 1 0 2852 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1635444444
transform 1 0 1380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1635444444
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1137_
timestamp 1635444444
transform 1 0 1472 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1138_
timestamp 1635444444
transform -1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1635444444
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_39
timestamp 1635444444
transform 1 0 4692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1635444444
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1132_
timestamp 1635444444
transform 1 0 3772 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_30_50
timestamp 1635444444
transform 1 0 5704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_54
timestamp 1635444444
transform 1 0 6072 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_65
timestamp 1635444444
transform 1 0 7084 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1283_
timestamp 1635444444
transform 1 0 6164 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1661_
timestamp 1635444444
transform 1 0 5428 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1635444444
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1635444444
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1292_
timestamp 1635444444
transform 1 0 8924 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1293_
timestamp 1635444444
transform -1 0 8280 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_102
timestamp 1635444444
transform 1 0 10488 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_109
timestamp 1635444444
transform 1 0 11132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_94
timestamp 1635444444
transform 1 0 9752 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0883_
timestamp 1635444444
transform 1 0 10764 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_122
timestamp 1635444444
transform 1 0 12328 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_130
timestamp 1635444444
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1105_
timestamp 1635444444
transform 1 0 12696 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1205_
timestamp 1635444444
transform 1 0 11500 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1635444444
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_141
timestamp 1635444444
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_145
timestamp 1635444444
transform 1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1635444444
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1635444444
transform 1 0 14168 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1767_
timestamp 1635444444
transform -1 0 15640 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_158
timestamp 1635444444
transform 1 0 15640 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_166
timestamp 1635444444
transform 1 0 16376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1542_
timestamp 1635444444
transform -1 0 16376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1563_
timestamp 1635444444
transform -1 0 17664 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_30_180
timestamp 1635444444
transform 1 0 17664 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_184
timestamp 1635444444
transform 1 0 18032 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1635444444
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1635444444
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1635444444
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1586_
timestamp 1635444444
transform -1 0 18492 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_200
timestamp 1635444444
transform 1 0 19504 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_204
timestamp 1635444444
transform 1 0 19872 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_214
timestamp 1635444444
transform 1 0 20792 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1583_
timestamp 1635444444
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1774_
timestamp 1635444444
transform 1 0 19964 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_222
timestamp 1635444444
transform 1 0 21528 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_232
timestamp 1635444444
transform 1 0 22448 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1788_
timestamp 1635444444
transform 1 0 21620 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 1635444444
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1635444444
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1635444444
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1635444444
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1635444444
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1635444444
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1635444444
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1635444444
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1635444444
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_316
timestamp 1635444444
transform 1 0 30176 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1635444444
transform -1 0 30820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1635444444
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1689_
timestamp 1635444444
transform 1 0 29900 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_6
timestamp 1635444444
transform 1 0 1656 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1635444444
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1635444444
transform 1 0 2208 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1635444444
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_28
timestamp 1635444444
transform 1 0 3680 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_34
timestamp 1635444444
transform 1 0 4232 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1635444444
transform 1 0 4324 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1635444444
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1635444444
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_60
timestamp 1635444444
transform 1 0 6624 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1635444444
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1710_
timestamp 1635444444
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_72
timestamp 1635444444
transform 1 0 7728 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_80
timestamp 1635444444
transform 1 0 8464 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_84
timestamp 1635444444
transform 1 0 8832 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1430_
timestamp 1635444444
transform -1 0 8832 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_100
timestamp 1635444444
transform 1 0 10304 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1635444444
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_91
timestamp 1635444444
transform 1 0 9476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0979_
timestamp 1635444444
transform -1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1635444444
transform 1 0 9844 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1389_
timestamp 1635444444
transform -1 0 9476 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1635444444
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1635444444
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 11868 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 1635444444
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1951_
timestamp 1635444444
transform -1 0 15548 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1635444444
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1635444444
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1635444444
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1635444444
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1179_
timestamp 1635444444
transform -1 0 17112 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1541_
timestamp 1635444444
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_178
timestamp 1635444444
transform 1 0 17480 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_188
timestamp 1635444444
transform 1 0 18400 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1771_
timestamp 1635444444
transform 1 0 17572 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1808_
timestamp 1635444444
transform 1 0 18768 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_201
timestamp 1635444444
transform 1 0 19596 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_212
timestamp 1635444444
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1627_
timestamp 1635444444
transform 1 0 20976 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_1  _1637_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 20608 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1635444444
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1635444444
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1635444444
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1635444444
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _1731_
timestamp 1635444444
transform 1 0 22172 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_241
timestamp 1635444444
transform 1 0 23276 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_253
timestamp 1635444444
transform 1 0 24380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_265
timestamp 1635444444
transform 1 0 25484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1635444444
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1635444444
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1635444444
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1635444444
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_305
timestamp 1635444444
transform 1 0 29164 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_311
timestamp 1635444444
transform 1 0 29716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_316
timestamp 1635444444
transform 1 0 30176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1635444444
transform -1 0 30820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1635444444
transform 1 0 29808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1635444444
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1635444444
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1635444444
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1635444444
transform 1 0 1840 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1635444444
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_29
timestamp 1635444444
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp 1635444444
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1635444444
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1131_
timestamp 1635444444
transform 1 0 4048 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_45
timestamp 1635444444
transform 1 0 5244 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_49
timestamp 1635444444
transform 1 0 5612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1284_
timestamp 1635444444
transform 1 0 6348 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1672_
timestamp 1635444444
transform 1 0 5336 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_66
timestamp 1635444444
transform 1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_76
timestamp 1635444444
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1635444444
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1635444444
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _1442_
timestamp 1635444444
transform -1 0 8096 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_109
timestamp 1635444444
transform 1 0 11132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1635444444
transform 1 0 9292 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1635444444
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1388_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 10396 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1390_
timestamp 1635444444
transform 1 0 9384 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_32_129
timestamp 1635444444
transform 1 0 12972 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1635444444
transform 1 0 11500 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1635444444
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_149
timestamp 1635444444
transform 1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1635444444
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1635444444
transform -1 0 13616 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_164
timestamp 1635444444
transform 1 0 16192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_168
timestamp 1635444444
transform 1 0 16560 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_172
timestamp 1635444444
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1525_
timestamp 1635444444
transform 1 0 16652 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 15548 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_32_185
timestamp 1635444444
transform 1 0 18124 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1635444444
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1635444444
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1772_
timestamp 1635444444
transform 1 0 17296 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_200
timestamp 1635444444
transform 1 0 19504 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_204
timestamp 1635444444
transform 1 0 19872 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_212
timestamp 1635444444
transform 1 0 20608 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1635444444
transform -1 0 19504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1635_
timestamp 1635444444
transform 1 0 19964 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_32_229
timestamp 1635444444
transform 1 0 22172 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _0913_
timestamp 1635444444
transform -1 0 22172 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_32_241
timestamp 1635444444
transform 1 0 23276 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1635444444
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1635444444
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1635444444
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1635444444
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1635444444
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1635444444
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1635444444
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1635444444
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp 1635444444
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_317
timestamp 1635444444
transform 1 0 30268 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1635444444
transform -1 0 30820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1635444444
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1136_
timestamp 1635444444
transform 1 0 1472 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1135_
timestamp 1635444444
transform 1 0 1564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1635444444
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1635444444
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1635444444
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1635444444
transform 1 0 1380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1635444444
transform 1 0 2668 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_14
timestamp 1635444444
transform 1 0 2392 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_13
timestamp 1635444444
transform 1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1684_
timestamp 1635444444
transform 1 0 3036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_20
timestamp 1635444444
transform 1 0 2944 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_20
timestamp 1635444444
transform 1 0 2944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_28
timestamp 1635444444
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1635444444
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_38
timestamp 1635444444
transform 1 0 4600 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1635444444
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1133_
timestamp 1635444444
transform 1 0 3772 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1635444444
transform 1 0 3772 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_33_45
timestamp 1635444444
transform 1 0 5244 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1635444444
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_57
timestamp 1635444444
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_46
timestamp 1635444444
transform 1 0 5336 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_63
timestamp 1635444444
transform 1 0 6900 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1635444444
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1699_
timestamp 1635444444
transform 1 0 5612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1635444444
transform 1 0 6624 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1635444444
transform -1 0 6900 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__or2b_1  _1425_
timestamp 1635444444
transform 1 0 7912 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 1635444444
transform -1 0 7544 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_70
timestamp 1635444444
transform 1 0 7544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_76
timestamp 1635444444
transform 1 0 8096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1303_
timestamp 1635444444
transform -1 0 10028 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _1278_
timestamp 1635444444
transform -1 0 8924 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1635444444
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1635444444
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1635444444
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_85
timestamp 1635444444
transform 1 0 8924 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_101
timestamp 1635444444
transform 1 0 10396 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1635444444
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_94
timestamp 1635444444
transform 1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1635444444
transform 1 0 10764 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1635444444
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1300_
timestamp 1635444444
transform -1 0 9752 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1301_
timestamp 1635444444
transform 1 0 10120 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1400_
timestamp 1635444444
transform -1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_117
timestamp 1635444444
transform 1 0 11868 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_125
timestamp 1635444444
transform 1 0 12604 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1635444444
transform 1 0 11868 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1635444444
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1635444444
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1188_
timestamp 1635444444
transform -1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1204_
timestamp 1635444444
transform -1 0 11868 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1529_
timestamp 1635444444
transform 1 0 13340 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 13984 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1635444444
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1635444444
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_140
timestamp 1635444444
transform 1 0 13984 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_133
timestamp 1635444444
transform 1 0 13340 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1766_
timestamp 1635444444
transform 1 0 14812 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1765_
timestamp 1635444444
transform -1 0 15456 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_34_141
timestamp 1635444444
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_146
timestamp 1635444444
transform 1 0 14536 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_156
timestamp 1635444444
transform 1 0 15456 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1635444444
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1635444444
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_158
timestamp 1635444444
transform 1 0 15640 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_171
timestamp 1635444444
transform 1 0 16836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1635444444
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1526_
timestamp 1635444444
transform -1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1764_
timestamp 1635444444
transform -1 0 16836 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1785_
timestamp 1635444444
transform 1 0 16836 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1784_
timestamp 1635444444
transform 1 0 17204 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1524_
timestamp 1635444444
transform 1 0 18032 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_34_184
timestamp 1635444444
transform 1 0 18032 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1635444444
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1773_
timestamp 1635444444
transform -1 0 19688 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1606_
timestamp 1635444444
transform 1 0 18400 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_191
timestamp 1635444444
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_189
timestamp 1635444444
transform 1 0 18492 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1635444444
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1635444444
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_202
timestamp 1635444444
transform 1 0 19688 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1635444444
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_204
timestamp 1635444444
transform 1 0 19872 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_210
timestamp 1635444444
transform 1 0 20424 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1620_
timestamp 1635444444
transform 1 0 19228 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1739_
timestamp 1635444444
transform 1 0 20516 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1762_
timestamp 1635444444
transform 1 0 20240 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1635444444
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_234
timestamp 1635444444
transform 1 0 22632 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_220
timestamp 1635444444
transform 1 0 21344 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_229
timestamp 1635444444
transform 1 0 22172 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1635444444
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1040_
timestamp 1635444444
transform -1 0 22172 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1794_
timestamp 1635444444
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_33_246
timestamp 1635444444
transform 1 0 23736 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_258
timestamp 1635444444
transform 1 0 24840 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_241
timestamp 1635444444
transform 1 0 23276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1635444444
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1635444444
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1635444444
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_270
timestamp 1635444444
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1635444444
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1635444444
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1635444444
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1635444444
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1635444444
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1635444444
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1635444444
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1635444444
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1635444444
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_317
timestamp 1635444444
transform 1 0 30268 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1635444444
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1635444444
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_317
timestamp 1635444444
transform 1 0 30268 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1635444444
transform -1 0 30820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1635444444
transform -1 0 30820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1635444444
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1635444444
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1635444444
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1635444444
transform 1 0 1932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_25
timestamp 1635444444
transform 1 0 3404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1635444444
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1635444444
transform 1 0 3772 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1635444444
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_65
timestamp 1635444444
transform 1 0 7084 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1635444444
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1281_
timestamp 1635444444
transform -1 0 7084 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_69
timestamp 1635444444
transform 1 0 7452 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_74
timestamp 1635444444
transform 1 0 7912 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_86
timestamp 1635444444
transform 1 0 9016 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1308_
timestamp 1635444444
transform 1 0 8280 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1397_
timestamp 1635444444
transform -1 0 7912 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_106
timestamp 1635444444
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1635444444
transform 1 0 9384 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_35_122
timestamp 1635444444
transform 1 0 12328 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1635444444
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1216_
timestamp 1635444444
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_35_134
timestamp 1635444444
transform 1 0 13432 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_146
timestamp 1635444444
transform 1 0 14536 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1763_
timestamp 1635444444
transform 1 0 14904 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1635444444
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1635444444
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1635444444
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1537_
timestamp 1635444444
transform 1 0 16652 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1635444444
transform 1 0 17480 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_191
timestamp 1635444444
transform 1 0 18676 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _1622_
timestamp 1635444444
transform 1 0 19044 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1798_
timestamp 1635444444
transform 1 0 17848 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1635444444
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_211
timestamp 1635444444
transform 1 0 20516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1635444444
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1635444444
transform -1 0 21160 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1636_
timestamp 1635444444
transform 1 0 20056 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1635444444
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1635444444
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1635444444
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1635444444
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1635444444
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1635444444
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1635444444
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1635444444
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1635444444
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1635444444
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_305
timestamp 1635444444
transform 1 0 29164 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_311
timestamp 1635444444
transform 1 0 29716 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_316
timestamp 1635444444
transform 1 0 30176 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1635444444
transform -1 0 30820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1635444444
transform 1 0 29808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1635444444
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1635444444
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1635444444
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1635444444
transform 1 0 1840 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1635444444
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp 1635444444
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_40
timestamp 1635444444
transform 1 0 4784 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1635444444
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1267_
timestamp 1635444444
transform -1 0 4784 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_52
timestamp 1635444444
transform 1 0 5888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_58
timestamp 1635444444
transform 1 0 6440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_62
timestamp 1635444444
transform 1 0 6808 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1386_
timestamp 1635444444
transform 1 0 6532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_66
timestamp 1635444444
transform 1 0 7176 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_71
timestamp 1635444444
transform 1 0 7636 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1635444444
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_85
timestamp 1635444444
transform 1 0 8924 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1635444444
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1635444444
transform -1 0 8464 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1387_
timestamp 1635444444
transform -1 0 9384 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_wb_clk_i
timestamp 1635444444
transform 1 0 7268 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_90
timestamp 1635444444
transform 1 0 9384 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1635444444
transform 1 0 9752 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1635444444
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_130
timestamp 1635444444
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1635444444
transform 1 0 11592 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1635444444
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1635444444
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_149
timestamp 1635444444
transform 1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1635444444
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_1  _1536_
timestamp 1635444444
transform 1 0 15088 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_158
timestamp 1635444444
transform 1 0 15640 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_166
timestamp 1635444444
transform 1 0 16376 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_174
timestamp 1635444444
transform 1 0 17112 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_1  _1538_
timestamp 1635444444
transform 1 0 16468 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_36_182
timestamp 1635444444
transform 1 0 17848 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1635444444
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1635444444
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1781_
timestamp 1635444444
transform 1 0 17940 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_206
timestamp 1635444444
transform 1 0 20056 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_216
timestamp 1635444444
transform 1 0 20976 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1041_
timestamp 1635444444
transform -1 0 20976 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1777_
timestamp 1635444444
transform 1 0 19228 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_36_222
timestamp 1635444444
transform 1 0 21528 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_228
timestamp 1635444444
transform 1 0 22080 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_235
timestamp 1635444444
transform 1 0 22724 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1635444444
transform 1 0 22448 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1035_
timestamp 1635444444
transform -1 0 22080 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_36_247
timestamp 1635444444
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1635444444
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1635444444
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1635444444
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1635444444
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1635444444
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1635444444
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1635444444
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1635444444
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_309
timestamp 1635444444
transform 1 0 29532 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_317
timestamp 1635444444
transform 1 0 30268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1635444444
transform -1 0 30820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1635444444
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_13
timestamp 1635444444
transform 1 0 2300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_20
timestamp 1635444444
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_6
timestamp 1635444444
transform 1 0 1656 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1635444444
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1635444444
transform -1 0 1656 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1635444444
transform 1 0 2024 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1635444444
transform -1 0 2944 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_32
timestamp 1635444444
transform 1 0 4048 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1268_
timestamp 1635444444
transform -1 0 5336 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_37_46
timestamp 1635444444
transform 1 0 5336 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1635444444
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1635444444
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1272_
timestamp 1635444444
transform 1 0 6348 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_37_67
timestamp 1635444444
transform 1 0 7268 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_80
timestamp 1635444444
transform 1 0 8464 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1391_
timestamp 1635444444
transform -1 0 8464 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_37_100
timestamp 1635444444
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_88
timestamp 1635444444
transform 1 0 9200 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1302_
timestamp 1635444444
transform -1 0 10304 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1635444444
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_121
timestamp 1635444444
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1635444444
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1635444444
transform 1 0 12420 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_37_139
timestamp 1635444444
transform 1 0 13892 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1635444444
transform -1 0 15732 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_37_159
timestamp 1635444444
transform 1 0 15732 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1635444444
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1635444444
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1812_
timestamp 1635444444
transform -1 0 17480 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_37_178
timestamp 1635444444
transform 1 0 17480 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_184
timestamp 1635444444
transform 1 0 18032 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_190
timestamp 1635444444
transform 1 0 18584 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1531_
timestamp 1635444444
transform 1 0 18952 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1621_
timestamp 1635444444
transform 1 0 18124 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_37_197
timestamp 1635444444
transform 1 0 19228 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_201
timestamp 1635444444
transform 1 0 19596 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_205
timestamp 1635444444
transform 1 0 19964 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1635444444
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1635444444
transform -1 0 19964 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1042_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 20976 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_37_230
timestamp 1635444444
transform 1 0 22264 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_239
timestamp 1635444444
transform 1 0 23092 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1635444444
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0911_
timestamp 1635444444
transform 1 0 21804 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1033_
timestamp 1635444444
transform -1 0 23092 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_37_251
timestamp 1635444444
transform 1 0 24196 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_263
timestamp 1635444444
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1635444444
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1635444444
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1635444444
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1635444444
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1635444444
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1635444444
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_317
timestamp 1635444444
transform 1 0 30268 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1635444444
transform -1 0 30820 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_13
timestamp 1635444444
transform 1 0 2300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_6
timestamp 1635444444
transform 1 0 1656 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1635444444
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1635444444
transform -1 0 1656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1635444444
transform -1 0 2300 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1635444444
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1635444444
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1635444444
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1635444444
transform 1 0 4048 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_48
timestamp 1635444444
transform 1 0 5520 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1635444444
transform 1 0 5888 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_68
timestamp 1635444444
transform 1 0 7360 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_75
timestamp 1635444444
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1635444444
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_85
timestamp 1635444444
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1635444444
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1385_
timestamp 1635444444
transform 1 0 7728 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_105
timestamp 1635444444
transform 1 0 10764 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_97
timestamp 1635444444
transform 1 0 10028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1218_
timestamp 1635444444
transform 1 0 10856 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1309_
timestamp 1635444444
transform 1 0 9200 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_115
timestamp 1635444444
transform 1 0 11684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_128
timestamp 1635444444
transform 1 0 12880 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _1202_
timestamp 1635444444
transform 1 0 12052 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1635444444
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_145
timestamp 1635444444
transform 1 0 14444 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_151
timestamp 1635444444
transform 1 0 14996 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1635444444
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1607_
timestamp 1635444444
transform 1 0 14536 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_38_158
timestamp 1635444444
transform 1 0 15640 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_171
timestamp 1635444444
transform 1 0 16836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1543_
timestamp 1635444444
transform 1 0 15364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1557_
timestamp 1635444444
transform 1 0 16008 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_38_183
timestamp 1635444444
transform 1 0 17940 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_188
timestamp 1635444444
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1635444444
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1530_
timestamp 1635444444
transform -1 0 18400 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1635444444
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1635444444
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_214
timestamp 1635444444
transform 1 0 20792 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_4  _0894_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 21988 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1635444444
transform 1 0 19412 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1039_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 20792 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_227
timestamp 1635444444
transform 1 0 21988 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_238
timestamp 1635444444
transform 1 0 23000 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0892_
timestamp 1635444444
transform -1 0 23000 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1635444444
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1635444444
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1635444444
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1635444444
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0912_
timestamp 1635444444
transform 1 0 23368 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1635444444
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1635444444
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1635444444
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1635444444
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1635444444
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_309
timestamp 1635444444
transform 1 0 29532 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_316
timestamp 1635444444
transform 1 0 30176 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1635444444
transform -1 0 30820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1635444444
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1635444444
transform 1 0 29808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1635444444
transform -1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1635444444
transform 1 0 1380 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1635444444
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1635444444
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_7
timestamp 1635444444
transform 1 0 1748 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1392_
timestamp 1635444444
transform -1 0 2944 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1635444444
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_15
timestamp 1635444444
transform 1 0 2484 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_17
timestamp 1635444444
transform 1 0 2668 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_13
timestamp 1635444444
transform 1 0 2300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1635444444
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1635444444
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_38
timestamp 1635444444
transform 1 0 4600 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1635444444
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1275_
timestamp 1635444444
transform -1 0 4600 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1276_
timestamp 1635444444
transform -1 0 5428 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1398_
timestamp 1635444444
transform 1 0 4968 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1635444444
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1635444444
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_45
timestamp 1635444444
transform 1 0 5244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_58
timestamp 1635444444
transform 1 0 6440 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1635444444
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1280_
timestamp 1635444444
transform 1 0 5612 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1282_
timestamp 1635444444
transform 1 0 6348 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1402_
timestamp 1635444444
transform 1 0 7360 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1401_
timestamp 1635444444
transform 1 0 7636 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_40_66
timestamp 1635444444
transform 1 0 7176 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_70
timestamp 1635444444
transform 1 0 7544 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_66
timestamp 1635444444
transform 1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1396_
timestamp 1635444444
transform -1 0 9200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1635444444
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1635444444
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1635444444
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_78
timestamp 1635444444
transform 1 0 8280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1306_
timestamp 1635444444
transform 1 0 9108 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_39_86
timestamp 1635444444
transform 1 0 9016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_103
timestamp 1635444444
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_96
timestamp 1635444444
transform 1 0 9936 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_88
timestamp 1635444444
transform 1 0 9200 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1208_
timestamp 1635444444
transform -1 0 10580 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1635444444
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_wb_clk_i
timestamp 1635444444
transform -1 0 12052 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1190_
timestamp 1635444444
transform 1 0 12052 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1635444444
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_118
timestamp 1635444444
transform 1 0 11960 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_110
timestamp 1635444444
transform 1 0 11224 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_119
timestamp 1635444444
transform 1 0 12052 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1635444444
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1635444444
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_127
timestamp 1635444444
transform 1 0 12788 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1635444444
transform 1 0 12880 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_40_128
timestamp 1635444444
transform 1 0 12880 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_144
timestamp 1635444444
transform 1 0 14352 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_151
timestamp 1635444444
transform 1 0 14996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_141
timestamp 1635444444
transform 1 0 14076 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_145
timestamp 1635444444
transform 1 0 14444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1635444444
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1544_
timestamp 1635444444
transform 1 0 14720 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 14444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1630_
timestamp 1635444444
transform 1 0 14812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1635444444
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_157
timestamp 1635444444
transform 1 0 15548 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_170
timestamp 1635444444
transform 1 0 16744 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1635444444
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_2  _1558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1769_
timestamp 1635444444
transform -1 0 17940 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1783_
timestamp 1635444444
transform -1 0 16192 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1813_
timestamp 1635444444
transform -1 0 16744 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_39_181
timestamp 1635444444
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_194
timestamp 1635444444
transform 1 0 18952 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_183
timestamp 1635444444
transform 1 0 17940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_187
timestamp 1635444444
transform 1 0 18308 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1635444444
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1635444444
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1635444444
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1533_
timestamp 1635444444
transform -1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1797_
timestamp 1635444444
transform 1 0 18124 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_39_211
timestamp 1635444444
transform 1 0 20516 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1635444444
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_201
timestamp 1635444444
transform 1 0 19596 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_205
timestamp 1635444444
transform 1 0 19964 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_212
timestamp 1635444444
transform 1 0 20608 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1635444444
transform 1 0 21068 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1037_
timestamp 1635444444
transform -1 0 20516 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1635444444
transform -1 0 19964 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1527_
timestamp 1635444444
transform 1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1635444444
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_225
timestamp 1635444444
transform 1 0 21804 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1635444444
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_224
timestamp 1635444444
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_234
timestamp 1635444444
transform 1 0 22632 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1635444444
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0886_
timestamp 1635444444
transform -1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0893_
timestamp 1635444444
transform 1 0 22632 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1795_
timestamp 1635444444
transform 1 0 21804 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_39_244
timestamp 1635444444
transform 1 0 23552 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_256
timestamp 1635444444
transform 1 0 24656 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1635444444
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1635444444
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1635444444
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_268
timestamp 1635444444
transform 1 0 25760 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1635444444
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1635444444
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1635444444
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1635444444
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1635444444
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1635444444
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1635444444
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1635444444
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_39_317
timestamp 1635444444
transform 1 0 30268 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1635444444
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_309
timestamp 1635444444
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_317
timestamp 1635444444
transform 1 0 30268 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1635444444
transform -1 0 30820 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1635444444
transform -1 0 30820 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1635444444
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_15
timestamp 1635444444
transform 1 0 2484 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_20
timestamp 1635444444
transform 1 0 2944 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_7
timestamp 1635444444
transform 1 0 1748 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1635444444
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1403_
timestamp 1635444444
transform -1 0 2944 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1635444444
transform -1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_41
timestamp 1635444444
transform 1 0 4876 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1273_
timestamp 1635444444
transform 1 0 4048 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_41_47
timestamp 1635444444
transform 1 0 5428 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1635444444
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1635444444
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_63
timestamp 1635444444
transform 1 0 6900 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1635444444
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1635444444
transform -1 0 6900 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_wb_clk_i
timestamp 1635444444
transform -1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_76
timestamp 1635444444
transform 1 0 8096 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_80
timestamp 1635444444
transform 1 0 8464 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1419_
timestamp 1635444444
transform 1 0 8556 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1787_
timestamp 1635444444
transform 1 0 7268 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1635444444
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_90
timestamp 1635444444
transform 1 0 9384 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_98
timestamp 1635444444
transform 1 0 10120 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1214_
timestamp 1635444444
transform 1 0 10212 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_41_129
timestamp 1635444444
transform 1 0 12972 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1635444444
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1635444444
transform 1 0 11500 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_41_141
timestamp 1635444444
transform 1 0 14076 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_147
timestamp 1635444444
transform 1 0 14628 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _1609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 15272 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_154
timestamp 1635444444
transform 1 0 15272 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1635444444
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1635444444
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1635444444
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1635444444
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1628_
timestamp 1635444444
transform 1 0 15640 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_177
timestamp 1635444444
transform 1 0 17388 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_187
timestamp 1635444444
transform 1 0 18308 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1532_
timestamp 1635444444
transform -1 0 19228 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1770_
timestamp 1635444444
transform -1 0 18308 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_41_197
timestamp 1635444444
transform 1 0 19228 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_205
timestamp 1635444444
transform 1 0 19964 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1635444444
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1050_
timestamp 1635444444
transform 1 0 19596 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1051_
timestamp 1635444444
transform 1 0 20332 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1635444444
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1635444444
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1635444444
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1635444444
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1635444444
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1635444444
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1635444444
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1635444444
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1635444444
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1635444444
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1635444444
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1635444444
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_317
timestamp 1635444444
transform 1 0 30268 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1635444444
transform -1 0 30820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1635444444
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1635444444
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1635444444
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1635444444
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_29
timestamp 1635444444
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_33
timestamp 1635444444
transform 1 0 4140 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1635444444
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1860_
timestamp 1635444444
transform 1 0 4232 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_42_51
timestamp 1635444444
transform 1 0 5796 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1635444444
transform 1 0 6164 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_42_71
timestamp 1635444444
transform 1 0 7636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_75
timestamp 1635444444
transform 1 0 8004 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_79
timestamp 1635444444
transform 1 0 8372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1635444444
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1635444444
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1399_
timestamp 1635444444
transform -1 0 8372 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1418_
timestamp 1635444444
transform 1 0 8924 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_42_100
timestamp 1635444444
transform 1 0 10304 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 1635444444
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_92
timestamp 1635444444
transform 1 0 9568 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1212_
timestamp 1635444444
transform -1 0 11132 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_42_117
timestamp 1635444444
transform 1 0 11868 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_128
timestamp 1635444444
transform 1 0 12880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1200_
timestamp 1635444444
transform 1 0 12052 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 1635444444
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1635444444
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1635444444
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_145
timestamp 1635444444
transform 1 0 14444 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_150
timestamp 1635444444
transform 1 0 14904 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1635444444
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1587_
timestamp 1635444444
transform 1 0 13248 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_wb_clk_i
timestamp 1635444444
transform 1 0 14536 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_157
timestamp 1635444444
transform 1 0 15548 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_165
timestamp 1635444444
transform 1 0 16284 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1629_
timestamp 1635444444
transform 1 0 15272 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1780_
timestamp 1635444444
transform -1 0 17388 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_177
timestamp 1635444444
transform 1 0 17388 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1635444444
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1635444444
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1809_
timestamp 1635444444
transform 1 0 17756 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_42_197
timestamp 1635444444
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_208
timestamp 1635444444
transform 1 0 20240 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1056_
timestamp 1635444444
transform 1 0 19504 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1058_
timestamp 1635444444
transform 1 0 20608 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_221
timestamp 1635444444
transform 1 0 21436 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1635444444
transform 1 0 21804 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_42_241
timestamp 1635444444
transform 1 0 23276 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1635444444
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1635444444
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1635444444
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1635444444
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1635444444
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1635444444
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1635444444
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1635444444
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_309
timestamp 1635444444
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_316
timestamp 1635444444
transform 1 0 30176 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1635444444
transform -1 0 30820 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1635444444
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1635444444
transform 1 0 29808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_15
timestamp 1635444444
transform 1 0 2484 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_20
timestamp 1635444444
transform 1 0 2944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_7
timestamp 1635444444
transform 1 0 1748 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1635444444
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1420_
timestamp 1635444444
transform -1 0 2944 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1635444444
transform -1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_28
timestamp 1635444444
transform 1 0 3680 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_37
timestamp 1635444444
transform 1 0 4508 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1274_
timestamp 1635444444
transform -1 0 4508 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1415_
timestamp 1635444444
transform 1 0 4876 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_44
timestamp 1635444444
transform 1 0 5152 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1635444444
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1635444444
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1635444444
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1793_
timestamp 1635444444
transform 1 0 6532 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_wb_clk_i
timestamp 1635444444
transform -1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_68
timestamp 1635444444
transform 1 0 7360 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_79
timestamp 1635444444
transform 1 0 8372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1409_
timestamp 1635444444
transform 1 0 7728 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1792_
timestamp 1635444444
transform 1 0 8924 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_43_101
timestamp 1635444444
transform 1 0 10396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1635444444
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_94
timestamp 1635444444
transform 1 0 9752 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1407_
timestamp 1635444444
transform -1 0 10396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1408_
timestamp 1635444444
transform -1 0 11040 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_122
timestamp 1635444444
transform 1 0 12328 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_126
timestamp 1635444444
transform 1 0 12696 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1635444444
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1199_
timestamp 1635444444
transform -1 0 12328 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1635444444
transform -1 0 14260 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_43_143
timestamp 1635444444
transform 1 0 14260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_152
timestamp 1635444444
transform 1 0 15088 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1567_
timestamp 1635444444
transform 1 0 14812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_158
timestamp 1635444444
transform 1 0 15640 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1635444444
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1635444444
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1556_
timestamp 1635444444
transform 1 0 15732 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1775_
timestamp 1635444444
transform 1 0 16652 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_43_178
timestamp 1635444444
transform 1 0 17480 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_186
timestamp 1635444444
transform 1 0 18216 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_196
timestamp 1635444444
transform 1 0 19136 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1806_
timestamp 1635444444
transform 1 0 18308 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_43_200
timestamp 1635444444
transform 1 0 19504 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_207
timestamp 1635444444
transform 1 0 20148 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1052_
timestamp 1635444444
transform 1 0 20516 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o211ai_1  _1057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 19596 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1635444444
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1635444444
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1952_
timestamp 1635444444
transform 1 0 21804 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_43_241
timestamp 1635444444
transform 1 0 23276 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_253
timestamp 1635444444
transform 1 0 24380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_265
timestamp 1635444444
transform 1 0 25484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1635444444
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1635444444
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1635444444
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1635444444
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1635444444
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_317
timestamp 1635444444
transform 1 0 30268 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1635444444
transform -1 0 30820 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_15
timestamp 1635444444
transform 1 0 2484 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1635444444
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_7
timestamp 1635444444
transform 1 0 1748 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1635444444
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1411_
timestamp 1635444444
transform -1 0 2944 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1635444444
transform -1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_29
timestamp 1635444444
transform 1 0 3772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_33
timestamp 1635444444
transform 1 0 4140 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_42
timestamp 1635444444
transform 1 0 4968 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1635444444
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1269_
timestamp 1635444444
transform 1 0 4232 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_50
timestamp 1635444444
transform 1 0 5704 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_58
timestamp 1635444444
transform 1 0 6440 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1196_
timestamp 1635444444
transform -1 0 6440 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1735_
timestamp 1635444444
transform 1 0 6992 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_73
timestamp 1635444444
transform 1 0 7820 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1635444444
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_85
timestamp 1635444444
transform 1 0 8924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1635444444
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1406_
timestamp 1635444444
transform -1 0 8464 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_104
timestamp 1635444444
transform 1 0 10672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_96
timestamp 1635444444
transform 1 0 9936 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1307_
timestamp 1635444444
transform 1 0 9200 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1414_
timestamp 1635444444
transform -1 0 11316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1635444444
transform -1 0 10672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_111
timestamp 1635444444
transform 1 0 11316 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_126
timestamp 1635444444
transform 1 0 12696 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1197_
timestamp 1635444444
transform 1 0 11868 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1635444444
transform -1 0 13432 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1635444444
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1635444444
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_148
timestamp 1635444444
transform 1 0 14720 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1635444444
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1545_
timestamp 1635444444
transform 1 0 15088 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1589_
timestamp 1635444444
transform 1 0 14260 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_44_155
timestamp 1635444444
transform 1 0 15364 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_162
timestamp 1635444444
transform 1 0 16008 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1546_
timestamp 1635444444
transform 1 0 15732 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1600_
timestamp 1635444444
transform 1 0 17112 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_44_179
timestamp 1635444444
transform 1 0 17572 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1635444444
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1635444444
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1807_
timestamp 1635444444
transform 1 0 17940 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_44_200
timestamp 1635444444
transform 1 0 19504 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_208
timestamp 1635444444
transform 1 0 20240 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_217
timestamp 1635444444
transform 1 0 21068 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1054_
timestamp 1635444444
transform -1 0 21068 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1588_
timestamp 1635444444
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_233
timestamp 1635444444
transform 1 0 22540 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_240
timestamp 1635444444
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1635444444
transform -1 0 23184 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0889_
timestamp 1635444444
transform 1 0 21620 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1635444444
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1635444444
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1635444444
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1635444444
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1635444444
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1635444444
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1635444444
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_309
timestamp 1635444444
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_317
timestamp 1635444444
transform 1 0 30268 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1635444444
transform -1 0 30820 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1635444444
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_19
timestamp 1635444444
transform 1 0 2852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_7
timestamp 1635444444
transform 1 0 1748 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1635444444
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1635444444
transform -1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_23
timestamp 1635444444
transform 1 0 3220 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_40
timestamp 1635444444
transform 1 0 4784 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1635444444
transform 1 0 3312 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_45_44
timestamp 1635444444
transform 1 0 5152 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1635444444
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_57
timestamp 1635444444
transform 1 0 6348 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_63
timestamp 1635444444
transform 1 0 6900 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1635444444
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1191_
timestamp 1635444444
transform 1 0 6624 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1198_
timestamp 1635444444
transform -1 0 5888 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_76
timestamp 1635444444
transform 1 0 8096 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_84
timestamp 1635444444
transform 1 0 8832 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1410_
timestamp 1635444444
transform -1 0 8096 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1635444444
transform -1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1635444444
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_90
timestamp 1635444444
transform 1 0 9384 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1841_
timestamp 1635444444
transform 1 0 9476 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_45_116
timestamp 1635444444
transform 1 0 11776 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1635444444
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1416_
timestamp 1635444444
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1635444444
transform 1 0 12512 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_45_140
timestamp 1635444444
transform 1 0 13984 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1568_
timestamp 1635444444
transform -1 0 15364 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_155
timestamp 1635444444
transform 1 0 15364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1635444444
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_172
timestamp 1635444444
transform 1 0 16928 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1635444444
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1569_
timestamp 1635444444
transform 1 0 15732 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1570_
timestamp 1635444444
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_179
timestamp 1635444444
transform 1 0 17572 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_191
timestamp 1635444444
transform 1 0 18676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1602_
timestamp 1635444444
transform 1 0 17940 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1603_
timestamp 1635444444
transform -1 0 17572 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_197
timestamp 1635444444
transform 1 0 19228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_202
timestamp 1635444444
transform 1 0 19688 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_212
timestamp 1635444444
transform 1 0 20608 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1045_
timestamp 1635444444
transform -1 0 20608 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1055_
timestamp 1635444444
transform 1 0 19320 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_230
timestamp 1635444444
transform 1 0 22264 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1635444444
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0888_
timestamp 1635444444
transform -1 0 22264 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_45_242
timestamp 1635444444
transform 1 0 23368 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_254
timestamp 1635444444
transform 1 0 24472 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_266
timestamp 1635444444
transform 1 0 25576 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1635444444
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1635444444
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1635444444
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1635444444
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1635444444
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_317
timestamp 1635444444
transform 1 0 30268 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1635444444
transform -1 0 30820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1635444444
transform -1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1635444444
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1635444444
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_7
timestamp 1635444444
transform 1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1433_
timestamp 1635444444
transform 1 0 2116 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1427_
timestamp 1635444444
transform -1 0 2852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1083_
timestamp 1635444444
transform -1 0 3128 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_14
timestamp 1635444444
transform 1 0 2392 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_19
timestamp 1635444444
transform 1 0 2852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_15
timestamp 1635444444
transform 1 0 2484 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1635444444
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1082_
timestamp 1635444444
transform -1 0 4232 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1635444444
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_22
timestamp 1635444444
transform 1 0 3128 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_29
timestamp 1635444444
transform 1 0 3772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1635444444
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1444_
timestamp 1635444444
transform -1 0 4876 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_41
timestamp 1635444444
transform 1 0 4876 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_34
timestamp 1635444444
transform 1 0 4232 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_35
timestamp 1635444444
transform 1 0 4324 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1861_
timestamp 1635444444
transform 1 0 4416 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_4  _0980_
timestamp 1635444444
transform 1 0 5336 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_45
timestamp 1635444444
transform 1 0 5244 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1635444444
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1635444444
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_52
timestamp 1635444444
transform 1 0 5888 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_53
timestamp 1635444444
transform 1 0 5980 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1635444444
transform -1 0 6900 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1438_
timestamp 1635444444
transform 1 0 6808 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_61
timestamp 1635444444
transform 1 0 6716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_63
timestamp 1635444444
transform 1 0 6900 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_65
timestamp 1635444444
transform 1 0 7084 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1437_
timestamp 1635444444
transform -1 0 7820 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1432_
timestamp 1635444444
transform 1 0 7452 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_46_73
timestamp 1635444444
transform 1 0 7820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1431_
timestamp 1635444444
transform -1 0 8464 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1426_
timestamp 1635444444
transform 1 0 8464 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1635444444
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_76
timestamp 1635444444
transform 1 0 8096 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1635444444
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1635444444
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1304_
timestamp 1635444444
transform 1 0 9108 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_103
timestamp 1635444444
transform 1 0 10580 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_108
timestamp 1635444444
transform 1 0 11040 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_95
timestamp 1635444444
transform 1 0 9844 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_101
timestamp 1635444444
transform 1 0 10396 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1635444444
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_89
timestamp 1635444444
transform 1 0 9292 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1192_
timestamp 1635444444
transform -1 0 11040 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1305_
timestamp 1635444444
transform 1 0 9660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1424_
timestamp 1635444444
transform -1 0 11040 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_128
timestamp 1635444444
transform 1 0 12880 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_116
timestamp 1635444444
transform 1 0 11776 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_124
timestamp 1635444444
transform 1 0 12512 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1635444444
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1195_
timestamp 1635444444
transform -1 0 12512 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1417_
timestamp 1635444444
transform 1 0 11500 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1635444444
transform 1 0 11408 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1635444444
transform 1 0 13064 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_46_141
timestamp 1635444444
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_150
timestamp 1635444444
transform 1 0 14904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_146
timestamp 1635444444
transform 1 0 14536 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1635444444
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1590_
timestamp 1635444444
transform 1 0 14904 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1591_
timestamp 1635444444
transform -1 0 14904 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1592_
timestamp 1635444444
transform 1 0 15272 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1580_
timestamp 1635444444
transform 1 0 15732 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_47_153
timestamp 1635444444
transform 1 0 15180 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_162
timestamp 1635444444
transform 1 0 16008 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_158
timestamp 1635444444
transform 1 0 15640 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1803_
timestamp 1635444444
transform 1 0 16100 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1635444444
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1635444444
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1635444444
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_172
timestamp 1635444444
transform 1 0 16928 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1796_
timestamp 1635444444
transform 1 0 17020 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_46_179
timestamp 1635444444
transform 1 0 17572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1635444444
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_182
timestamp 1635444444
transform 1 0 17848 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_195
timestamp 1635444444
transform 1 0 19044 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1635444444
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1565_
timestamp 1635444444
transform 1 0 17296 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1599_
timestamp 1635444444
transform 1 0 18400 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1601_
timestamp 1635444444
transform 1 0 17940 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_46_206
timestamp 1635444444
transform 1 0 20056 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_218
timestamp 1635444444
transform 1 0 21160 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_207
timestamp 1635444444
transform 1 0 20148 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_216
timestamp 1635444444
transform 1 0 20976 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1047_
timestamp 1635444444
transform -1 0 21160 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_1  _1048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 20332 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1811_
timestamp 1635444444
transform 1 0 19228 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_46_225
timestamp 1635444444
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1635444444
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_230
timestamp 1635444444
transform 1 0 22264 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1635444444
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1031_
timestamp 1635444444
transform -1 0 22264 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1635444444
transform 1 0 21528 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1635444444
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1635444444
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_242
timestamp 1635444444
transform 1 0 23368 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_254
timestamp 1635444444
transform 1 0 24472 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1635444444
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1635444444
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1635444444
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_266
timestamp 1635444444
transform 1 0 25576 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1635444444
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1635444444
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1635444444
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1635444444
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1635444444
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1635444444
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_305
timestamp 1635444444
transform 1 0 29164 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1635444444
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1635444444
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1635444444
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1635444444
transform 1 0 29808 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1363_
timestamp 1635444444
transform 1 0 29808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_311
timestamp 1635444444
transform 1 0 29716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1635444444
transform -1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1635444444
transform -1 0 30820 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_316
timestamp 1635444444
transform 1 0 30176 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_316
timestamp 1635444444
transform 1 0 30176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_15
timestamp 1635444444
transform 1 0 2484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1635444444
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_7
timestamp 1635444444
transform 1 0 1748 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1635444444
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1439_
timestamp 1635444444
transform -1 0 2852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1635444444
transform -1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1635444444
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_32
timestamp 1635444444
transform 1 0 4048 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_40
timestamp 1635444444
transform 1 0 4784 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1635444444
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3772 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1635444444
transform -1 0 5244 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_45
timestamp 1635444444
transform 1 0 5244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_52
timestamp 1635444444
transform 1 0 5888 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_56
timestamp 1635444444
transform 1 0 6256 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1635444444
transform -1 0 5888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1789_
timestamp 1635444444
transform 1 0 6348 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_66
timestamp 1635444444
transform 1 0 7176 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_79
timestamp 1635444444
transform 1 0 8372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1635444444
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1635444444
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1423_
timestamp 1635444444
transform -1 0 9200 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1786_
timestamp 1635444444
transform 1 0 7544 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_48_88
timestamp 1635444444
transform 1 0 9200 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1635444444
transform 1 0 9936 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_112
timestamp 1635444444
transform 1 0 11408 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_120
timestamp 1635444444
transform 1 0 12144 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1194_
timestamp 1635444444
transform 1 0 12696 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1635444444
transform 1 0 11776 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_134
timestamp 1635444444
transform 1 0 13432 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1635444444
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_149
timestamp 1635444444
transform 1 0 14812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1635444444
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0900_
timestamp 1635444444
transform 1 0 14444 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_158
timestamp 1635444444
transform 1 0 15640 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_166
timestamp 1635444444
transform 1 0 16376 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1635444444
transform 1 0 15180 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1799_
timestamp 1635444444
transform 1 0 16468 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_48_176
timestamp 1635444444
transform 1 0 17296 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_182
timestamp 1635444444
transform 1 0 17848 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1635444444
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1635444444
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1760_
timestamp 1635444444
transform -1 0 18768 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1635444444
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_201
timestamp 1635444444
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_206
timestamp 1635444444
transform 1 0 20056 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_214
timestamp 1635444444
transform 1 0 20792 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_218
timestamp 1635444444
transform 1 0 21160 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1032_
timestamp 1635444444
transform 1 0 19688 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1365_
timestamp 1635444444
transform 1 0 20424 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_236
timestamp 1635444444
transform 1 0 22816 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _1954_
timestamp 1635444444
transform 1 0 21252 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1635444444
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1635444444
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1635444444
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1635444444
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1635444444
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1635444444
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1635444444
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1635444444
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_309
timestamp 1635444444
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_317
timestamp 1635444444
transform 1 0 30268 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1635444444
transform -1 0 30820 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1635444444
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_15
timestamp 1635444444
transform 1 0 2484 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_7
timestamp 1635444444
transform 1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1635444444
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1635444444
transform -1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1635444444
transform 1 0 2116 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_23
timestamp 1635444444
transform 1 0 3220 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_28
timestamp 1635444444
transform 1 0 3680 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_35
timestamp 1635444444
transform 1 0 4324 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1330_
timestamp 1635444444
transform -1 0 3680 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1332_
timestamp 1635444444
transform -1 0 4324 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1338_
timestamp 1635444444
transform 1 0 5060 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_46
timestamp 1635444444
transform 1 0 5336 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1635444444
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_57
timestamp 1635444444
transform 1 0 6348 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1635444444
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1790_
timestamp 1635444444
transform 1 0 6624 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_69
timestamp 1635444444
transform 1 0 7452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_76
timestamp 1635444444
transform 1 0 8096 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_82
timestamp 1635444444
transform 1 0 8648 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1405_
timestamp 1635444444
transform 1 0 7820 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1791_
timestamp 1635444444
transform 1 0 8740 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_92
timestamp 1635444444
transform 1 0 9568 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_99
timestamp 1635444444
transform 1 0 10212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1429_
timestamp 1635444444
transform 1 0 9936 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1635444444
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_113
timestamp 1635444444
transform 1 0 11500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_119
timestamp 1635444444
transform 1 0 12052 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_127
timestamp 1635444444
transform 1 0 12788 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1635444444
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1635444444
transform -1 0 12052 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1187_
timestamp 1635444444
transform -1 0 12788 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1201_
timestamp 1635444444
transform -1 0 13892 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_139
timestamp 1635444444
transform 1 0 13892 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_145
timestamp 1635444444
transform 1 0 14444 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_150
timestamp 1635444444
transform 1 0 14904 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0916_
timestamp 1635444444
transform -1 0 14904 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_158
timestamp 1635444444
transform 1 0 15640 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1635444444
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1635444444
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1566_
timestamp 1635444444
transform 1 0 15916 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1581_
timestamp 1635444444
transform 1 0 16652 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_178
timestamp 1635444444
transform 1 0 17480 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_188
timestamp 1635444444
transform 1 0 18400 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__o211ai_1  _1582_
timestamp 1635444444
transform -1 0 18400 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_200
timestamp 1635444444
transform 1 0 19504 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_208
timestamp 1635444444
transform 1 0 20240 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1635444444
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1366_
timestamp 1635444444
transform -1 0 21068 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1635444444
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_225
timestamp 1635444444
transform 1 0 21804 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_232
timestamp 1635444444
transform 1 0 22448 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1635444444
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1368_
timestamp 1635444444
transform -1 0 22448 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1825_
timestamp 1635444444
transform 1 0 22816 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_49_253
timestamp 1635444444
transform 1 0 24380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_265
timestamp 1635444444
transform 1 0 25484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1635444444
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1635444444
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1635444444
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1635444444
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_305
timestamp 1635444444
transform 1 0 29164 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_311
timestamp 1635444444
transform 1 0 29716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_316
timestamp 1635444444
transform 1 0 30176 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1635444444
transform -1 0 30820 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1635444444
transform 1 0 29808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_17
timestamp 1635444444
transform 1 0 2668 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_6
timestamp 1635444444
transform 1 0 1656 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1635444444
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1329_
timestamp 1635444444
transform 1 0 3036 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1447_
timestamp 1635444444
transform -1 0 1656 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1450_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2024 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1635444444
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_29
timestamp 1635444444
transform 1 0 3772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1635444444
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1635444444
transform 1 0 4140 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_49
timestamp 1635444444
transform 1 0 5612 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_56
timestamp 1635444444
transform 1 0 6256 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_64
timestamp 1635444444
transform 1 0 6992 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1339_
timestamp 1635444444
transform 1 0 5980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_70
timestamp 1635444444
transform 1 0 7544 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_74
timestamp 1635444444
transform 1 0 7912 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_78
timestamp 1635444444
transform 1 0 8280 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_85
timestamp 1635444444
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1635444444
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1395_
timestamp 1635444444
transform 1 0 8004 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_wb_clk_i
timestamp 1635444444
transform 1 0 7176 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_102
timestamp 1635444444
transform 1 0 10488 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_109
timestamp 1635444444
transform 1 0 11132 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_94
timestamp 1635444444
transform 1 0 9752 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1209_
timestamp 1635444444
transform -1 0 11132 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1422_
timestamp 1635444444
transform 1 0 9476 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_121
timestamp 1635444444
transform 1 0 12236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1193_
timestamp 1635444444
transform 1 0 12604 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1203_
timestamp 1635444444
transform -1 0 12236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_135
timestamp 1635444444
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1635444444
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1635444444
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1635444444
transform 1 0 14076 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_50_157
timestamp 1635444444
transform 1 0 15548 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_166
timestamp 1635444444
transform 1 0 16376 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1564_
timestamp 1635444444
transform -1 0 16376 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1801_
timestamp 1635444444
transform -1 0 17572 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_179
timestamp 1635444444
transform 1 0 17572 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_187
timestamp 1635444444
transform 1 0 18308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1635444444
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1635444444
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0901_
timestamp 1635444444
transform 1 0 17940 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_197
timestamp 1635444444
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_210
timestamp 1635444444
transform 1 0 20424 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_2  _1030_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 19780 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _1373_
timestamp 1635444444
transform -1 0 21436 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_50_221
timestamp 1635444444
transform 1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1635444444
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_1  _1367_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 21804 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1635444444
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1635444444
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1635444444
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1635444444
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1635444444
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1635444444
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1635444444
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1635444444
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1635444444
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_309
timestamp 1635444444
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_317
timestamp 1635444444
transform 1 0 30268 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1635444444
transform -1 0 30820 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1635444444
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_16
timestamp 1635444444
transform 1 0 2576 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_3
timestamp 1635444444
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1635444444
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1446_
timestamp 1635444444
transform 1 0 1932 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_51_22
timestamp 1635444444
transform 1 0 3128 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_39
timestamp 1635444444
transform 1 0 4692 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1635444444
transform 1 0 3220 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_51_47
timestamp 1635444444
transform 1 0 5428 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1635444444
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1635444444
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1436_
timestamp 1635444444
transform -1 0 5888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1635444444
transform 1 0 6348 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_73
timestamp 1635444444
transform 1 0 7820 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_83
timestamp 1635444444
transform 1 0 8740 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1404_
timestamp 1635444444
transform -1 0 8740 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 1635444444
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_91
timestamp 1635444444
transform 1 0 9476 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1635444444
transform 1 0 9568 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_51_113
timestamp 1635444444
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_118
timestamp 1635444444
transform 1 0 11960 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1635444444
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1181_
timestamp 1635444444
transform -1 0 11960 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1185_
timestamp 1635444444
transform 1 0 12328 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_51_132
timestamp 1635444444
transform 1 0 13248 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_140
timestamp 1635444444
transform 1 0 13984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1635444444
transform 1 0 14168 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_51_158
timestamp 1635444444
transform 1 0 15640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1635444444
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1635444444
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1800_
timestamp 1635444444
transform 1 0 16652 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_178
timestamp 1635444444
transform 1 0 17480 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_191
timestamp 1635444444
transform 1 0 18676 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0923_
timestamp 1635444444
transform 1 0 19044 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1805_
timestamp 1635444444
transform 1 0 17848 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_51_199
timestamp 1635444444
transform 1 0 19412 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_215
timestamp 1635444444
transform 1 0 20884 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0972_
timestamp 1635444444
transform 1 0 19964 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1635444444
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_230
timestamp 1635444444
transform 1 0 22264 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1635444444
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1635444444
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0890_
timestamp 1635444444
transform -1 0 22264 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1635444444
transform 1 0 22632 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1635444444
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1635444444
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1635444444
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1635444444
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1635444444
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1635444444
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1635444444
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1635444444
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_317
timestamp 1635444444
transform 1 0 30268 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1635444444
transform -1 0 30820 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1453_
timestamp 1635444444
transform 1 0 1380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1449_
timestamp 1635444444
transform -1 0 1656 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1635444444
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1635444444
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_6
timestamp 1635444444
transform 1 0 1656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_6
timestamp 1635444444
transform 1 0 1656 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1452_
timestamp 1635444444
transform 1 0 2024 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1448_
timestamp 1635444444
transform 1 0 2024 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1454_
timestamp 1635444444
transform 1 0 3036 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1451_
timestamp 1635444444
transform 1 0 3036 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_17
timestamp 1635444444
transform 1 0 2668 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_17
timestamp 1635444444
transform 1 0 2668 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1635444444
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_33
timestamp 1635444444
transform 1 0 4140 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_24
timestamp 1635444444
transform 1 0 3312 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_37
timestamp 1635444444
transform 1 0 4508 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1635444444
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1316_
timestamp 1635444444
transform -1 0 5796 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1331_
timestamp 1635444444
transform -1 0 4508 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1334_
timestamp 1635444444
transform -1 0 5520 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1635444444
transform 1 0 3772 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_48
timestamp 1635444444
transform 1 0 5520 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_61
timestamp 1635444444
transform 1 0 6716 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1635444444
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1635444444
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1635444444
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1337_
timestamp 1635444444
transform -1 0 6716 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1340_
timestamp 1635444444
transform -1 0 7912 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1635444444
transform -1 0 7820 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_52_74
timestamp 1635444444
transform 1 0 7912 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1635444444
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_73
timestamp 1635444444
transform 1 0 7820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_77
timestamp 1635444444
transform 1 0 8188 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_84
timestamp 1635444444
transform 1 0 8832 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1635444444
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _1394_
timestamp 1635444444
transform -1 0 9476 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1428_
timestamp 1635444444
transform 1 0 8280 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1412_
timestamp 1635444444
transform 1 0 9476 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_90
timestamp 1635444444
transform 1 0 9384 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_91
timestamp 1635444444
transform 1 0 9476 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1393_
timestamp 1635444444
transform 1 0 9844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_97
timestamp 1635444444
transform 1 0 10028 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_98
timestamp 1635444444
transform 1 0 10120 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_wb_clk_i
timestamp 1635444444
transform -1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1413_
timestamp 1635444444
transform 1 0 10488 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_103
timestamp 1635444444
transform 1 0 10580 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_105
timestamp 1635444444
transform 1 0 10764 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1635444444
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_109
timestamp 1635444444
transform 1 0 11132 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_119
timestamp 1635444444
transform 1 0 12052 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_122
timestamp 1635444444
transform 1 0 12328 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_128
timestamp 1635444444
transform 1 0 12880 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1635444444
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1182_
timestamp 1635444444
transform -1 0 13340 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1186_
timestamp 1635444444
transform 1 0 12972 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1206_
timestamp 1635444444
transform 1 0 11224 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1213_
timestamp 1635444444
transform 1 0 11500 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1635444444
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1635444444
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_149
timestamp 1635444444
transform 1 0 14812 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_137
timestamp 1635444444
transform 1 0 13708 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_149
timestamp 1635444444
transform 1 0 14812 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1635444444
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1207_
timestamp 1635444444
transform -1 0 14812 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1215_
timestamp 1635444444
transform 1 0 14076 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_wb_clk_i
timestamp 1635444444
transform 1 0 15916 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1635444444
transform 1 0 15180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1741_
timestamp 1635444444
transform 1 0 15364 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_52_157
timestamp 1635444444
transform 1 0 15548 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1579_
timestamp 1635444444
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1578_
timestamp 1635444444
transform 1 0 16928 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1635444444
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_172
timestamp 1635444444
transform 1 0 16928 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1635444444
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_171
timestamp 1635444444
transform 1 0 16836 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_165
timestamp 1635444444
transform 1 0 16284 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_179
timestamp 1635444444
transform 1 0 17572 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_187
timestamp 1635444444
transform 1 0 18308 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1635444444
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_187
timestamp 1635444444
transform 1 0 18308 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1635444444
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1343_
timestamp 1635444444
transform -1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1355_
timestamp 1635444444
transform 1 0 18676 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1740_
timestamp 1635444444
transform -1 0 18308 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_52_197
timestamp 1635444444
transform 1 0 19228 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_208
timestamp 1635444444
transform 1 0 20240 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_200
timestamp 1635444444
transform 1 0 19504 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_207
timestamp 1635444444
transform 1 0 20148 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1635444444
transform 1 0 19872 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_4  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 22080 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__and3_1  _1312_
timestamp 1635444444
transform 1 0 19780 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _1313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 21344 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_52_228
timestamp 1635444444
transform 1 0 22080 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_236
timestamp 1635444444
transform 1 0 22816 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1635444444
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_235
timestamp 1635444444
transform 1 0 22724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1635444444
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0922_
timestamp 1635444444
transform -1 0 22816 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0948_
timestamp 1635444444
transform 1 0 21804 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1635444444
transform 1 0 23184 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_243
timestamp 1635444444
transform 1 0 23460 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1635444444
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1635444444
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_247
timestamp 1635444444
transform 1 0 23828 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_259
timestamp 1635444444
transform 1 0 24932 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1635444444
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1635444444
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1635444444
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1635444444
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1635444444
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1635444444
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1635444444
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1635444444
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1635444444
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1635444444
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_305
timestamp 1635444444
transform 1 0 29164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1635444444
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_309
timestamp 1635444444
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_317
timestamp 1635444444
transform 1 0 30268 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_316
timestamp 1635444444
transform 1 0 30176 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1635444444
transform -1 0 30820 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1635444444
transform -1 0 30820 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1635444444
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1635444444
transform -1 0 30176 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_54_15
timestamp 1635444444
transform 1 0 2484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 1635444444
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_7
timestamp 1635444444
transform 1 0 1748 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1635444444
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1326_
timestamp 1635444444
transform 1 0 2576 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1635444444
transform -1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1635444444
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_38
timestamp 1635444444
transform 1 0 4600 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1635444444
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1314_
timestamp 1635444444
transform -1 0 5888 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1327_
timestamp 1635444444
transform -1 0 4600 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_54_52
timestamp 1635444444
transform 1 0 5888 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_59
timestamp 1635444444
transform 1 0 6532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1315_
timestamp 1635444444
transform -1 0 6532 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1335_
timestamp 1635444444
transform 1 0 6900 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_66
timestamp 1635444444
transform 1 0 7176 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_73
timestamp 1635444444
transform 1 0 7820 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1635444444
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1635444444
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1635444444
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1336_
timestamp 1635444444
transform 1 0 7544 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1342_
timestamp 1635444444
transform 1 0 8188 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_100
timestamp 1635444444
transform 1 0 10304 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_105
timestamp 1635444444
transform 1 0 10764 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_89
timestamp 1635444444
transform 1 0 9292 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_96
timestamp 1635444444
transform 1 0 9936 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1062_
timestamp 1635444444
transform -1 0 11684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1217_
timestamp 1635444444
transform 1 0 10396 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1421_
timestamp 1635444444
transform -1 0 9936 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_115
timestamp 1635444444
transform 1 0 11684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_127
timestamp 1635444444
transform 1 0 12788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1635444444
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1635444444
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1635444444
transform 1 0 14076 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_157
timestamp 1635444444
transform 1 0 15548 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_164
timestamp 1635444444
transform 1 0 16192 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_172
timestamp 1635444444
transform 1 0 16928 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1635444444
transform 1 0 15916 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_180
timestamp 1635444444
transform 1 0 17664 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_188
timestamp 1635444444
transform 1 0 18400 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1635444444
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1635444444
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1635444444
transform -1 0 17664 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1344_
timestamp 1635444444
transform 1 0 18492 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_206
timestamp 1635444444
transform 1 0 20056 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_214
timestamp 1635444444
transform 1 0 20792 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0920_
timestamp 1635444444
transform -1 0 22080 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0921_
timestamp 1635444444
transform 1 0 20424 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1345_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 19228 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_54_228
timestamp 1635444444
transform 1 0 22080 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_240
timestamp 1635444444
transform 1 0 23184 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1635444444
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1635444444
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1635444444
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1635444444
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1635444444
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1635444444
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1635444444
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_309
timestamp 1635444444
transform 1 0 29532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_317
timestamp 1635444444
transform 1 0 30268 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1635444444
transform -1 0 30820 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1635444444
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_15
timestamp 1635444444
transform 1 0 2484 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1635444444
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_7
timestamp 1635444444
transform 1 0 1748 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1635444444
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1455_
timestamp 1635444444
transform 1 0 1840 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1635444444
transform 1 0 2852 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_35
timestamp 1635444444
transform 1 0 4324 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_39
timestamp 1635444444
transform 1 0 4692 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1320_
timestamp 1635444444
transform -1 0 5704 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_55_50
timestamp 1635444444
transform 1 0 5704 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1635444444
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_64
timestamp 1635444444
transform 1 0 6992 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1635444444
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0961_
timestamp 1635444444
transform 1 0 6716 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_84
timestamp 1635444444
transform 1 0 8832 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1965_
timestamp 1635444444
transform 1 0 7360 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1635444444
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1967_
timestamp 1635444444
transform -1 0 11040 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_55_113
timestamp 1635444444
transform 1 0 11500 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_131
timestamp 1635444444
transform 1 0 13156 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1635444444
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1874_
timestamp 1635444444
transform 1 0 11592 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_55_143
timestamp 1635444444
transform 1 0 14260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_151
timestamp 1635444444
transform 1 0 14996 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _0917_
timestamp 1635444444
transform 1 0 15088 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_160
timestamp 1635444444
transform 1 0 15824 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_169
timestamp 1635444444
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1635444444
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_184
timestamp 1635444444
transform 1 0 18032 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0924_
timestamp 1635444444
transform 1 0 17204 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1742_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 19228 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_55_197
timestamp 1635444444
transform 1 0 19228 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_204
timestamp 1635444444
transform 1 0 19872 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_208
timestamp 1635444444
transform 1 0 20240 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_214
timestamp 1635444444
transform 1 0 20792 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0973_
timestamp 1635444444
transform 1 0 20332 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1354_
timestamp 1635444444
transform 1 0 19596 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1635444444
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1635444444
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1635444444
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1635444444
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1635444444
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1635444444
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1635444444
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1635444444
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1635444444
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1635444444
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1635444444
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1635444444
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_317
timestamp 1635444444
transform 1 0 30268 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1635444444
transform -1 0 30820 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_14
timestamp 1635444444
transform 1 0 2392 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_7
timestamp 1635444444
transform 1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1635444444
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1325_
timestamp 1635444444
transform -1 0 3220 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1635444444
transform 1 0 2116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1635444444
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_23
timestamp 1635444444
transform 1 0 3220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1635444444
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_29
timestamp 1635444444
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_35
timestamp 1635444444
transform 1 0 4324 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_42
timestamp 1635444444
transform 1 0 4968 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1635444444
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1311_
timestamp 1635444444
transform -1 0 4968 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1341_
timestamp 1635444444
transform 1 0 4048 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_46
timestamp 1635444444
transform 1 0 5336 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_51
timestamp 1635444444
transform 1 0 5796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_60
timestamp 1635444444
transform 1 0 6624 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0957_
timestamp 1635444444
transform 1 0 6348 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1240_
timestamp 1635444444
transform 1 0 5428 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1964_
timestamp 1635444444
transform 1 0 6992 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1635444444
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_85
timestamp 1635444444
transform 1 0 8924 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1635444444
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0946_
timestamp 1635444444
transform 1 0 9016 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_103
timestamp 1635444444
transform 1 0 10580 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_89
timestamp 1635444444
transform 1 0 9292 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_93
timestamp 1635444444
transform 1 0 9660 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0947_
timestamp 1635444444
transform -1 0 11224 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0955_
timestamp 1635444444
transform 1 0 9752 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_56_110
timestamp 1635444444
transform 1 0 11224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_130
timestamp 1635444444
transform 1 0 13064 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1635444444
transform 1 0 11592 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1635444444
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_141
timestamp 1635444444
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_149
timestamp 1635444444
transform 1 0 14812 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1635444444
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1972_
timestamp 1635444444
transform 1 0 15088 0 1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_56_169
timestamp 1635444444
transform 1 0 16652 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1971_
timestamp 1635444444
transform 1 0 17020 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1635444444
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1635444444
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1635444444
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_197
timestamp 1635444444
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_201
timestamp 1635444444
transform 1 0 19596 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_205
timestamp 1635444444
transform 1 0 19964 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_214
timestamp 1635444444
transform 1 0 20792 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1635444444
transform 1 0 19688 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0928_
timestamp 1635444444
transform 1 0 20332 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_56_226
timestamp 1635444444
transform 1 0 21896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1635444444
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _0966_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 22540 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1635444444
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1635444444
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1635444444
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1635444444
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1635444444
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1635444444
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1635444444
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1635444444
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1635444444
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_309
timestamp 1635444444
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_317
timestamp 1635444444
transform 1 0 30268 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1635444444
transform -1 0 30820 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1635444444
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_13
timestamp 1635444444
transform 1 0 2300 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_17
timestamp 1635444444
transform 1 0 2668 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_7
timestamp 1635444444
transform 1 0 1748 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1635444444
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1322_
timestamp 1635444444
transform -1 0 3312 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1323_
timestamp 1635444444
transform 1 0 2392 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1635444444
transform -1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_24
timestamp 1635444444
transform 1 0 3312 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_28
timestamp 1635444444
transform 1 0 3680 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_38
timestamp 1635444444
transform 1 0 4600 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1324_
timestamp 1635444444
transform -1 0 4600 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_57_46
timestamp 1635444444
transform 1 0 5336 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1635444444
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1635444444
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_57
timestamp 1635444444
transform 1 0 6348 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_61
timestamp 1635444444
transform 1 0 6716 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1635444444
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0956_
timestamp 1635444444
transform -1 0 7360 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0960_
timestamp 1635444444
transform 1 0 6440 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1248_
timestamp 1635444444
transform -1 0 5796 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_68
timestamp 1635444444
transform 1 0 7360 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_83
timestamp 1635444444
transform 1 0 8740 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0959_
timestamp 1635444444
transform -1 0 8740 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_101
timestamp 1635444444
transform 1 0 10396 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1635444444
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_91
timestamp 1635444444
transform 1 0 9476 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0951_
timestamp 1635444444
transform -1 0 10396 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0953_
timestamp 1635444444
transform 1 0 10764 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_120
timestamp 1635444444
transform 1 0 12144 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_128
timestamp 1635444444
transform 1 0 12880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1635444444
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__o221ai_1  _1211_
timestamp 1635444444
transform -1 0 12144 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1635444444
transform -1 0 14628 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_57_147
timestamp 1635444444
transform 1 0 14628 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_155
timestamp 1635444444
transform 1 0 15364 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_159
timestamp 1635444444
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1635444444
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_172
timestamp 1635444444
transform 1 0 16928 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1635444444
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0918_
timestamp 1635444444
transform 1 0 15456 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0919_
timestamp 1635444444
transform 1 0 16652 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_184
timestamp 1635444444
transform 1 0 18032 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_189
timestamp 1635444444
transform 1 0 18492 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1346_
timestamp 1635444444
transform 1 0 18860 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1351_
timestamp 1635444444
transform -1 0 18492 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_201
timestamp 1635444444
transform 1 0 19596 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_209
timestamp 1635444444
transform 1 0 20332 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1737_
timestamp 1635444444
transform -1 0 21344 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1635444444
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_225
timestamp 1635444444
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_234
timestamp 1635444444
transform 1 0 22632 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1635444444
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1362_
timestamp 1635444444
transform 1 0 22356 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_246
timestamp 1635444444
transform 1 0 23736 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_258
timestamp 1635444444
transform 1 0 24840 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_270
timestamp 1635444444
transform 1 0 25944 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1635444444
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1635444444
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1635444444
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1635444444
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_305
timestamp 1635444444
transform 1 0 29164 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_316
timestamp 1635444444
transform 1 0 30176 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1635444444
transform -1 0 30820 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1635444444
transform 1 0 29900 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_15
timestamp 1635444444
transform 1 0 2484 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1635444444
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_7
timestamp 1635444444
transform 1 0 1748 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1635444444
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1458_
timestamp 1635444444
transform 1 0 1840 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1635444444
transform -1 0 3220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_23
timestamp 1635444444
transform 1 0 3220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1635444444
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1635444444
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1635444444
transform 1 0 3772 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_45
timestamp 1635444444
transform 1 0 5244 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_58
timestamp 1635444444
transform 1 0 6440 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0964_
timestamp 1635444444
transform 1 0 6992 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1317_
timestamp 1635444444
transform -1 0 6440 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_58_67
timestamp 1635444444
transform 1 0 7268 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_80
timestamp 1635444444
transform 1 0 8464 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1635444444
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1635444444
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0963_
timestamp 1635444444
transform -1 0 8464 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_58_92
timestamp 1635444444
transform 1 0 9568 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0952_
timestamp 1635444444
transform 1 0 9292 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1966_
timestamp 1635444444
transform -1 0 11408 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_112
timestamp 1635444444
transform 1 0 11408 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_126
timestamp 1635444444
transform 1 0 12696 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0950_
timestamp 1635444444
transform 1 0 11776 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1635444444
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1635444444
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1888_
timestamp 1635444444
transform 1 0 14076 0 1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_58_158
timestamp 1635444444
transform 1 0 15640 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_170
timestamp 1635444444
transform 1 0 16744 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_185
timestamp 1635444444
transform 1 0 18124 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1635444444
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1635444444
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1635444444
transform -1 0 18768 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1347_
timestamp 1635444444
transform -1 0 18124 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_197
timestamp 1635444444
transform 1 0 19228 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_209
timestamp 1635444444
transform 1 0 20332 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_2  _0930_
timestamp 1635444444
transform 1 0 20700 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1734_
timestamp 1635444444
transform 1 0 19504 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_58_220
timestamp 1635444444
transform 1 0 21344 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_227
timestamp 1635444444
transform 1 0 21988 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_234
timestamp 1635444444
transform 1 0 22632 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1635444444
transform 1 0 21712 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1361_
timestamp 1635444444
transform 1 0 22356 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_246
timestamp 1635444444
transform 1 0 23736 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1635444444
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1635444444
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1635444444
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1635444444
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1635444444
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1635444444
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1635444444
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_309
timestamp 1635444444
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_317
timestamp 1635444444
transform 1 0 30268 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1635444444
transform -1 0 30820 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1635444444
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _1462_
timestamp 1635444444
transform 1 0 1840 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1460_
timestamp 1635444444
transform 1 0 1840 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1635444444
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1635444444
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_7
timestamp 1635444444
transform 1 0 1748 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_3
timestamp 1635444444
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_7
timestamp 1635444444
transform 1 0 1748 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1635444444
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_15
timestamp 1635444444
transform 1 0 2484 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_15
timestamp 1635444444
transform 1 0 2484 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1635444444
transform 1 0 2852 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_32
timestamp 1635444444
transform 1 0 4048 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_23
timestamp 1635444444
transform 1 0 3220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1635444444
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1635444444
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1321_
timestamp 1635444444
transform 1 0 3220 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1635444444
transform 1 0 3772 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1635444444
transform -1 0 5888 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _0944_
timestamp 1635444444
transform -1 0 6072 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_45
timestamp 1635444444
transform 1 0 5244 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_52
timestamp 1635444444
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1328_
timestamp 1635444444
transform -1 0 6624 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906__1
timestamp 1635444444
transform -1 0 6716 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1635444444
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_61
timestamp 1635444444
transform 1 0 6716 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_54
timestamp 1635444444
transform 1 0 6072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_60
timestamp 1635444444
transform 1 0 6624 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0907_
timestamp 1635444444
transform -1 0 7268 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0967_
timestamp 1635444444
transform 1 0 7636 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0945_
timestamp 1635444444
transform -1 0 7912 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_69
timestamp 1635444444
transform 1 0 7452 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_74
timestamp 1635444444
transform 1 0 7912 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_67
timestamp 1635444444
transform 1 0 7268 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1635444444
transform 1 0 8648 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1635444444
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_85
timestamp 1635444444
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1635444444
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_85
timestamp 1635444444
transform 1 0 8924 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1635444444
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_93
timestamp 1635444444
transform 1 0 9660 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_106
timestamp 1635444444
transform 1 0 10856 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_99
timestamp 1635444444
transform 1 0 10212 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0932_
timestamp 1635444444
transform 1 0 9292 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0933_
timestamp 1635444444
transform 1 0 9844 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0940_
timestamp 1635444444
transform -1 0 10856 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1635444444
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_116
timestamp 1635444444
transform 1 0 11776 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_114
timestamp 1635444444
transform 1 0 11592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1635444444
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1875_
timestamp 1635444444
transform 1 0 11684 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1887_
timestamp 1635444444
transform 1 0 12328 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  net99_2
timestamp 1635444444
transform 1 0 11500 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_139
timestamp 1635444444
transform 1 0 13892 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_132
timestamp 1635444444
transform 1 0 13248 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_60_141
timestamp 1635444444
transform 1 0 14076 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_147
timestamp 1635444444
transform 1 0 14628 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1635444444
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14720 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1823_
timestamp 1635444444
transform 1 0 14260 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1635444444
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1635444444
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_174
timestamp 1635444444
transform 1 0 17112 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_169
timestamp 1635444444
transform 1 0 16652 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1635444444
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1577_
timestamp 1635444444
transform -1 0 17112 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1804_
timestamp 1635444444
transform -1 0 17848 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_59_194
timestamp 1635444444
transform 1 0 18952 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_182
timestamp 1635444444
transform 1 0 17848 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_191
timestamp 1635444444
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1635444444
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1635444444
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1576_
timestamp 1635444444
transform 1 0 18216 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1635444444
transform 1 0 17480 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_59_206
timestamp 1635444444
transform 1 0 20056 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1635444444
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_197
timestamp 1635444444
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_205
timestamp 1635444444
transform 1 0 19964 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_212
timestamp 1635444444
transform 1 0 20608 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1222_
timestamp 1635444444
transform -1 0 21252 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1223_
timestamp 1635444444
transform 1 0 20424 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1350_
timestamp 1635444444
transform 1 0 19320 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1523_
timestamp 1635444444
transform 1 0 20056 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1635444444
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1635444444
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1635444444
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_219
timestamp 1635444444
transform 1 0 21252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_231
timestamp 1635444444
transform 1 0 22356 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1635444444
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0962_
timestamp 1635444444
transform -1 0 22356 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1635444444
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1635444444
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_243
timestamp 1635444444
transform 1 0 23460 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1635444444
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1635444444
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1635444444
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1635444444
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1635444444
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1635444444
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1635444444
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1635444444
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1635444444
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1635444444
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1635444444
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1635444444
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1635444444
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_59_317
timestamp 1635444444
transform 1 0 30268 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1635444444
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_309
timestamp 1635444444
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_316
timestamp 1635444444
transform 1 0 30176 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1635444444
transform -1 0 30820 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1635444444
transform -1 0 30820 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1635444444
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1635444444
transform 1 0 29900 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_15
timestamp 1635444444
transform 1 0 2484 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1635444444
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_7
timestamp 1635444444
transform 1 0 1748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1635444444
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1318_
timestamp 1635444444
transform 1 0 2852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1464_
timestamp 1635444444
transform 1 0 1840 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_61_22
timestamp 1635444444
transform 1 0 3128 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_29
timestamp 1635444444
transform 1 0 3772 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_37
timestamp 1635444444
transform 1 0 4508 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_42
timestamp 1635444444
transform 1 0 4968 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1310_
timestamp 1635444444
transform -1 0 4968 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1319_
timestamp 1635444444
transform 1 0 3496 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1635444444
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1635444444
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_63
timestamp 1635444444
transform 1 0 6900 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1635444444
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1249_
timestamp 1635444444
transform -1 0 5796 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1382_
timestamp 1635444444
transform 1 0 6348 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_71
timestamp 1635444444
transform 1 0 7636 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1635444444
transform 1 0 7820 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1635444444
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_89
timestamp 1635444444
transform 1 0 9292 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_95
timestamp 1635444444
transform 1 0 9844 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0943_
timestamp 1635444444
transform 1 0 9936 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1635444444
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1635444444
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_121
timestamp 1635444444
transform 1 0 12236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1635444444
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _0904_
timestamp 1635444444
transform 1 0 11684 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1183_
timestamp 1635444444
transform 1 0 12604 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_133
timestamp 1635444444
transform 1 0 13340 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_145
timestamp 1635444444
transform 1 0 14444 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_157
timestamp 1635444444
transform 1 0 15548 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 1635444444
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1635444444
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1810_
timestamp 1635444444
transform -1 0 17480 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_61_178
timestamp 1635444444
transform 1 0 17480 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_184
timestamp 1635444444
transform 1 0 18032 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1635444444
transform 1 0 18124 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_61_201
timestamp 1635444444
transform 1 0 19596 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_207
timestamp 1635444444
transform 1 0 20148 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_211
timestamp 1635444444
transform 1 0 20516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1221_
timestamp 1635444444
transform -1 0 20516 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1635444444
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1635444444
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1635444444
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1635444444
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1635444444
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1635444444
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1635444444
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1635444444
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1635444444
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1635444444
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1635444444
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1635444444
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_317
timestamp 1635444444
transform 1 0 30268 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1635444444
transform -1 0 30820 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_15
timestamp 1635444444
transform 1 0 2484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_7
timestamp 1635444444
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1635444444
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1456_
timestamp 1635444444
transform 1 0 2852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1635444444
transform -1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1635444444
transform -1 0 2484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_22
timestamp 1635444444
transform 1 0 3128 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_32
timestamp 1635444444
transform 1 0 4048 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_39
timestamp 1635444444
transform 1 0 4692 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1635444444
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0992_
timestamp 1635444444
transform 1 0 3772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1250_
timestamp 1635444444
transform 1 0 5060 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1459_
timestamp 1635444444
transform 1 0 4416 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_46
timestamp 1635444444
transform 1 0 5336 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_60
timestamp 1635444444
transform 1 0 6624 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1434_
timestamp 1635444444
transform 1 0 5704 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _1435_
timestamp 1635444444
transform -1 0 7544 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_70
timestamp 1635444444
transform 1 0 7544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1635444444
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1635444444
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1635444444
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0965_
timestamp 1635444444
transform -1 0 8188 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1465_
timestamp 1635444444
transform 1 0 8924 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_88
timestamp 1635444444
transform 1 0 9200 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_95
timestamp 1635444444
transform 1 0 9844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0941_
timestamp 1635444444
transform 1 0 9568 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1968_
timestamp 1635444444
transform 1 0 10212 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_115
timestamp 1635444444
transform 1 0 11684 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_123
timestamp 1635444444
transform 1 0 12420 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__a221o_1  _1184_
timestamp 1635444444
transform -1 0 13340 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1635444444
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1635444444
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_141
timestamp 1635444444
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_149
timestamp 1635444444
transform 1 0 14812 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1635444444
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1817_
timestamp 1635444444
transform 1 0 15088 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_62_173
timestamp 1635444444
transform 1 0 17020 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_182
timestamp 1635444444
transform 1 0 17848 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1635444444
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1635444444
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1635444444
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1348_
timestamp 1635444444
transform 1 0 17572 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1349_
timestamp 1635444444
transform -1 0 18492 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_197
timestamp 1635444444
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_210
timestamp 1635444444
transform 1 0 20424 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1522_
timestamp 1635444444
transform -1 0 21344 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1758_
timestamp 1635444444
transform 1 0 19596 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_220
timestamp 1635444444
transform 1 0 21344 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_232
timestamp 1635444444
transform 1 0 22448 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_244
timestamp 1635444444
transform 1 0 23552 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1635444444
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1635444444
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1635444444
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1635444444
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1635444444
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1635444444
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1635444444
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_309
timestamp 1635444444
transform 1 0 29532 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_317
timestamp 1635444444
transform 1 0 30268 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1635444444
transform -1 0 30820 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1635444444
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_17
timestamp 1635444444
transform 1 0 2668 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_6
timestamp 1635444444
transform 1 0 1656 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1635444444
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1635444444
transform -1 0 1656 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1472_
timestamp 1635444444
transform 1 0 2024 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_63_28
timestamp 1635444444
transform 1 0 3680 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_41
timestamp 1635444444
transform 1 0 4876 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0990_
timestamp 1635444444
transform 1 0 3404 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0994_
timestamp 1635444444
transform -1 0 4876 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_63_50
timestamp 1635444444
transform 1 0 5704 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_57
timestamp 1635444444
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1635444444
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0968_
timestamp 1635444444
transform -1 0 5704 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1440_
timestamp 1635444444
transform -1 0 7452 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_69
timestamp 1635444444
transform 1 0 7452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_76
timestamp 1635444444
transform 1 0 8096 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_84
timestamp 1635444444
transform 1 0 8832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0908_
timestamp 1635444444
transform 1 0 9016 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1383_
timestamp 1635444444
transform 1 0 7820 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_107
timestamp 1635444444
transform 1 0 10948 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_89
timestamp 1635444444
transform 1 0 9292 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_97
timestamp 1635444444
transform 1 0 10028 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0935_
timestamp 1635444444
transform 1 0 10120 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1635444444
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_116
timestamp 1635444444
transform 1 0 11776 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_122
timestamp 1635444444
transform 1 0 12328 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_127
timestamp 1635444444
transform 1 0 12788 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1635444444
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0936_
timestamp 1635444444
transform -1 0 11776 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0998_
timestamp 1635444444
transform 1 0 12420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1210_
timestamp 1635444444
transform 1 0 13156 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_134
timestamp 1635444444
transform 1 0 13432 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_145
timestamp 1635444444
transform 1 0 14444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_152
timestamp 1635444444
transform 1 0 15088 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1571_
timestamp 1635444444
transform -1 0 15088 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1594_
timestamp 1635444444
transform -1 0 14444 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1635444444
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1635444444
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1635444444
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1761_
timestamp 1635444444
transform -1 0 17664 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_63_180
timestamp 1635444444
transform 1 0 17664 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_188
timestamp 1635444444
transform 1 0 18400 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_193
timestamp 1635444444
transform 1 0 18860 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1352_
timestamp 1635444444
transform 1 0 18584 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1635444444
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1828_
timestamp 1635444444
transform 1 0 19228 0 -1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1635444444
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_231
timestamp 1635444444
transform 1 0 22356 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1635444444
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0958_
timestamp 1635444444
transform -1 0 22356 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_243
timestamp 1635444444
transform 1 0 23460 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_255
timestamp 1635444444
transform 1 0 24564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_267
timestamp 1635444444
transform 1 0 25668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1635444444
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1635444444
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1635444444
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1635444444
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1635444444
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_317
timestamp 1635444444
transform 1 0 30268 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1635444444
transform -1 0 30820 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_16
timestamp 1635444444
transform 1 0 2576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_3
timestamp 1635444444
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1635444444
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1467_
timestamp 1635444444
transform 1 0 1932 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1635444444
transform 1 0 2944 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1635444444
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_32
timestamp 1635444444
transform 1 0 4048 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1635444444
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0981_
timestamp 1635444444
transform -1 0 5704 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0989_
timestamp 1635444444
transform -1 0 4048 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_50
timestamp 1635444444
transform 1 0 5704 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1635444444
transform 1 0 6072 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_64_70
timestamp 1635444444
transform 1 0 7544 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_76
timestamp 1635444444
transform 1 0 8096 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 1635444444
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1635444444
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1003_
timestamp 1635444444
transform -1 0 8464 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1005_
timestamp 1635444444
transform -1 0 9752 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_64_102
timestamp 1635444444
transform 1 0 10488 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_94
timestamp 1635444444
transform 1 0 9752 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1635444444
transform 1 0 10580 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_64_119
timestamp 1635444444
transform 1 0 12052 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_125
timestamp 1635444444
transform 1 0 12604 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_131
timestamp 1635444444
transform 1 0 13156 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1610_
timestamp 1635444444
transform -1 0 13156 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1635444444
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_148
timestamp 1635444444
transform 1 0 14720 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1635444444
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_2  _1572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14076 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1816_
timestamp 1635444444
transform 1 0 15088 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_64_173
timestamp 1635444444
transform 1 0 17020 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_190
timestamp 1635444444
transform 1 0 18584 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1635444444
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1759_
timestamp 1635444444
transform -1 0 18584 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_200
timestamp 1635444444
transform 1 0 19504 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_212
timestamp 1635444444
transform 1 0 20608 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1353_
timestamp 1635444444
transform -1 0 19504 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_224
timestamp 1635444444
transform 1 0 21712 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_236
timestamp 1635444444
transform 1 0 22816 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1635444444
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1635444444
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1635444444
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1635444444
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1635444444
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1635444444
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1635444444
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1635444444
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_309
timestamp 1635444444
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_316
timestamp 1635444444
transform 1 0 30176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1635444444
transform -1 0 30820 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1635444444
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1635444444
transform 1 0 29900 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_7
timestamp 1635444444
transform 1 0 1748 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1635444444
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1635444444
transform -1 0 3772 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1635444444
transform -1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_29
timestamp 1635444444
transform 1 0 3772 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1958_
timestamp 1635444444
transform 1 0 4140 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_65_49
timestamp 1635444444
transform 1 0 5612 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1635444444
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1635444444
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1251_
timestamp 1635444444
transform -1 0 7176 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_65_66
timestamp 1635444444
transform 1 0 7176 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_73
timestamp 1635444444
transform 1 0 7820 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1468_
timestamp 1635444444
transform 1 0 7544 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1635444444
transform 1 0 8188 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_65_106
timestamp 1635444444
transform 1 0 10856 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_93
timestamp 1635444444
transform 1 0 9660 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0939_
timestamp 1635444444
transform 1 0 10028 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_65_129
timestamp 1635444444
transform 1 0 12972 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1635444444
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1970_
timestamp 1635444444
transform 1 0 11500 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_137
timestamp 1635444444
transform 1 0 13708 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_147
timestamp 1635444444
transform 1 0 14628 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1593_
timestamp 1635444444
transform 1 0 14996 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1596_
timestamp 1635444444
transform -1 0 14628 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1612_
timestamp 1635444444
transform -1 0 13708 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_154
timestamp 1635444444
transform 1 0 15272 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1635444444
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_169
timestamp 1635444444
transform 1 0 16652 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1635444444
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_177
timestamp 1635444444
transform 1 0 17388 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_185
timestamp 1635444444
transform 1 0 18124 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_192
timestamp 1635444444
transform 1 0 18768 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1597_
timestamp 1635444444
transform 1 0 17664 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1598_
timestamp 1635444444
transform 1 0 18492 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_204
timestamp 1635444444
transform 1 0 19872 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_216
timestamp 1635444444
transform 1 0 20976 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1635444444
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1635444444
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1635444444
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1635444444
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1635444444
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1635444444
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1635444444
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1635444444
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1635444444
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1635444444
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1635444444
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_317
timestamp 1635444444
transform 1 0 30268 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1635444444
transform -1 0 30820 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1635444444
transform -1 0 1656 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1635444444
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1635444444
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_6
timestamp 1635444444
transform 1 0 1656 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_3
timestamp 1635444444
transform 1 0 1380 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1474_
timestamp 1635444444
transform 1 0 2024 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1470_
timestamp 1635444444
transform 1 0 1932 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1635444444
transform 1 0 2944 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1635444444
transform 1 0 3036 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_17
timestamp 1635444444
transform 1 0 2668 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_16
timestamp 1635444444
transform 1 0 2576 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1635444444
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_38
timestamp 1635444444
transform 1 0 4600 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_24
timestamp 1635444444
transform 1 0 3312 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_30
timestamp 1635444444
transform 1 0 3864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_34
timestamp 1635444444
transform 1 0 4232 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1635444444
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0991_
timestamp 1635444444
transform -1 0 4600 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0993_
timestamp 1635444444
transform 1 0 3956 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1231_
timestamp 1635444444
transform 1 0 4968 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1635444444
transform 1 0 5612 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0976_
timestamp 1635444444
transform 1 0 5428 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_67_52
timestamp 1635444444
transform 1 0 5888 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_45
timestamp 1635444444
transform 1 0 5244 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_46
timestamp 1635444444
transform 1 0 5336 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0978_
timestamp 1635444444
transform 1 0 6716 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1635444444
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_57
timestamp 1635444444
transform 1 0 6348 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_57
timestamp 1635444444
transform 1 0 6348 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1635444444
transform 1 0 6532 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_66_71
timestamp 1635444444
transform 1 0 7636 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_80
timestamp 1635444444
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_75
timestamp 1635444444
transform 1 0 8004 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1635444444
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0995_
timestamp 1635444444
transform 1 0 8188 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0999_
timestamp 1635444444
transform 1 0 8556 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1002_
timestamp 1635444444
transform 1 0 8924 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_66_100
timestamp 1635444444
transform 1 0 10304 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_104
timestamp 1635444444
transform 1 0 10672 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_94
timestamp 1635444444
transform 1 0 9752 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_103
timestamp 1635444444
transform 1 0 10580 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_90
timestamp 1635444444
transform 1 0 9384 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_98
timestamp 1635444444
transform 1 0 10120 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0925_
timestamp 1635444444
transform 1 0 10396 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0926_
timestamp 1635444444
transform 1 0 11040 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0937_
timestamp 1635444444
transform 1 0 10304 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1611_
timestamp 1635444444
transform -1 0 12420 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1635444444
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_113
timestamp 1635444444
transform 1 0 11500 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1635444444
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_119
timestamp 1635444444
transform 1 0 12052 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_111
timestamp 1635444444
transform 1 0 11316 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_2  _1617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 12788 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_67_121
timestamp 1635444444
transform 1 0 12236 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_123
timestamp 1635444444
transform 1 0 12420 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1815_
timestamp 1635444444
transform 1 0 12512 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_66_136
timestamp 1635444444
transform 1 0 13616 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_146
timestamp 1635444444
transform 1 0 14536 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_145
timestamp 1635444444
transform 1 0 14444 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_151
timestamp 1635444444
transform 1 0 14996 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1635444444
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1547_
timestamp 1635444444
transform 1 0 15088 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1595_
timestamp 1635444444
transform 1 0 14904 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1613_
timestamp 1635444444
transform -1 0 14536 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1635444444
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1635444444
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_155
timestamp 1635444444
transform 1 0 15364 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_164
timestamp 1635444444
transform 1 0 16192 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_172
timestamp 1635444444
transform 1 0 16928 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1635444444
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1548_
timestamp 1635444444
transform 1 0 15732 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1552_
timestamp 1635444444
transform -1 0 16928 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_177
timestamp 1635444444
transform 1 0 17388 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_181
timestamp 1635444444
transform 1 0 17756 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_187
timestamp 1635444444
transform 1 0 18308 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1635444444
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_185
timestamp 1635444444
transform 1 0 18124 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1635444444
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1554_
timestamp 1635444444
transform 1 0 17848 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1776_
timestamp 1635444444
transform -1 0 19320 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1779_
timestamp 1635444444
transform 1 0 17296 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_66_202
timestamp 1635444444
transform 1 0 19688 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1635444444
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_198
timestamp 1635444444
transform 1 0 19320 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_211
timestamp 1635444444
transform 1 0 20516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1618_
timestamp 1635444444
transform 1 0 19228 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1635444444
transform 1 0 20056 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1738_
timestamp 1635444444
transform -1 0 20516 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1635444444
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1635444444
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1635444444
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_231
timestamp 1635444444
transform 1 0 22356 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1635444444
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0954_
timestamp 1635444444
transform -1 0 22356 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1635444444
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1635444444
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1635444444
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_243
timestamp 1635444444
transform 1 0 23460 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_255
timestamp 1635444444
transform 1 0 24564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1635444444
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1635444444
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1635444444
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_267
timestamp 1635444444
transform 1 0 25668 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1635444444
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1635444444
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1635444444
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1635444444
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1635444444
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1635444444
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1635444444
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1635444444
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_309
timestamp 1635444444
transform 1 0 29532 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_317
timestamp 1635444444
transform 1 0 30268 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_317
timestamp 1635444444
transform 1 0 30268 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1635444444
transform -1 0 30820 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1635444444
transform -1 0 30820 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1635444444
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_16
timestamp 1635444444
transform 1 0 2576 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_20
timestamp 1635444444
transform 1 0 2944 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_3
timestamp 1635444444
transform 1 0 1380 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1635444444
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0986_
timestamp 1635444444
transform -1 0 3312 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1476_
timestamp 1635444444
transform 1 0 1932 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_68_24
timestamp 1635444444
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_38
timestamp 1635444444
transform 1 0 4600 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1635444444
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0988_
timestamp 1635444444
transform -1 0 4600 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1466_
timestamp 1635444444
transform 1 0 4968 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_45
timestamp 1635444444
transform 1 0 5244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_49
timestamp 1635444444
transform 1 0 5612 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_53
timestamp 1635444444
transform 1 0 5980 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1245_
timestamp 1635444444
transform -1 0 5980 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1247_
timestamp 1635444444
transform 1 0 6348 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_68_66
timestamp 1635444444
transform 1 0 7176 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_73
timestamp 1635444444
transform 1 0 7820 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_80
timestamp 1635444444
transform 1 0 8464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_85
timestamp 1635444444
transform 1 0 8924 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1635444444
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1004_
timestamp 1635444444
transform -1 0 8464 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1635444444
transform -1 0 7820 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1635444444
transform 1 0 9016 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_102
timestamp 1635444444
transform 1 0 10488 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_114
timestamp 1635444444
transform 1 0 11592 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_121
timestamp 1635444444
transform 1 0 12236 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_130
timestamp 1635444444
transform 1 0 13064 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1614_
timestamp 1635444444
transform -1 0 12236 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1615_
timestamp 1635444444
transform 1 0 12604 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_68_138
timestamp 1635444444
transform 1 0 13800 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_141
timestamp 1635444444
transform 1 0 14076 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1635444444
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1819_
timestamp 1635444444
transform 1 0 14444 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_68_166
timestamp 1635444444
transform 1 0 16376 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1778_
timestamp 1635444444
transform -1 0 17572 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_68_179
timestamp 1635444444
transform 1 0 17572 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_186
timestamp 1635444444
transform 1 0 18216 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_194
timestamp 1635444444
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1635444444
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1635444444
transform 1 0 17940 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_197
timestamp 1635444444
transform 1 0 19228 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_206
timestamp 1635444444
transform 1 0 20056 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_218
timestamp 1635444444
transform 1 0 21160 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1633_
timestamp 1635444444
transform 1 0 19596 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_68_230
timestamp 1635444444
transform 1 0 22264 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_242
timestamp 1635444444
transform 1 0 23368 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1635444444
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1635444444
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1635444444
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1635444444
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1635444444
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1635444444
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1635444444
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1635444444
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_309
timestamp 1635444444
transform 1 0 29532 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_316
timestamp 1635444444
transform 1 0 30176 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1635444444
transform -1 0 30820 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1635444444
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1635444444
transform 1 0 29900 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_18
timestamp 1635444444
transform 1 0 2760 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_7
timestamp 1635444444
transform 1 0 1748 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1635444444
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0987_
timestamp 1635444444
transform 1 0 2484 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1635444444
transform -1 0 1748 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_38
timestamp 1635444444
transform 1 0 4600 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0970_
timestamp 1635444444
transform 1 0 4968 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1635444444
transform 1 0 3128 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_45
timestamp 1635444444
transform 1 0 5244 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_52
timestamp 1635444444
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1635444444
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1244_
timestamp 1635444444
transform 1 0 6348 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1246_
timestamp 1635444444
transform 1 0 5612 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_66
timestamp 1635444444
transform 1 0 7176 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_75
timestamp 1635444444
transform 1 0 8004 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_82
timestamp 1635444444
transform 1 0 8648 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0997_
timestamp 1635444444
transform 1 0 8372 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1000_
timestamp 1635444444
transform 1 0 7728 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1635444444
transform -1 0 10488 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_69_102
timestamp 1635444444
transform 1 0 10488 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_110
timestamp 1635444444
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_113
timestamp 1635444444
transform 1 0 11500 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_117
timestamp 1635444444
transform 1 0 11868 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_121
timestamp 1635444444
transform 1 0 12236 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1635444444
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1631_
timestamp 1635444444
transform -1 0 12236 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1814_
timestamp 1635444444
transform 1 0 12604 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_69_146
timestamp 1635444444
transform 1 0 14536 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1736_
timestamp 1635444444
transform -1 0 15732 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_69_159
timestamp 1635444444
transform 1 0 15732 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1635444444
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1635444444
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1818_
timestamp 1635444444
transform 1 0 16652 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_69_190
timestamp 1635444444
transform 1 0 18584 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1619_
timestamp 1635444444
transform 1 0 18952 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_197
timestamp 1635444444
transform 1 0 19228 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_209
timestamp 1635444444
transform 1 0 20332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_221
timestamp 1635444444
transform 1 0 21436 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_232
timestamp 1635444444
transform 1 0 22448 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1635444444
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0949_
timestamp 1635444444
transform -1 0 22448 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_69_244
timestamp 1635444444
transform 1 0 23552 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_256
timestamp 1635444444
transform 1 0 24656 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_268
timestamp 1635444444
transform 1 0 25760 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1635444444
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1635444444
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1635444444
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1635444444
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_317
timestamp 1635444444
transform 1 0 30268 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1635444444
transform -1 0 30820 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_18
timestamp 1635444444
transform 1 0 2760 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_7
timestamp 1635444444
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1635444444
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1482_
timestamp 1635444444
transform 1 0 2116 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1635444444
transform -1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_26
timestamp 1635444444
transform 1 0 3496 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_29
timestamp 1635444444
transform 1 0 3772 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1635444444
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0982_
timestamp 1635444444
transform -1 0 5152 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_70_44
timestamp 1635444444
transform 1 0 5152 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_58
timestamp 1635444444
transform 1 0 6440 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_62
timestamp 1635444444
transform 1 0 6808 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1225_
timestamp 1635444444
transform 1 0 6900 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1381_
timestamp 1635444444
transform -1 0 6440 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_70_73
timestamp 1635444444
transform 1 0 7820 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_81
timestamp 1635444444
transform 1 0 8556 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1635444444
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0996_
timestamp 1635444444
transform -1 0 9200 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_107
timestamp 1635444444
transform 1 0 10948 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_88
timestamp 1635444444
transform 1 0 9200 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_95
timestamp 1635444444
transform 1 0 9844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1001_
timestamp 1635444444
transform 1 0 9568 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_119
timestamp 1635444444
transform 1 0 12052 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_125
timestamp 1635444444
transform 1 0 12604 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1616_
timestamp 1635444444
transform -1 0 13248 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1632_
timestamp 1635444444
transform -1 0 12604 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_132
timestamp 1635444444
transform 1 0 13248 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_141
timestamp 1635444444
transform 1 0 14076 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1635444444
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1820_
timestamp 1635444444
transform 1 0 14444 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_70_166
timestamp 1635444444
transform 1 0 16376 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1551_
timestamp 1635444444
transform 1 0 16744 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_70_175
timestamp 1635444444
transform 1 0 17204 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_183
timestamp 1635444444
transform 1 0 17940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1635444444
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1635444444
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1553_
timestamp 1635444444
transform -1 0 17940 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1635444444
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1635444444
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1635444444
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1635444444
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1635444444
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1635444444
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1635444444
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1635444444
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1635444444
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1635444444
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1635444444
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1635444444
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1635444444
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_309
timestamp 1635444444
transform 1 0 29532 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_317
timestamp 1635444444
transform 1 0 30268 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1635444444
transform -1 0 30820 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1635444444
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_16
timestamp 1635444444
transform 1 0 2576 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_71_3
timestamp 1635444444
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1635444444
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1479_
timestamp 1635444444
transform 1 0 1932 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_71_22
timestamp 1635444444
transform 1 0 3128 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_32
timestamp 1635444444
transform 1 0 4048 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0985_
timestamp 1635444444
transform 1 0 3220 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1962_
timestamp 1635444444
transform -1 0 5888 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_52
timestamp 1635444444
transform 1 0 5888 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_57
timestamp 1635444444
transform 1 0 6348 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1635444444
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1635444444
transform -1 0 8188 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_77
timestamp 1635444444
transform 1 0 8188 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1226_
timestamp 1635444444
transform 1 0 8556 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_71_103
timestamp 1635444444
transform 1 0 10580 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_91
timestamp 1635444444
transform 1 0 9476 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1635444444
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1635444444
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1635444444
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1635444444
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1635444444
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1635444444
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_164
timestamp 1635444444
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_173
timestamp 1635444444
transform 1 0 17020 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1635444444
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1549_
timestamp 1635444444
transform -1 0 16192 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1550_
timestamp 1635444444
transform -1 0 17020 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_185
timestamp 1635444444
transform 1 0 18124 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_197
timestamp 1635444444
transform 1 0 19228 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_209
timestamp 1635444444
transform 1 0 20332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_221
timestamp 1635444444
transform 1 0 21436 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1635444444
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1635444444
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1635444444
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1635444444
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1635444444
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1635444444
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1635444444
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1635444444
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1635444444
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1635444444
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_305
timestamp 1635444444
transform 1 0 29164 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_316
timestamp 1635444444
transform 1 0 30176 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1635444444
transform -1 0 30820 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1635444444
transform 1 0 29900 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1635444444
transform -1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1635444444
transform -1 0 1748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1635444444
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1635444444
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_7
timestamp 1635444444
transform 1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_7
timestamp 1635444444
transform 1 0 1748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1486_
timestamp 1635444444
transform 1 0 2116 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1484_
timestamp 1635444444
transform 1 0 2116 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_73_18
timestamp 1635444444
transform 1 0 2760 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_18
timestamp 1635444444
transform 1 0 2760 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_26
timestamp 1635444444
transform 1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_29
timestamp 1635444444
transform 1 0 3772 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_37
timestamp 1635444444
transform 1 0 4508 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_42
timestamp 1635444444
transform 1 0 4968 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1635444444
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1635444444
transform 1 0 4692 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0983_
timestamp 1635444444
transform 1 0 3496 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1961_
timestamp 1635444444
transform 1 0 3772 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1481_
timestamp 1635444444
transform 1 0 5612 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _1238_
timestamp 1635444444
transform 1 0 5612 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_52
timestamp 1635444444
transform 1 0 5888 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_48
timestamp 1635444444
transform 1 0 5520 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_45
timestamp 1635444444
transform 1 0 5244 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1241_
timestamp 1635444444
transform 1 0 6716 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1635444444
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_57
timestamp 1635444444
transform 1 0 6348 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_63
timestamp 1635444444
transform 1 0 6900 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_59
timestamp 1635444444
transform 1 0 6532 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1635444444
transform -1 0 8464 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_72_80
timestamp 1635444444
transform 1 0 8464 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_70
timestamp 1635444444
transform 1 0 7544 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_77
timestamp 1635444444
transform 1 0 8188 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1635444444
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1239_
timestamp 1635444444
transform 1 0 7912 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1243_
timestamp 1635444444
transform -1 0 9200 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_100
timestamp 1635444444
transform 1 0 10304 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_88
timestamp 1635444444
transform 1 0 9200 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_101
timestamp 1635444444
transform 1 0 10396 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_109
timestamp 1635444444
transform 1 0 11132 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_89
timestamp 1635444444
transform 1 0 9292 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_112
timestamp 1635444444
transform 1 0 11408 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_124
timestamp 1635444444
transform 1 0 12512 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1635444444
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1635444444
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1635444444
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_136
timestamp 1635444444
transform 1 0 13616 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1635444444
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1635444444
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1635444444
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1635444444
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1635444444
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1635444444
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1635444444
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1635444444
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1635444444
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1635444444
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1635444444
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1635444444
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1635444444
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1635444444
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1635444444
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1635444444
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1635444444
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1635444444
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1635444444
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1635444444
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1635444444
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1635444444
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1635444444
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1635444444
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1635444444
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1635444444
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1635444444
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1635444444
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1635444444
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1635444444
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1635444444
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1635444444
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1635444444
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1635444444
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1635444444
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1635444444
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1635444444
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1635444444
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1635444444
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1635444444
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1635444444
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1635444444
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1635444444
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_309
timestamp 1635444444
transform 1 0 29532 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_317
timestamp 1635444444
transform 1 0 30268 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_73_317
timestamp 1635444444
transform 1 0 30268 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1635444444
transform -1 0 30820 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1635444444
transform -1 0 30820 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1635444444
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_18
timestamp 1635444444
transform 1 0 2760 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_7
timestamp 1635444444
transform 1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1635444444
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1488_
timestamp 1635444444
transform 1 0 2116 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1635444444
transform -1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_26
timestamp 1635444444
transform 1 0 3496 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_32
timestamp 1635444444
transform 1 0 4048 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_36
timestamp 1635444444
transform 1 0 4416 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1635444444
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0984_
timestamp 1635444444
transform -1 0 4048 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1491_
timestamp 1635444444
transform -1 0 5152 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_74_44
timestamp 1635444444
transform 1 0 5152 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_52
timestamp 1635444444
transform 1 0 5888 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_56
timestamp 1635444444
transform 1 0 6256 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1234_
timestamp 1635444444
transform -1 0 7452 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1242_
timestamp 1635444444
transform 1 0 5980 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_69
timestamp 1635444444
transform 1 0 7452 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_80
timestamp 1635444444
transform 1 0 8464 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1635444444
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1219_
timestamp 1635444444
transform -1 0 9200 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1220_
timestamp 1635444444
transform 1 0 8188 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_100
timestamp 1635444444
transform 1 0 10304 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_88
timestamp 1635444444
transform 1 0 9200 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_112
timestamp 1635444444
transform 1 0 11408 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_124
timestamp 1635444444
transform 1 0 12512 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_136
timestamp 1635444444
transform 1 0 13616 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1635444444
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1635444444
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1635444444
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1635444444
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1635444444
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1635444444
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1635444444
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1635444444
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_197
timestamp 1635444444
transform 1 0 19228 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_206
timestamp 1635444444
transform 1 0 20056 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_218
timestamp 1635444444
transform 1 0 21160 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _0942_
timestamp 1635444444
transform -1 0 20056 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_230
timestamp 1635444444
transform 1 0 22264 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_242
timestamp 1635444444
transform 1 0 23368 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1635444444
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1635444444
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1635444444
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1635444444
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1635444444
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1635444444
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1635444444
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1635444444
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_309
timestamp 1635444444
transform 1 0 29532 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_317
timestamp 1635444444
transform 1 0 30268 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1635444444
transform -1 0 30820 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1635444444
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_14
timestamp 1635444444
transform 1 0 2392 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_21
timestamp 1635444444
transform 1 0 3036 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_7
timestamp 1635444444
transform 1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1635444444
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1469_
timestamp 1635444444
transform 1 0 2116 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1473_
timestamp 1635444444
transform -1 0 3036 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1635444444
transform -1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_28
timestamp 1635444444
transform 1 0 3680 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_35
timestamp 1635444444
transform 1 0 4324 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_42
timestamp 1635444444
transform 1 0 4968 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1475_
timestamp 1635444444
transform 1 0 3404 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1480_
timestamp 1635444444
transform 1 0 4048 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1487_
timestamp 1635444444
transform 1 0 4692 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_75_48
timestamp 1635444444
transform 1 0 5520 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_52
timestamp 1635444444
transform 1 0 5888 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_60
timestamp 1635444444
transform 1 0 6624 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1635444444
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1232_
timestamp 1635444444
transform -1 0 6624 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1235_
timestamp 1635444444
transform 1 0 5612 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_77
timestamp 1635444444
transform 1 0 8188 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1230_
timestamp 1635444444
transform 1 0 7360 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1635444444
transform 1 0 8556 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_75_104
timestamp 1635444444
transform 1 0 10672 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_97
timestamp 1635444444
transform 1 0 10028 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1228_
timestamp 1635444444
transform -1 0 10672 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1635444444
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1635444444
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1635444444
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1635444444
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1635444444
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1635444444
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1635444444
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1635444444
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1635444444
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1635444444
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1635444444
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1635444444
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1635444444
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1635444444
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1635444444
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1635444444
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1635444444
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1635444444
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1635444444
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1635444444
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1635444444
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1635444444
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1635444444
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1635444444
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_305
timestamp 1635444444
transform 1 0 29164 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_316
timestamp 1635444444
transform 1 0 30176 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1635444444
transform -1 0 30820 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1635444444
transform 1 0 29900 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_14
timestamp 1635444444
transform 1 0 2392 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_21
timestamp 1635444444
transform 1 0 3036 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_7
timestamp 1635444444
transform 1 0 1748 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1635444444
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1471_
timestamp 1635444444
transform -1 0 2392 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1478_
timestamp 1635444444
transform 1 0 2760 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1635444444
transform -1 0 1748 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1635444444
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_32
timestamp 1635444444
transform 1 0 4048 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_40
timestamp 1635444444
transform 1 0 4784 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1635444444
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1485_
timestamp 1635444444
transform 1 0 3772 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1495_
timestamp 1635444444
transform 1 0 4876 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_76_48
timestamp 1635444444
transform 1 0 5520 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1635444444
transform 1 0 5888 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_76_68
timestamp 1635444444
transform 1 0 7360 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_76
timestamp 1635444444
transform 1 0 8096 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_80
timestamp 1635444444
transform 1 0 8464 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1635444444
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1229_
timestamp 1635444444
transform 1 0 8188 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1635444444
transform 1 0 8924 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_101
timestamp 1635444444
transform 1 0 10396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_113
timestamp 1635444444
transform 1 0 11500 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_125
timestamp 1635444444
transform 1 0 12604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_137
timestamp 1635444444
transform 1 0 13708 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1635444444
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1635444444
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1635444444
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1635444444
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1635444444
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1635444444
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1635444444
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1635444444
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_197
timestamp 1635444444
transform 1 0 19228 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_211
timestamp 1635444444
transform 1 0 20516 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _0934_
timestamp 1635444444
transform -1 0 20516 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0938_
timestamp 1635444444
transform -1 0 21436 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1635444444
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1635444444
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1635444444
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1635444444
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1635444444
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1635444444
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1635444444
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1635444444
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1635444444
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1635444444
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1635444444
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_309
timestamp 1635444444
transform 1 0 29532 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_317
timestamp 1635444444
transform 1 0 30268 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1635444444
transform -1 0 30820 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1635444444
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_14
timestamp 1635444444
transform 1 0 2392 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_21
timestamp 1635444444
transform 1 0 3036 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_7
timestamp 1635444444
transform 1 0 1748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1635444444
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1477_
timestamp 1635444444
transform 1 0 2116 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1483_
timestamp 1635444444
transform 1 0 2760 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1635444444
transform -1 0 1748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_29
timestamp 1635444444
transform 1 0 3772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_37
timestamp 1635444444
transform 1 0 4508 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1493_
timestamp 1635444444
transform -1 0 5520 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1499_
timestamp 1635444444
transform 1 0 3864 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_77_48
timestamp 1635444444
transform 1 0 5520 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_57
timestamp 1635444444
transform 1 0 6348 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1635444444
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1635444444
transform 1 0 6716 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_77_77
timestamp 1635444444
transform 1 0 8188 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1227_
timestamp 1635444444
transform -1 0 9384 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_77_102
timestamp 1635444444
transform 1 0 10488 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_90
timestamp 1635444444
transform 1 0 9384 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_110
timestamp 1635444444
transform 1 0 11224 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1635444444
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1635444444
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1635444444
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1635444444
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1635444444
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1635444444
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1635444444
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1635444444
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1635444444
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1635444444
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1635444444
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1635444444
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1635444444
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1635444444
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1635444444
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1635444444
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1635444444
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1635444444
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1635444444
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1635444444
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1635444444
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1635444444
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1635444444
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1635444444
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1635444444
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_317
timestamp 1635444444
transform 1 0 30268 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1635444444
transform -1 0 30820 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_15
timestamp 1635444444
transform 1 0 2484 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_7
timestamp 1635444444
transform 1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1635444444
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1489_
timestamp 1635444444
transform 1 0 2852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1635444444
transform -1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1635444444
transform -1 0 2484 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_22
timestamp 1635444444
transform 1 0 3128 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_78_29
timestamp 1635444444
transform 1 0 3772 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_35
timestamp 1635444444
transform 1 0 4324 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1635444444
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1490_
timestamp 1635444444
transform -1 0 4324 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1497_
timestamp 1635444444
transform 1 0 4692 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_78_46
timestamp 1635444444
transform 1 0 5336 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_53
timestamp 1635444444
transform 1 0 5980 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_61
timestamp 1635444444
transform 1 0 6716 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1233_
timestamp 1635444444
transform 1 0 5704 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1237_
timestamp 1635444444
transform -1 0 7636 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_78_71
timestamp 1635444444
transform 1 0 7636 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_78
timestamp 1635444444
transform 1 0 8280 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1635444444
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1635444444
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1635444444
transform 1 0 8004 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1635444444
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1635444444
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1635444444
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1635444444
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1635444444
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1635444444
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1635444444
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1635444444
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1635444444
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1635444444
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1635444444
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1635444444
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1635444444
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1635444444
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1635444444
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1635444444
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1635444444
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1635444444
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1635444444
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1635444444
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1635444444
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1635444444
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1635444444
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1635444444
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1635444444
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1635444444
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_309
timestamp 1635444444
transform 1 0 29532 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_316
timestamp 1635444444
transform 1 0 30176 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1635444444
transform -1 0 30820 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1635444444
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1635444444
transform 1 0 29900 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_15
timestamp 1635444444
transform 1 0 2484 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_7
timestamp 1635444444
transform 1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1635444444
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1635444444
transform -1 0 2484 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1635444444
transform -1 0 3220 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1635444444
transform -1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_23
timestamp 1635444444
transform 1 0 3220 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_27
timestamp 1635444444
transform 1 0 3588 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_32
timestamp 1635444444
transform 1 0 4048 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_39
timestamp 1635444444
transform 1 0 4692 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1635444444
transform 1 0 3680 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1635444444
transform 1 0 3772 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1494_
timestamp 1635444444
transform 1 0 4416 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1635444444
transform 1 0 5060 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_46
timestamp 1635444444
transform 1 0 5336 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_54
timestamp 1635444444
transform 1 0 6072 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_57
timestamp 1635444444
transform 1 0 6348 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_61
timestamp 1635444444
transform 1 0 6716 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1635444444
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1236_
timestamp 1635444444
transform 1 0 6440 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 1635444444
transform 1 0 7084 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_68
timestamp 1635444444
transform 1 0 7360 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_80
timestamp 1635444444
transform 1 0 8464 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_85
timestamp 1635444444
transform 1 0 8924 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1635444444
transform 1 0 8832 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_109
timestamp 1635444444
transform 1 0 11132 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_97
timestamp 1635444444
transform 1 0 10028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1635444444
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1635444444
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1635444444
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_137
timestamp 1635444444
transform 1 0 13708 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_141
timestamp 1635444444
transform 1 0 14076 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1635444444
transform 1 0 13984 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_153
timestamp 1635444444
transform 1 0 15180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_165
timestamp 1635444444
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1635444444
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1635444444
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1635444444
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_193
timestamp 1635444444
transform 1 0 18860 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1635444444
transform 1 0 19136 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_197
timestamp 1635444444
transform 1 0 19228 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_209
timestamp 1635444444
transform 1 0 20332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_221
timestamp 1635444444
transform 1 0 21436 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1635444444
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1635444444
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1635444444
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_249
timestamp 1635444444
transform 1 0 24012 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_253
timestamp 1635444444
transform 1 0 24380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1635444444
transform 1 0 24288 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_265
timestamp 1635444444
transform 1 0 25484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_277
timestamp 1635444444
transform 1 0 26588 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1635444444
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1635444444
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1635444444
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_305
timestamp 1635444444
transform 1 0 29164 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_309
timestamp 1635444444
transform 1 0 29532 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_316
timestamp 1635444444
transform 1 0 30176 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1635444444
transform -1 0 30820 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1635444444
transform 1 0 29440 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1635444444
transform 1 0 29900 0 -1 45696
box -38 -48 314 592
<< labels >>
rlabel metal3 s 31200 4904 32000 5024 6 hb_clk_o
port 0 nsew signal tristate
rlabel metal3 s 31200 6944 32000 7064 6 hb_clkn_o
port 1 nsew signal tristate
rlabel metal3 s 31200 2864 32000 2984 6 hb_csn_o
port 2 nsew signal tristate
rlabel metal3 s 31200 32920 32000 33040 6 hb_dq_i[0]
port 3 nsew signal input
rlabel metal3 s 31200 34960 32000 35080 6 hb_dq_i[1]
port 4 nsew signal input
rlabel metal3 s 31200 36864 32000 36984 6 hb_dq_i[2]
port 5 nsew signal input
rlabel metal3 s 31200 38904 32000 39024 6 hb_dq_i[3]
port 6 nsew signal input
rlabel metal3 s 31200 40944 32000 41064 6 hb_dq_i[4]
port 7 nsew signal input
rlabel metal3 s 31200 42848 32000 42968 6 hb_dq_i[5]
port 8 nsew signal input
rlabel metal3 s 31200 44888 32000 45008 6 hb_dq_i[6]
port 9 nsew signal input
rlabel metal3 s 31200 46928 32000 47048 6 hb_dq_i[7]
port 10 nsew signal input
rlabel metal3 s 31200 14832 32000 14952 6 hb_dq_o[0]
port 11 nsew signal tristate
rlabel metal3 s 31200 16872 32000 16992 6 hb_dq_o[1]
port 12 nsew signal tristate
rlabel metal3 s 31200 18912 32000 19032 6 hb_dq_o[2]
port 13 nsew signal tristate
rlabel metal3 s 31200 20952 32000 21072 6 hb_dq_o[3]
port 14 nsew signal tristate
rlabel metal3 s 31200 22856 32000 22976 6 hb_dq_o[4]
port 15 nsew signal tristate
rlabel metal3 s 31200 24896 32000 25016 6 hb_dq_o[5]
port 16 nsew signal tristate
rlabel metal3 s 31200 26936 32000 27056 6 hb_dq_o[6]
port 17 nsew signal tristate
rlabel metal3 s 31200 28840 32000 28960 6 hb_dq_o[7]
port 18 nsew signal tristate
rlabel metal3 s 31200 12928 32000 13048 6 hb_dq_oen
port 19 nsew signal tristate
rlabel metal3 s 31200 960 32000 1080 6 hb_rstn_o
port 20 nsew signal tristate
rlabel metal3 s 31200 30880 32000 31000 6 hb_rwds_i
port 21 nsew signal input
rlabel metal3 s 31200 8848 32000 8968 6 hb_rwds_o
port 22 nsew signal tristate
rlabel metal3 s 31200 10888 32000 11008 6 hb_rwds_oen
port 23 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 rst_i
port 24 nsew signal input
rlabel metal4 s 5909 2128 6229 45744 6 vccd1
port 25 nsew power input
rlabel metal4 s 15839 2128 16159 45744 6 vccd1
port 25 nsew power input
rlabel metal4 s 25770 2128 26090 45744 6 vccd1
port 25 nsew power input
rlabel metal4 s 10874 2128 11194 45744 6 vssd1
port 26 nsew ground input
rlabel metal4 s 20805 2128 21125 45744 6 vssd1
port 26 nsew ground input
rlabel metal2 s 1122 0 1178 800 6 wb_clk_i
port 27 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wb_rst_i
port 28 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 wbs_ack_o
port 29 nsew signal tristate
rlabel metal2 s 7930 0 7986 800 6 wbs_adr_i[0]
port 30 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[10]
port 31 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[11]
port 32 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_adr_i[12]
port 33 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[13]
port 34 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[14]
port 35 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[15]
port 36 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[16]
port 37 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[17]
port 38 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_adr_i[18]
port 39 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[19]
port 40 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[1]
port 41 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_adr_i[20]
port 42 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[21]
port 43 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[22]
port 44 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[23]
port 45 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[24]
port 46 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_adr_i[25]
port 47 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_adr_i[26]
port 48 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[27]
port 49 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[28]
port 50 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[29]
port 51 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_adr_i[2]
port 52 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[30]
port 53 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_adr_i[31]
port 54 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[3]
port 55 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_adr_i[4]
port 56 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_adr_i[5]
port 57 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[6]
port 58 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[7]
port 59 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_adr_i[8]
port 60 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[9]
port 61 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_cyc_i
port 62 nsew signal input
rlabel metal3 s 0 280 800 400 6 wbs_dat_i[0]
port 63 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 wbs_dat_i[10]
port 64 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 wbs_dat_i[11]
port 65 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 wbs_dat_i[12]
port 66 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 wbs_dat_i[13]
port 67 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 wbs_dat_i[14]
port 68 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 wbs_dat_i[15]
port 69 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 wbs_dat_i[16]
port 70 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 wbs_dat_i[17]
port 71 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 wbs_dat_i[18]
port 72 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 wbs_dat_i[19]
port 73 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wbs_dat_i[1]
port 74 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 wbs_dat_i[20]
port 75 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 wbs_dat_i[21]
port 76 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 wbs_dat_i[22]
port 77 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 wbs_dat_i[23]
port 78 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 wbs_dat_i[24]
port 79 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 wbs_dat_i[25]
port 80 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wbs_dat_i[26]
port 81 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 wbs_dat_i[27]
port 82 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 wbs_dat_i[28]
port 83 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 wbs_dat_i[29]
port 84 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 wbs_dat_i[2]
port 85 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 wbs_dat_i[30]
port 86 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wbs_dat_i[31]
port 87 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 wbs_dat_i[3]
port 88 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 wbs_dat_i[4]
port 89 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 wbs_dat_i[5]
port 90 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 wbs_dat_i[6]
port 91 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 wbs_dat_i[7]
port 92 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wbs_dat_i[8]
port 93 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wbs_dat_i[9]
port 94 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 wbs_dat_o[0]
port 95 nsew signal tristate
rlabel metal3 s 0 31288 800 31408 6 wbs_dat_o[10]
port 96 nsew signal tristate
rlabel metal3 s 0 31968 800 32088 6 wbs_dat_o[11]
port 97 nsew signal tristate
rlabel metal3 s 0 32648 800 32768 6 wbs_dat_o[12]
port 98 nsew signal tristate
rlabel metal3 s 0 33464 800 33584 6 wbs_dat_o[13]
port 99 nsew signal tristate
rlabel metal3 s 0 34144 800 34264 6 wbs_dat_o[14]
port 100 nsew signal tristate
rlabel metal3 s 0 34960 800 35080 6 wbs_dat_o[15]
port 101 nsew signal tristate
rlabel metal3 s 0 35640 800 35760 6 wbs_dat_o[16]
port 102 nsew signal tristate
rlabel metal3 s 0 36456 800 36576 6 wbs_dat_o[17]
port 103 nsew signal tristate
rlabel metal3 s 0 37136 800 37256 6 wbs_dat_o[18]
port 104 nsew signal tristate
rlabel metal3 s 0 37816 800 37936 6 wbs_dat_o[19]
port 105 nsew signal tristate
rlabel metal3 s 0 24624 800 24744 6 wbs_dat_o[1]
port 106 nsew signal tristate
rlabel metal3 s 0 38632 800 38752 6 wbs_dat_o[20]
port 107 nsew signal tristate
rlabel metal3 s 0 39312 800 39432 6 wbs_dat_o[21]
port 108 nsew signal tristate
rlabel metal3 s 0 40128 800 40248 6 wbs_dat_o[22]
port 109 nsew signal tristate
rlabel metal3 s 0 40808 800 40928 6 wbs_dat_o[23]
port 110 nsew signal tristate
rlabel metal3 s 0 41624 800 41744 6 wbs_dat_o[24]
port 111 nsew signal tristate
rlabel metal3 s 0 42304 800 42424 6 wbs_dat_o[25]
port 112 nsew signal tristate
rlabel metal3 s 0 42984 800 43104 6 wbs_dat_o[26]
port 113 nsew signal tristate
rlabel metal3 s 0 43800 800 43920 6 wbs_dat_o[27]
port 114 nsew signal tristate
rlabel metal3 s 0 44480 800 44600 6 wbs_dat_o[28]
port 115 nsew signal tristate
rlabel metal3 s 0 45296 800 45416 6 wbs_dat_o[29]
port 116 nsew signal tristate
rlabel metal3 s 0 25304 800 25424 6 wbs_dat_o[2]
port 117 nsew signal tristate
rlabel metal3 s 0 45976 800 46096 6 wbs_dat_o[30]
port 118 nsew signal tristate
rlabel metal3 s 0 46792 800 46912 6 wbs_dat_o[31]
port 119 nsew signal tristate
rlabel metal3 s 0 26120 800 26240 6 wbs_dat_o[3]
port 120 nsew signal tristate
rlabel metal3 s 0 26800 800 26920 6 wbs_dat_o[4]
port 121 nsew signal tristate
rlabel metal3 s 0 27480 800 27600 6 wbs_dat_o[5]
port 122 nsew signal tristate
rlabel metal3 s 0 28296 800 28416 6 wbs_dat_o[6]
port 123 nsew signal tristate
rlabel metal3 s 0 28976 800 29096 6 wbs_dat_o[7]
port 124 nsew signal tristate
rlabel metal3 s 0 29792 800 29912 6 wbs_dat_o[8]
port 125 nsew signal tristate
rlabel metal3 s 0 30472 800 30592 6 wbs_dat_o[9]
port 126 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 wbs_sel_i[0]
port 127 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_sel_i[1]
port 128 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_sel_i[2]
port 129 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_sel_i[3]
port 130 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_stb_i
port 131 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_we_i
port 132 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32000 48000
<< end >>
