magic
tech sky130A
magscale 1 2
timestamp 1636594562
<< locali >>
rect 7573 43775 7607 43945
rect 3801 38199 3835 38369
rect 13737 37655 13771 37757
rect 19533 33439 19567 33609
rect 20177 29699 20211 29801
rect 7849 23715 7883 23817
rect 17601 23103 17635 23205
rect 17417 13311 17451 13481
rect 8769 10999 8803 11169
rect 9137 10455 9171 10625
rect 19073 8959 19107 9129
rect 3893 5083 3927 5253
<< viali >>
rect 1685 45441 1719 45475
rect 2421 45441 2455 45475
rect 3157 45441 3191 45475
rect 3985 45441 4019 45475
rect 4629 45441 4663 45475
rect 30113 45441 30147 45475
rect 2237 45305 2271 45339
rect 2973 45305 3007 45339
rect 3801 45305 3835 45339
rect 1501 45237 1535 45271
rect 4445 45237 4479 45271
rect 29929 45237 29963 45271
rect 2237 45033 2271 45067
rect 4445 45033 4479 45067
rect 5457 45033 5491 45067
rect 1685 44829 1719 44863
rect 2421 44829 2455 44863
rect 3065 44829 3099 44863
rect 3985 44829 4019 44863
rect 4629 44829 4663 44863
rect 5825 44829 5859 44863
rect 6653 44829 6687 44863
rect 9137 44829 9171 44863
rect 30113 44829 30147 44863
rect 6920 44761 6954 44795
rect 1501 44693 1535 44727
rect 2881 44693 2915 44727
rect 3801 44693 3835 44727
rect 5273 44693 5307 44727
rect 5457 44693 5491 44727
rect 8033 44693 8067 44727
rect 8953 44693 8987 44727
rect 29929 44693 29963 44727
rect 4813 44489 4847 44523
rect 5273 44489 5307 44523
rect 6561 44489 6595 44523
rect 7021 44489 7055 44523
rect 4629 44421 4663 44455
rect 5457 44421 5491 44455
rect 1685 44353 1719 44387
rect 2329 44353 2363 44387
rect 2973 44353 3007 44387
rect 3617 44353 3651 44387
rect 6377 44353 6411 44387
rect 7205 44353 7239 44387
rect 7573 44353 7607 44387
rect 7757 44353 7791 44387
rect 8217 44353 8251 44387
rect 8401 44353 8435 44387
rect 8585 44353 8619 44387
rect 8769 44353 8803 44387
rect 9413 44353 9447 44387
rect 18337 44353 18371 44387
rect 30113 44353 30147 44387
rect 7389 44285 7423 44319
rect 7481 44285 7515 44319
rect 8493 44285 8527 44319
rect 18521 44285 18555 44319
rect 4261 44217 4295 44251
rect 5825 44217 5859 44251
rect 8953 44217 8987 44251
rect 1501 44149 1535 44183
rect 2145 44149 2179 44183
rect 2789 44149 2823 44183
rect 3433 44149 3467 44183
rect 4629 44149 4663 44183
rect 5457 44149 5491 44183
rect 9597 44149 9631 44183
rect 18153 44149 18187 44183
rect 29929 44149 29963 44183
rect 5273 43945 5307 43979
rect 5457 43945 5491 43979
rect 6561 43945 6595 43979
rect 7573 43945 7607 43979
rect 18153 43945 18187 43979
rect 2513 43877 2547 43911
rect 10333 43877 10367 43911
rect 8033 43809 8067 43843
rect 8953 43809 8987 43843
rect 1869 43741 1903 43775
rect 2329 43741 2363 43775
rect 3157 43741 3191 43775
rect 3801 43741 3835 43775
rect 5825 43741 5859 43775
rect 6745 43741 6779 43775
rect 7573 43741 7607 43775
rect 7665 43741 7699 43775
rect 7849 43741 7883 43775
rect 7941 43741 7975 43775
rect 8217 43741 8251 43775
rect 18337 43741 18371 43775
rect 18521 43741 18555 43775
rect 8401 43673 8435 43707
rect 9198 43673 9232 43707
rect 1685 43605 1719 43639
rect 2973 43605 3007 43639
rect 3985 43605 4019 43639
rect 5457 43605 5491 43639
rect 8125 43401 8159 43435
rect 8861 43401 8895 43435
rect 18153 43401 18187 43435
rect 9974 43333 10008 43367
rect 1685 43265 1719 43299
rect 2513 43265 2547 43299
rect 3893 43265 3927 43299
rect 4537 43265 4571 43299
rect 4997 43265 5031 43299
rect 5641 43265 5675 43299
rect 7012 43265 7046 43299
rect 10241 43265 10275 43299
rect 18337 43265 18371 43299
rect 6745 43197 6779 43231
rect 18521 43197 18555 43231
rect 1501 43061 1535 43095
rect 2697 43061 2731 43095
rect 3709 43061 3743 43095
rect 4353 43061 4387 43095
rect 5181 43061 5215 43095
rect 5825 43061 5859 43095
rect 6193 42857 6227 42891
rect 7021 42857 7055 42891
rect 1685 42653 1719 42687
rect 2145 42653 2179 42687
rect 3065 42653 3099 42687
rect 4169 42653 4203 42687
rect 6561 42653 6595 42687
rect 7205 42653 7239 42687
rect 7389 42653 7423 42687
rect 7478 42653 7512 42687
rect 7573 42653 7607 42687
rect 7757 42653 7791 42687
rect 8217 42653 8251 42687
rect 8953 42653 8987 42687
rect 30113 42653 30147 42687
rect 4436 42585 4470 42619
rect 1501 42517 1535 42551
rect 2329 42517 2363 42551
rect 3249 42517 3283 42551
rect 5549 42517 5583 42551
rect 6009 42517 6043 42551
rect 6193 42517 6227 42551
rect 8401 42517 8435 42551
rect 9137 42517 9171 42551
rect 29929 42517 29963 42551
rect 5273 42313 5307 42347
rect 6745 42313 6779 42347
rect 7941 42313 7975 42347
rect 5457 42245 5491 42279
rect 1685 42177 1719 42211
rect 2329 42177 2363 42211
rect 2789 42177 2823 42211
rect 3056 42177 3090 42211
rect 4813 42177 4847 42211
rect 5825 42177 5859 42211
rect 6929 42177 6963 42211
rect 9054 42177 9088 42211
rect 9321 42109 9355 42143
rect 4629 42041 4663 42075
rect 1501 41973 1535 42007
rect 2145 41973 2179 42007
rect 4169 41973 4203 42007
rect 5457 41973 5491 42007
rect 2881 41769 2915 41803
rect 4445 41769 4479 41803
rect 5641 41769 5675 41803
rect 5825 41769 5859 41803
rect 8125 41769 8159 41803
rect 9137 41769 9171 41803
rect 6193 41701 6227 41735
rect 6929 41701 6963 41735
rect 4905 41633 4939 41667
rect 21373 41633 21407 41667
rect 1869 41565 1903 41599
rect 3065 41565 3099 41599
rect 3985 41565 4019 41599
rect 4629 41565 4663 41599
rect 4813 41565 4847 41599
rect 4997 41565 5031 41599
rect 5181 41565 5215 41599
rect 6745 41565 6779 41599
rect 7389 41565 7423 41599
rect 7573 41565 7607 41599
rect 7665 41565 7699 41599
rect 7757 41565 7791 41599
rect 7941 41565 7975 41599
rect 8953 41565 8987 41599
rect 13001 41565 13035 41599
rect 15945 41565 15979 41599
rect 21833 41565 21867 41599
rect 21925 41565 21959 41599
rect 5825 41497 5859 41531
rect 1685 41429 1719 41463
rect 3801 41429 3835 41463
rect 12817 41429 12851 41463
rect 16129 41429 16163 41463
rect 2421 41225 2455 41259
rect 3433 41225 3467 41259
rect 5273 41225 5307 41259
rect 6561 41225 6595 41259
rect 21925 41225 21959 41259
rect 2605 41157 2639 41191
rect 5457 41157 5491 41191
rect 1685 41089 1719 41123
rect 3617 41089 3651 41123
rect 3985 41089 4019 41123
rect 4169 41089 4203 41123
rect 4629 41089 4663 41123
rect 7674 41089 7708 41123
rect 8677 41089 8711 41123
rect 15025 41089 15059 41123
rect 15117 41089 15151 41123
rect 15669 41089 15703 41123
rect 15853 41089 15887 41123
rect 16681 41089 16715 41123
rect 17417 41089 17451 41123
rect 22109 41089 22143 41123
rect 30113 41089 30147 41123
rect 3801 41021 3835 41055
rect 3893 41021 3927 41055
rect 7941 41021 7975 41055
rect 8401 41021 8435 41055
rect 12633 41021 12667 41055
rect 12817 41021 12851 41055
rect 13553 41021 13587 41055
rect 13691 41021 13725 41055
rect 13829 41021 13863 41055
rect 22293 41021 22327 41055
rect 2973 40953 3007 40987
rect 5825 40953 5859 40987
rect 13277 40953 13311 40987
rect 29929 40953 29963 40987
rect 1501 40885 1535 40919
rect 2605 40885 2639 40919
rect 4813 40885 4847 40919
rect 5457 40885 5491 40919
rect 14473 40885 14507 40919
rect 16037 40885 16071 40919
rect 16681 40885 16715 40919
rect 17417 40885 17451 40919
rect 6653 40681 6687 40715
rect 9597 40681 9631 40715
rect 12541 40681 12575 40715
rect 4997 40613 5031 40647
rect 4261 40545 4295 40579
rect 6285 40545 6319 40579
rect 7389 40545 7423 40579
rect 14565 40545 14599 40579
rect 14749 40545 14783 40579
rect 16129 40545 16163 40579
rect 16773 40545 16807 40579
rect 17049 40545 17083 40579
rect 17187 40545 17221 40579
rect 1685 40477 1719 40511
rect 2605 40477 2639 40511
rect 3985 40477 4019 40511
rect 4169 40477 4203 40511
rect 4353 40477 4387 40511
rect 4537 40477 4571 40511
rect 5181 40477 5215 40511
rect 5917 40477 5951 40511
rect 6101 40477 6135 40511
rect 6193 40477 6227 40511
rect 6469 40477 6503 40511
rect 7113 40477 7147 40511
rect 8953 40477 8987 40511
rect 9781 40477 9815 40511
rect 12357 40477 12391 40511
rect 13001 40477 13035 40511
rect 16313 40477 16347 40511
rect 17325 40477 17359 40511
rect 18613 40477 18647 40511
rect 1501 40341 1535 40375
rect 2789 40341 2823 40375
rect 3801 40341 3835 40375
rect 9137 40341 9171 40375
rect 13185 40341 13219 40375
rect 14841 40341 14875 40375
rect 15209 40341 15243 40375
rect 17969 40341 18003 40375
rect 18429 40341 18463 40375
rect 2237 40137 2271 40171
rect 4261 40137 4295 40171
rect 7665 40137 7699 40171
rect 8585 40137 8619 40171
rect 9229 40137 9263 40171
rect 14657 40137 14691 40171
rect 16865 40137 16899 40171
rect 17509 40137 17543 40171
rect 17877 40137 17911 40171
rect 3148 40069 3182 40103
rect 5457 40069 5491 40103
rect 15577 40069 15611 40103
rect 17969 40069 18003 40103
rect 18889 40069 18923 40103
rect 19809 40069 19843 40103
rect 19993 40069 20027 40103
rect 1869 40001 1903 40035
rect 5825 40001 5859 40035
rect 6837 40001 6871 40035
rect 7481 40001 7515 40035
rect 8401 40001 8435 40035
rect 9045 40001 9079 40035
rect 9873 40001 9907 40035
rect 12817 40001 12851 40035
rect 13001 40001 13035 40035
rect 15761 40001 15795 40035
rect 16681 40001 16715 40035
rect 18705 40001 18739 40035
rect 2881 39933 2915 39967
rect 13737 39933 13771 39967
rect 13854 39933 13888 39967
rect 14013 39933 14047 39967
rect 18061 39933 18095 39967
rect 5273 39865 5307 39899
rect 13461 39865 13495 39899
rect 15945 39865 15979 39899
rect 2237 39797 2271 39831
rect 2421 39797 2455 39831
rect 5457 39797 5491 39831
rect 6929 39797 6963 39831
rect 9689 39797 9723 39831
rect 19073 39797 19107 39831
rect 20177 39797 20211 39831
rect 2881 39593 2915 39627
rect 5825 39593 5859 39627
rect 8217 39593 8251 39627
rect 13001 39593 13035 39627
rect 18521 39593 18555 39627
rect 15301 39525 15335 39559
rect 20545 39525 20579 39559
rect 9413 39457 9447 39491
rect 14657 39457 14691 39491
rect 15694 39457 15728 39491
rect 17049 39457 17083 39491
rect 1685 39389 1719 39423
rect 2421 39389 2455 39423
rect 3065 39389 3099 39423
rect 3801 39389 3835 39423
rect 4537 39389 4571 39423
rect 5365 39389 5399 39423
rect 6009 39389 6043 39423
rect 6469 39389 6503 39423
rect 6653 39389 6687 39423
rect 6745 39389 6779 39423
rect 6883 39389 6917 39423
rect 7021 39389 7055 39423
rect 8401 39389 8435 39423
rect 12633 39389 12667 39423
rect 14841 39389 14875 39423
rect 15577 39389 15611 39423
rect 15853 39389 15887 39423
rect 18153 39389 18187 39423
rect 19441 39389 19475 39423
rect 21741 39389 21775 39423
rect 21925 39389 21959 39423
rect 30113 39389 30147 39423
rect 9680 39321 9714 39355
rect 12817 39321 12851 39355
rect 16497 39321 16531 39355
rect 17325 39321 17359 39355
rect 18337 39321 18371 39355
rect 19993 39321 20027 39355
rect 20269 39321 20303 39355
rect 1501 39253 1535 39287
rect 2237 39253 2271 39287
rect 3985 39253 4019 39287
rect 4721 39253 4755 39287
rect 5181 39253 5215 39287
rect 7205 39253 7239 39287
rect 10793 39253 10827 39287
rect 17233 39253 17267 39287
rect 17693 39253 17727 39287
rect 19257 39253 19291 39287
rect 20085 39253 20119 39287
rect 21557 39253 21591 39287
rect 29929 39253 29963 39287
rect 2421 39049 2455 39083
rect 8217 39049 8251 39083
rect 13553 39049 13587 39083
rect 16129 39049 16163 39083
rect 19165 39049 19199 39083
rect 20269 39049 20303 39083
rect 2237 38981 2271 39015
rect 7104 38981 7138 39015
rect 13829 38981 13863 39015
rect 19073 38981 19107 39015
rect 2881 38913 2915 38947
rect 4077 38913 4111 38947
rect 4445 38913 4479 38947
rect 4629 38913 4663 38947
rect 5825 38913 5859 38947
rect 6837 38913 6871 38947
rect 9229 38913 9263 38947
rect 9496 38913 9530 38947
rect 13277 38913 13311 38947
rect 14289 38913 14323 38947
rect 15326 38913 15360 38947
rect 20085 38913 20119 38947
rect 1869 38845 1903 38879
rect 4261 38845 4295 38879
rect 4353 38845 4387 38879
rect 13185 38845 13219 38879
rect 14473 38845 14507 38879
rect 14933 38845 14967 38879
rect 15209 38845 15243 38879
rect 15485 38845 15519 38879
rect 18889 38845 18923 38879
rect 2237 38709 2271 38743
rect 3065 38709 3099 38743
rect 3893 38709 3927 38743
rect 5733 38709 5767 38743
rect 10609 38709 10643 38743
rect 19533 38709 19567 38743
rect 1869 38505 1903 38539
rect 2053 38505 2087 38539
rect 5365 38505 5399 38539
rect 12541 38505 12575 38539
rect 14289 38505 14323 38539
rect 17417 38505 17451 38539
rect 1501 38437 1535 38471
rect 18613 38437 18647 38471
rect 2881 38369 2915 38403
rect 3801 38369 3835 38403
rect 3985 38369 4019 38403
rect 6101 38369 6135 38403
rect 7481 38369 7515 38403
rect 9229 38369 9263 38403
rect 13001 38369 13035 38403
rect 2697 38301 2731 38335
rect 2973 38301 3007 38335
rect 3065 38301 3099 38335
rect 3249 38301 3283 38335
rect 1869 38233 1903 38267
rect 4252 38301 4286 38335
rect 5825 38301 5859 38335
rect 7297 38301 7331 38335
rect 7573 38301 7607 38335
rect 7665 38301 7699 38335
rect 7849 38301 7883 38335
rect 8953 38301 8987 38335
rect 9137 38301 9171 38335
rect 9321 38301 9355 38335
rect 9505 38301 9539 38335
rect 9689 38301 9723 38335
rect 10885 38301 10919 38335
rect 12357 38301 12391 38335
rect 13185 38301 13219 38335
rect 13369 38301 13403 38335
rect 14105 38301 14139 38335
rect 17601 38301 17635 38335
rect 18429 38301 18463 38335
rect 19441 38301 19475 38335
rect 30113 38301 30147 38335
rect 2513 38165 2547 38199
rect 3801 38165 3835 38199
rect 7113 38165 7147 38199
rect 10701 38165 10735 38199
rect 19257 38165 19291 38199
rect 29929 38165 29963 38199
rect 1961 37961 1995 37995
rect 2145 37961 2179 37995
rect 3065 37961 3099 37995
rect 9413 37961 9447 37995
rect 12725 37961 12759 37995
rect 13829 37961 13863 37995
rect 21925 37961 21959 37995
rect 4178 37893 4212 37927
rect 17693 37893 17727 37927
rect 5549 37825 5583 37859
rect 5825 37825 5859 37859
rect 8033 37825 8067 37859
rect 8677 37825 8711 37859
rect 8861 37825 8895 37859
rect 9229 37825 9263 37859
rect 9965 37825 9999 37859
rect 10609 37825 10643 37859
rect 11713 37825 11747 37859
rect 12909 37825 12943 37859
rect 13093 37825 13127 37859
rect 14013 37825 14047 37859
rect 14933 37825 14967 37859
rect 16865 37825 16899 37859
rect 17509 37825 17543 37859
rect 17877 37825 17911 37859
rect 18337 37825 18371 37859
rect 18981 37825 19015 37859
rect 19248 37825 19282 37859
rect 22109 37825 22143 37859
rect 2513 37757 2547 37791
rect 4445 37757 4479 37791
rect 6377 37757 6411 37791
rect 6653 37757 6687 37791
rect 8953 37757 8987 37791
rect 9045 37757 9079 37791
rect 13737 37757 13771 37791
rect 14289 37757 14323 37791
rect 14841 37757 14875 37791
rect 22293 37757 22327 37791
rect 10793 37689 10827 37723
rect 2145 37621 2179 37655
rect 8217 37621 8251 37655
rect 10149 37621 10183 37655
rect 11529 37621 11563 37655
rect 13093 37621 13127 37655
rect 13737 37621 13771 37655
rect 14197 37621 14231 37655
rect 17049 37621 17083 37655
rect 18521 37621 18555 37655
rect 20361 37621 20395 37655
rect 2237 37417 2271 37451
rect 6929 37417 6963 37451
rect 7481 37417 7515 37451
rect 12909 37417 12943 37451
rect 14105 37417 14139 37451
rect 12817 37349 12851 37383
rect 10885 37281 10919 37315
rect 13001 37281 13035 37315
rect 15577 37281 15611 37315
rect 15853 37281 15887 37315
rect 15991 37281 16025 37315
rect 17693 37281 17727 37315
rect 17877 37281 17911 37315
rect 1869 37213 1903 37247
rect 2881 37213 2915 37247
rect 3985 37213 4019 37247
rect 4629 37213 4663 37247
rect 5549 37213 5583 37247
rect 5816 37213 5850 37247
rect 7389 37213 7423 37247
rect 10333 37213 10367 37247
rect 12725 37213 12759 37247
rect 14105 37213 14139 37247
rect 14289 37213 14323 37247
rect 14933 37213 14967 37247
rect 15117 37213 15151 37247
rect 16129 37213 16163 37247
rect 17969 37213 18003 37247
rect 19441 37213 19475 37247
rect 20269 37213 20303 37247
rect 20453 37213 20487 37247
rect 2237 37145 2271 37179
rect 10066 37145 10100 37179
rect 11152 37145 11186 37179
rect 2421 37077 2455 37111
rect 3065 37077 3099 37111
rect 3801 37077 3835 37111
rect 4445 37077 4479 37111
rect 7849 37077 7883 37111
rect 8953 37077 8987 37111
rect 12265 37077 12299 37111
rect 16773 37077 16807 37111
rect 18337 37077 18371 37111
rect 19257 37077 19291 37111
rect 20361 37077 20395 37111
rect 3709 36873 3743 36907
rect 4997 36873 5031 36907
rect 8953 36873 8987 36907
rect 12909 36873 12943 36907
rect 13461 36873 13495 36907
rect 15761 36873 15795 36907
rect 17141 36873 17175 36907
rect 17509 36873 17543 36907
rect 10977 36805 11011 36839
rect 11774 36805 11808 36839
rect 1685 36737 1719 36771
rect 2145 36737 2179 36771
rect 2881 36737 2915 36771
rect 3525 36737 3559 36771
rect 4353 36737 4387 36771
rect 4813 36737 4847 36771
rect 5641 36737 5675 36771
rect 6837 36737 6871 36771
rect 8217 36737 8251 36771
rect 8401 36737 8435 36771
rect 8769 36737 8803 36771
rect 9597 36737 9631 36771
rect 10241 36737 10275 36771
rect 10425 36737 10459 36771
rect 10517 36737 10551 36771
rect 10793 36737 10827 36771
rect 11529 36737 11563 36771
rect 13369 36737 13403 36771
rect 14197 36737 14231 36771
rect 14565 36737 14599 36771
rect 15209 36737 15243 36771
rect 15485 36737 15519 36771
rect 15577 36737 15611 36771
rect 18337 36737 18371 36771
rect 18604 36737 18638 36771
rect 20545 36737 20579 36771
rect 22109 36737 22143 36771
rect 30113 36737 30147 36771
rect 6561 36669 6595 36703
rect 8493 36669 8527 36703
rect 8585 36669 8619 36703
rect 10609 36669 10643 36703
rect 14749 36669 14783 36703
rect 15301 36669 15335 36703
rect 16865 36669 16899 36703
rect 17049 36669 17083 36703
rect 20637 36669 20671 36703
rect 20729 36669 20763 36703
rect 22293 36669 22327 36703
rect 3065 36601 3099 36635
rect 5457 36601 5491 36635
rect 14289 36601 14323 36635
rect 19717 36601 19751 36635
rect 29929 36601 29963 36635
rect 1501 36533 1535 36567
rect 2329 36533 2363 36567
rect 4169 36533 4203 36567
rect 9781 36533 9815 36567
rect 20177 36533 20211 36567
rect 21925 36533 21959 36567
rect 5181 36329 5215 36363
rect 7205 36329 7239 36363
rect 9781 36329 9815 36363
rect 11069 36329 11103 36363
rect 14197 36329 14231 36363
rect 16773 36329 16807 36363
rect 18613 36329 18647 36363
rect 20545 36329 20579 36363
rect 3801 36261 3835 36295
rect 4721 36261 4755 36295
rect 11529 36261 11563 36295
rect 6377 36193 6411 36227
rect 6653 36193 6687 36227
rect 10609 36193 10643 36227
rect 10701 36193 10735 36227
rect 14933 36193 14967 36227
rect 15117 36193 15151 36227
rect 15577 36193 15611 36227
rect 15853 36193 15887 36227
rect 15991 36193 16025 36227
rect 21373 36193 21407 36227
rect 1685 36125 1719 36159
rect 2329 36125 2363 36159
rect 2789 36125 2823 36159
rect 3985 36125 4019 36159
rect 4537 36125 4571 36159
rect 5365 36125 5399 36159
rect 7113 36125 7147 36159
rect 8033 36125 8067 36159
rect 9137 36125 9171 36159
rect 9597 36125 9631 36159
rect 10333 36125 10367 36159
rect 10517 36125 10551 36159
rect 10885 36125 10919 36159
rect 11713 36125 11747 36159
rect 14105 36125 14139 36159
rect 14289 36125 14323 36159
rect 16129 36125 16163 36159
rect 17509 36125 17543 36159
rect 18429 36125 18463 36159
rect 18613 36125 18647 36159
rect 20085 36125 20119 36159
rect 20361 36125 20395 36159
rect 21097 36125 21131 36159
rect 1501 35989 1535 36023
rect 2145 35989 2179 36023
rect 2973 35989 3007 36023
rect 7573 35989 7607 36023
rect 8217 35989 8251 36023
rect 8953 35989 8987 36023
rect 17325 35989 17359 36023
rect 20177 35989 20211 36023
rect 2421 35785 2455 35819
rect 7021 35785 7055 35819
rect 8217 35785 8251 35819
rect 18245 35785 18279 35819
rect 18981 35785 19015 35819
rect 19165 35785 19199 35819
rect 20913 35785 20947 35819
rect 2237 35717 2271 35751
rect 1869 35649 1903 35683
rect 3157 35649 3191 35683
rect 3424 35649 3458 35683
rect 5181 35649 5215 35683
rect 5825 35649 5859 35683
rect 6837 35649 6871 35683
rect 8033 35649 8067 35683
rect 9413 35649 9447 35683
rect 9781 35649 9815 35683
rect 9965 35649 9999 35683
rect 10793 35649 10827 35683
rect 11529 35649 11563 35683
rect 17049 35649 17083 35683
rect 17877 35649 17911 35683
rect 18061 35649 18095 35683
rect 19162 35649 19196 35683
rect 20085 35649 20119 35683
rect 20269 35649 20303 35683
rect 20821 35649 20855 35683
rect 9597 35581 9631 35615
rect 9689 35581 9723 35615
rect 16773 35581 16807 35615
rect 16957 35581 16991 35615
rect 19625 35581 19659 35615
rect 2237 35445 2271 35479
rect 4537 35445 4571 35479
rect 4997 35445 5031 35479
rect 5641 35445 5675 35479
rect 9229 35445 9263 35479
rect 10609 35445 10643 35479
rect 11713 35445 11747 35479
rect 17417 35445 17451 35479
rect 19533 35445 19567 35479
rect 20177 35445 20211 35479
rect 2237 35241 2271 35275
rect 4445 35241 4479 35275
rect 10793 35241 10827 35275
rect 13093 35241 13127 35275
rect 16405 35241 16439 35275
rect 21005 35241 21039 35275
rect 1869 35173 1903 35207
rect 2421 35173 2455 35207
rect 15209 35173 15243 35207
rect 18705 35173 18739 35207
rect 4905 35105 4939 35139
rect 8401 35105 8435 35139
rect 8953 35105 8987 35139
rect 11713 35105 11747 35139
rect 14749 35105 14783 35139
rect 15602 35105 15636 35139
rect 17325 35105 17359 35139
rect 20361 35105 20395 35139
rect 3157 35037 3191 35071
rect 4261 35037 4295 35071
rect 9220 35037 9254 35071
rect 10977 35037 11011 35071
rect 14565 35037 14599 35071
rect 15485 35037 15519 35071
rect 15761 35037 15795 35071
rect 20913 35037 20947 35071
rect 21189 35037 21223 35071
rect 2237 34969 2271 35003
rect 5150 34969 5184 35003
rect 8134 34969 8168 35003
rect 11980 34969 12014 35003
rect 17592 34969 17626 35003
rect 2973 34901 3007 34935
rect 6285 34901 6319 34935
rect 7021 34901 7055 34935
rect 10333 34901 10367 34935
rect 19717 34901 19751 34935
rect 20085 34901 20119 34935
rect 20177 34901 20211 34935
rect 21373 34901 21407 34935
rect 1869 34697 1903 34731
rect 3525 34697 3559 34731
rect 4721 34697 4755 34731
rect 7573 34697 7607 34731
rect 11621 34697 11655 34731
rect 16129 34697 16163 34731
rect 16957 34697 16991 34731
rect 17325 34697 17359 34731
rect 17417 34697 17451 34731
rect 18245 34697 18279 34731
rect 18889 34697 18923 34731
rect 19073 34697 19107 34731
rect 2053 34629 2087 34663
rect 20269 34629 20303 34663
rect 2421 34561 2455 34595
rect 2881 34561 2915 34595
rect 3709 34561 3743 34595
rect 4077 34561 4111 34595
rect 4261 34561 4295 34595
rect 4905 34561 4939 34595
rect 5089 34561 5123 34595
rect 5273 34561 5307 34595
rect 5457 34561 5491 34595
rect 6377 34561 6411 34595
rect 7757 34561 7791 34595
rect 8125 34561 8159 34595
rect 8309 34561 8343 34595
rect 9229 34561 9263 34595
rect 10241 34561 10275 34595
rect 10425 34561 10459 34595
rect 10609 34561 10643 34595
rect 10793 34561 10827 34595
rect 11805 34561 11839 34595
rect 12357 34561 12391 34595
rect 12624 34561 12658 34595
rect 14473 34561 14507 34595
rect 15326 34561 15360 34595
rect 18153 34561 18187 34595
rect 18337 34561 18371 34595
rect 19070 34561 19104 34595
rect 20177 34561 20211 34595
rect 30113 34561 30147 34595
rect 3893 34493 3927 34527
rect 3985 34493 4019 34527
rect 5181 34493 5215 34527
rect 6837 34493 6871 34527
rect 7941 34493 7975 34527
rect 8033 34493 8067 34527
rect 8953 34493 8987 34527
rect 10517 34493 10551 34527
rect 14289 34493 14323 34527
rect 15209 34493 15243 34527
rect 15485 34493 15519 34527
rect 17601 34493 17635 34527
rect 19441 34493 19475 34527
rect 19533 34493 19567 34527
rect 29837 34493 29871 34527
rect 14933 34425 14967 34459
rect 2053 34357 2087 34391
rect 3065 34357 3099 34391
rect 6469 34357 6503 34391
rect 10977 34357 11011 34391
rect 13737 34357 13771 34391
rect 2237 34153 2271 34187
rect 6101 34153 6135 34187
rect 7573 34153 7607 34187
rect 1869 34085 1903 34119
rect 14105 34085 14139 34119
rect 15669 34085 15703 34119
rect 18613 34085 18647 34119
rect 20453 34085 20487 34119
rect 3801 34017 3835 34051
rect 9781 34017 9815 34051
rect 9873 34017 9907 34051
rect 10609 34017 10643 34051
rect 3157 33949 3191 33983
rect 6285 33949 6319 33983
rect 6929 33949 6963 33983
rect 7389 33949 7423 33983
rect 8217 33949 8251 33983
rect 9597 33949 9631 33983
rect 9965 33949 9999 33983
rect 10149 33949 10183 33983
rect 10876 33949 10910 33983
rect 12449 33949 12483 33983
rect 12542 33949 12576 33983
rect 12953 33949 12987 33983
rect 14243 33949 14277 33983
rect 14601 33949 14635 33983
rect 14749 33949 14783 33983
rect 15485 33949 15519 33983
rect 16129 33949 16163 33983
rect 17877 33949 17911 33983
rect 18061 33949 18095 33983
rect 18521 33949 18555 33983
rect 19993 33949 20027 33983
rect 20637 33949 20671 33983
rect 21741 33949 21775 33983
rect 2237 33881 2271 33915
rect 4046 33881 4080 33915
rect 12725 33881 12759 33915
rect 12817 33881 12851 33915
rect 14381 33881 14415 33915
rect 14473 33881 14507 33915
rect 17969 33881 18003 33915
rect 21005 33881 21039 33915
rect 2421 33813 2455 33847
rect 2973 33813 3007 33847
rect 5181 33813 5215 33847
rect 6837 33813 6871 33847
rect 8309 33813 8343 33847
rect 9413 33813 9447 33847
rect 11989 33813 12023 33847
rect 13093 33813 13127 33847
rect 16313 33813 16347 33847
rect 19901 33813 19935 33847
rect 20729 33813 20763 33847
rect 20821 33813 20855 33847
rect 21925 33813 21959 33847
rect 2973 33609 3007 33643
rect 3617 33609 3651 33643
rect 6377 33609 6411 33643
rect 14289 33609 14323 33643
rect 19533 33609 19567 33643
rect 19993 33609 20027 33643
rect 20729 33609 20763 33643
rect 15393 33541 15427 33575
rect 17325 33541 17359 33575
rect 18337 33541 18371 33575
rect 18521 33541 18555 33575
rect 1685 33473 1719 33507
rect 2329 33473 2363 33507
rect 3157 33473 3191 33507
rect 3801 33473 3835 33507
rect 4077 33473 4111 33507
rect 4169 33473 4203 33507
rect 4353 33473 4387 33507
rect 5549 33473 5583 33507
rect 6561 33473 6595 33507
rect 7757 33473 7791 33507
rect 8033 33473 8067 33507
rect 8125 33473 8159 33507
rect 8309 33473 8343 33507
rect 8769 33473 8803 33507
rect 9597 33473 9631 33507
rect 10333 33473 10367 33507
rect 11805 33473 11839 33507
rect 13176 33473 13210 33507
rect 15025 33473 15059 33507
rect 15118 33473 15152 33507
rect 15301 33473 15335 33507
rect 15490 33473 15524 33507
rect 17509 33473 17543 33507
rect 20637 33541 20671 33575
rect 20839 33541 20873 33575
rect 21005 33541 21039 33575
rect 21925 33541 21959 33575
rect 19625 33473 19659 33507
rect 19717 33473 19751 33507
rect 21833 33473 21867 33507
rect 22661 33473 22695 33507
rect 29837 33473 29871 33507
rect 3985 33405 4019 33439
rect 7941 33405 7975 33439
rect 10057 33405 10091 33439
rect 11529 33405 11563 33439
rect 12909 33405 12943 33439
rect 17141 33405 17175 33439
rect 18245 33405 18279 33439
rect 19533 33405 19567 33439
rect 5365 33337 5399 33371
rect 8953 33337 8987 33371
rect 20453 33337 20487 33371
rect 1501 33269 1535 33303
rect 2145 33269 2179 33303
rect 7573 33269 7607 33303
rect 9413 33269 9447 33303
rect 15669 33269 15703 33303
rect 18797 33269 18831 33303
rect 19809 33269 19843 33303
rect 22477 33269 22511 33303
rect 30021 33269 30055 33303
rect 2237 33065 2271 33099
rect 5733 33065 5767 33099
rect 10701 33065 10735 33099
rect 12081 33065 12115 33099
rect 19257 33065 19291 33099
rect 19809 33065 19843 33099
rect 21557 33065 21591 33099
rect 22201 33065 22235 33099
rect 1869 32997 1903 33031
rect 16405 32997 16439 33031
rect 7941 32929 7975 32963
rect 8033 32929 8067 32963
rect 9321 32929 9355 32963
rect 11621 32929 11655 32963
rect 15025 32929 15059 32963
rect 16957 32929 16991 32963
rect 19717 32929 19751 32963
rect 20913 32929 20947 32963
rect 2881 32861 2915 32895
rect 3801 32861 3835 32895
rect 7021 32861 7055 32895
rect 7665 32861 7699 32895
rect 7849 32861 7883 32895
rect 8217 32861 8251 32895
rect 9577 32861 9611 32895
rect 11529 32861 11563 32895
rect 11805 32861 11839 32895
rect 11897 32861 11931 32895
rect 12081 32861 12115 32895
rect 15292 32861 15326 32895
rect 19533 32861 19567 32895
rect 19625 32861 19659 32895
rect 19993 32861 20027 32895
rect 2237 32793 2271 32827
rect 4046 32793 4080 32827
rect 5825 32793 5859 32827
rect 17224 32793 17258 32827
rect 21189 32793 21223 32827
rect 22385 32793 22419 32827
rect 2421 32725 2455 32759
rect 3065 32725 3099 32759
rect 5181 32725 5215 32759
rect 6837 32725 6871 32759
rect 8401 32725 8435 32759
rect 18337 32725 18371 32759
rect 21097 32725 21131 32759
rect 22017 32725 22051 32759
rect 22185 32725 22219 32759
rect 3341 32521 3375 32555
rect 3801 32521 3835 32555
rect 8217 32521 8251 32555
rect 10057 32521 10091 32555
rect 15485 32521 15519 32555
rect 17877 32521 17911 32555
rect 19257 32521 19291 32555
rect 21991 32521 22025 32555
rect 7104 32453 7138 32487
rect 13706 32453 13740 32487
rect 19993 32453 20027 32487
rect 22201 32453 22235 32487
rect 1685 32385 1719 32419
rect 2421 32385 2455 32419
rect 3157 32385 3191 32419
rect 3985 32385 4019 32419
rect 4261 32385 4295 32419
rect 4353 32385 4387 32419
rect 4537 32385 4571 32419
rect 5365 32385 5399 32419
rect 8933 32385 8967 32419
rect 10885 32385 10919 32419
rect 11796 32385 11830 32419
rect 13461 32385 13495 32419
rect 15393 32385 15427 32419
rect 17141 32385 17175 32419
rect 17325 32385 17359 32419
rect 17693 32385 17727 32419
rect 18521 32385 18555 32419
rect 18705 32385 18739 32419
rect 18889 32385 18923 32419
rect 19073 32385 19107 32419
rect 20545 32385 20579 32419
rect 20913 32385 20947 32419
rect 21281 32385 21315 32419
rect 4169 32317 4203 32351
rect 5549 32317 5583 32351
rect 6837 32317 6871 32351
rect 8677 32317 8711 32351
rect 11529 32317 11563 32351
rect 17417 32317 17451 32351
rect 17509 32317 17543 32351
rect 18797 32317 18831 32351
rect 20637 32317 20671 32351
rect 21097 32317 21131 32351
rect 1501 32181 1535 32215
rect 2237 32181 2271 32215
rect 10609 32181 10643 32215
rect 12909 32181 12943 32215
rect 14841 32181 14875 32215
rect 21833 32181 21867 32215
rect 22017 32181 22051 32215
rect 2329 31977 2363 32011
rect 2973 31977 3007 32011
rect 6377 31977 6411 32011
rect 7021 31977 7055 32011
rect 9689 31977 9723 32011
rect 18521 31977 18555 32011
rect 20545 31977 20579 32011
rect 1961 31909 1995 31943
rect 2513 31909 2547 31943
rect 4077 31909 4111 31943
rect 7481 31909 7515 31943
rect 8125 31909 8159 31943
rect 10609 31909 10643 31943
rect 12633 31909 12667 31943
rect 13093 31909 13127 31943
rect 19625 31909 19659 31943
rect 5641 31841 5675 31875
rect 9505 31841 9539 31875
rect 18429 31841 18463 31875
rect 18613 31841 18647 31875
rect 20913 31841 20947 31875
rect 3157 31773 3191 31807
rect 5365 31773 5399 31807
rect 6193 31773 6227 31807
rect 6837 31773 6871 31807
rect 7665 31773 7699 31807
rect 8309 31773 8343 31807
rect 9965 31773 9999 31807
rect 10425 31773 10459 31807
rect 11253 31773 11287 31807
rect 13277 31773 13311 31807
rect 14105 31773 14139 31807
rect 18705 31773 18739 31807
rect 20637 31773 20671 31807
rect 20821 31773 20855 31807
rect 21006 31773 21040 31807
rect 21189 31773 21223 31807
rect 29837 31773 29871 31807
rect 4261 31705 4295 31739
rect 11520 31705 11554 31739
rect 14350 31705 14384 31739
rect 19809 31705 19843 31739
rect 2329 31637 2363 31671
rect 15485 31637 15519 31671
rect 30021 31637 30055 31671
rect 2513 31433 2547 31467
rect 8309 31433 8343 31467
rect 11805 31433 11839 31467
rect 13553 31433 13587 31467
rect 15393 31433 15427 31467
rect 17233 31433 17267 31467
rect 18705 31433 18739 31467
rect 19073 31433 19107 31467
rect 21925 31433 21959 31467
rect 2329 31365 2363 31399
rect 20085 31365 20119 31399
rect 1961 31297 1995 31331
rect 3617 31297 3651 31331
rect 3801 31297 3835 31331
rect 3985 31297 4019 31331
rect 4169 31297 4203 31331
rect 5089 31297 5123 31331
rect 6561 31297 6595 31331
rect 6745 31297 6779 31331
rect 6929 31297 6963 31331
rect 7113 31297 7147 31331
rect 7757 31297 7791 31331
rect 8401 31297 8435 31331
rect 9045 31297 9079 31331
rect 9505 31297 9539 31331
rect 10425 31297 10459 31331
rect 11984 31297 12018 31331
rect 12081 31297 12115 31331
rect 12173 31297 12207 31331
rect 12356 31297 12390 31331
rect 12449 31297 12483 31331
rect 12909 31297 12943 31331
rect 13002 31297 13036 31331
rect 13185 31297 13219 31331
rect 13277 31297 13311 31331
rect 13413 31297 13447 31331
rect 15761 31297 15795 31331
rect 17325 31297 17359 31331
rect 18613 31297 18647 31331
rect 20913 31297 20947 31331
rect 21833 31297 21867 31331
rect 3893 31229 3927 31263
rect 4813 31229 4847 31263
rect 6837 31229 6871 31263
rect 15853 31229 15887 31263
rect 16037 31229 16071 31263
rect 17141 31229 17175 31263
rect 18429 31229 18463 31263
rect 20269 31161 20303 31195
rect 2329 31093 2363 31127
rect 3433 31093 3467 31127
rect 6377 31093 6411 31127
rect 7573 31093 7607 31127
rect 8861 31093 8895 31127
rect 9597 31093 9631 31127
rect 9965 31093 9999 31127
rect 10517 31093 10551 31127
rect 10885 31093 10919 31127
rect 17693 31093 17727 31127
rect 20821 31093 20855 31127
rect 2329 30889 2363 30923
rect 8309 30889 8343 30923
rect 9137 30889 9171 30923
rect 11897 30889 11931 30923
rect 29929 30889 29963 30923
rect 1961 30821 1995 30855
rect 3985 30821 4019 30855
rect 21005 30821 21039 30855
rect 4905 30753 4939 30787
rect 5641 30753 5675 30787
rect 11529 30753 11563 30787
rect 13185 30753 13219 30787
rect 16865 30753 16899 30787
rect 17969 30753 18003 30787
rect 20269 30753 20303 30787
rect 20545 30753 20579 30787
rect 2973 30685 3007 30719
rect 3801 30685 3835 30719
rect 4629 30685 4663 30719
rect 4813 30685 4847 30719
rect 4997 30685 5031 30719
rect 5181 30685 5215 30719
rect 5908 30685 5942 30719
rect 8401 30685 8435 30719
rect 9413 30685 9447 30719
rect 10057 30685 10091 30719
rect 10701 30685 10735 30719
rect 11161 30685 11195 30719
rect 11345 30685 11379 30719
rect 11437 30685 11471 30719
rect 11713 30685 11747 30719
rect 12909 30685 12943 30719
rect 14289 30685 14323 30719
rect 16957 30685 16991 30719
rect 17877 30685 17911 30719
rect 18153 30685 18187 30719
rect 18245 30685 18279 30719
rect 29929 30685 29963 30719
rect 30113 30685 30147 30719
rect 2329 30617 2363 30651
rect 14556 30617 14590 30651
rect 21189 30617 21223 30651
rect 21373 30617 21407 30651
rect 2513 30549 2547 30583
rect 3157 30549 3191 30583
rect 4445 30549 4479 30583
rect 7021 30549 7055 30583
rect 7941 30549 7975 30583
rect 8953 30549 8987 30583
rect 9873 30549 9907 30583
rect 10517 30549 10551 30583
rect 15669 30549 15703 30583
rect 17049 30549 17083 30583
rect 17417 30549 17451 30583
rect 18429 30549 18463 30583
rect 2237 30345 2271 30379
rect 4261 30345 4295 30379
rect 4721 30345 4755 30379
rect 14749 30345 14783 30379
rect 18981 30345 19015 30379
rect 19809 30345 19843 30379
rect 3148 30277 3182 30311
rect 10977 30277 11011 30311
rect 12265 30277 12299 30311
rect 15301 30277 15335 30311
rect 15485 30277 15519 30311
rect 18899 30277 18933 30311
rect 19890 30277 19924 30311
rect 19993 30277 20027 30311
rect 1869 30209 1903 30243
rect 4905 30209 4939 30243
rect 5365 30209 5399 30243
rect 6561 30209 6595 30243
rect 6837 30209 6871 30243
rect 6929 30209 6963 30243
rect 7113 30209 7147 30243
rect 7941 30209 7975 30243
rect 8585 30209 8619 30243
rect 9137 30209 9171 30243
rect 10793 30209 10827 30243
rect 11529 30209 11563 30243
rect 11713 30209 11747 30243
rect 12081 30209 12115 30243
rect 13093 30209 13127 30243
rect 14105 30209 14139 30243
rect 14198 30209 14232 30243
rect 14381 30209 14415 30243
rect 14473 30209 14507 30243
rect 14611 30209 14645 30243
rect 15945 30209 15979 30243
rect 17049 30209 17083 30243
rect 17877 30209 17911 30243
rect 18797 30209 18831 30243
rect 19165 30209 19199 30243
rect 19625 30209 19659 30243
rect 20913 30209 20947 30243
rect 22937 30209 22971 30243
rect 29193 30209 29227 30243
rect 29837 30209 29871 30243
rect 2881 30141 2915 30175
rect 5457 30141 5491 30175
rect 6745 30141 6779 30175
rect 10517 30141 10551 30175
rect 11805 30141 11839 30175
rect 11897 30141 11931 30175
rect 12817 30141 12851 30175
rect 17141 30141 17175 30175
rect 17325 30141 17359 30175
rect 16037 30073 16071 30107
rect 18613 30073 18647 30107
rect 20177 30073 20211 30107
rect 29377 30073 29411 30107
rect 30021 30073 30055 30107
rect 2237 30005 2271 30039
rect 2421 30005 2455 30039
rect 6377 30005 6411 30039
rect 7757 30005 7791 30039
rect 8401 30005 8435 30039
rect 9321 30005 9355 30039
rect 10609 30005 10643 30039
rect 16681 30005 16715 30039
rect 18061 30005 18095 30039
rect 21005 30005 21039 30039
rect 22753 30005 22787 30039
rect 1501 29801 1535 29835
rect 2973 29801 3007 29835
rect 5089 29801 5123 29835
rect 11069 29801 11103 29835
rect 15577 29801 15611 29835
rect 19625 29801 19659 29835
rect 20177 29801 20211 29835
rect 2145 29733 2179 29767
rect 3801 29733 3835 29767
rect 11805 29733 11839 29767
rect 21925 29733 21959 29767
rect 12541 29665 12575 29699
rect 16865 29665 16899 29699
rect 18061 29665 18095 29699
rect 18245 29665 18279 29699
rect 19441 29665 19475 29699
rect 20177 29665 20211 29699
rect 20545 29665 20579 29699
rect 20637 29665 20671 29699
rect 22385 29665 22419 29699
rect 1685 29597 1719 29631
rect 2329 29597 2363 29631
rect 3157 29597 3191 29631
rect 3985 29597 4019 29631
rect 4629 29597 4663 29631
rect 6469 29597 6503 29631
rect 7849 29597 7883 29631
rect 9689 29597 9723 29631
rect 11621 29597 11655 29631
rect 12265 29597 12299 29631
rect 14197 29597 14231 29631
rect 16589 29597 16623 29631
rect 16773 29597 16807 29631
rect 16957 29597 16991 29631
rect 17141 29597 17175 29631
rect 18337 29597 18371 29631
rect 19349 29597 19383 29631
rect 19717 29597 19751 29631
rect 20361 29597 20395 29631
rect 20453 29597 20487 29631
rect 21741 29597 21775 29631
rect 22652 29597 22686 29631
rect 6224 29529 6258 29563
rect 7021 29529 7055 29563
rect 9934 29529 9968 29563
rect 14442 29529 14476 29563
rect 16405 29529 16439 29563
rect 21557 29529 21591 29563
rect 4445 29461 4479 29495
rect 7113 29461 7147 29495
rect 7665 29461 7699 29495
rect 18705 29461 18739 29495
rect 19349 29461 19383 29495
rect 20821 29461 20855 29495
rect 23765 29461 23799 29495
rect 2789 29257 2823 29291
rect 5181 29257 5215 29291
rect 5825 29257 5859 29291
rect 7297 29257 7331 29291
rect 8125 29257 8159 29291
rect 9505 29257 9539 29291
rect 10885 29257 10919 29291
rect 14013 29257 14047 29291
rect 16037 29257 16071 29291
rect 16681 29257 16715 29291
rect 17141 29257 17175 29291
rect 21005 29257 21039 29291
rect 23213 29257 23247 29291
rect 4068 29189 4102 29223
rect 9597 29189 9631 29223
rect 12633 29189 12667 29223
rect 13645 29189 13679 29223
rect 15025 29189 15059 29223
rect 1685 29121 1719 29155
rect 2145 29121 2179 29155
rect 2973 29121 3007 29155
rect 5641 29121 5675 29155
rect 8309 29121 8343 29155
rect 10977 29121 11011 29155
rect 13369 29121 13403 29155
rect 13462 29121 13496 29155
rect 13737 29121 13771 29155
rect 13834 29121 13868 29155
rect 15209 29121 15243 29155
rect 15393 29121 15427 29155
rect 15853 29121 15887 29155
rect 17049 29121 17083 29155
rect 18429 29121 18463 29155
rect 18521 29121 18555 29155
rect 18797 29121 18831 29155
rect 19441 29121 19475 29155
rect 19717 29121 19751 29155
rect 20913 29121 20947 29155
rect 3801 29053 3835 29087
rect 7389 29053 7423 29087
rect 7573 29053 7607 29087
rect 9689 29053 9723 29087
rect 17325 29053 17359 29087
rect 21833 29053 21867 29087
rect 22109 29053 22143 29087
rect 1501 28985 1535 29019
rect 2329 28985 2363 29019
rect 9137 28985 9171 29019
rect 12449 28985 12483 29019
rect 6929 28917 6963 28951
rect 18245 28917 18279 28951
rect 18705 28917 18739 28951
rect 2421 28713 2455 28747
rect 3801 28713 3835 28747
rect 4813 28713 4847 28747
rect 6193 28713 6227 28747
rect 11897 28713 11931 28747
rect 14197 28713 14231 28747
rect 15669 28713 15703 28747
rect 16865 28713 16899 28747
rect 22477 28713 22511 28747
rect 6653 28645 6687 28679
rect 18153 28645 18187 28679
rect 3157 28577 3191 28611
rect 7297 28577 7331 28611
rect 9505 28577 9539 28611
rect 11253 28577 11287 28611
rect 15025 28577 15059 28611
rect 20729 28577 20763 28611
rect 21833 28577 21867 28611
rect 22318 28577 22352 28611
rect 1685 28509 1719 28543
rect 2421 28509 2455 28543
rect 2605 28509 2639 28543
rect 3065 28509 3099 28543
rect 3249 28509 3283 28543
rect 3985 28509 4019 28543
rect 4629 28509 4663 28543
rect 6009 28509 6043 28543
rect 7021 28509 7055 28543
rect 8401 28509 8435 28543
rect 9321 28509 9355 28543
rect 10333 28509 10367 28543
rect 11069 28509 11103 28543
rect 11805 28509 11839 28543
rect 12771 28509 12805 28543
rect 13184 28509 13218 28543
rect 13277 28509 13311 28543
rect 14289 28509 14323 28543
rect 15577 28509 15611 28543
rect 16957 28509 16991 28543
rect 18061 28509 18095 28543
rect 18245 28509 18279 28543
rect 18337 28509 18371 28543
rect 18521 28509 18555 28543
rect 20177 28509 20211 28543
rect 20269 28509 20303 28543
rect 20453 28509 20487 28543
rect 20637 28509 20671 28543
rect 22109 28509 22143 28543
rect 29837 28509 29871 28543
rect 12909 28441 12943 28475
rect 13001 28441 13035 28475
rect 14841 28441 14875 28475
rect 20545 28441 20579 28475
rect 1501 28373 1535 28407
rect 7113 28373 7147 28407
rect 8309 28373 8343 28407
rect 8953 28373 8987 28407
rect 9413 28373 9447 28407
rect 10241 28373 10275 28407
rect 12633 28373 12667 28407
rect 17877 28373 17911 28407
rect 22201 28373 22235 28407
rect 30021 28373 30055 28407
rect 2145 28169 2179 28203
rect 6745 28169 6779 28203
rect 8493 28169 8527 28203
rect 14289 28169 14323 28203
rect 17049 28169 17083 28203
rect 18613 28169 18647 28203
rect 19073 28169 19107 28203
rect 20913 28169 20947 28203
rect 21925 28169 21959 28203
rect 30021 28169 30055 28203
rect 3709 28101 3743 28135
rect 12357 28101 12391 28135
rect 14749 28101 14783 28135
rect 1685 28033 1719 28067
rect 2329 28033 2363 28067
rect 2881 28033 2915 28067
rect 3617 28033 3651 28067
rect 3801 28033 3835 28067
rect 6561 28033 6595 28067
rect 7665 28033 7699 28067
rect 8677 28033 8711 28067
rect 8769 28033 8803 28067
rect 9045 28033 9079 28067
rect 9597 28033 9631 28067
rect 9864 28033 9898 28067
rect 11621 28033 11655 28067
rect 11713 28033 11747 28067
rect 12909 28033 12943 28067
rect 13176 28033 13210 28067
rect 14933 28033 14967 28067
rect 15485 28033 15519 28067
rect 16681 28033 16715 28067
rect 16865 28033 16899 28067
rect 17877 28033 17911 28067
rect 18061 28033 18095 28067
rect 18153 28033 18187 28067
rect 18429 28033 18463 28067
rect 19441 28033 19475 28067
rect 20269 28033 20303 28067
rect 20453 28033 20487 28067
rect 20729 28033 20763 28067
rect 21833 28033 21867 28067
rect 29929 28033 29963 28067
rect 30113 28033 30147 28067
rect 7205 27965 7239 27999
rect 18245 27965 18279 27999
rect 19533 27965 19567 27999
rect 19625 27965 19659 27999
rect 12173 27897 12207 27931
rect 20545 27897 20579 27931
rect 20637 27897 20671 27931
rect 1501 27829 1535 27863
rect 3065 27829 3099 27863
rect 7573 27829 7607 27863
rect 8953 27829 8987 27863
rect 10977 27829 11011 27863
rect 15577 27829 15611 27863
rect 16957 27625 16991 27659
rect 17969 27625 18003 27659
rect 19441 27625 19475 27659
rect 20453 27625 20487 27659
rect 4261 27557 4295 27591
rect 5825 27557 5859 27591
rect 6653 27557 6687 27591
rect 9689 27557 9723 27591
rect 10701 27557 10735 27591
rect 15485 27557 15519 27591
rect 20085 27557 20119 27591
rect 7665 27489 7699 27523
rect 9229 27489 9263 27523
rect 10609 27489 10643 27523
rect 11345 27489 11379 27523
rect 14841 27489 14875 27523
rect 15393 27489 15427 27523
rect 15577 27489 15611 27523
rect 16405 27489 16439 27523
rect 18521 27489 18555 27523
rect 19993 27489 20027 27523
rect 3065 27421 3099 27455
rect 3249 27421 3283 27455
rect 5641 27421 5675 27455
rect 5733 27421 5767 27455
rect 5917 27421 5951 27455
rect 6561 27421 6595 27455
rect 7389 27421 7423 27455
rect 7481 27421 7515 27455
rect 7757 27421 7791 27455
rect 8309 27421 8343 27455
rect 8401 27421 8435 27455
rect 8953 27421 8987 27455
rect 9141 27421 9175 27455
rect 9321 27421 9355 27455
rect 9505 27421 9539 27455
rect 10793 27421 10827 27455
rect 10885 27421 10919 27455
rect 14381 27421 14415 27455
rect 14473 27421 14507 27455
rect 14657 27421 14691 27455
rect 15301 27421 15335 27455
rect 16589 27421 16623 27455
rect 18337 27421 18371 27455
rect 19349 27421 19383 27455
rect 20269 27421 20303 27455
rect 21373 27421 21407 27455
rect 21649 27421 21683 27455
rect 29837 27421 29871 27455
rect 4445 27353 4479 27387
rect 6101 27353 6135 27387
rect 11590 27353 11624 27387
rect 3157 27285 3191 27319
rect 7205 27285 7239 27319
rect 12725 27285 12759 27319
rect 16497 27285 16531 27319
rect 18429 27285 18463 27319
rect 30021 27285 30055 27319
rect 6469 27081 6503 27115
rect 10977 27081 11011 27115
rect 16865 27081 16899 27115
rect 17233 27081 17267 27115
rect 18153 27081 18187 27115
rect 19533 27081 19567 27115
rect 29929 27081 29963 27115
rect 8401 27013 8435 27047
rect 11989 27013 12023 27047
rect 12173 27013 12207 27047
rect 1685 26945 1719 26979
rect 5558 26945 5592 26979
rect 6561 26945 6595 26979
rect 7113 26945 7147 26979
rect 7297 26945 7331 26979
rect 7665 26945 7699 26979
rect 8585 26945 8619 26979
rect 9137 26945 9171 26979
rect 9230 26945 9264 26979
rect 9413 26945 9447 26979
rect 9505 26945 9539 26979
rect 9602 26945 9636 26979
rect 10241 26945 10275 26979
rect 10425 26945 10459 26979
rect 10517 26945 10551 26979
rect 10793 26945 10827 26979
rect 12633 26945 12667 26979
rect 12889 26945 12923 26979
rect 14657 26945 14691 26979
rect 14933 26945 14967 26979
rect 15025 26945 15059 26979
rect 15209 26945 15243 26979
rect 15669 26945 15703 26979
rect 15853 26945 15887 26979
rect 18521 26945 18555 26979
rect 19717 26945 19751 26979
rect 19901 26945 19935 26979
rect 20821 26945 20855 26979
rect 22100 26945 22134 26979
rect 30113 26945 30147 26979
rect 5825 26877 5859 26911
rect 7389 26877 7423 26911
rect 7481 26877 7515 26911
rect 10609 26877 10643 26911
rect 14749 26877 14783 26911
rect 17325 26877 17359 26911
rect 17509 26877 17543 26911
rect 18613 26877 18647 26911
rect 18705 26877 18739 26911
rect 20729 26877 20763 26911
rect 21833 26877 21867 26911
rect 1501 26809 1535 26843
rect 4445 26741 4479 26775
rect 7849 26741 7883 26775
rect 9781 26741 9815 26775
rect 14013 26741 14047 26775
rect 16037 26741 16071 26775
rect 20453 26741 20487 26775
rect 20821 26741 20855 26775
rect 23213 26741 23247 26775
rect 7021 26537 7055 26571
rect 8309 26537 8343 26571
rect 9689 26537 9723 26571
rect 12633 26537 12667 26571
rect 14381 26537 14415 26571
rect 15117 26537 15151 26571
rect 16497 26537 16531 26571
rect 17785 26537 17819 26571
rect 19625 26537 19659 26571
rect 3801 26469 3835 26503
rect 5641 26469 5675 26503
rect 7481 26401 7515 26435
rect 7665 26401 7699 26435
rect 12173 26401 12207 26435
rect 14289 26401 14323 26435
rect 20821 26401 20855 26435
rect 20913 26401 20947 26435
rect 21741 26401 21775 26435
rect 1685 26333 1719 26367
rect 3065 26333 3099 26367
rect 3249 26333 3283 26367
rect 4925 26333 4959 26367
rect 5181 26333 5215 26367
rect 5779 26333 5813 26367
rect 6009 26333 6043 26367
rect 6137 26333 6171 26367
rect 6285 26333 6319 26367
rect 7389 26333 7423 26367
rect 8401 26333 8435 26367
rect 9045 26333 9079 26367
rect 9193 26333 9227 26367
rect 9321 26333 9355 26367
rect 9510 26333 9544 26367
rect 10333 26333 10367 26367
rect 11897 26333 11931 26367
rect 12081 26333 12115 26367
rect 12265 26333 12299 26367
rect 12449 26333 12483 26367
rect 14197 26333 14231 26367
rect 15025 26333 15059 26367
rect 15669 26333 15703 26367
rect 15853 26333 15887 26367
rect 16313 26333 16347 26367
rect 17417 26333 17451 26367
rect 18245 26333 18279 26367
rect 19533 26333 19567 26367
rect 19809 26333 19843 26367
rect 19901 26333 19935 26367
rect 20545 26333 20579 26367
rect 20729 26333 20763 26367
rect 21097 26333 21131 26367
rect 5917 26265 5951 26299
rect 9413 26265 9447 26299
rect 10241 26265 10275 26299
rect 17601 26265 17635 26299
rect 18337 26265 18371 26299
rect 21281 26265 21315 26299
rect 21986 26265 22020 26299
rect 1501 26197 1535 26231
rect 3157 26197 3191 26231
rect 14565 26197 14599 26231
rect 15761 26197 15795 26231
rect 19993 26197 20027 26231
rect 23121 26197 23155 26231
rect 3249 25993 3283 26027
rect 4537 25993 4571 26027
rect 10885 25993 10919 26027
rect 15669 25993 15703 26027
rect 17601 25993 17635 26027
rect 20085 25993 20119 26027
rect 21925 25993 21959 26027
rect 4905 25925 4939 25959
rect 5733 25925 5767 25959
rect 7573 25925 7607 25959
rect 7757 25925 7791 25959
rect 8677 25925 8711 25959
rect 13369 25925 13403 25959
rect 14841 25925 14875 25959
rect 19441 25925 19475 25959
rect 1685 25857 1719 25891
rect 3157 25857 3191 25891
rect 3341 25857 3375 25891
rect 4716 25857 4750 25891
rect 4813 25857 4847 25891
rect 5088 25857 5122 25891
rect 5181 25857 5215 25891
rect 5825 25857 5859 25891
rect 6469 25857 6503 25891
rect 6745 25857 6779 25891
rect 9505 25857 9539 25891
rect 9772 25857 9806 25891
rect 11989 25857 12023 25891
rect 12173 25857 12207 25891
rect 12265 25857 12299 25891
rect 12541 25857 12575 25891
rect 14749 25857 14783 25891
rect 15761 25857 15795 25891
rect 16957 25857 16991 25891
rect 17969 25857 18003 25891
rect 19901 25857 19935 25891
rect 20545 25857 20579 25891
rect 20729 25857 20763 25891
rect 20821 25857 20855 25891
rect 21097 25857 21131 25891
rect 22017 25857 22051 25891
rect 29837 25857 29871 25891
rect 8769 25789 8803 25823
rect 8861 25789 8895 25823
rect 12357 25789 12391 25823
rect 15577 25789 15611 25823
rect 18061 25789 18095 25823
rect 18153 25789 18187 25823
rect 19809 25789 19843 25823
rect 20913 25789 20947 25823
rect 21281 25789 21315 25823
rect 6561 25721 6595 25755
rect 6653 25721 6687 25755
rect 8309 25721 8343 25755
rect 13185 25721 13219 25755
rect 1501 25653 1535 25687
rect 6929 25653 6963 25687
rect 12725 25653 12759 25687
rect 16129 25653 16163 25687
rect 17049 25653 17083 25687
rect 19625 25653 19659 25687
rect 30021 25653 30055 25687
rect 6377 25449 6411 25483
rect 10333 25449 10367 25483
rect 14197 25449 14231 25483
rect 19717 25449 19751 25483
rect 20637 25449 20671 25483
rect 20913 25449 20947 25483
rect 6929 25381 6963 25415
rect 12633 25381 12667 25415
rect 15025 25381 15059 25415
rect 7481 25313 7515 25347
rect 9413 25313 9447 25347
rect 16865 25313 16899 25347
rect 19809 25313 19843 25347
rect 20545 25313 20579 25347
rect 6285 25245 6319 25279
rect 8125 25245 8159 25279
rect 8953 25245 8987 25279
rect 9137 25245 9171 25279
rect 9321 25245 9355 25279
rect 9505 25245 9539 25279
rect 9689 25245 9723 25279
rect 10425 25245 10459 25279
rect 11253 25245 11287 25279
rect 14105 25245 14139 25279
rect 15945 25245 15979 25279
rect 16957 25245 16991 25279
rect 19533 25245 19567 25279
rect 19625 25245 19659 25279
rect 20269 25245 20303 25279
rect 20729 25245 20763 25279
rect 21649 25245 21683 25279
rect 5733 25177 5767 25211
rect 7297 25177 7331 25211
rect 11520 25177 11554 25211
rect 14841 25177 14875 25211
rect 16129 25177 16163 25211
rect 17049 25177 17083 25211
rect 18613 25177 18647 25211
rect 21741 25177 21775 25211
rect 5641 25109 5675 25143
rect 7389 25109 7423 25143
rect 8217 25109 8251 25143
rect 15761 25109 15795 25143
rect 17417 25109 17451 25143
rect 18521 25109 18555 25143
rect 6929 24905 6963 24939
rect 9689 24905 9723 24939
rect 12265 24905 12299 24939
rect 12909 24905 12943 24939
rect 17693 24905 17727 24939
rect 19441 24905 19475 24939
rect 22201 24905 22235 24939
rect 9413 24837 9447 24871
rect 23029 24837 23063 24871
rect 23213 24837 23247 24871
rect 1685 24769 1719 24803
rect 3157 24769 3191 24803
rect 3341 24769 3375 24803
rect 5558 24769 5592 24803
rect 5825 24769 5859 24803
rect 7113 24769 7147 24803
rect 7389 24769 7423 24803
rect 7481 24769 7515 24803
rect 7665 24767 7699 24801
rect 8125 24769 8159 24803
rect 9045 24769 9079 24803
rect 9193 24769 9227 24803
rect 9321 24769 9355 24803
rect 9510 24769 9544 24803
rect 10425 24769 10459 24803
rect 10517 24769 10551 24803
rect 10701 24769 10735 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 12081 24769 12115 24803
rect 14022 24769 14056 24803
rect 14289 24769 14323 24803
rect 14749 24769 14783 24803
rect 15393 24769 15427 24803
rect 16681 24769 16715 24803
rect 18889 24769 18923 24803
rect 19533 24769 19567 24803
rect 19993 24769 20027 24803
rect 20913 24769 20947 24803
rect 21005 24769 21039 24803
rect 3249 24701 3283 24735
rect 7297 24701 7331 24735
rect 8217 24701 8251 24735
rect 10609 24701 10643 24735
rect 11805 24701 11839 24735
rect 11897 24701 11931 24735
rect 17417 24701 17451 24735
rect 17601 24701 17635 24735
rect 22293 24701 22327 24735
rect 22385 24701 22419 24735
rect 1501 24633 1535 24667
rect 10885 24633 10919 24667
rect 14841 24633 14875 24667
rect 4445 24565 4479 24599
rect 15485 24565 15519 24599
rect 16773 24565 16807 24599
rect 18061 24565 18095 24599
rect 18705 24565 18739 24599
rect 20085 24565 20119 24599
rect 21833 24565 21867 24599
rect 23397 24565 23431 24599
rect 5733 24361 5767 24395
rect 8217 24361 8251 24395
rect 9505 24361 9539 24395
rect 9965 24361 9999 24395
rect 13185 24361 13219 24395
rect 15485 24361 15519 24395
rect 19901 24361 19935 24395
rect 20085 24361 20119 24395
rect 11069 24293 11103 24327
rect 22845 24293 22879 24327
rect 6193 24225 6227 24259
rect 7481 24225 7515 24259
rect 9045 24225 9079 24259
rect 10425 24225 10459 24259
rect 12173 24225 12207 24259
rect 16313 24225 16347 24259
rect 17601 24225 17635 24259
rect 17785 24225 17819 24259
rect 20177 24225 20211 24259
rect 21097 24225 21131 24259
rect 1685 24157 1719 24191
rect 3065 24157 3099 24191
rect 3249 24157 3283 24191
rect 3801 24157 3835 24191
rect 5917 24157 5951 24191
rect 6101 24157 6135 24191
rect 6285 24157 6319 24191
rect 6469 24157 6503 24191
rect 7297 24157 7331 24191
rect 8309 24157 8343 24191
rect 8953 24157 8987 24191
rect 9229 24157 9263 24191
rect 9321 24157 9355 24191
rect 10149 24157 10183 24191
rect 10241 24157 10275 24191
rect 10517 24157 10551 24191
rect 11161 24157 11195 24191
rect 11897 24157 11931 24191
rect 12081 24157 12115 24191
rect 12265 24157 12299 24191
rect 12449 24157 12483 24191
rect 13093 24157 13127 24191
rect 14197 24157 14231 24191
rect 14381 24157 14415 24191
rect 14841 24157 14875 24191
rect 14934 24157 14968 24191
rect 15117 24157 15151 24191
rect 15209 24157 15243 24191
rect 15306 24157 15340 24191
rect 16037 24157 16071 24191
rect 16221 24157 16255 24191
rect 16405 24157 16439 24191
rect 16589 24157 16623 24191
rect 19257 24157 19291 24191
rect 20269 24157 20303 24191
rect 21005 24157 21039 24191
rect 21557 24157 21591 24191
rect 23029 24157 23063 24191
rect 23765 24157 23799 24191
rect 29837 24157 29871 24191
rect 3157 24089 3191 24123
rect 4068 24089 4102 24123
rect 17877 24089 17911 24123
rect 22017 24089 22051 24123
rect 22201 24089 22235 24123
rect 1501 24021 1535 24055
rect 5181 24021 5215 24055
rect 6929 24021 6963 24055
rect 7389 24021 7423 24055
rect 12633 24021 12667 24055
rect 14289 24021 14323 24055
rect 16773 24021 16807 24055
rect 18245 24021 18279 24055
rect 19349 24021 19383 24055
rect 21373 24021 21407 24055
rect 22385 24021 22419 24055
rect 23673 24021 23707 24055
rect 30021 24021 30055 24055
rect 3985 23817 4019 23851
rect 7849 23817 7883 23851
rect 14105 23817 14139 23851
rect 14933 23817 14967 23851
rect 16129 23817 16163 23851
rect 18613 23817 18647 23851
rect 29929 23817 29963 23851
rect 5549 23749 5583 23783
rect 7297 23749 7331 23783
rect 8217 23749 8251 23783
rect 8309 23749 8343 23783
rect 10793 23749 10827 23783
rect 12970 23749 13004 23783
rect 14565 23749 14599 23783
rect 15761 23749 15795 23783
rect 19625 23749 19659 23783
rect 4169 23681 4203 23715
rect 4537 23681 4571 23715
rect 4721 23681 4755 23715
rect 5733 23681 5767 23715
rect 6377 23681 6411 23715
rect 7849 23681 7883 23715
rect 8120 23681 8154 23715
rect 8492 23681 8526 23715
rect 8585 23681 8619 23715
rect 9045 23681 9079 23715
rect 9229 23681 9263 23715
rect 9597 23681 9631 23715
rect 11529 23681 11563 23715
rect 11713 23681 11747 23715
rect 11805 23681 11839 23715
rect 12081 23681 12115 23715
rect 12725 23681 12759 23715
rect 14749 23681 14783 23715
rect 16681 23681 16715 23715
rect 17141 23681 17175 23715
rect 17509 23681 17543 23715
rect 18521 23681 18555 23715
rect 19717 23681 19751 23715
rect 20407 23681 20441 23715
rect 20542 23681 20576 23715
rect 20637 23681 20671 23715
rect 20821 23681 20855 23715
rect 22201 23681 22235 23715
rect 23489 23681 23523 23715
rect 30113 23681 30147 23715
rect 1409 23613 1443 23647
rect 1685 23613 1719 23647
rect 4353 23613 4387 23647
rect 4445 23613 4479 23647
rect 9321 23613 9355 23647
rect 9413 23613 9447 23647
rect 11897 23613 11931 23647
rect 15485 23613 15519 23647
rect 15669 23613 15703 23647
rect 17233 23613 17267 23647
rect 17417 23613 17451 23647
rect 18705 23613 18739 23647
rect 22477 23613 22511 23647
rect 6469 23477 6503 23511
rect 7205 23477 7239 23511
rect 7941 23477 7975 23511
rect 9781 23477 9815 23511
rect 10885 23477 10919 23511
rect 12265 23477 12299 23511
rect 16773 23477 16807 23511
rect 18153 23477 18187 23511
rect 20177 23477 20211 23511
rect 23581 23477 23615 23511
rect 7205 23273 7239 23307
rect 9045 23273 9079 23307
rect 11161 23273 11195 23307
rect 13553 23273 13587 23307
rect 15761 23273 15795 23307
rect 17141 23273 17175 23307
rect 17877 23273 17911 23307
rect 19349 23273 19383 23307
rect 20637 23273 20671 23307
rect 6745 23205 6779 23239
rect 17601 23205 17635 23239
rect 21925 23205 21959 23239
rect 4537 23137 4571 23171
rect 4629 23137 4663 23171
rect 7665 23137 7699 23171
rect 16589 23137 16623 23171
rect 1409 23069 1443 23103
rect 4353 23069 4387 23103
rect 4721 23069 4755 23103
rect 4905 23069 4939 23103
rect 5365 23069 5399 23103
rect 7389 23069 7423 23103
rect 7573 23069 7607 23103
rect 7757 23069 7791 23103
rect 7941 23069 7975 23103
rect 8953 23069 8987 23103
rect 9781 23069 9815 23103
rect 10037 23069 10071 23103
rect 12173 23069 12207 23103
rect 14749 23069 14783 23103
rect 14841 23069 14875 23103
rect 15025 23069 15059 23103
rect 15669 23069 15703 23103
rect 16681 23069 16715 23103
rect 17601 23069 17635 23103
rect 17693 23069 17727 23103
rect 17877 23069 17911 23103
rect 18337 23069 18371 23103
rect 19257 23069 19291 23103
rect 19533 23069 19567 23103
rect 20361 23069 20395 23103
rect 20545 23069 20579 23103
rect 20729 23069 20763 23103
rect 22293 23069 22327 23103
rect 22937 23069 22971 23103
rect 23121 23069 23155 23103
rect 5632 23001 5666 23035
rect 12440 23001 12474 23035
rect 15209 23001 15243 23035
rect 19717 23001 19751 23035
rect 22109 23001 22143 23035
rect 22753 23001 22787 23035
rect 1593 22933 1627 22967
rect 4169 22933 4203 22967
rect 16773 22933 16807 22967
rect 18521 22933 18555 22967
rect 5457 22729 5491 22763
rect 6377 22729 6411 22763
rect 9137 22729 9171 22763
rect 9597 22729 9631 22763
rect 14841 22729 14875 22763
rect 16681 22729 16715 22763
rect 18705 22729 18739 22763
rect 20085 22729 20119 22763
rect 23121 22729 23155 22763
rect 4322 22661 4356 22695
rect 12970 22661 13004 22695
rect 17141 22661 17175 22695
rect 21005 22661 21039 22695
rect 1409 22593 1443 22627
rect 2053 22593 2087 22627
rect 2697 22593 2731 22627
rect 4077 22593 4111 22627
rect 6561 22593 6595 22627
rect 6929 22593 6963 22627
rect 7113 22593 7147 22627
rect 7757 22593 7791 22627
rect 8024 22593 8058 22627
rect 10710 22593 10744 22627
rect 10977 22593 11011 22627
rect 11529 22593 11563 22627
rect 11713 22593 11747 22627
rect 11805 22593 11839 22627
rect 12081 22593 12115 22627
rect 12725 22593 12759 22627
rect 14749 22593 14783 22627
rect 17049 22593 17083 22627
rect 18797 22593 18831 22627
rect 19993 22593 20027 22627
rect 21189 22593 21223 22627
rect 29837 22593 29871 22627
rect 6745 22525 6779 22559
rect 6837 22525 6871 22559
rect 11897 22525 11931 22559
rect 17233 22525 17267 22559
rect 18521 22525 18555 22559
rect 20177 22525 20211 22559
rect 24133 22525 24167 22559
rect 2237 22457 2271 22491
rect 20821 22457 20855 22491
rect 1593 22389 1627 22423
rect 2881 22389 2915 22423
rect 12265 22389 12299 22423
rect 14105 22389 14139 22423
rect 19165 22389 19199 22423
rect 19625 22389 19659 22423
rect 30021 22389 30055 22423
rect 10977 22185 11011 22219
rect 17141 22185 17175 22219
rect 16681 22117 16715 22151
rect 5273 22049 5307 22083
rect 6193 22049 6227 22083
rect 8953 22049 8987 22083
rect 9229 22049 9263 22083
rect 10609 22049 10643 22083
rect 11897 22049 11931 22083
rect 12357 22049 12391 22083
rect 15669 22049 15703 22083
rect 18153 22049 18187 22083
rect 18245 22049 18279 22083
rect 21189 22049 21223 22083
rect 22385 22049 22419 22083
rect 1869 21981 1903 22015
rect 5549 21981 5583 22015
rect 8125 21981 8159 22015
rect 10241 21981 10275 22015
rect 10425 21981 10459 22015
rect 10517 21981 10551 22015
rect 10793 21981 10827 22015
rect 11621 21981 11655 22015
rect 11805 21981 11839 22015
rect 11989 21981 12023 22015
rect 12173 21981 12207 22015
rect 15393 21981 15427 22015
rect 15766 21981 15800 22015
rect 16681 21981 16715 22015
rect 16865 21981 16899 22015
rect 16957 21981 16991 22015
rect 17233 21981 17267 22015
rect 19441 21981 19475 22015
rect 19625 21981 19659 22015
rect 21097 21981 21131 22015
rect 22293 21981 22327 22015
rect 2136 21913 2170 21947
rect 6460 21913 6494 21947
rect 8309 21913 8343 21947
rect 15577 21913 15611 21947
rect 15669 21913 15703 21947
rect 21005 21913 21039 21947
rect 22201 21913 22235 21947
rect 3249 21845 3283 21879
rect 7573 21845 7607 21879
rect 17693 21845 17727 21879
rect 18061 21845 18095 21879
rect 19257 21845 19291 21879
rect 20637 21845 20671 21879
rect 21833 21845 21867 21879
rect 4905 21641 4939 21675
rect 5733 21641 5767 21675
rect 13001 21641 13035 21675
rect 15485 21641 15519 21675
rect 15945 21641 15979 21675
rect 17417 21641 17451 21675
rect 19073 21641 19107 21675
rect 7941 21573 7975 21607
rect 10793 21573 10827 21607
rect 11888 21573 11922 21607
rect 20085 21573 20119 21607
rect 21833 21573 21867 21607
rect 22017 21573 22051 21607
rect 22201 21573 22235 21607
rect 1685 21505 1719 21539
rect 1952 21505 1986 21539
rect 3709 21505 3743 21539
rect 4997 21505 5031 21539
rect 5825 21505 5859 21539
rect 6929 21505 6963 21539
rect 7205 21505 7239 21539
rect 8125 21505 8159 21539
rect 8677 21505 8711 21539
rect 8953 21505 8987 21539
rect 10149 21505 10183 21539
rect 15577 21505 15611 21539
rect 16681 21505 16715 21539
rect 16865 21505 16899 21539
rect 17233 21505 17267 21539
rect 18245 21505 18279 21539
rect 19073 21505 19107 21539
rect 19257 21505 19291 21539
rect 19349 21505 19383 21539
rect 19625 21505 19659 21539
rect 20269 21505 20303 21539
rect 11621 21437 11655 21471
rect 15301 21437 15335 21471
rect 16957 21437 16991 21471
rect 17049 21437 17083 21471
rect 18337 21437 18371 21471
rect 18521 21437 18555 21471
rect 19533 21437 19567 21471
rect 3525 21369 3559 21403
rect 10977 21369 11011 21403
rect 17877 21369 17911 21403
rect 3065 21301 3099 21335
rect 10057 21301 10091 21335
rect 20453 21301 20487 21335
rect 2237 21097 2271 21131
rect 6745 21097 6779 21131
rect 8953 21097 8987 21131
rect 10425 21097 10459 21131
rect 11161 21097 11195 21131
rect 19257 21097 19291 21131
rect 19717 21097 19751 21131
rect 20545 21097 20579 21131
rect 8125 21029 8159 21063
rect 13185 21029 13219 21063
rect 17601 21029 17635 21063
rect 6285 20961 6319 20995
rect 6377 20961 6411 20995
rect 7389 20961 7423 20995
rect 15025 20961 15059 20995
rect 16497 20961 16531 20995
rect 18245 20961 18279 20995
rect 21005 20961 21039 20995
rect 21097 20961 21131 20995
rect 1501 20893 1535 20927
rect 1685 20893 1719 20927
rect 1777 20893 1811 20927
rect 1869 20893 1903 20927
rect 2053 20893 2087 20927
rect 3065 20893 3099 20927
rect 3801 20893 3835 20927
rect 4629 20893 4663 20927
rect 6009 20893 6043 20927
rect 6193 20893 6227 20927
rect 6561 20893 6595 20927
rect 7573 20893 7607 20927
rect 14105 20893 14139 20927
rect 15209 20893 15243 20927
rect 18061 20893 18095 20927
rect 19441 20893 19475 20927
rect 19533 20893 19567 20927
rect 19809 20893 19843 20927
rect 29837 20893 29871 20927
rect 3893 20825 3927 20859
rect 8309 20825 8343 20859
rect 9137 20825 9171 20859
rect 9321 20825 9355 20859
rect 10517 20825 10551 20859
rect 11253 20825 11287 20859
rect 13369 20825 13403 20859
rect 13553 20825 13587 20859
rect 14197 20825 14231 20859
rect 16681 20825 16715 20859
rect 17969 20825 18003 20859
rect 20913 20825 20947 20859
rect 3157 20757 3191 20791
rect 4445 20757 4479 20791
rect 15117 20757 15151 20791
rect 15577 20757 15611 20791
rect 16773 20757 16807 20791
rect 17141 20757 17175 20791
rect 30021 20757 30055 20791
rect 2421 20553 2455 20587
rect 8125 20553 8159 20587
rect 8953 20553 8987 20587
rect 15393 20553 15427 20587
rect 15485 20553 15519 20587
rect 16865 20553 16899 20587
rect 19533 20553 19567 20587
rect 22293 20553 22327 20587
rect 29929 20553 29963 20587
rect 8309 20485 8343 20519
rect 22201 20485 22235 20519
rect 1685 20417 1719 20451
rect 1869 20417 1903 20451
rect 2237 20417 2271 20451
rect 3065 20417 3099 20451
rect 3976 20417 4010 20451
rect 5549 20417 5583 20451
rect 6469 20417 6503 20451
rect 6562 20417 6596 20451
rect 6745 20417 6779 20451
rect 6837 20417 6871 20451
rect 6975 20417 7009 20451
rect 8493 20417 8527 20451
rect 9413 20417 9447 20451
rect 9873 20417 9907 20451
rect 9965 20417 9999 20451
rect 10609 20417 10643 20451
rect 11529 20417 11563 20451
rect 11713 20417 11747 20451
rect 11805 20417 11839 20451
rect 12081 20417 12115 20451
rect 13461 20417 13495 20451
rect 14105 20417 14139 20451
rect 14565 20417 14599 20451
rect 16681 20417 16715 20451
rect 18521 20417 18555 20451
rect 18705 20417 18739 20451
rect 20361 20417 20395 20451
rect 20545 20417 20579 20451
rect 20637 20417 20671 20451
rect 20913 20417 20947 20451
rect 30113 20417 30147 20451
rect 1961 20349 1995 20383
rect 2053 20349 2087 20383
rect 3709 20349 3743 20383
rect 11897 20349 11931 20383
rect 15577 20349 15611 20383
rect 19625 20349 19659 20383
rect 19717 20349 19751 20383
rect 22385 20349 22419 20383
rect 13553 20281 13587 20315
rect 14427 20281 14461 20315
rect 21833 20281 21867 20315
rect 2881 20213 2915 20247
rect 5089 20213 5123 20247
rect 5641 20213 5675 20247
rect 7113 20213 7147 20247
rect 9137 20213 9171 20247
rect 10701 20213 10735 20247
rect 12265 20213 12299 20247
rect 14197 20213 14231 20247
rect 14289 20213 14323 20247
rect 15025 20213 15059 20247
rect 18521 20213 18555 20247
rect 19165 20213 19199 20247
rect 20361 20213 20395 20247
rect 20821 20213 20855 20247
rect 4537 20009 4571 20043
rect 5641 20009 5675 20043
rect 9413 20009 9447 20043
rect 12909 20009 12943 20043
rect 13461 20009 13495 20043
rect 16681 20009 16715 20043
rect 20177 20009 20211 20043
rect 20637 20009 20671 20043
rect 7573 19941 7607 19975
rect 9873 19941 9907 19975
rect 10425 19941 10459 19975
rect 4169 19873 4203 19907
rect 6463 19873 6497 19907
rect 10609 19873 10643 19907
rect 11529 19873 11563 19907
rect 14473 19873 14507 19907
rect 15853 19873 15887 19907
rect 16037 19873 16071 19907
rect 17877 19873 17911 19907
rect 1777 19805 1811 19839
rect 3801 19805 3835 19839
rect 3985 19805 4019 19839
rect 4077 19805 4111 19839
rect 4353 19805 4387 19839
rect 5733 19805 5767 19839
rect 6193 19805 6227 19839
rect 6377 19805 6411 19839
rect 6561 19805 6595 19839
rect 6745 19805 6779 19839
rect 7757 19805 7791 19839
rect 9597 19805 9631 19839
rect 9689 19805 9723 19839
rect 9965 19805 9999 19839
rect 10701 19805 10735 19839
rect 10977 19805 11011 19839
rect 11796 19805 11830 19839
rect 13553 19805 13587 19839
rect 14105 19805 14139 19839
rect 14289 19805 14323 19839
rect 14381 19805 14415 19839
rect 14565 19805 14599 19839
rect 15761 19805 15795 19839
rect 15945 19805 15979 19839
rect 16773 19805 16807 19839
rect 17693 19805 17727 19839
rect 19441 19805 19475 19839
rect 20361 19805 20395 19839
rect 20453 19805 20487 19839
rect 20729 19805 20763 19839
rect 21189 19805 21223 19839
rect 21373 19805 21407 19839
rect 2044 19737 2078 19771
rect 7941 19737 7975 19771
rect 11069 19737 11103 19771
rect 19349 19737 19383 19771
rect 3157 19669 3191 19703
rect 6929 19669 6963 19703
rect 14749 19669 14783 19703
rect 15577 19669 15611 19703
rect 17325 19669 17359 19703
rect 17785 19669 17819 19703
rect 21281 19669 21315 19703
rect 8217 19465 8251 19499
rect 13185 19465 13219 19499
rect 14105 19465 14139 19499
rect 16681 19465 16715 19499
rect 17601 19465 17635 19499
rect 18797 19465 18831 19499
rect 19165 19465 19199 19499
rect 20729 19465 20763 19499
rect 30021 19465 30055 19499
rect 2237 19397 2271 19431
rect 11897 19397 11931 19431
rect 15218 19397 15252 19431
rect 18061 19397 18095 19431
rect 20637 19397 20671 19431
rect 1501 19329 1535 19363
rect 1685 19329 1719 19363
rect 1869 19329 1903 19363
rect 2053 19329 2087 19363
rect 3525 19329 3559 19363
rect 4261 19329 4295 19363
rect 4528 19329 4562 19363
rect 6837 19329 6871 19363
rect 7104 19329 7138 19363
rect 9229 19329 9263 19363
rect 10241 19329 10275 19363
rect 10425 19329 10459 19363
rect 15485 19329 15519 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 17969 19329 18003 19363
rect 19257 19329 19291 19363
rect 29837 19329 29871 19363
rect 1777 19261 1811 19295
rect 3801 19261 3835 19295
rect 8769 19261 8803 19295
rect 10057 19261 10091 19295
rect 18245 19261 18279 19295
rect 19349 19261 19383 19295
rect 20821 19261 20855 19295
rect 5641 19125 5675 19159
rect 8953 19125 8987 19159
rect 20269 19125 20303 19159
rect 4813 18921 4847 18955
rect 5917 18921 5951 18955
rect 18153 18921 18187 18955
rect 19257 18921 19291 18955
rect 21097 18921 21131 18955
rect 1869 18785 1903 18819
rect 4445 18785 4479 18819
rect 9229 18785 9263 18819
rect 15025 18785 15059 18819
rect 16681 18785 16715 18819
rect 19809 18785 19843 18819
rect 21649 18785 21683 18819
rect 4077 18717 4111 18751
rect 4261 18717 4295 18751
rect 4353 18717 4387 18751
rect 4629 18717 4663 18751
rect 5273 18717 5307 18751
rect 7297 18717 7331 18751
rect 8953 18717 8987 18751
rect 9137 18717 9171 18751
rect 9321 18717 9355 18751
rect 9505 18717 9539 18751
rect 10793 18717 10827 18751
rect 11253 18717 11287 18751
rect 12541 18717 12575 18751
rect 12725 18717 12759 18751
rect 14381 18717 14415 18751
rect 16221 18717 16255 18751
rect 18337 18717 18371 18751
rect 19625 18717 19659 18751
rect 20453 18717 20487 18751
rect 2136 18649 2170 18683
rect 7030 18649 7064 18683
rect 14105 18649 14139 18683
rect 15209 18649 15243 18683
rect 21465 18649 21499 18683
rect 3249 18581 3283 18615
rect 5365 18581 5399 18615
rect 9689 18581 9723 18615
rect 10609 18581 10643 18615
rect 11437 18581 11471 18615
rect 12633 18581 12667 18615
rect 15117 18581 15151 18615
rect 15577 18581 15611 18615
rect 19717 18581 19751 18615
rect 20637 18581 20671 18615
rect 21557 18581 21591 18615
rect 2513 18377 2547 18411
rect 10241 18377 10275 18411
rect 12909 18377 12943 18411
rect 15485 18377 15519 18411
rect 18981 18377 19015 18411
rect 19533 18377 19567 18411
rect 20913 18377 20947 18411
rect 21925 18377 21959 18411
rect 4721 18309 4755 18343
rect 13921 18309 13955 18343
rect 15393 18309 15427 18343
rect 1777 18241 1811 18275
rect 1961 18241 1995 18275
rect 2145 18241 2179 18275
rect 2329 18241 2363 18275
rect 3525 18241 3559 18275
rect 3709 18241 3743 18275
rect 4077 18241 4111 18275
rect 4905 18241 4939 18275
rect 5641 18241 5675 18275
rect 6377 18241 6411 18275
rect 7021 18241 7055 18275
rect 8953 18241 8987 18275
rect 9137 18241 9171 18275
rect 9229 18241 9263 18275
rect 9505 18241 9539 18275
rect 10333 18241 10367 18275
rect 11785 18241 11819 18275
rect 13645 18241 13679 18275
rect 17233 18241 17267 18275
rect 18337 18241 18371 18275
rect 19073 18241 19107 18275
rect 19718 18241 19752 18275
rect 19809 18241 19843 18275
rect 20085 18241 20119 18275
rect 20545 18241 20579 18275
rect 20729 18241 20763 18275
rect 22017 18241 22051 18275
rect 29837 18241 29871 18275
rect 2053 18173 2087 18207
rect 3801 18173 3835 18207
rect 3893 18173 3927 18207
rect 5457 18173 5491 18207
rect 9321 18173 9355 18207
rect 9689 18173 9723 18207
rect 11529 18173 11563 18207
rect 15577 18173 15611 18207
rect 17509 18173 17543 18207
rect 18061 18173 18095 18207
rect 13737 18105 13771 18139
rect 4261 18037 4295 18071
rect 6469 18037 6503 18071
rect 7113 18037 7147 18071
rect 13829 18037 13863 18071
rect 15025 18037 15059 18071
rect 19993 18037 20027 18071
rect 30021 18037 30055 18071
rect 2973 17833 3007 17867
rect 11161 17833 11195 17867
rect 13001 17833 13035 17867
rect 14749 17833 14783 17867
rect 15301 17833 15335 17867
rect 15393 17833 15427 17867
rect 16681 17833 16715 17867
rect 17141 17833 17175 17867
rect 19349 17833 19383 17867
rect 20269 17833 20303 17867
rect 29929 17833 29963 17867
rect 14473 17765 14507 17799
rect 18337 17765 18371 17799
rect 20177 17765 20211 17799
rect 2053 17697 2087 17731
rect 3801 17697 3835 17731
rect 6653 17697 6687 17731
rect 7941 17697 7975 17731
rect 9781 17697 9815 17731
rect 14289 17697 14323 17731
rect 14381 17697 14415 17731
rect 15485 17697 15519 17731
rect 16129 17697 16163 17731
rect 17325 17697 17359 17731
rect 17785 17697 17819 17731
rect 20361 17697 20395 17731
rect 1777 17629 1811 17663
rect 1961 17629 1995 17663
rect 2145 17629 2179 17663
rect 2329 17629 2363 17663
rect 2789 17629 2823 17663
rect 4077 17629 4111 17663
rect 5365 17629 5399 17663
rect 6377 17629 6411 17663
rect 7665 17629 7699 17663
rect 7849 17629 7883 17663
rect 8033 17629 8067 17663
rect 8217 17629 8251 17663
rect 10037 17629 10071 17663
rect 11621 17629 11655 17663
rect 14105 17629 14139 17663
rect 14565 17629 14599 17663
rect 15209 17629 15243 17663
rect 16221 17629 16255 17663
rect 16313 17629 16347 17663
rect 17417 17629 17451 17663
rect 18245 17629 18279 17663
rect 19441 17629 19475 17663
rect 20085 17629 20119 17663
rect 21005 17629 21039 17663
rect 30113 17629 30147 17663
rect 11866 17561 11900 17595
rect 20913 17561 20947 17595
rect 1593 17493 1627 17527
rect 5457 17493 5491 17527
rect 8401 17493 8435 17527
rect 8677 17289 8711 17323
rect 9873 17289 9907 17323
rect 15853 17289 15887 17323
rect 16773 17289 16807 17323
rect 17693 17289 17727 17323
rect 6837 17221 6871 17255
rect 7564 17221 7598 17255
rect 12256 17221 12290 17255
rect 17325 17221 17359 17255
rect 1676 17153 1710 17187
rect 3249 17153 3283 17187
rect 4077 17153 4111 17187
rect 4344 17153 4378 17187
rect 6653 17153 6687 17187
rect 9137 17153 9171 17187
rect 9321 17153 9355 17187
rect 9689 17153 9723 17187
rect 13829 17153 13863 17187
rect 14565 17153 14599 17187
rect 14749 17153 14783 17187
rect 15117 17153 15151 17187
rect 15945 17153 15979 17187
rect 16681 17153 16715 17187
rect 17509 17153 17543 17187
rect 19073 17153 19107 17187
rect 19533 17153 19567 17187
rect 19717 17153 19751 17187
rect 20085 17153 20119 17187
rect 1409 17085 1443 17119
rect 7297 17085 7331 17119
rect 9413 17085 9447 17119
rect 9505 17085 9539 17119
rect 11989 17085 12023 17119
rect 14841 17085 14875 17119
rect 14933 17085 14967 17119
rect 19809 17085 19843 17119
rect 19901 17085 19935 17119
rect 2789 17017 2823 17051
rect 3433 16949 3467 16983
rect 5457 16949 5491 16983
rect 13369 16949 13403 16983
rect 13921 16949 13955 16983
rect 15301 16949 15335 16983
rect 18981 16949 19015 16983
rect 20269 16949 20303 16983
rect 6285 16745 6319 16779
rect 18337 16745 18371 16779
rect 19257 16745 19291 16779
rect 13277 16677 13311 16711
rect 2145 16609 2179 16643
rect 4353 16609 4387 16643
rect 6837 16609 6871 16643
rect 9229 16609 9263 16643
rect 13185 16609 13219 16643
rect 13406 16609 13440 16643
rect 14841 16609 14875 16643
rect 16957 16609 16991 16643
rect 19625 16609 19659 16643
rect 1409 16541 1443 16575
rect 2421 16541 2455 16575
rect 4609 16541 4643 16575
rect 6193 16541 6227 16575
rect 8953 16541 8987 16575
rect 11989 16541 12023 16575
rect 12357 16541 12391 16575
rect 15117 16541 15151 16575
rect 16497 16541 16531 16575
rect 17233 16541 17267 16575
rect 19441 16541 19475 16575
rect 19714 16541 19748 16575
rect 19805 16541 19839 16575
rect 19993 16541 20027 16575
rect 20637 16541 20671 16575
rect 20893 16541 20927 16575
rect 29837 16541 29871 16575
rect 7104 16473 7138 16507
rect 12817 16473 12851 16507
rect 13553 16473 13587 16507
rect 1593 16405 1627 16439
rect 5733 16405 5767 16439
rect 8217 16405 8251 16439
rect 22017 16405 22051 16439
rect 30021 16405 30055 16439
rect 7205 16201 7239 16235
rect 13461 16201 13495 16235
rect 14473 16201 14507 16235
rect 17417 16201 17451 16235
rect 18521 16133 18555 16167
rect 20146 16133 20180 16167
rect 1409 16065 1443 16099
rect 2596 16065 2630 16099
rect 4445 16065 4479 16099
rect 5457 16065 5491 16099
rect 6561 16065 6595 16099
rect 7389 16065 7423 16099
rect 7757 16065 7791 16099
rect 7941 16065 7975 16099
rect 9045 16065 9079 16099
rect 10057 16065 10091 16099
rect 10241 16065 10275 16099
rect 10609 16065 10643 16099
rect 12357 16065 12391 16099
rect 12541 16065 12575 16099
rect 13645 16065 13679 16099
rect 13829 16065 13863 16099
rect 13921 16065 13955 16099
rect 14657 16065 14691 16099
rect 14841 16065 14875 16099
rect 16681 16065 16715 16099
rect 16865 16065 16899 16099
rect 17049 16065 17083 16099
rect 17233 16065 17267 16099
rect 18245 16065 18279 16099
rect 18383 16065 18417 16099
rect 18613 16065 18647 16099
rect 18751 16065 18785 16099
rect 2329 15997 2363 16031
rect 4169 15997 4203 16031
rect 7573 15997 7607 16031
rect 7671 15997 7705 16031
rect 8769 15997 8803 16031
rect 10333 15997 10367 16031
rect 10425 15997 10459 16031
rect 16957 15997 16991 16031
rect 19901 15997 19935 16031
rect 3709 15929 3743 15963
rect 13737 15929 13771 15963
rect 1593 15861 1627 15895
rect 5549 15861 5583 15895
rect 6653 15861 6687 15895
rect 10793 15861 10827 15895
rect 12357 15861 12391 15895
rect 18889 15861 18923 15895
rect 21281 15861 21315 15895
rect 4537 15657 4571 15691
rect 11437 15657 11471 15691
rect 13369 15657 13403 15691
rect 16129 15657 16163 15691
rect 17141 15657 17175 15691
rect 17693 15657 17727 15691
rect 21097 15657 21131 15691
rect 29929 15657 29963 15691
rect 20269 15589 20303 15623
rect 2421 15521 2455 15555
rect 2881 15521 2915 15555
rect 4077 15521 4111 15555
rect 14841 15521 14875 15555
rect 17785 15521 17819 15555
rect 1409 15453 1443 15487
rect 2145 15453 2179 15487
rect 2333 15453 2367 15487
rect 2513 15453 2547 15487
rect 2697 15453 2731 15487
rect 3801 15453 3835 15487
rect 3985 15453 4019 15487
rect 4169 15453 4203 15487
rect 4353 15453 4387 15487
rect 4997 15453 5031 15487
rect 5641 15453 5675 15487
rect 5825 15453 5859 15487
rect 5911 15453 5945 15487
rect 6009 15453 6043 15487
rect 6193 15453 6227 15487
rect 6837 15453 6871 15487
rect 7481 15453 7515 15487
rect 8125 15453 8159 15487
rect 8953 15453 8987 15487
rect 9101 15453 9135 15487
rect 9229 15453 9263 15487
rect 9418 15453 9452 15487
rect 10057 15453 10091 15487
rect 11989 15453 12023 15487
rect 12256 15453 12290 15487
rect 14473 15453 14507 15487
rect 14657 15453 14691 15487
rect 14749 15453 14783 15487
rect 15025 15453 15059 15487
rect 16221 15453 16255 15487
rect 17693 15453 17727 15487
rect 19625 15453 19659 15487
rect 19809 15453 19843 15487
rect 21281 15453 21315 15487
rect 22017 15453 22051 15487
rect 29929 15453 29963 15487
rect 30113 15453 30147 15487
rect 9321 15385 9355 15419
rect 10302 15385 10336 15419
rect 17049 15385 17083 15419
rect 20453 15385 20487 15419
rect 1593 15317 1627 15351
rect 5089 15317 5123 15351
rect 6377 15317 6411 15351
rect 6929 15317 6963 15351
rect 7573 15317 7607 15351
rect 8217 15317 8251 15351
rect 9597 15317 9631 15351
rect 15209 15317 15243 15351
rect 18061 15317 18095 15351
rect 19441 15317 19475 15351
rect 21833 15317 21867 15351
rect 5273 15113 5307 15147
rect 8861 15113 8895 15147
rect 14013 15113 14047 15147
rect 19073 15113 19107 15147
rect 29285 15113 29319 15147
rect 3433 15045 3467 15079
rect 4138 15045 4172 15079
rect 12081 15045 12115 15079
rect 14740 15045 14774 15079
rect 16865 15045 16899 15079
rect 17049 15045 17083 15079
rect 18061 15045 18095 15079
rect 18245 15045 18279 15079
rect 18981 15045 19015 15079
rect 21833 15045 21867 15079
rect 1409 14977 1443 15011
rect 2237 14977 2271 15011
rect 2697 14977 2731 15011
rect 2881 14977 2915 15011
rect 3249 14977 3283 15011
rect 6377 14977 6411 15011
rect 6561 14977 6595 15011
rect 6745 14977 6779 15011
rect 6929 14977 6963 15011
rect 8769 14977 8803 15011
rect 10710 14977 10744 15011
rect 10977 14977 11011 15011
rect 12541 14977 12575 15011
rect 12725 14977 12759 15011
rect 13553 14977 13587 15011
rect 13829 14977 13863 15011
rect 16681 14977 16715 15011
rect 20545 14977 20579 15011
rect 20637 14977 20671 15011
rect 22017 14977 22051 15011
rect 29193 14977 29227 15011
rect 29377 14977 29411 15011
rect 29837 14977 29871 15011
rect 2973 14909 3007 14943
rect 3065 14909 3099 14943
rect 3893 14909 3927 14943
rect 6653 14909 6687 14943
rect 12817 14909 12851 14943
rect 14473 14909 14507 14943
rect 20269 14909 20303 14943
rect 7113 14841 7147 14875
rect 17877 14841 17911 14875
rect 20821 14841 20855 14875
rect 1593 14773 1627 14807
rect 2053 14773 2087 14807
rect 9597 14773 9631 14807
rect 13645 14773 13679 14807
rect 15853 14773 15887 14807
rect 20361 14773 20395 14807
rect 22201 14773 22235 14807
rect 30021 14773 30055 14807
rect 2881 14569 2915 14603
rect 6469 14569 6503 14603
rect 7665 14569 7699 14603
rect 11989 14569 12023 14603
rect 14565 14569 14599 14603
rect 16129 14569 16163 14603
rect 22109 14569 22143 14603
rect 29009 14569 29043 14603
rect 10333 14501 10367 14535
rect 19809 14501 19843 14535
rect 20269 14501 20303 14535
rect 5181 14433 5215 14467
rect 7297 14433 7331 14467
rect 12725 14433 12759 14467
rect 16129 14433 16163 14467
rect 18153 14433 18187 14467
rect 30021 14433 30055 14467
rect 1501 14365 1535 14399
rect 5733 14365 5767 14399
rect 5917 14365 5951 14399
rect 6009 14365 6043 14399
rect 6101 14365 6135 14399
rect 6285 14365 6319 14399
rect 6929 14365 6963 14399
rect 7113 14365 7147 14399
rect 7205 14365 7239 14399
rect 7481 14365 7515 14399
rect 8953 14365 8987 14399
rect 11805 14365 11839 14399
rect 13369 14365 13403 14399
rect 13553 14365 13587 14399
rect 14657 14365 14691 14399
rect 15393 14365 15427 14399
rect 16037 14365 16071 14399
rect 16957 14365 16991 14399
rect 17141 14365 17175 14399
rect 17325 14365 17359 14399
rect 17509 14365 17543 14399
rect 18061 14365 18095 14399
rect 18337 14365 18371 14399
rect 18429 14365 18463 14399
rect 19717 14365 19751 14399
rect 19993 14365 20027 14399
rect 20085 14365 20119 14399
rect 20729 14365 20763 14399
rect 21005 14365 21039 14399
rect 22017 14365 22051 14399
rect 22293 14365 22327 14399
rect 22385 14365 22419 14399
rect 28825 14365 28859 14399
rect 29929 14365 29963 14399
rect 30113 14365 30147 14399
rect 1746 14297 1780 14331
rect 4914 14297 4948 14331
rect 8217 14297 8251 14331
rect 9198 14297 9232 14331
rect 12541 14297 12575 14331
rect 16313 14297 16347 14331
rect 22569 14297 22603 14331
rect 3801 14229 3835 14263
rect 8309 14229 8343 14263
rect 13185 14229 13219 14263
rect 15301 14229 15335 14263
rect 15853 14229 15887 14263
rect 17325 14229 17359 14263
rect 18613 14229 18647 14263
rect 1409 14025 1443 14059
rect 4629 14025 4663 14059
rect 7573 14025 7607 14059
rect 30021 14025 30055 14059
rect 8309 13957 8343 13991
rect 9137 13957 9171 13991
rect 14749 13957 14783 13991
rect 1593 13889 1627 13923
rect 1961 13889 1995 13923
rect 2145 13889 2179 13923
rect 3893 13889 3927 13923
rect 4077 13889 4111 13923
rect 4261 13889 4295 13923
rect 4445 13889 4479 13923
rect 5181 13889 5215 13923
rect 6837 13889 6871 13923
rect 7021 13889 7055 13923
rect 7113 13889 7147 13923
rect 7389 13889 7423 13923
rect 8033 13889 8067 13923
rect 8153 13889 8187 13923
rect 8401 13889 8435 13923
rect 8498 13889 8532 13923
rect 9321 13889 9355 13923
rect 9505 13889 9539 13923
rect 10241 13889 10275 13923
rect 12633 13889 12667 13923
rect 13369 13889 13403 13923
rect 13737 13889 13771 13923
rect 14565 13889 14599 13923
rect 15577 13889 15611 13923
rect 16773 13889 16807 13923
rect 16957 13889 16991 13923
rect 17509 13889 17543 13923
rect 19542 13889 19576 13923
rect 19809 13889 19843 13923
rect 20729 13889 20763 13923
rect 22293 13889 22327 13923
rect 29929 13889 29963 13923
rect 30113 13889 30147 13923
rect 1777 13821 1811 13855
rect 1869 13821 1903 13855
rect 2605 13821 2639 13855
rect 2881 13821 2915 13855
rect 4169 13821 4203 13855
rect 5273 13821 5307 13855
rect 7205 13821 7239 13855
rect 12449 13821 12483 13855
rect 14381 13821 14415 13855
rect 20453 13821 20487 13855
rect 22569 13821 22603 13855
rect 8677 13753 8711 13787
rect 16681 13753 16715 13787
rect 18429 13753 18463 13787
rect 10425 13685 10459 13719
rect 15301 13685 15335 13719
rect 4261 13481 4295 13515
rect 4997 13481 5031 13515
rect 6561 13481 6595 13515
rect 12081 13481 12115 13515
rect 16221 13481 16255 13515
rect 17417 13481 17451 13515
rect 19349 13481 19383 13515
rect 1869 13413 1903 13447
rect 11621 13413 11655 13447
rect 6193 13345 6227 13379
rect 8401 13345 8435 13379
rect 12449 13345 12483 13379
rect 16313 13345 16347 13379
rect 17601 13345 17635 13379
rect 20361 13345 20395 13379
rect 1961 13277 1995 13311
rect 2421 13277 2455 13311
rect 2697 13277 2731 13311
rect 4905 13277 4939 13311
rect 5825 13277 5859 13311
rect 6009 13277 6043 13311
rect 6104 13277 6138 13311
rect 6377 13277 6411 13311
rect 8125 13277 8159 13311
rect 10241 13277 10275 13311
rect 12265 13277 12299 13311
rect 13461 13277 13495 13311
rect 13553 13277 13587 13311
rect 15393 13277 15427 13311
rect 16221 13277 16255 13311
rect 17417 13277 17451 13311
rect 17509 13277 17543 13311
rect 17785 13277 17819 13311
rect 17877 13277 17911 13311
rect 19533 13277 19567 13311
rect 20269 13277 20303 13311
rect 20545 13277 20579 13311
rect 20637 13277 20671 13311
rect 20821 13277 20855 13311
rect 29837 13277 29871 13311
rect 4353 13209 4387 13243
rect 9413 13209 9447 13243
rect 10508 13209 10542 13243
rect 14473 13209 14507 13243
rect 15025 13209 15059 13243
rect 15209 13209 15243 13243
rect 18061 13209 18095 13243
rect 9505 13141 9539 13175
rect 14381 13141 14415 13175
rect 16589 13141 16623 13175
rect 30021 13141 30055 13175
rect 2881 12937 2915 12971
rect 4629 12937 4663 12971
rect 9137 12937 9171 12971
rect 11621 12937 11655 12971
rect 12817 12937 12851 12971
rect 18061 12937 18095 12971
rect 30021 12937 30055 12971
rect 5457 12869 5491 12903
rect 8769 12869 8803 12903
rect 8969 12869 9003 12903
rect 13461 12869 13495 12903
rect 14749 12869 14783 12903
rect 15669 12869 15703 12903
rect 17233 12869 17267 12903
rect 19165 12869 19199 12903
rect 1757 12801 1791 12835
rect 3341 12801 3375 12835
rect 3525 12801 3559 12835
rect 3893 12801 3927 12835
rect 4721 12801 4755 12835
rect 5273 12801 5307 12835
rect 5549 12801 5583 12835
rect 5677 12801 5711 12835
rect 7297 12801 7331 12835
rect 7573 12801 7607 12835
rect 8125 12801 8159 12835
rect 10057 12801 10091 12835
rect 10793 12801 10827 12835
rect 11529 12801 11563 12835
rect 11713 12801 11747 12835
rect 12633 12801 12667 12835
rect 13645 12801 13679 12835
rect 15393 12801 15427 12835
rect 16681 12801 16715 12835
rect 16957 12801 16991 12835
rect 17049 12801 17083 12835
rect 17693 12801 17727 12835
rect 18521 12801 18555 12835
rect 18613 12801 18647 12835
rect 19349 12801 19383 12835
rect 19993 12801 20027 12835
rect 20269 12801 20303 12835
rect 20361 12801 20395 12835
rect 29929 12801 29963 12835
rect 30113 12801 30147 12835
rect 1501 12733 1535 12767
rect 3617 12733 3651 12767
rect 3709 12733 3743 12767
rect 17785 12733 17819 12767
rect 20085 12733 20119 12767
rect 8309 12665 8343 12699
rect 9689 12665 9723 12699
rect 10977 12665 11011 12699
rect 20545 12665 20579 12699
rect 4077 12597 4111 12631
rect 5273 12597 5307 12631
rect 8953 12597 8987 12631
rect 14841 12597 14875 12631
rect 16773 12597 16807 12631
rect 17693 12597 17727 12631
rect 19533 12597 19567 12631
rect 1593 12393 1627 12427
rect 6653 12393 6687 12427
rect 17877 12393 17911 12427
rect 1961 12257 1995 12291
rect 6285 12257 6319 12291
rect 7389 12257 7423 12291
rect 7481 12257 7515 12291
rect 13277 12257 13311 12291
rect 14105 12257 14139 12291
rect 18521 12257 18555 12291
rect 1777 12189 1811 12223
rect 2053 12189 2087 12223
rect 2145 12189 2179 12223
rect 2329 12189 2363 12223
rect 2789 12189 2823 12223
rect 3801 12189 3835 12223
rect 5917 12189 5951 12223
rect 6101 12189 6135 12223
rect 6193 12189 6227 12223
rect 6469 12189 6503 12223
rect 7113 12189 7147 12223
rect 7297 12189 7331 12223
rect 7665 12189 7699 12223
rect 9413 12189 9447 12223
rect 9597 12189 9631 12223
rect 10333 12189 10367 12223
rect 10977 12189 11011 12223
rect 12817 12189 12851 12223
rect 13001 12189 13035 12223
rect 13185 12189 13219 12223
rect 13369 12189 13403 12223
rect 13553 12189 13587 12223
rect 15945 12189 15979 12223
rect 16221 12189 16255 12223
rect 18002 12189 18036 12223
rect 18429 12189 18463 12223
rect 20545 12189 20579 12223
rect 29929 12189 29963 12223
rect 30113 12189 30147 12223
rect 4068 12121 4102 12155
rect 9229 12121 9263 12155
rect 11244 12121 11278 12155
rect 14372 12121 14406 12155
rect 19257 12121 19291 12155
rect 19441 12121 19475 12155
rect 20085 12121 20119 12155
rect 2973 12053 3007 12087
rect 5181 12053 5215 12087
rect 7849 12053 7883 12087
rect 10149 12053 10183 12087
rect 12357 12053 12391 12087
rect 15485 12053 15519 12087
rect 18061 12053 18095 12087
rect 19625 12053 19659 12087
rect 30021 12053 30055 12087
rect 4997 11849 5031 11883
rect 10977 11849 11011 11883
rect 13829 11849 13863 11883
rect 15669 11849 15703 11883
rect 17877 11849 17911 11883
rect 18337 11849 18371 11883
rect 18521 11849 18555 11883
rect 20545 11849 20579 11883
rect 21189 11849 21223 11883
rect 12716 11781 12750 11815
rect 1409 11713 1443 11747
rect 2421 11713 2455 11747
rect 2605 11713 2639 11747
rect 2973 11713 3007 11747
rect 3617 11713 3651 11747
rect 3873 11713 3907 11747
rect 5641 11713 5675 11747
rect 6377 11713 6411 11747
rect 7021 11713 7055 11747
rect 7205 11713 7239 11747
rect 7389 11713 7423 11747
rect 7573 11713 7607 11747
rect 8217 11713 8251 11747
rect 8484 11713 8518 11747
rect 10241 11713 10275 11747
rect 10425 11713 10459 11747
rect 10609 11713 10643 11747
rect 10793 11713 10827 11747
rect 14289 11713 14323 11747
rect 14545 11713 14579 11747
rect 17141 11713 17175 11747
rect 17325 11713 17359 11747
rect 17509 11713 17543 11747
rect 17693 11713 17727 11747
rect 18462 11713 18496 11747
rect 18889 11713 18923 11747
rect 19809 11713 19843 11747
rect 19993 11713 20027 11747
rect 20177 11713 20211 11747
rect 20361 11713 20395 11747
rect 21189 11713 21223 11747
rect 29193 11713 29227 11747
rect 29837 11713 29871 11747
rect 2697 11645 2731 11679
rect 2789 11645 2823 11679
rect 3157 11645 3191 11679
rect 7297 11645 7331 11679
rect 10517 11645 10551 11679
rect 12449 11645 12483 11679
rect 17417 11645 17451 11679
rect 18981 11645 19015 11679
rect 20085 11645 20119 11679
rect 1593 11577 1627 11611
rect 5825 11577 5859 11611
rect 29377 11577 29411 11611
rect 6469 11509 6503 11543
rect 7757 11509 7791 11543
rect 9597 11509 9631 11543
rect 30021 11509 30055 11543
rect 6929 11305 6963 11339
rect 9413 11305 9447 11339
rect 13553 11305 13587 11339
rect 14841 11305 14875 11339
rect 16405 11305 16439 11339
rect 18613 11305 18647 11339
rect 20545 11305 20579 11339
rect 21097 11237 21131 11271
rect 5365 11169 5399 11203
rect 8769 11169 8803 11203
rect 11161 11169 11195 11203
rect 11253 11169 11287 11203
rect 12357 11169 12391 11203
rect 13093 11169 13127 11203
rect 14381 11169 14415 11203
rect 16865 11169 16899 11203
rect 17785 11169 17819 11203
rect 20177 11169 20211 11203
rect 1409 11101 1443 11135
rect 5181 11101 5215 11135
rect 5457 11101 5491 11135
rect 5585 11101 5619 11135
rect 8042 11101 8076 11135
rect 8309 11101 8343 11135
rect 5365 11033 5399 11067
rect 8953 11101 8987 11135
rect 9321 11101 9355 11135
rect 9505 11101 9539 11135
rect 10885 11101 10919 11135
rect 11069 11101 11103 11135
rect 11420 11101 11454 11135
rect 12817 11101 12851 11135
rect 13001 11101 13035 11135
rect 13185 11101 13219 11135
rect 13369 11101 13403 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 14473 11101 14507 11135
rect 14668 11101 14702 11135
rect 15669 11101 15703 11135
rect 15853 11101 15887 11135
rect 15945 11101 15979 11135
rect 16037 11101 16071 11135
rect 16221 11101 16255 11135
rect 17269 11095 17303 11129
rect 17969 11101 18003 11135
rect 18521 11101 18555 11135
rect 19809 11101 19843 11135
rect 19993 11101 20027 11135
rect 20085 11101 20119 11135
rect 20361 11101 20395 11135
rect 21189 11101 21223 11135
rect 10149 11033 10183 11067
rect 12173 11033 12207 11067
rect 16865 11033 16899 11067
rect 17049 11033 17083 11067
rect 17141 11033 17175 11067
rect 1593 10965 1627 10999
rect 8769 10965 8803 10999
rect 9137 10965 9171 10999
rect 10241 10965 10275 10999
rect 11621 10965 11655 10999
rect 2881 10761 2915 10795
rect 6837 10761 6871 10795
rect 15117 10761 15151 10795
rect 17509 10761 17543 10795
rect 18061 10761 18095 10795
rect 20453 10761 20487 10795
rect 21005 10761 21039 10795
rect 5089 10693 5123 10727
rect 5365 10693 5399 10727
rect 7389 10693 7423 10727
rect 8585 10693 8619 10727
rect 11713 10693 11747 10727
rect 14289 10693 14323 10727
rect 1501 10625 1535 10659
rect 1768 10625 1802 10659
rect 5273 10625 5307 10659
rect 5462 10625 5496 10659
rect 6929 10625 6963 10659
rect 7573 10625 7607 10659
rect 8401 10625 8435 10659
rect 9137 10625 9171 10659
rect 9229 10625 9263 10659
rect 9413 10625 9447 10659
rect 10149 10625 10183 10659
rect 10333 10625 10367 10659
rect 10701 10625 10735 10659
rect 12357 10625 12391 10659
rect 12633 10625 12667 10659
rect 14197 10625 14231 10659
rect 15209 10625 15243 10659
rect 15669 10625 15703 10659
rect 15853 10625 15887 10659
rect 15945 10625 15979 10659
rect 16073 10625 16107 10659
rect 16773 10625 16807 10659
rect 16957 10625 16991 10659
rect 17049 10625 17083 10659
rect 17325 10625 17359 10659
rect 17969 10625 18003 10659
rect 18797 10625 18831 10659
rect 19717 10625 19751 10659
rect 19901 10625 19935 10659
rect 20085 10625 20119 10659
rect 20269 10625 20303 10659
rect 21097 10625 21131 10659
rect 5089 10489 5123 10523
rect 9597 10557 9631 10591
rect 10425 10557 10459 10591
rect 10517 10557 10551 10591
rect 15761 10557 15795 10591
rect 17141 10557 17175 10591
rect 19257 10557 19291 10591
rect 19993 10557 20027 10591
rect 11897 10489 11931 10523
rect 9137 10421 9171 10455
rect 10885 10421 10919 10455
rect 19073 10421 19107 10455
rect 2237 10217 2271 10251
rect 9321 10217 9355 10251
rect 11621 10217 11655 10251
rect 13461 10217 13495 10251
rect 17509 10217 17543 10251
rect 20361 10217 20395 10251
rect 18521 10149 18555 10183
rect 1777 10081 1811 10115
rect 3801 10081 3835 10115
rect 6285 10081 6319 10115
rect 10241 10081 10275 10115
rect 14473 10081 14507 10115
rect 16681 10081 16715 10115
rect 1501 10013 1535 10047
rect 1685 10013 1719 10047
rect 1869 10013 1903 10047
rect 2053 10013 2087 10047
rect 2697 10013 2731 10047
rect 6193 10013 6227 10047
rect 6382 9991 6416 10025
rect 7113 10013 7147 10047
rect 7849 10013 7883 10047
rect 10508 10013 10542 10047
rect 12081 10013 12115 10047
rect 12337 10013 12371 10047
rect 14105 10013 14139 10047
rect 14289 10013 14323 10047
rect 14381 10013 14415 10047
rect 14657 10013 14691 10047
rect 16589 10013 16623 10047
rect 16793 10013 16827 10047
rect 17417 10013 17451 10047
rect 18337 10013 18371 10047
rect 18613 10013 18647 10047
rect 20453 10013 20487 10047
rect 22477 10013 22511 10047
rect 29837 10013 29871 10047
rect 4046 9945 4080 9979
rect 6009 9945 6043 9979
rect 6285 9945 6319 9979
rect 6929 9945 6963 9979
rect 7665 9945 7699 9979
rect 9505 9945 9539 9979
rect 9689 9945 9723 9979
rect 15393 9945 15427 9979
rect 15577 9945 15611 9979
rect 16405 9945 16439 9979
rect 16681 9945 16715 9979
rect 22232 9945 22266 9979
rect 2881 9877 2915 9911
rect 5181 9877 5215 9911
rect 14841 9877 14875 9911
rect 18153 9877 18187 9911
rect 21097 9877 21131 9911
rect 30021 9877 30055 9911
rect 3341 9673 3375 9707
rect 19257 9673 19291 9707
rect 19809 9673 19843 9707
rect 6929 9605 6963 9639
rect 10701 9605 10735 9639
rect 10885 9605 10919 9639
rect 14044 9605 14078 9639
rect 1409 9537 1443 9571
rect 2605 9537 2639 9571
rect 2789 9537 2823 9571
rect 3157 9537 3191 9571
rect 4077 9537 4111 9571
rect 4261 9537 4295 9571
rect 4445 9537 4479 9571
rect 4629 9537 4663 9571
rect 5457 9537 5491 9571
rect 6556 9559 6590 9593
rect 6653 9537 6687 9571
rect 6745 9537 6779 9571
rect 9965 9537 9999 9571
rect 14922 9537 14956 9571
rect 15117 9537 15151 9571
rect 15301 9537 15335 9571
rect 15485 9537 15519 9571
rect 15937 9537 15971 9571
rect 18144 9537 18178 9571
rect 19717 9537 19751 9571
rect 22089 9537 22123 9571
rect 2881 9469 2915 9503
rect 2973 9469 3007 9503
rect 4353 9469 4387 9503
rect 5273 9469 5307 9503
rect 8309 9469 8343 9503
rect 8585 9469 8619 9503
rect 12173 9469 12207 9503
rect 12449 9469 12483 9503
rect 14289 9469 14323 9503
rect 15209 9469 15243 9503
rect 16037 9469 16071 9503
rect 17877 9469 17911 9503
rect 21833 9469 21867 9503
rect 6929 9401 6963 9435
rect 1593 9333 1627 9367
rect 4813 9333 4847 9367
rect 12909 9333 12943 9367
rect 14749 9333 14783 9367
rect 23213 9333 23247 9367
rect 5181 9129 5215 9163
rect 6837 9129 6871 9163
rect 9689 9129 9723 9163
rect 10241 9129 10275 9163
rect 19073 9129 19107 9163
rect 19625 9129 19659 9163
rect 20269 9129 20303 9163
rect 21925 9129 21959 9163
rect 16129 9061 16163 9095
rect 2697 8993 2731 9027
rect 9229 8993 9263 9027
rect 12725 8993 12759 9027
rect 21465 8993 21499 9027
rect 1409 8925 1443 8959
rect 2329 8925 2363 8959
rect 2513 8925 2547 8959
rect 2605 8925 2639 8959
rect 2881 8925 2915 8959
rect 3801 8925 3835 8959
rect 8217 8925 8251 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9321 8925 9355 8959
rect 9505 8925 9539 8959
rect 10149 8925 10183 8959
rect 10977 8925 11011 8959
rect 11437 8925 11471 8959
rect 11621 8925 11655 8959
rect 13001 8925 13035 8959
rect 14289 8925 14323 8959
rect 16313 8925 16347 8959
rect 16957 8925 16991 8959
rect 17877 8925 17911 8959
rect 18061 8925 18095 8959
rect 18147 8925 18181 8959
rect 18245 8925 18279 8959
rect 18429 8925 18463 8959
rect 19073 8925 19107 8959
rect 19533 8925 19567 8959
rect 20177 8925 20211 8959
rect 21189 8925 21223 8959
rect 21373 8925 21407 8959
rect 21557 8925 21591 8959
rect 21741 8925 21775 8959
rect 4057 8857 4091 8891
rect 5825 8857 5859 8891
rect 7950 8857 7984 8891
rect 14534 8857 14568 8891
rect 1593 8789 1627 8823
rect 3065 8789 3099 8823
rect 5733 8789 5767 8823
rect 10885 8789 10919 8823
rect 11529 8789 11563 8823
rect 15669 8789 15703 8823
rect 17049 8789 17083 8823
rect 18613 8789 18647 8823
rect 2789 8585 2823 8619
rect 5733 8585 5767 8619
rect 10241 8585 10275 8619
rect 10609 8585 10643 8619
rect 14105 8585 14139 8619
rect 19901 8585 19935 8619
rect 22569 8585 22603 8619
rect 3617 8517 3651 8551
rect 7205 8517 7239 8551
rect 7849 8517 7883 8551
rect 11989 8517 12023 8551
rect 1409 8449 1443 8483
rect 1676 8449 1710 8483
rect 3801 8449 3835 8483
rect 4353 8449 4387 8483
rect 4620 8449 4654 8483
rect 6469 8449 6503 8483
rect 6653 8449 6687 8483
rect 7021 8449 7055 8483
rect 8401 8449 8435 8483
rect 8677 8449 8711 8483
rect 11897 8449 11931 8483
rect 13369 8449 13403 8483
rect 13553 8449 13587 8483
rect 13921 8449 13955 8483
rect 14832 8449 14866 8483
rect 16681 8449 16715 8483
rect 16937 8449 16971 8483
rect 18521 8449 18555 8483
rect 18797 8449 18831 8483
rect 21833 8449 21867 8483
rect 22017 8449 22051 8483
rect 22385 8449 22419 8483
rect 29837 8449 29871 8483
rect 6745 8381 6779 8415
rect 6837 8381 6871 8415
rect 10701 8381 10735 8415
rect 10885 8381 10919 8415
rect 12081 8381 12115 8415
rect 13645 8381 13679 8415
rect 13737 8381 13771 8415
rect 14565 8381 14599 8415
rect 22109 8381 22143 8415
rect 22201 8381 22235 8415
rect 7665 8313 7699 8347
rect 11529 8313 11563 8347
rect 15945 8313 15979 8347
rect 30021 8313 30055 8347
rect 18061 8245 18095 8279
rect 2651 8041 2685 8075
rect 9045 8041 9079 8075
rect 9413 8041 9447 8075
rect 10333 8041 10367 8075
rect 10793 8041 10827 8075
rect 12541 8041 12575 8075
rect 16405 8041 16439 8075
rect 21097 8041 21131 8075
rect 8401 7973 8435 8007
rect 9873 7973 9907 8007
rect 2421 7905 2455 7939
rect 9321 7905 9355 7939
rect 10241 7905 10275 7939
rect 11989 7905 12023 7939
rect 15945 7905 15979 7939
rect 21833 7905 21867 7939
rect 1409 7837 1443 7871
rect 3985 7837 4019 7871
rect 4261 7837 4295 7871
rect 5733 7837 5767 7871
rect 6009 7837 6043 7871
rect 9413 7837 9447 7871
rect 10057 7837 10091 7871
rect 10977 7837 11011 7871
rect 13001 7837 13035 7871
rect 13093 7837 13127 7871
rect 13277 7837 13311 7871
rect 15669 7837 15703 7871
rect 15853 7837 15887 7871
rect 16037 7837 16071 7871
rect 16221 7837 16255 7871
rect 17049 7837 17083 7871
rect 17693 7837 17727 7871
rect 17969 7837 18003 7871
rect 19717 7837 19751 7871
rect 21557 7837 21591 7871
rect 21741 7837 21775 7871
rect 21925 7837 21959 7871
rect 22109 7837 22143 7871
rect 7113 7769 7147 7803
rect 7297 7769 7331 7803
rect 8217 7769 8251 7803
rect 10333 7769 10367 7803
rect 11161 7769 11195 7803
rect 12081 7769 12115 7803
rect 17233 7769 17267 7803
rect 19984 7769 20018 7803
rect 1593 7701 1627 7735
rect 12173 7701 12207 7735
rect 13461 7701 13495 7735
rect 22293 7701 22327 7735
rect 2237 7497 2271 7531
rect 10149 7497 10183 7531
rect 11621 7497 11655 7531
rect 13461 7497 13495 7531
rect 13829 7497 13863 7531
rect 23213 7497 23247 7531
rect 5549 7429 5583 7463
rect 5733 7429 5767 7463
rect 14381 7429 14415 7463
rect 22100 7429 22134 7463
rect 1501 7361 1535 7395
rect 1685 7361 1719 7395
rect 1777 7361 1811 7395
rect 2053 7361 2087 7395
rect 3525 7361 3559 7395
rect 3801 7361 3835 7395
rect 4537 7361 4571 7395
rect 6745 7361 6779 7395
rect 6929 7361 6963 7395
rect 7297 7361 7331 7395
rect 8493 7361 8527 7395
rect 8677 7361 8711 7395
rect 8769 7361 8803 7395
rect 9045 7361 9079 7395
rect 10333 7361 10367 7395
rect 10609 7361 10643 7395
rect 11529 7361 11563 7395
rect 11713 7361 11747 7395
rect 12173 7361 12207 7395
rect 12449 7361 12483 7395
rect 14289 7361 14323 7395
rect 14473 7361 14507 7395
rect 15301 7361 15335 7395
rect 15485 7361 15519 7395
rect 15577 7361 15611 7395
rect 15853 7361 15887 7395
rect 17969 7361 18003 7395
rect 18613 7361 18647 7395
rect 20913 7361 20947 7395
rect 29837 7361 29871 7395
rect 1869 7293 1903 7327
rect 4261 7293 4295 7327
rect 7021 7293 7055 7327
rect 7113 7293 7147 7327
rect 8861 7293 8895 7327
rect 10517 7293 10551 7327
rect 12265 7293 12299 7327
rect 13185 7293 13219 7327
rect 13369 7293 13403 7327
rect 15669 7293 15703 7327
rect 17693 7293 17727 7327
rect 19441 7293 19475 7327
rect 19717 7293 19751 7327
rect 21833 7293 21867 7327
rect 7481 7157 7515 7191
rect 9229 7157 9263 7191
rect 10517 7157 10551 7191
rect 12633 7157 12667 7191
rect 16037 7157 16071 7191
rect 18521 7157 18555 7191
rect 20821 7157 20855 7191
rect 30021 7157 30055 7191
rect 7021 6953 7055 6987
rect 10333 6953 10367 6987
rect 20085 6953 20119 6987
rect 29929 6953 29963 6987
rect 18153 6885 18187 6919
rect 2053 6817 2087 6851
rect 4077 6817 4111 6851
rect 4169 6817 4203 6851
rect 5181 6817 5215 6851
rect 6101 6817 6135 6851
rect 12265 6817 12299 6851
rect 14841 6817 14875 6851
rect 16957 6817 16991 6851
rect 19625 6817 19659 6851
rect 20545 6817 20579 6851
rect 1685 6749 1719 6783
rect 1869 6749 1903 6783
rect 1961 6749 1995 6783
rect 2237 6749 2271 6783
rect 3801 6749 3835 6783
rect 3985 6749 4019 6783
rect 4353 6749 4387 6783
rect 5273 6749 5307 6783
rect 5825 6749 5859 6783
rect 5917 6749 5951 6783
rect 6193 6749 6227 6783
rect 6469 6749 6503 6783
rect 8134 6749 8168 6783
rect 8401 6749 8435 6783
rect 8953 6749 8987 6783
rect 9220 6749 9254 6783
rect 12541 6749 12575 6783
rect 14565 6749 14599 6783
rect 16037 6749 16071 6783
rect 16589 6749 16623 6783
rect 16773 6749 16807 6783
rect 16865 6749 16899 6783
rect 17141 6749 17175 6783
rect 19349 6749 19383 6783
rect 19533 6749 19567 6783
rect 19717 6749 19751 6783
rect 19901 6749 19935 6783
rect 29929 6749 29963 6783
rect 30113 6749 30147 6783
rect 3157 6681 3191 6715
rect 10977 6681 11011 6715
rect 17969 6681 18003 6715
rect 20812 6681 20846 6715
rect 2421 6613 2455 6647
rect 3065 6613 3099 6647
rect 4537 6613 4571 6647
rect 10885 6613 10919 6647
rect 12449 6613 12483 6647
rect 12909 6613 12943 6647
rect 15853 6613 15887 6647
rect 17325 6613 17359 6647
rect 21925 6613 21959 6647
rect 2973 6409 3007 6443
rect 5365 6409 5399 6443
rect 11897 6409 11931 6443
rect 15761 6409 15795 6443
rect 16681 6409 16715 6443
rect 18521 6409 18555 6443
rect 21097 6409 21131 6443
rect 4252 6341 4286 6375
rect 6561 6341 6595 6375
rect 6791 6341 6825 6375
rect 8585 6341 8619 6375
rect 1593 6273 1627 6307
rect 1860 6273 1894 6307
rect 3985 6273 4019 6307
rect 6464 6273 6498 6307
rect 6653 6273 6687 6307
rect 7353 6273 7387 6307
rect 7481 6273 7515 6307
rect 7573 6273 7607 6307
rect 7757 6273 7791 6307
rect 10057 6273 10091 6307
rect 10333 6273 10367 6307
rect 12081 6273 12115 6307
rect 12357 6273 12391 6307
rect 14381 6273 14415 6307
rect 14648 6273 14682 6307
rect 17794 6273 17828 6307
rect 18061 6273 18095 6307
rect 19634 6273 19668 6307
rect 19901 6273 19935 6307
rect 20361 6273 20395 6307
rect 20545 6273 20579 6307
rect 20637 6273 20671 6307
rect 20913 6273 20947 6307
rect 13645 6205 13679 6239
rect 13921 6205 13955 6239
rect 20729 6205 20763 6239
rect 7757 6137 7791 6171
rect 6837 6069 6871 6103
rect 8677 6069 8711 6103
rect 12265 6069 12299 6103
rect 3249 5865 3283 5899
rect 5549 5865 5583 5899
rect 13185 5865 13219 5899
rect 13553 5865 13587 5899
rect 15025 5865 15059 5899
rect 17049 5865 17083 5899
rect 18245 5865 18279 5899
rect 20637 5865 20671 5899
rect 29837 5865 29871 5899
rect 11989 5797 12023 5831
rect 1869 5729 1903 5763
rect 4169 5729 4203 5763
rect 6561 5729 6595 5763
rect 12633 5729 12667 5763
rect 14105 5729 14139 5763
rect 15669 5729 15703 5763
rect 17877 5729 17911 5763
rect 19257 5729 19291 5763
rect 6285 5661 6319 5695
rect 6469 5661 6503 5695
rect 6653 5661 6687 5695
rect 6837 5661 6871 5695
rect 13369 5661 13403 5695
rect 13553 5661 13587 5695
rect 14197 5661 14231 5695
rect 14381 5661 14415 5695
rect 15209 5661 15243 5695
rect 15925 5661 15959 5695
rect 17509 5661 17543 5695
rect 17693 5661 17727 5695
rect 17785 5661 17819 5695
rect 18061 5661 18095 5695
rect 19533 5661 19567 5695
rect 20729 5661 20763 5695
rect 29837 5661 29871 5695
rect 2136 5593 2170 5627
rect 4436 5593 4470 5627
rect 10241 5593 10275 5627
rect 10609 5593 10643 5627
rect 10977 5593 11011 5627
rect 11069 5593 11103 5627
rect 12449 5593 12483 5627
rect 7021 5525 7055 5559
rect 10057 5525 10091 5559
rect 11345 5525 11379 5559
rect 12357 5525 12391 5559
rect 14565 5525 14599 5559
rect 2697 5321 2731 5355
rect 4721 5321 4755 5355
rect 6653 5321 6687 5355
rect 11621 5321 11655 5355
rect 13001 5321 13035 5355
rect 13369 5321 13403 5355
rect 15117 5321 15151 5355
rect 19901 5321 19935 5355
rect 30021 5321 30055 5355
rect 3893 5253 3927 5287
rect 7766 5253 7800 5287
rect 21036 5253 21070 5287
rect 2881 5185 2915 5219
rect 3157 5185 3191 5219
rect 3249 5185 3283 5219
rect 3433 5185 3467 5219
rect 1409 5117 1443 5151
rect 1685 5117 1719 5151
rect 3065 5117 3099 5151
rect 3985 5185 4019 5219
rect 4169 5185 4203 5219
rect 4261 5185 4295 5219
rect 4537 5185 4571 5219
rect 5365 5185 5399 5219
rect 8749 5185 8783 5219
rect 10793 5185 10827 5219
rect 11805 5185 11839 5219
rect 11989 5185 12023 5219
rect 14381 5185 14415 5219
rect 15301 5185 15335 5219
rect 15485 5185 15519 5219
rect 15669 5185 15703 5219
rect 15853 5185 15887 5219
rect 17325 5185 17359 5219
rect 18337 5185 18371 5219
rect 21281 5185 21315 5219
rect 29837 5185 29871 5219
rect 4353 5117 4387 5151
rect 8033 5117 8067 5151
rect 8493 5117 8527 5151
rect 12081 5117 12115 5151
rect 13461 5117 13495 5151
rect 13553 5117 13587 5151
rect 15577 5117 15611 5151
rect 17601 5117 17635 5151
rect 18061 5117 18095 5151
rect 3893 5049 3927 5083
rect 5181 5049 5215 5083
rect 10977 5049 11011 5083
rect 14197 5049 14231 5083
rect 17509 5049 17543 5083
rect 18153 5049 18187 5083
rect 9873 4981 9907 5015
rect 17141 4981 17175 5015
rect 18521 4981 18555 5015
rect 2881 4777 2915 4811
rect 8401 4777 8435 4811
rect 11345 4777 11379 4811
rect 15117 4777 15151 4811
rect 14657 4709 14691 4743
rect 17233 4709 17267 4743
rect 1409 4641 1443 4675
rect 1685 4641 1719 4675
rect 5549 4641 5583 4675
rect 6745 4641 6779 4675
rect 7941 4641 7975 4675
rect 13277 4641 13311 4675
rect 15761 4641 15795 4675
rect 18245 4641 18279 4675
rect 19625 4641 19659 4675
rect 2697 4573 2731 4607
rect 5365 4573 5399 4607
rect 5641 4573 5675 4607
rect 5733 4573 5767 4607
rect 5917 4573 5951 4607
rect 6377 4573 6411 4607
rect 6561 4573 6595 4607
rect 6653 4573 6687 4607
rect 6929 4573 6963 4607
rect 7665 4573 7699 4607
rect 7849 4573 7883 4607
rect 8033 4573 8067 4607
rect 8217 4573 8251 4607
rect 8953 4573 8987 4607
rect 9137 4573 9171 4607
rect 9229 4573 9263 4607
rect 9321 4573 9355 4607
rect 9505 4573 9539 4607
rect 10701 4573 10735 4607
rect 13553 4573 13587 4607
rect 14473 4573 14507 4607
rect 16497 4573 16531 4607
rect 16681 4573 16715 4607
rect 16773 4573 16807 4607
rect 17417 4573 17451 4607
rect 17969 4573 18003 4607
rect 18157 4573 18191 4607
rect 18337 4573 18371 4607
rect 18521 4573 18555 4607
rect 30113 4573 30147 4607
rect 11529 4505 11563 4539
rect 11713 4505 11747 4539
rect 15485 4505 15519 4539
rect 19892 4505 19926 4539
rect 5181 4437 5215 4471
rect 7113 4437 7147 4471
rect 9689 4437 9723 4471
rect 10793 4437 10827 4471
rect 15577 4437 15611 4471
rect 16313 4437 16347 4471
rect 18705 4437 18739 4471
rect 21005 4437 21039 4471
rect 29929 4437 29963 4471
rect 7757 4233 7791 4267
rect 12449 4233 12483 4267
rect 13185 4233 13219 4267
rect 15025 4233 15059 4267
rect 16681 4233 16715 4267
rect 19809 4233 19843 4267
rect 21005 4233 21039 4267
rect 1869 4165 1903 4199
rect 2237 4165 2271 4199
rect 15393 4165 15427 4199
rect 17049 4165 17083 4199
rect 18696 4165 18730 4199
rect 2697 4097 2731 4131
rect 3433 4097 3467 4131
rect 4261 4097 4295 4131
rect 4445 4097 4479 4131
rect 4813 4097 4847 4131
rect 6377 4097 6411 4131
rect 6644 4097 6678 4131
rect 8861 4097 8895 4131
rect 9045 4097 9079 4131
rect 9137 4097 9171 4131
rect 9229 4097 9263 4131
rect 9413 4097 9447 4131
rect 10149 4097 10183 4131
rect 10793 4097 10827 4131
rect 12081 4097 12115 4131
rect 13185 4097 13219 4131
rect 14565 4097 14599 4131
rect 15485 4097 15519 4131
rect 17141 4097 17175 4131
rect 20269 4097 20303 4131
rect 20453 4097 20487 4131
rect 20821 4097 20855 4131
rect 28549 4097 28583 4131
rect 29193 4097 29227 4131
rect 29837 4097 29871 4131
rect 4537 4029 4571 4063
rect 4629 4029 4663 4063
rect 10885 4029 10919 4063
rect 12173 4029 12207 4063
rect 12909 4029 12943 4063
rect 14289 4029 14323 4063
rect 15669 4029 15703 4063
rect 17233 4029 17267 4063
rect 18429 4029 18463 4063
rect 20545 4029 20579 4063
rect 20637 4029 20671 4063
rect 2881 3961 2915 3995
rect 3617 3961 3651 3995
rect 13093 3961 13127 3995
rect 4997 3893 5031 3927
rect 9597 3893 9631 3927
rect 10241 3893 10275 3927
rect 12081 3893 12115 3927
rect 28733 3893 28767 3927
rect 29377 3893 29411 3927
rect 30021 3893 30055 3927
rect 2145 3689 2179 3723
rect 3985 3689 4019 3723
rect 10885 3689 10919 3723
rect 11621 3689 11655 3723
rect 15669 3689 15703 3723
rect 16865 3689 16899 3723
rect 18153 3689 18187 3723
rect 18521 3689 18555 3723
rect 20177 3689 20211 3723
rect 20821 3689 20855 3723
rect 22293 3689 22327 3723
rect 22937 3689 22971 3723
rect 3065 3621 3099 3655
rect 13093 3621 13127 3655
rect 11713 3553 11747 3587
rect 14105 3553 14139 3587
rect 16221 3553 16255 3587
rect 17325 3553 17359 3587
rect 17417 3553 17451 3587
rect 18061 3553 18095 3587
rect 19717 3553 19751 3587
rect 19809 3553 19843 3587
rect 1869 3485 1903 3519
rect 3801 3485 3835 3519
rect 5089 3485 5123 3519
rect 9505 3485 9539 3519
rect 9772 3485 9806 3519
rect 11805 3485 11839 3519
rect 12265 3485 12299 3519
rect 12725 3485 12759 3519
rect 13093 3485 13127 3519
rect 14381 3485 14415 3519
rect 16037 3485 16071 3519
rect 17233 3485 17267 3519
rect 18337 3485 18371 3519
rect 19441 3485 19475 3519
rect 19625 3485 19659 3519
rect 19993 3485 20027 3519
rect 20913 3485 20947 3519
rect 21005 3485 21039 3519
rect 22477 3485 22511 3519
rect 23121 3485 23155 3519
rect 28089 3485 28123 3519
rect 28825 3485 28859 3519
rect 29745 3485 29779 3519
rect 2789 3417 2823 3451
rect 5334 3417 5368 3451
rect 16129 3417 16163 3451
rect 21465 3417 21499 3451
rect 21649 3417 21683 3451
rect 21833 3417 21867 3451
rect 6469 3349 6503 3383
rect 11437 3349 11471 3383
rect 20637 3349 20671 3383
rect 27905 3349 27939 3383
rect 28641 3349 28675 3383
rect 29561 3349 29595 3383
rect 5365 3145 5399 3179
rect 7481 3145 7515 3179
rect 10793 3145 10827 3179
rect 11529 3145 11563 3179
rect 13829 3145 13863 3179
rect 17601 3145 17635 3179
rect 19165 3145 19199 3179
rect 19257 3145 19291 3179
rect 21833 3145 21867 3179
rect 22937 3145 22971 3179
rect 23581 3145 23615 3179
rect 27261 3145 27295 3179
rect 29377 3145 29411 3179
rect 1869 3077 1903 3111
rect 12725 3077 12759 3111
rect 14289 3077 14323 3111
rect 15485 3077 15519 3111
rect 16681 3077 16715 3111
rect 27721 3077 27755 3111
rect 28181 3077 28215 3111
rect 28365 3077 28399 3111
rect 2789 3009 2823 3043
rect 3985 3009 4019 3043
rect 4252 3009 4286 3043
rect 6561 3009 6595 3043
rect 7297 3009 7331 3043
rect 8401 3009 8435 3043
rect 8585 3009 8619 3043
rect 8953 3009 8987 3043
rect 9413 3009 9447 3043
rect 9680 3009 9714 3043
rect 11713 3009 11747 3043
rect 11989 3009 12023 3043
rect 13185 3009 13219 3043
rect 13277 3009 13311 3043
rect 14197 3009 14231 3043
rect 15209 3009 15243 3043
rect 15945 3009 15979 3043
rect 16895 3009 16929 3043
rect 17141 3009 17175 3043
rect 17969 3009 18003 3043
rect 20177 3009 20211 3043
rect 20453 3009 20487 3043
rect 20637 3009 20671 3043
rect 22017 3009 22051 3043
rect 22109 3009 22143 3043
rect 22477 3009 22511 3043
rect 23121 3009 23155 3043
rect 23765 3009 23799 3043
rect 24409 3009 24443 3043
rect 27445 3009 27479 3043
rect 29561 3009 29595 3043
rect 29929 3009 29963 3043
rect 30021 3009 30055 3043
rect 11897 2941 11931 2975
rect 14381 2941 14415 2975
rect 15393 2941 15427 2975
rect 18061 2941 18095 2975
rect 18153 2941 18187 2975
rect 19349 2941 19383 2975
rect 27629 2941 27663 2975
rect 2145 2873 2179 2907
rect 15025 2873 15059 2907
rect 16129 2873 16163 2907
rect 17049 2873 17083 2907
rect 20821 2873 20855 2907
rect 28549 2873 28583 2907
rect 3065 2805 3099 2839
rect 6745 2805 6779 2839
rect 11897 2805 11931 2839
rect 15209 2805 15243 2839
rect 18797 2805 18831 2839
rect 20269 2805 20303 2839
rect 22385 2805 22419 2839
rect 24225 2805 24259 2839
rect 27721 2805 27755 2839
rect 29561 2805 29595 2839
rect 4445 2601 4479 2635
rect 6561 2601 6595 2635
rect 8217 2601 8251 2635
rect 9137 2601 9171 2635
rect 14105 2601 14139 2635
rect 14473 2601 14507 2635
rect 15117 2601 15151 2635
rect 15485 2601 15519 2635
rect 16129 2601 16163 2635
rect 16681 2601 16715 2635
rect 17785 2601 17819 2635
rect 18245 2601 18279 2635
rect 19257 2601 19291 2635
rect 20269 2601 20303 2635
rect 20729 2601 20763 2635
rect 21833 2601 21867 2635
rect 22109 2601 22143 2635
rect 24409 2601 24443 2635
rect 25697 2601 25731 2635
rect 27169 2601 27203 2635
rect 27629 2601 27663 2635
rect 3065 2533 3099 2567
rect 7573 2533 7607 2567
rect 17325 2533 17359 2567
rect 2237 2465 2271 2499
rect 9873 2465 9907 2499
rect 11805 2465 11839 2499
rect 14565 2465 14599 2499
rect 15025 2465 15059 2499
rect 20453 2465 20487 2499
rect 1961 2397 1995 2431
rect 2881 2397 2915 2431
rect 4997 2397 5031 2431
rect 5273 2397 5307 2431
rect 6377 2397 6411 2431
rect 7389 2397 7423 2431
rect 8033 2397 8067 2431
rect 8953 2397 8987 2431
rect 9597 2397 9631 2431
rect 11529 2397 11563 2431
rect 12817 2397 12851 2431
rect 14289 2397 14323 2431
rect 15301 2397 15335 2431
rect 15945 2397 15979 2431
rect 16865 2397 16899 2431
rect 17509 2397 17543 2431
rect 17601 2397 17635 2431
rect 17785 2397 17819 2431
rect 18429 2397 18463 2431
rect 18613 2397 18647 2431
rect 18705 2397 18739 2431
rect 19441 2397 19475 2431
rect 20545 2397 20579 2431
rect 22017 2397 22051 2431
rect 22201 2397 22235 2431
rect 22845 2397 22879 2431
rect 23489 2397 23523 2431
rect 24593 2397 24627 2431
rect 25237 2397 25271 2431
rect 25881 2397 25915 2431
rect 26985 2397 27019 2431
rect 27813 2397 27847 2431
rect 28733 2397 28767 2431
rect 29837 2397 29871 2431
rect 4169 2329 4203 2363
rect 20269 2329 20303 2363
rect 13001 2261 13035 2295
rect 22661 2261 22695 2295
rect 23305 2261 23339 2295
rect 25053 2261 25087 2295
rect 28917 2261 28951 2295
rect 30021 2261 30055 2295
<< metal1 >>
rect 1104 45722 30820 45744
rect 1104 45670 10880 45722
rect 10932 45670 10944 45722
rect 10996 45670 11008 45722
rect 11060 45670 11072 45722
rect 11124 45670 11136 45722
rect 11188 45670 20811 45722
rect 20863 45670 20875 45722
rect 20927 45670 20939 45722
rect 20991 45670 21003 45722
rect 21055 45670 21067 45722
rect 21119 45670 30820 45722
rect 1104 45648 30820 45670
rect 1394 45432 1400 45484
rect 1452 45472 1458 45484
rect 1673 45475 1731 45481
rect 1673 45472 1685 45475
rect 1452 45444 1685 45472
rect 1452 45432 1458 45444
rect 1673 45441 1685 45444
rect 1719 45441 1731 45475
rect 1673 45435 1731 45441
rect 2409 45475 2467 45481
rect 2409 45441 2421 45475
rect 2455 45441 2467 45475
rect 2409 45435 2467 45441
rect 2424 45404 2452 45435
rect 2866 45432 2872 45484
rect 2924 45472 2930 45484
rect 3050 45472 3056 45484
rect 2924 45444 3056 45472
rect 2924 45432 2930 45444
rect 3050 45432 3056 45444
rect 3108 45432 3114 45484
rect 3142 45432 3148 45484
rect 3200 45472 3206 45484
rect 3973 45475 4031 45481
rect 3200 45444 3245 45472
rect 3200 45432 3206 45444
rect 3973 45441 3985 45475
rect 4019 45441 4031 45475
rect 3973 45435 4031 45441
rect 4617 45475 4675 45481
rect 4617 45441 4629 45475
rect 4663 45472 4675 45475
rect 4798 45472 4804 45484
rect 4663 45444 4804 45472
rect 4663 45441 4675 45444
rect 4617 45435 4675 45441
rect 3988 45404 4016 45435
rect 4798 45432 4804 45444
rect 4856 45432 4862 45484
rect 30098 45472 30104 45484
rect 30059 45444 30104 45472
rect 30098 45432 30104 45444
rect 30156 45432 30162 45484
rect 5258 45404 5264 45416
rect 2424 45376 3832 45404
rect 3988 45376 5264 45404
rect 2222 45336 2228 45348
rect 2183 45308 2228 45336
rect 2222 45296 2228 45308
rect 2280 45296 2286 45348
rect 2958 45336 2964 45348
rect 2919 45308 2964 45336
rect 2958 45296 2964 45308
rect 3016 45296 3022 45348
rect 3804 45345 3832 45376
rect 5258 45364 5264 45376
rect 5316 45364 5322 45416
rect 3789 45339 3847 45345
rect 3789 45305 3801 45339
rect 3835 45305 3847 45339
rect 3789 45299 3847 45305
rect 1489 45271 1547 45277
rect 1489 45237 1501 45271
rect 1535 45268 1547 45271
rect 2774 45268 2780 45280
rect 1535 45240 2780 45268
rect 1535 45237 1547 45240
rect 1489 45231 1547 45237
rect 2774 45228 2780 45240
rect 2832 45228 2838 45280
rect 2866 45228 2872 45280
rect 2924 45268 2930 45280
rect 4433 45271 4491 45277
rect 4433 45268 4445 45271
rect 2924 45240 4445 45268
rect 2924 45228 2930 45240
rect 4433 45237 4445 45240
rect 4479 45237 4491 45271
rect 29914 45268 29920 45280
rect 29875 45240 29920 45268
rect 4433 45231 4491 45237
rect 29914 45228 29920 45240
rect 29972 45228 29978 45280
rect 1104 45178 30820 45200
rect 1104 45126 5915 45178
rect 5967 45126 5979 45178
rect 6031 45126 6043 45178
rect 6095 45126 6107 45178
rect 6159 45126 6171 45178
rect 6223 45126 15846 45178
rect 15898 45126 15910 45178
rect 15962 45126 15974 45178
rect 16026 45126 16038 45178
rect 16090 45126 16102 45178
rect 16154 45126 25776 45178
rect 25828 45126 25840 45178
rect 25892 45126 25904 45178
rect 25956 45126 25968 45178
rect 26020 45126 26032 45178
rect 26084 45126 30820 45178
rect 1104 45104 30820 45126
rect 2225 45067 2283 45073
rect 2225 45033 2237 45067
rect 2271 45064 2283 45067
rect 3050 45064 3056 45076
rect 2271 45036 3056 45064
rect 2271 45033 2283 45036
rect 2225 45027 2283 45033
rect 3050 45024 3056 45036
rect 3108 45024 3114 45076
rect 3142 45024 3148 45076
rect 3200 45064 3206 45076
rect 4433 45067 4491 45073
rect 4433 45064 4445 45067
rect 3200 45036 4445 45064
rect 3200 45024 3206 45036
rect 4433 45033 4445 45036
rect 4479 45033 4491 45067
rect 4433 45027 4491 45033
rect 5166 45024 5172 45076
rect 5224 45064 5230 45076
rect 5445 45067 5503 45073
rect 5445 45064 5457 45067
rect 5224 45036 5457 45064
rect 5224 45024 5230 45036
rect 5445 45033 5457 45036
rect 5491 45033 5503 45067
rect 5445 45027 5503 45033
rect 5718 44928 5724 44940
rect 3068 44900 5724 44928
rect 1673 44863 1731 44869
rect 1673 44829 1685 44863
rect 1719 44829 1731 44863
rect 1673 44823 1731 44829
rect 2409 44863 2467 44869
rect 2409 44829 2421 44863
rect 2455 44860 2467 44863
rect 2866 44860 2872 44872
rect 2455 44832 2872 44860
rect 2455 44829 2467 44832
rect 2409 44823 2467 44829
rect 1688 44792 1716 44823
rect 2866 44820 2872 44832
rect 2924 44820 2930 44872
rect 3068 44869 3096 44900
rect 5718 44888 5724 44900
rect 5776 44888 5782 44940
rect 3053 44863 3111 44869
rect 3053 44829 3065 44863
rect 3099 44829 3111 44863
rect 3053 44823 3111 44829
rect 3973 44863 4031 44869
rect 3973 44829 3985 44863
rect 4019 44860 4031 44863
rect 4522 44860 4528 44872
rect 4019 44832 4528 44860
rect 4019 44829 4031 44832
rect 3973 44823 4031 44829
rect 4522 44820 4528 44832
rect 4580 44820 4586 44872
rect 4617 44863 4675 44869
rect 4617 44829 4629 44863
rect 4663 44860 4675 44863
rect 4663 44832 5304 44860
rect 4663 44829 4675 44832
rect 4617 44823 4675 44829
rect 1688 44764 3832 44792
rect 1486 44724 1492 44736
rect 1447 44696 1492 44724
rect 1486 44684 1492 44696
rect 1544 44684 1550 44736
rect 2866 44724 2872 44736
rect 2827 44696 2872 44724
rect 2866 44684 2872 44696
rect 2924 44684 2930 44736
rect 3804 44733 3832 44764
rect 5276 44733 5304 44832
rect 5534 44820 5540 44872
rect 5592 44860 5598 44872
rect 5813 44863 5871 44869
rect 5813 44860 5825 44863
rect 5592 44832 5825 44860
rect 5592 44820 5598 44832
rect 5813 44829 5825 44832
rect 5859 44829 5871 44863
rect 5813 44823 5871 44829
rect 6546 44820 6552 44872
rect 6604 44860 6610 44872
rect 6641 44863 6699 44869
rect 6641 44860 6653 44863
rect 6604 44832 6653 44860
rect 6604 44820 6610 44832
rect 6641 44829 6653 44832
rect 6687 44829 6699 44863
rect 6641 44823 6699 44829
rect 8386 44820 8392 44872
rect 8444 44860 8450 44872
rect 9125 44863 9183 44869
rect 9125 44860 9137 44863
rect 8444 44832 9137 44860
rect 8444 44820 8450 44832
rect 9125 44829 9137 44832
rect 9171 44829 9183 44863
rect 9125 44823 9183 44829
rect 30101 44863 30159 44869
rect 30101 44829 30113 44863
rect 30147 44860 30159 44863
rect 30190 44860 30196 44872
rect 30147 44832 30196 44860
rect 30147 44829 30159 44832
rect 30101 44823 30159 44829
rect 30190 44820 30196 44832
rect 30248 44820 30254 44872
rect 6908 44795 6966 44801
rect 6908 44761 6920 44795
rect 6954 44792 6966 44795
rect 7006 44792 7012 44804
rect 6954 44764 7012 44792
rect 6954 44761 6966 44764
rect 6908 44755 6966 44761
rect 7006 44752 7012 44764
rect 7064 44752 7070 44804
rect 3789 44727 3847 44733
rect 3789 44693 3801 44727
rect 3835 44693 3847 44727
rect 3789 44687 3847 44693
rect 5261 44727 5319 44733
rect 5261 44693 5273 44727
rect 5307 44693 5319 44727
rect 5261 44687 5319 44693
rect 5445 44727 5503 44733
rect 5445 44693 5457 44727
rect 5491 44724 5503 44727
rect 6270 44724 6276 44736
rect 5491 44696 6276 44724
rect 5491 44693 5503 44696
rect 5445 44687 5503 44693
rect 6270 44684 6276 44696
rect 6328 44684 6334 44736
rect 7190 44684 7196 44736
rect 7248 44724 7254 44736
rect 8021 44727 8079 44733
rect 8021 44724 8033 44727
rect 7248 44696 8033 44724
rect 7248 44684 7254 44696
rect 8021 44693 8033 44696
rect 8067 44693 8079 44727
rect 8938 44724 8944 44736
rect 8899 44696 8944 44724
rect 8021 44687 8079 44693
rect 8938 44684 8944 44696
rect 8996 44684 9002 44736
rect 28994 44684 29000 44736
rect 29052 44724 29058 44736
rect 29917 44727 29975 44733
rect 29917 44724 29929 44727
rect 29052 44696 29929 44724
rect 29052 44684 29058 44696
rect 29917 44693 29929 44696
rect 29963 44693 29975 44727
rect 29917 44687 29975 44693
rect 1104 44634 30820 44656
rect 1104 44582 10880 44634
rect 10932 44582 10944 44634
rect 10996 44582 11008 44634
rect 11060 44582 11072 44634
rect 11124 44582 11136 44634
rect 11188 44582 20811 44634
rect 20863 44582 20875 44634
rect 20927 44582 20939 44634
rect 20991 44582 21003 44634
rect 21055 44582 21067 44634
rect 21119 44582 30820 44634
rect 1104 44560 30820 44582
rect 4798 44520 4804 44532
rect 4759 44492 4804 44520
rect 4798 44480 4804 44492
rect 4856 44480 4862 44532
rect 5258 44520 5264 44532
rect 5219 44492 5264 44520
rect 5258 44480 5264 44492
rect 5316 44480 5322 44532
rect 6546 44520 6552 44532
rect 6507 44492 6552 44520
rect 6546 44480 6552 44492
rect 6604 44480 6610 44532
rect 7006 44520 7012 44532
rect 6967 44492 7012 44520
rect 7006 44480 7012 44492
rect 7064 44480 7070 44532
rect 7558 44480 7564 44532
rect 7616 44520 7622 44532
rect 7616 44492 8708 44520
rect 7616 44480 7622 44492
rect 2866 44452 2872 44464
rect 1688 44424 2872 44452
rect 1688 44393 1716 44424
rect 2866 44412 2872 44424
rect 2924 44412 2930 44464
rect 4617 44455 4675 44461
rect 4617 44421 4629 44455
rect 4663 44421 4675 44455
rect 4617 44415 4675 44421
rect 5445 44455 5503 44461
rect 5445 44421 5457 44455
rect 5491 44452 5503 44455
rect 8680 44452 8708 44492
rect 8754 44480 8760 44532
rect 8812 44520 8818 44532
rect 10502 44520 10508 44532
rect 8812 44492 10508 44520
rect 8812 44480 8818 44492
rect 10502 44480 10508 44492
rect 10560 44520 10566 44532
rect 18138 44520 18144 44532
rect 10560 44492 18144 44520
rect 10560 44480 10566 44492
rect 18138 44480 18144 44492
rect 18196 44480 18202 44532
rect 5491 44424 6914 44452
rect 5491 44421 5503 44424
rect 5445 44415 5503 44421
rect 1673 44387 1731 44393
rect 1673 44353 1685 44387
rect 1719 44353 1731 44387
rect 2314 44384 2320 44396
rect 2275 44356 2320 44384
rect 1673 44347 1731 44353
rect 2314 44344 2320 44356
rect 2372 44344 2378 44396
rect 2961 44387 3019 44393
rect 2961 44353 2973 44387
rect 3007 44353 3019 44387
rect 2961 44347 3019 44353
rect 3605 44387 3663 44393
rect 3605 44353 3617 44387
rect 3651 44384 3663 44387
rect 4246 44384 4252 44396
rect 3651 44356 4252 44384
rect 3651 44353 3663 44356
rect 3605 44347 3663 44353
rect 2976 44316 3004 44347
rect 4246 44344 4252 44356
rect 4304 44344 4310 44396
rect 3970 44316 3976 44328
rect 2976 44288 3976 44316
rect 3970 44276 3976 44288
rect 4028 44276 4034 44328
rect 4632 44316 4660 44415
rect 6362 44384 6368 44396
rect 6323 44356 6368 44384
rect 6362 44344 6368 44356
rect 6420 44344 6426 44396
rect 6886 44384 6914 44424
rect 7392 44424 8616 44452
rect 8680 44424 16574 44452
rect 7190 44384 7196 44396
rect 6886 44356 7196 44384
rect 7190 44344 7196 44356
rect 7248 44344 7254 44396
rect 7392 44328 7420 44424
rect 7558 44384 7564 44396
rect 7519 44356 7564 44384
rect 7558 44344 7564 44356
rect 7616 44344 7622 44396
rect 7742 44384 7748 44396
rect 7703 44356 7748 44384
rect 7742 44344 7748 44356
rect 7800 44384 7806 44396
rect 8205 44387 8263 44393
rect 8205 44384 8217 44387
rect 7800 44356 8217 44384
rect 7800 44344 7806 44356
rect 8205 44353 8217 44356
rect 8251 44353 8263 44387
rect 8205 44347 8263 44353
rect 8294 44344 8300 44396
rect 8352 44384 8358 44396
rect 8588 44393 8616 44424
rect 8389 44387 8447 44393
rect 8389 44384 8401 44387
rect 8352 44356 8401 44384
rect 8352 44344 8358 44356
rect 8389 44353 8401 44356
rect 8435 44353 8447 44387
rect 8389 44347 8447 44353
rect 8573 44387 8631 44393
rect 8573 44353 8585 44387
rect 8619 44353 8631 44387
rect 8573 44347 8631 44353
rect 8757 44387 8815 44393
rect 8757 44353 8769 44387
rect 8803 44353 8815 44387
rect 8757 44347 8815 44353
rect 7374 44316 7380 44328
rect 4632 44288 6914 44316
rect 7335 44288 7380 44316
rect 4249 44251 4307 44257
rect 4249 44217 4261 44251
rect 4295 44248 4307 44251
rect 5534 44248 5540 44260
rect 4295 44220 5540 44248
rect 4295 44217 4307 44220
rect 4249 44211 4307 44217
rect 5534 44208 5540 44220
rect 5592 44248 5598 44260
rect 5813 44251 5871 44257
rect 5813 44248 5825 44251
rect 5592 44220 5825 44248
rect 5592 44208 5598 44220
rect 5813 44217 5825 44220
rect 5859 44217 5871 44251
rect 6886 44248 6914 44288
rect 7374 44276 7380 44288
rect 7432 44276 7438 44328
rect 7469 44319 7527 44325
rect 7469 44285 7481 44319
rect 7515 44316 7527 44319
rect 7834 44316 7840 44328
rect 7515 44288 7840 44316
rect 7515 44285 7527 44288
rect 7469 44279 7527 44285
rect 7834 44276 7840 44288
rect 7892 44316 7898 44328
rect 8481 44319 8539 44325
rect 8481 44316 8493 44319
rect 7892 44288 8493 44316
rect 7892 44276 7898 44288
rect 8481 44285 8493 44288
rect 8527 44285 8539 44319
rect 8481 44279 8539 44285
rect 8772 44248 8800 44347
rect 9122 44344 9128 44396
rect 9180 44384 9186 44396
rect 9401 44387 9459 44393
rect 9401 44384 9413 44387
rect 9180 44356 9413 44384
rect 9180 44344 9186 44356
rect 9401 44353 9413 44356
rect 9447 44353 9459 44387
rect 9401 44347 9459 44353
rect 8846 44248 8852 44260
rect 6886 44220 8852 44248
rect 5813 44211 5871 44217
rect 8846 44208 8852 44220
rect 8904 44208 8910 44260
rect 8941 44251 8999 44257
rect 8941 44217 8953 44251
rect 8987 44248 8999 44251
rect 9950 44248 9956 44260
rect 8987 44220 9956 44248
rect 8987 44217 8999 44220
rect 8941 44211 8999 44217
rect 9950 44208 9956 44220
rect 10008 44208 10014 44260
rect 16546 44248 16574 44424
rect 18322 44384 18328 44396
rect 18283 44356 18328 44384
rect 18322 44344 18328 44356
rect 18380 44344 18386 44396
rect 30098 44384 30104 44396
rect 30059 44356 30104 44384
rect 30098 44344 30104 44356
rect 30156 44344 30162 44396
rect 18509 44319 18567 44325
rect 18509 44285 18521 44319
rect 18555 44316 18567 44319
rect 29914 44316 29920 44328
rect 18555 44288 29920 44316
rect 18555 44285 18567 44288
rect 18509 44279 18567 44285
rect 29914 44276 29920 44288
rect 29972 44276 29978 44328
rect 18046 44248 18052 44260
rect 16546 44220 18052 44248
rect 18046 44208 18052 44220
rect 18104 44208 18110 44260
rect 1486 44180 1492 44192
rect 1447 44152 1492 44180
rect 1486 44140 1492 44152
rect 1544 44140 1550 44192
rect 1946 44140 1952 44192
rect 2004 44180 2010 44192
rect 2133 44183 2191 44189
rect 2133 44180 2145 44183
rect 2004 44152 2145 44180
rect 2004 44140 2010 44152
rect 2133 44149 2145 44152
rect 2179 44149 2191 44183
rect 2133 44143 2191 44149
rect 2777 44183 2835 44189
rect 2777 44149 2789 44183
rect 2823 44180 2835 44183
rect 2958 44180 2964 44192
rect 2823 44152 2964 44180
rect 2823 44149 2835 44152
rect 2777 44143 2835 44149
rect 2958 44140 2964 44152
rect 3016 44140 3022 44192
rect 3418 44180 3424 44192
rect 3379 44152 3424 44180
rect 3418 44140 3424 44152
rect 3476 44140 3482 44192
rect 4617 44183 4675 44189
rect 4617 44149 4629 44183
rect 4663 44180 4675 44183
rect 5166 44180 5172 44192
rect 4663 44152 5172 44180
rect 4663 44149 4675 44152
rect 4617 44143 4675 44149
rect 5166 44140 5172 44152
rect 5224 44180 5230 44192
rect 5445 44183 5503 44189
rect 5445 44180 5457 44183
rect 5224 44152 5457 44180
rect 5224 44140 5230 44152
rect 5445 44149 5457 44152
rect 5491 44149 5503 44183
rect 5445 44143 5503 44149
rect 8294 44140 8300 44192
rect 8352 44180 8358 44192
rect 8754 44180 8760 44192
rect 8352 44152 8760 44180
rect 8352 44140 8358 44152
rect 8754 44140 8760 44152
rect 8812 44140 8818 44192
rect 9585 44183 9643 44189
rect 9585 44149 9597 44183
rect 9631 44180 9643 44183
rect 10226 44180 10232 44192
rect 9631 44152 10232 44180
rect 9631 44149 9643 44152
rect 9585 44143 9643 44149
rect 10226 44140 10232 44152
rect 10284 44140 10290 44192
rect 17954 44140 17960 44192
rect 18012 44180 18018 44192
rect 18141 44183 18199 44189
rect 18141 44180 18153 44183
rect 18012 44152 18153 44180
rect 18012 44140 18018 44152
rect 18141 44149 18153 44152
rect 18187 44149 18199 44183
rect 29914 44180 29920 44192
rect 29875 44152 29920 44180
rect 18141 44143 18199 44149
rect 29914 44140 29920 44152
rect 29972 44140 29978 44192
rect 1104 44090 30820 44112
rect 1104 44038 5915 44090
rect 5967 44038 5979 44090
rect 6031 44038 6043 44090
rect 6095 44038 6107 44090
rect 6159 44038 6171 44090
rect 6223 44038 15846 44090
rect 15898 44038 15910 44090
rect 15962 44038 15974 44090
rect 16026 44038 16038 44090
rect 16090 44038 16102 44090
rect 16154 44038 25776 44090
rect 25828 44038 25840 44090
rect 25892 44038 25904 44090
rect 25956 44038 25968 44090
rect 26020 44038 26032 44090
rect 26084 44038 30820 44090
rect 1104 44016 30820 44038
rect 4522 43936 4528 43988
rect 4580 43976 4586 43988
rect 5261 43979 5319 43985
rect 5261 43976 5273 43979
rect 4580 43948 5273 43976
rect 4580 43936 4586 43948
rect 5261 43945 5273 43948
rect 5307 43945 5319 43979
rect 5261 43939 5319 43945
rect 5445 43979 5503 43985
rect 5445 43945 5457 43979
rect 5491 43945 5503 43979
rect 5445 43939 5503 43945
rect 2501 43911 2559 43917
rect 2501 43877 2513 43911
rect 2547 43908 2559 43911
rect 3142 43908 3148 43920
rect 2547 43880 3148 43908
rect 2547 43877 2559 43880
rect 2501 43871 2559 43877
rect 3142 43868 3148 43880
rect 3200 43868 3206 43920
rect 5166 43868 5172 43920
rect 5224 43908 5230 43920
rect 5460 43908 5488 43939
rect 6362 43936 6368 43988
rect 6420 43976 6426 43988
rect 6549 43979 6607 43985
rect 6549 43976 6561 43979
rect 6420 43948 6561 43976
rect 6420 43936 6426 43948
rect 6549 43945 6561 43948
rect 6595 43945 6607 43979
rect 6549 43939 6607 43945
rect 7561 43979 7619 43985
rect 7561 43945 7573 43979
rect 7607 43976 7619 43979
rect 7742 43976 7748 43988
rect 7607 43948 7748 43976
rect 7607 43945 7619 43948
rect 7561 43939 7619 43945
rect 7742 43936 7748 43948
rect 7800 43936 7806 43988
rect 18138 43976 18144 43988
rect 18099 43948 18144 43976
rect 18138 43936 18144 43948
rect 18196 43936 18202 43988
rect 5224 43880 5488 43908
rect 5224 43868 5230 43880
rect 6270 43868 6276 43920
rect 6328 43908 6334 43920
rect 10321 43911 10379 43917
rect 6328 43880 8248 43908
rect 6328 43868 6334 43880
rect 7374 43800 7380 43852
rect 7432 43840 7438 43852
rect 8021 43843 8079 43849
rect 8021 43840 8033 43843
rect 7432 43812 8033 43840
rect 7432 43800 7438 43812
rect 8021 43809 8033 43812
rect 8067 43809 8079 43843
rect 8021 43803 8079 43809
rect 1854 43772 1860 43784
rect 1815 43744 1860 43772
rect 1854 43732 1860 43744
rect 1912 43732 1918 43784
rect 2317 43775 2375 43781
rect 2317 43741 2329 43775
rect 2363 43772 2375 43775
rect 2498 43772 2504 43784
rect 2363 43744 2504 43772
rect 2363 43741 2375 43744
rect 2317 43735 2375 43741
rect 2498 43732 2504 43744
rect 2556 43732 2562 43784
rect 3145 43775 3203 43781
rect 3145 43741 3157 43775
rect 3191 43741 3203 43775
rect 3145 43735 3203 43741
rect 3789 43775 3847 43781
rect 3789 43741 3801 43775
rect 3835 43772 3847 43775
rect 5074 43772 5080 43784
rect 3835 43744 5080 43772
rect 3835 43741 3847 43744
rect 3789 43735 3847 43741
rect 3160 43704 3188 43735
rect 5074 43732 5080 43744
rect 5132 43732 5138 43784
rect 5534 43732 5540 43784
rect 5592 43772 5598 43784
rect 5813 43775 5871 43781
rect 5813 43772 5825 43775
rect 5592 43744 5825 43772
rect 5592 43732 5598 43744
rect 5813 43741 5825 43744
rect 5859 43741 5871 43775
rect 5813 43735 5871 43741
rect 5902 43732 5908 43784
rect 5960 43772 5966 43784
rect 6638 43772 6644 43784
rect 5960 43744 6644 43772
rect 5960 43732 5966 43744
rect 6638 43732 6644 43744
rect 6696 43772 6702 43784
rect 6733 43775 6791 43781
rect 6733 43772 6745 43775
rect 6696 43744 6745 43772
rect 6696 43732 6702 43744
rect 6733 43741 6745 43744
rect 6779 43741 6791 43775
rect 6733 43735 6791 43741
rect 7561 43775 7619 43781
rect 7561 43741 7573 43775
rect 7607 43772 7619 43775
rect 7653 43775 7711 43781
rect 7653 43772 7665 43775
rect 7607 43744 7665 43772
rect 7607 43741 7619 43744
rect 7561 43735 7619 43741
rect 7653 43741 7665 43744
rect 7699 43741 7711 43775
rect 7653 43735 7711 43741
rect 7837 43775 7895 43781
rect 7837 43741 7849 43775
rect 7883 43741 7895 43775
rect 7837 43735 7895 43741
rect 5626 43704 5632 43716
rect 3160 43676 5632 43704
rect 5626 43664 5632 43676
rect 5684 43664 5690 43716
rect 7668 43704 7696 43735
rect 7742 43704 7748 43716
rect 7668 43676 7748 43704
rect 7742 43664 7748 43676
rect 7800 43664 7806 43716
rect 1578 43596 1584 43648
rect 1636 43636 1642 43648
rect 1673 43639 1731 43645
rect 1673 43636 1685 43639
rect 1636 43608 1685 43636
rect 1636 43596 1642 43608
rect 1673 43605 1685 43608
rect 1719 43605 1731 43639
rect 1673 43599 1731 43605
rect 2961 43639 3019 43645
rect 2961 43605 2973 43639
rect 3007 43636 3019 43639
rect 3234 43636 3240 43648
rect 3007 43608 3240 43636
rect 3007 43605 3019 43608
rect 2961 43599 3019 43605
rect 3234 43596 3240 43608
rect 3292 43596 3298 43648
rect 3973 43639 4031 43645
rect 3973 43605 3985 43639
rect 4019 43636 4031 43639
rect 5350 43636 5356 43648
rect 4019 43608 5356 43636
rect 4019 43605 4031 43608
rect 3973 43599 4031 43605
rect 5350 43596 5356 43608
rect 5408 43596 5414 43648
rect 5445 43639 5503 43645
rect 5445 43605 5457 43639
rect 5491 43636 5503 43639
rect 7190 43636 7196 43648
rect 5491 43608 7196 43636
rect 5491 43605 5503 43608
rect 5445 43599 5503 43605
rect 7190 43596 7196 43608
rect 7248 43596 7254 43648
rect 7282 43596 7288 43648
rect 7340 43636 7346 43648
rect 7852 43636 7880 43735
rect 7926 43732 7932 43784
rect 7984 43772 7990 43784
rect 8220 43781 8248 43880
rect 10321 43877 10333 43911
rect 10367 43877 10379 43911
rect 10321 43871 10379 43877
rect 8938 43840 8944 43852
rect 8899 43812 8944 43840
rect 8938 43800 8944 43812
rect 8996 43800 9002 43852
rect 8205 43775 8263 43781
rect 7984 43744 8029 43772
rect 7984 43732 7990 43744
rect 8205 43741 8217 43775
rect 8251 43772 8263 43775
rect 10336 43772 10364 43871
rect 18322 43772 18328 43784
rect 8251 43744 10364 43772
rect 18283 43744 18328 43772
rect 8251 43741 8263 43744
rect 8205 43735 8263 43741
rect 18322 43732 18328 43744
rect 18380 43732 18386 43784
rect 18509 43775 18567 43781
rect 18509 43741 18521 43775
rect 18555 43772 18567 43775
rect 28994 43772 29000 43784
rect 18555 43744 29000 43772
rect 18555 43741 18567 43744
rect 18509 43735 18567 43741
rect 28994 43732 29000 43744
rect 29052 43732 29058 43784
rect 8389 43707 8447 43713
rect 8389 43673 8401 43707
rect 8435 43704 8447 43707
rect 9186 43707 9244 43713
rect 9186 43704 9198 43707
rect 8435 43676 9198 43704
rect 8435 43673 8447 43676
rect 8389 43667 8447 43673
rect 9186 43673 9198 43676
rect 9232 43673 9244 43707
rect 10686 43704 10692 43716
rect 9186 43667 9244 43673
rect 9324 43676 10692 43704
rect 9324 43636 9352 43676
rect 10686 43664 10692 43676
rect 10744 43704 10750 43716
rect 17954 43704 17960 43716
rect 10744 43676 17960 43704
rect 10744 43664 10750 43676
rect 17954 43664 17960 43676
rect 18012 43664 18018 43716
rect 7340 43608 9352 43636
rect 7340 43596 7346 43608
rect 1104 43546 30820 43568
rect 1104 43494 10880 43546
rect 10932 43494 10944 43546
rect 10996 43494 11008 43546
rect 11060 43494 11072 43546
rect 11124 43494 11136 43546
rect 11188 43494 20811 43546
rect 20863 43494 20875 43546
rect 20927 43494 20939 43546
rect 20991 43494 21003 43546
rect 21055 43494 21067 43546
rect 21119 43494 30820 43546
rect 1104 43472 30820 43494
rect 7190 43392 7196 43444
rect 7248 43432 7254 43444
rect 8113 43435 8171 43441
rect 8113 43432 8125 43435
rect 7248 43404 8125 43432
rect 7248 43392 7254 43404
rect 8113 43401 8125 43404
rect 8159 43401 8171 43435
rect 8846 43432 8852 43444
rect 8807 43404 8852 43432
rect 8113 43395 8171 43401
rect 8846 43392 8852 43404
rect 8904 43392 8910 43444
rect 18046 43392 18052 43444
rect 18104 43432 18110 43444
rect 18141 43435 18199 43441
rect 18141 43432 18153 43435
rect 18104 43404 18153 43432
rect 18104 43392 18110 43404
rect 18141 43401 18153 43404
rect 18187 43401 18199 43435
rect 18141 43395 18199 43401
rect 3418 43364 3424 43376
rect 1688 43336 3424 43364
rect 1688 43305 1716 43336
rect 3418 43324 3424 43336
rect 3476 43324 3482 43376
rect 9950 43324 9956 43376
rect 10008 43373 10014 43376
rect 10008 43364 10020 43373
rect 10008 43336 10053 43364
rect 10008 43327 10020 43336
rect 10008 43324 10014 43327
rect 1673 43299 1731 43305
rect 1673 43265 1685 43299
rect 1719 43265 1731 43299
rect 1673 43259 1731 43265
rect 2501 43299 2559 43305
rect 2501 43265 2513 43299
rect 2547 43296 2559 43299
rect 2866 43296 2872 43308
rect 2547 43268 2872 43296
rect 2547 43265 2559 43268
rect 2501 43259 2559 43265
rect 2866 43256 2872 43268
rect 2924 43256 2930 43308
rect 3878 43296 3884 43308
rect 3839 43268 3884 43296
rect 3878 43256 3884 43268
rect 3936 43256 3942 43308
rect 4522 43296 4528 43308
rect 4483 43268 4528 43296
rect 4522 43256 4528 43268
rect 4580 43256 4586 43308
rect 4985 43299 5043 43305
rect 4985 43265 4997 43299
rect 5031 43296 5043 43299
rect 5074 43296 5080 43308
rect 5031 43268 5080 43296
rect 5031 43265 5043 43268
rect 4985 43259 5043 43265
rect 5074 43256 5080 43268
rect 5132 43256 5138 43308
rect 5629 43299 5687 43305
rect 5629 43265 5641 43299
rect 5675 43296 5687 43299
rect 5902 43296 5908 43308
rect 5675 43268 5908 43296
rect 5675 43265 5687 43268
rect 5629 43259 5687 43265
rect 5902 43256 5908 43268
rect 5960 43256 5966 43308
rect 7006 43305 7012 43308
rect 7000 43259 7012 43305
rect 7064 43296 7070 43308
rect 10226 43296 10232 43308
rect 7064 43268 7100 43296
rect 10187 43268 10232 43296
rect 7006 43256 7012 43259
rect 7064 43256 7070 43268
rect 10226 43256 10232 43268
rect 10284 43256 10290 43308
rect 18322 43296 18328 43308
rect 18235 43268 18328 43296
rect 18322 43256 18328 43268
rect 18380 43296 18386 43308
rect 19058 43296 19064 43308
rect 18380 43268 19064 43296
rect 18380 43256 18386 43268
rect 19058 43256 19064 43268
rect 19116 43256 19122 43308
rect 6730 43228 6736 43240
rect 6691 43200 6736 43228
rect 6730 43188 6736 43200
rect 6788 43188 6794 43240
rect 18509 43231 18567 43237
rect 18509 43197 18521 43231
rect 18555 43228 18567 43231
rect 29914 43228 29920 43240
rect 18555 43200 29920 43228
rect 18555 43197 18567 43200
rect 18509 43191 18567 43197
rect 29914 43188 29920 43200
rect 29972 43188 29978 43240
rect 1486 43092 1492 43104
rect 1447 43064 1492 43092
rect 1486 43052 1492 43064
rect 1544 43052 1550 43104
rect 2685 43095 2743 43101
rect 2685 43061 2697 43095
rect 2731 43092 2743 43095
rect 2774 43092 2780 43104
rect 2731 43064 2780 43092
rect 2731 43061 2743 43064
rect 2685 43055 2743 43061
rect 2774 43052 2780 43064
rect 2832 43052 2838 43104
rect 3050 43052 3056 43104
rect 3108 43092 3114 43104
rect 3697 43095 3755 43101
rect 3697 43092 3709 43095
rect 3108 43064 3709 43092
rect 3108 43052 3114 43064
rect 3697 43061 3709 43064
rect 3743 43061 3755 43095
rect 4338 43092 4344 43104
rect 4299 43064 4344 43092
rect 3697 43055 3755 43061
rect 4338 43052 4344 43064
rect 4396 43052 4402 43104
rect 5166 43092 5172 43104
rect 5127 43064 5172 43092
rect 5166 43052 5172 43064
rect 5224 43052 5230 43104
rect 5813 43095 5871 43101
rect 5813 43061 5825 43095
rect 5859 43092 5871 43095
rect 6914 43092 6920 43104
rect 5859 43064 6920 43092
rect 5859 43061 5871 43064
rect 5813 43055 5871 43061
rect 6914 43052 6920 43064
rect 6972 43052 6978 43104
rect 1104 43002 30820 43024
rect 1104 42950 5915 43002
rect 5967 42950 5979 43002
rect 6031 42950 6043 43002
rect 6095 42950 6107 43002
rect 6159 42950 6171 43002
rect 6223 42950 15846 43002
rect 15898 42950 15910 43002
rect 15962 42950 15974 43002
rect 16026 42950 16038 43002
rect 16090 42950 16102 43002
rect 16154 42950 25776 43002
rect 25828 42950 25840 43002
rect 25892 42950 25904 43002
rect 25956 42950 25968 43002
rect 26020 42950 26032 43002
rect 26084 42950 30820 43002
rect 1104 42928 30820 42950
rect 5166 42848 5172 42900
rect 5224 42888 5230 42900
rect 6181 42891 6239 42897
rect 6181 42888 6193 42891
rect 5224 42860 6193 42888
rect 5224 42848 5230 42860
rect 6181 42857 6193 42860
rect 6227 42857 6239 42891
rect 7006 42888 7012 42900
rect 6967 42860 7012 42888
rect 6181 42851 6239 42857
rect 7006 42848 7012 42860
rect 7064 42848 7070 42900
rect 7834 42820 7840 42832
rect 7484 42792 7840 42820
rect 2958 42752 2964 42764
rect 1688 42724 2964 42752
rect 1688 42693 1716 42724
rect 2958 42712 2964 42724
rect 3016 42712 3022 42764
rect 1673 42687 1731 42693
rect 1673 42653 1685 42687
rect 1719 42653 1731 42687
rect 2130 42684 2136 42696
rect 2091 42656 2136 42684
rect 1673 42647 1731 42653
rect 2130 42644 2136 42656
rect 2188 42644 2194 42696
rect 3050 42684 3056 42696
rect 3011 42656 3056 42684
rect 3050 42644 3056 42656
rect 3108 42644 3114 42696
rect 4157 42687 4215 42693
rect 4157 42684 4169 42687
rect 3252 42656 4169 42684
rect 1486 42548 1492 42560
rect 1447 42520 1492 42548
rect 1486 42508 1492 42520
rect 1544 42508 1550 42560
rect 2317 42551 2375 42557
rect 2317 42517 2329 42551
rect 2363 42548 2375 42551
rect 2590 42548 2596 42560
rect 2363 42520 2596 42548
rect 2363 42517 2375 42520
rect 2317 42511 2375 42517
rect 2590 42508 2596 42520
rect 2648 42508 2654 42560
rect 3252 42557 3280 42656
rect 4157 42653 4169 42656
rect 4203 42653 4215 42687
rect 4157 42647 4215 42653
rect 5902 42644 5908 42696
rect 5960 42684 5966 42696
rect 6549 42687 6607 42693
rect 6549 42684 6561 42687
rect 5960 42656 6561 42684
rect 5960 42644 5966 42656
rect 6549 42653 6561 42656
rect 6595 42653 6607 42687
rect 7190 42684 7196 42696
rect 7151 42656 7196 42684
rect 6549 42647 6607 42653
rect 7190 42644 7196 42656
rect 7248 42644 7254 42696
rect 7374 42684 7380 42696
rect 7335 42656 7380 42684
rect 7374 42644 7380 42656
rect 7432 42644 7438 42696
rect 7484 42693 7512 42792
rect 7834 42780 7840 42792
rect 7892 42780 7898 42832
rect 7466 42687 7524 42693
rect 7466 42653 7478 42687
rect 7512 42653 7524 42687
rect 7466 42647 7524 42653
rect 7561 42687 7619 42693
rect 7561 42653 7573 42687
rect 7607 42684 7619 42687
rect 7650 42684 7656 42696
rect 7607 42656 7656 42684
rect 7607 42653 7619 42656
rect 7561 42647 7619 42653
rect 7650 42644 7656 42656
rect 7708 42644 7714 42696
rect 7742 42644 7748 42696
rect 7800 42684 7806 42696
rect 7800 42656 7893 42684
rect 7800 42644 7806 42656
rect 8018 42644 8024 42696
rect 8076 42684 8082 42696
rect 8205 42687 8263 42693
rect 8205 42684 8217 42687
rect 8076 42656 8217 42684
rect 8076 42644 8082 42656
rect 8205 42653 8217 42656
rect 8251 42684 8263 42687
rect 8941 42687 8999 42693
rect 8941 42684 8953 42687
rect 8251 42656 8953 42684
rect 8251 42653 8263 42656
rect 8205 42647 8263 42653
rect 8941 42653 8953 42656
rect 8987 42653 8999 42687
rect 30098 42684 30104 42696
rect 30059 42656 30104 42684
rect 8941 42647 8999 42653
rect 30098 42644 30104 42656
rect 30156 42644 30162 42696
rect 4430 42625 4436 42628
rect 4424 42579 4436 42625
rect 4488 42616 4494 42628
rect 4488 42588 4524 42616
rect 4430 42576 4436 42579
rect 4488 42576 4494 42588
rect 5718 42576 5724 42628
rect 5776 42616 5782 42628
rect 7760 42616 7788 42644
rect 10318 42616 10324 42628
rect 5776 42588 6040 42616
rect 7760 42588 10324 42616
rect 5776 42576 5782 42588
rect 3237 42551 3295 42557
rect 3237 42517 3249 42551
rect 3283 42517 3295 42551
rect 3237 42511 3295 42517
rect 5537 42551 5595 42557
rect 5537 42517 5549 42551
rect 5583 42548 5595 42551
rect 5810 42548 5816 42560
rect 5583 42520 5816 42548
rect 5583 42517 5595 42520
rect 5537 42511 5595 42517
rect 5810 42508 5816 42520
rect 5868 42508 5874 42560
rect 6012 42557 6040 42588
rect 10318 42576 10324 42588
rect 10376 42576 10382 42628
rect 5997 42551 6055 42557
rect 5997 42517 6009 42551
rect 6043 42517 6055 42551
rect 5997 42511 6055 42517
rect 6181 42551 6239 42557
rect 6181 42517 6193 42551
rect 6227 42548 6239 42551
rect 7926 42548 7932 42560
rect 6227 42520 7932 42548
rect 6227 42517 6239 42520
rect 6181 42511 6239 42517
rect 7926 42508 7932 42520
rect 7984 42508 7990 42560
rect 8386 42548 8392 42560
rect 8347 42520 8392 42548
rect 8386 42508 8392 42520
rect 8444 42508 8450 42560
rect 9122 42548 9128 42560
rect 9083 42520 9128 42548
rect 9122 42508 9128 42520
rect 9180 42508 9186 42560
rect 29914 42548 29920 42560
rect 29875 42520 29920 42548
rect 29914 42508 29920 42520
rect 29972 42508 29978 42560
rect 1104 42458 30820 42480
rect 1104 42406 10880 42458
rect 10932 42406 10944 42458
rect 10996 42406 11008 42458
rect 11060 42406 11072 42458
rect 11124 42406 11136 42458
rect 11188 42406 20811 42458
rect 20863 42406 20875 42458
rect 20927 42406 20939 42458
rect 20991 42406 21003 42458
rect 21055 42406 21067 42458
rect 21119 42406 30820 42458
rect 1104 42384 30820 42406
rect 4246 42304 4252 42356
rect 4304 42344 4310 42356
rect 5261 42347 5319 42353
rect 5261 42344 5273 42347
rect 4304 42316 5273 42344
rect 4304 42304 4310 42316
rect 5261 42313 5273 42316
rect 5307 42313 5319 42347
rect 6730 42344 6736 42356
rect 6691 42316 6736 42344
rect 5261 42307 5319 42313
rect 6730 42304 6736 42316
rect 6788 42304 6794 42356
rect 7374 42304 7380 42356
rect 7432 42344 7438 42356
rect 7742 42344 7748 42356
rect 7432 42316 7748 42344
rect 7432 42304 7438 42316
rect 7742 42304 7748 42316
rect 7800 42304 7806 42356
rect 7926 42344 7932 42356
rect 7887 42316 7932 42344
rect 7926 42304 7932 42316
rect 7984 42304 7990 42356
rect 4338 42276 4344 42288
rect 1688 42248 4344 42276
rect 1688 42217 1716 42248
rect 4338 42236 4344 42248
rect 4396 42236 4402 42288
rect 5445 42279 5503 42285
rect 5445 42245 5457 42279
rect 5491 42276 5503 42279
rect 6546 42276 6552 42288
rect 5491 42248 6552 42276
rect 5491 42245 5503 42248
rect 5445 42239 5503 42245
rect 6546 42236 6552 42248
rect 6604 42236 6610 42288
rect 1673 42211 1731 42217
rect 1673 42177 1685 42211
rect 1719 42177 1731 42211
rect 1673 42171 1731 42177
rect 2317 42211 2375 42217
rect 2317 42177 2329 42211
rect 2363 42208 2375 42211
rect 2406 42208 2412 42220
rect 2363 42180 2412 42208
rect 2363 42177 2375 42180
rect 2317 42171 2375 42177
rect 2406 42168 2412 42180
rect 2464 42168 2470 42220
rect 2774 42208 2780 42220
rect 2735 42180 2780 42208
rect 2774 42168 2780 42180
rect 2832 42168 2838 42220
rect 3044 42211 3102 42217
rect 3044 42177 3056 42211
rect 3090 42208 3102 42211
rect 3418 42208 3424 42220
rect 3090 42180 3424 42208
rect 3090 42177 3102 42180
rect 3044 42171 3102 42177
rect 3418 42168 3424 42180
rect 3476 42168 3482 42220
rect 3510 42168 3516 42220
rect 3568 42208 3574 42220
rect 4801 42211 4859 42217
rect 4801 42208 4813 42211
rect 3568 42180 4813 42208
rect 3568 42168 3574 42180
rect 4801 42177 4813 42180
rect 4847 42177 4859 42211
rect 4801 42171 4859 42177
rect 5813 42211 5871 42217
rect 5813 42177 5825 42211
rect 5859 42208 5871 42211
rect 5902 42208 5908 42220
rect 5859 42180 5908 42208
rect 5859 42177 5871 42180
rect 5813 42171 5871 42177
rect 5902 42168 5908 42180
rect 5960 42208 5966 42220
rect 6270 42208 6276 42220
rect 5960 42180 6276 42208
rect 5960 42168 5966 42180
rect 6270 42168 6276 42180
rect 6328 42168 6334 42220
rect 6914 42168 6920 42220
rect 6972 42208 6978 42220
rect 6972 42180 7017 42208
rect 6972 42168 6978 42180
rect 8110 42168 8116 42220
rect 8168 42208 8174 42220
rect 9042 42211 9100 42217
rect 9042 42208 9054 42211
rect 8168 42180 9054 42208
rect 8168 42168 8174 42180
rect 9042 42177 9054 42180
rect 9088 42177 9100 42211
rect 9042 42171 9100 42177
rect 5258 42100 5264 42152
rect 5316 42140 5322 42152
rect 8294 42140 8300 42152
rect 5316 42112 8300 42140
rect 5316 42100 5322 42112
rect 8294 42100 8300 42112
rect 8352 42100 8358 42152
rect 9306 42140 9312 42152
rect 9267 42112 9312 42140
rect 9306 42100 9312 42112
rect 9364 42100 9370 42152
rect 4062 42032 4068 42084
rect 4120 42072 4126 42084
rect 4617 42075 4675 42081
rect 4617 42072 4629 42075
rect 4120 42044 4629 42072
rect 4120 42032 4126 42044
rect 4617 42041 4629 42044
rect 4663 42041 4675 42075
rect 4617 42035 4675 42041
rect 1486 42004 1492 42016
rect 1447 41976 1492 42004
rect 1486 41964 1492 41976
rect 1544 41964 1550 42016
rect 2038 41964 2044 42016
rect 2096 42004 2102 42016
rect 2133 42007 2191 42013
rect 2133 42004 2145 42007
rect 2096 41976 2145 42004
rect 2096 41964 2102 41976
rect 2133 41973 2145 41976
rect 2179 41973 2191 42007
rect 2133 41967 2191 41973
rect 3694 41964 3700 42016
rect 3752 42004 3758 42016
rect 4157 42007 4215 42013
rect 4157 42004 4169 42007
rect 3752 41976 4169 42004
rect 3752 41964 3758 41976
rect 4157 41973 4169 41976
rect 4203 41973 4215 42007
rect 4157 41967 4215 41973
rect 5350 41964 5356 42016
rect 5408 42004 5414 42016
rect 5445 42007 5503 42013
rect 5445 42004 5457 42007
rect 5408 41976 5457 42004
rect 5408 41964 5414 41976
rect 5445 41973 5457 41976
rect 5491 41973 5503 42007
rect 5445 41967 5503 41973
rect 1104 41914 30820 41936
rect 1104 41862 5915 41914
rect 5967 41862 5979 41914
rect 6031 41862 6043 41914
rect 6095 41862 6107 41914
rect 6159 41862 6171 41914
rect 6223 41862 15846 41914
rect 15898 41862 15910 41914
rect 15962 41862 15974 41914
rect 16026 41862 16038 41914
rect 16090 41862 16102 41914
rect 16154 41862 25776 41914
rect 25828 41862 25840 41914
rect 25892 41862 25904 41914
rect 25956 41862 25968 41914
rect 26020 41862 26032 41914
rect 26084 41862 30820 41914
rect 1104 41840 30820 41862
rect 2866 41800 2872 41812
rect 2827 41772 2872 41800
rect 2866 41760 2872 41772
rect 2924 41760 2930 41812
rect 4430 41800 4436 41812
rect 4391 41772 4436 41800
rect 4430 41760 4436 41772
rect 4488 41760 4494 41812
rect 5626 41800 5632 41812
rect 5587 41772 5632 41800
rect 5626 41760 5632 41772
rect 5684 41760 5690 41812
rect 5813 41803 5871 41809
rect 5813 41769 5825 41803
rect 5859 41769 5871 41803
rect 8110 41800 8116 41812
rect 8071 41772 8116 41800
rect 5813 41763 5871 41769
rect 5350 41692 5356 41744
rect 5408 41732 5414 41744
rect 5828 41732 5856 41763
rect 8110 41760 8116 41772
rect 8168 41760 8174 41812
rect 9125 41803 9183 41809
rect 9125 41769 9137 41803
rect 9171 41800 9183 41803
rect 9306 41800 9312 41812
rect 9171 41772 9312 41800
rect 9171 41769 9183 41772
rect 9125 41763 9183 41769
rect 9306 41760 9312 41772
rect 9364 41760 9370 41812
rect 5408 41704 5856 41732
rect 6181 41735 6239 41741
rect 5408 41692 5414 41704
rect 6181 41701 6193 41735
rect 6227 41732 6239 41735
rect 6270 41732 6276 41744
rect 6227 41704 6276 41732
rect 6227 41701 6239 41704
rect 6181 41695 6239 41701
rect 6270 41692 6276 41704
rect 6328 41692 6334 41744
rect 6917 41735 6975 41741
rect 6917 41701 6929 41735
rect 6963 41701 6975 41735
rect 6917 41695 6975 41701
rect 4338 41624 4344 41676
rect 4396 41664 4402 41676
rect 4893 41667 4951 41673
rect 4893 41664 4905 41667
rect 4396 41636 4905 41664
rect 4396 41624 4402 41636
rect 4893 41633 4905 41636
rect 4939 41633 4951 41667
rect 5258 41664 5264 41676
rect 4893 41627 4951 41633
rect 5000 41636 5264 41664
rect 1762 41556 1768 41608
rect 1820 41596 1826 41608
rect 1857 41599 1915 41605
rect 1857 41596 1869 41599
rect 1820 41568 1869 41596
rect 1820 41556 1826 41568
rect 1857 41565 1869 41568
rect 1903 41565 1915 41599
rect 1857 41559 1915 41565
rect 2774 41556 2780 41608
rect 2832 41596 2838 41608
rect 3053 41599 3111 41605
rect 3053 41596 3065 41599
rect 2832 41568 3065 41596
rect 2832 41556 2838 41568
rect 3053 41565 3065 41568
rect 3099 41596 3111 41599
rect 3878 41596 3884 41608
rect 3099 41568 3884 41596
rect 3099 41565 3111 41568
rect 3053 41559 3111 41565
rect 3878 41556 3884 41568
rect 3936 41556 3942 41608
rect 3973 41599 4031 41605
rect 3973 41565 3985 41599
rect 4019 41596 4031 41599
rect 4430 41596 4436 41608
rect 4019 41568 4436 41596
rect 4019 41565 4031 41568
rect 3973 41559 4031 41565
rect 4430 41556 4436 41568
rect 4488 41556 4494 41608
rect 4617 41599 4675 41605
rect 4617 41565 4629 41599
rect 4663 41565 4675 41599
rect 4617 41559 4675 41565
rect 4632 41528 4660 41559
rect 4706 41556 4712 41608
rect 4764 41596 4770 41608
rect 5000 41605 5028 41636
rect 5258 41624 5264 41636
rect 5316 41624 5322 41676
rect 6932 41664 6960 41695
rect 7006 41692 7012 41744
rect 7064 41732 7070 41744
rect 7650 41732 7656 41744
rect 7064 41704 7656 41732
rect 7064 41692 7070 41704
rect 7650 41692 7656 41704
rect 7708 41732 7714 41744
rect 10226 41732 10232 41744
rect 7708 41704 10232 41732
rect 7708 41692 7714 41704
rect 10226 41692 10232 41704
rect 10284 41732 10290 41744
rect 10284 41704 16574 41732
rect 10284 41692 10290 41704
rect 16546 41664 16574 41704
rect 21361 41667 21419 41673
rect 21361 41664 21373 41667
rect 6932 41636 8984 41664
rect 16546 41636 21373 41664
rect 4801 41599 4859 41605
rect 4801 41596 4813 41599
rect 4764 41568 4813 41596
rect 4764 41556 4770 41568
rect 4801 41565 4813 41568
rect 4847 41565 4859 41599
rect 4801 41559 4859 41565
rect 4985 41599 5043 41605
rect 4985 41565 4997 41599
rect 5031 41565 5043 41599
rect 5166 41596 5172 41608
rect 5127 41568 5172 41596
rect 4985 41559 5043 41565
rect 5166 41556 5172 41568
rect 5224 41556 5230 41608
rect 6638 41556 6644 41608
rect 6696 41596 6702 41608
rect 6733 41599 6791 41605
rect 6733 41596 6745 41599
rect 6696 41568 6745 41596
rect 6696 41556 6702 41568
rect 6733 41565 6745 41568
rect 6779 41565 6791 41599
rect 7377 41599 7435 41605
rect 7377 41596 7389 41599
rect 6733 41559 6791 41565
rect 6886 41568 7389 41596
rect 5810 41528 5816 41540
rect 4632 41500 5816 41528
rect 5810 41488 5816 41500
rect 5868 41488 5874 41540
rect 6362 41488 6368 41540
rect 6420 41528 6426 41540
rect 6886 41528 6914 41568
rect 7377 41565 7389 41568
rect 7423 41565 7435 41599
rect 7377 41559 7435 41565
rect 7561 41599 7619 41605
rect 7561 41565 7573 41599
rect 7607 41565 7619 41599
rect 7561 41559 7619 41565
rect 7653 41599 7711 41605
rect 7653 41565 7665 41599
rect 7699 41565 7711 41599
rect 7653 41559 7711 41565
rect 6420 41500 6914 41528
rect 6420 41488 6426 41500
rect 1670 41460 1676 41472
rect 1631 41432 1676 41460
rect 1670 41420 1676 41432
rect 1728 41420 1734 41472
rect 2958 41420 2964 41472
rect 3016 41460 3022 41472
rect 3789 41463 3847 41469
rect 3789 41460 3801 41463
rect 3016 41432 3801 41460
rect 3016 41420 3022 41432
rect 3789 41429 3801 41432
rect 3835 41429 3847 41463
rect 3789 41423 3847 41429
rect 7466 41420 7472 41472
rect 7524 41460 7530 41472
rect 7576 41460 7604 41559
rect 7668 41528 7696 41559
rect 7742 41556 7748 41608
rect 7800 41596 7806 41608
rect 7926 41596 7932 41608
rect 7800 41568 7845 41596
rect 7887 41568 7932 41596
rect 7800 41556 7806 41568
rect 7926 41556 7932 41568
rect 7984 41556 7990 41608
rect 8956 41605 8984 41636
rect 21361 41633 21373 41636
rect 21407 41633 21419 41667
rect 21361 41627 21419 41633
rect 8941 41599 8999 41605
rect 8941 41565 8953 41599
rect 8987 41565 8999 41599
rect 12986 41596 12992 41608
rect 12947 41568 12992 41596
rect 8941 41559 8999 41565
rect 12986 41556 12992 41568
rect 13044 41556 13050 41608
rect 15746 41556 15752 41608
rect 15804 41596 15810 41608
rect 15933 41599 15991 41605
rect 15933 41596 15945 41599
rect 15804 41568 15945 41596
rect 15804 41556 15810 41568
rect 15933 41565 15945 41568
rect 15979 41565 15991 41599
rect 15933 41559 15991 41565
rect 21821 41599 21879 41605
rect 21821 41565 21833 41599
rect 21867 41565 21879 41599
rect 21821 41559 21879 41565
rect 21913 41599 21971 41605
rect 21913 41565 21925 41599
rect 21959 41596 21971 41599
rect 29914 41596 29920 41608
rect 21959 41568 29920 41596
rect 21959 41565 21971 41568
rect 21913 41559 21971 41565
rect 7834 41528 7840 41540
rect 7668 41500 7840 41528
rect 7834 41488 7840 41500
rect 7892 41488 7898 41540
rect 10134 41528 10140 41540
rect 7944 41500 10140 41528
rect 7944 41460 7972 41500
rect 10134 41488 10140 41500
rect 10192 41528 10198 41540
rect 21836 41528 21864 41559
rect 29914 41556 29920 41568
rect 29972 41556 29978 41608
rect 22002 41528 22008 41540
rect 10192 41500 16574 41528
rect 21836 41500 22008 41528
rect 10192 41488 10198 41500
rect 7524 41432 7972 41460
rect 7524 41420 7530 41432
rect 12618 41420 12624 41472
rect 12676 41460 12682 41472
rect 12805 41463 12863 41469
rect 12805 41460 12817 41463
rect 12676 41432 12817 41460
rect 12676 41420 12682 41432
rect 12805 41429 12817 41432
rect 12851 41429 12863 41463
rect 12805 41423 12863 41429
rect 16117 41463 16175 41469
rect 16117 41429 16129 41463
rect 16163 41460 16175 41463
rect 16298 41460 16304 41472
rect 16163 41432 16304 41460
rect 16163 41429 16175 41432
rect 16117 41423 16175 41429
rect 16298 41420 16304 41432
rect 16356 41420 16362 41472
rect 16546 41460 16574 41500
rect 22002 41488 22008 41500
rect 22060 41488 22066 41540
rect 21910 41460 21916 41472
rect 16546 41432 21916 41460
rect 21910 41420 21916 41432
rect 21968 41420 21974 41472
rect 1104 41370 30820 41392
rect 1104 41318 10880 41370
rect 10932 41318 10944 41370
rect 10996 41318 11008 41370
rect 11060 41318 11072 41370
rect 11124 41318 11136 41370
rect 11188 41318 20811 41370
rect 20863 41318 20875 41370
rect 20927 41318 20939 41370
rect 20991 41318 21003 41370
rect 21055 41318 21067 41370
rect 21119 41318 30820 41370
rect 1104 41296 30820 41318
rect 2314 41216 2320 41268
rect 2372 41256 2378 41268
rect 2409 41259 2467 41265
rect 2409 41256 2421 41259
rect 2372 41228 2421 41256
rect 2372 41216 2378 41228
rect 2409 41225 2421 41228
rect 2455 41225 2467 41259
rect 3418 41256 3424 41268
rect 3379 41228 3424 41256
rect 2409 41219 2467 41225
rect 3418 41216 3424 41228
rect 3476 41216 3482 41268
rect 3970 41216 3976 41268
rect 4028 41256 4034 41268
rect 5261 41259 5319 41265
rect 5261 41256 5273 41259
rect 4028 41228 5273 41256
rect 4028 41216 4034 41228
rect 5261 41225 5273 41228
rect 5307 41225 5319 41259
rect 6546 41256 6552 41268
rect 6507 41228 6552 41256
rect 5261 41219 5319 41225
rect 6546 41216 6552 41228
rect 6604 41216 6610 41268
rect 21910 41256 21916 41268
rect 21871 41228 21916 41256
rect 21910 41216 21916 41228
rect 21968 41216 21974 41268
rect 2593 41191 2651 41197
rect 2593 41157 2605 41191
rect 2639 41157 2651 41191
rect 5166 41188 5172 41200
rect 2593 41151 2651 41157
rect 4448 41160 5172 41188
rect 1673 41123 1731 41129
rect 1673 41089 1685 41123
rect 1719 41089 1731 41123
rect 2608 41120 2636 41151
rect 4448 41132 4476 41160
rect 5166 41148 5172 41160
rect 5224 41148 5230 41200
rect 5445 41191 5503 41197
rect 5445 41157 5457 41191
rect 5491 41188 5503 41191
rect 6362 41188 6368 41200
rect 5491 41160 6368 41188
rect 5491 41157 5503 41160
rect 5445 41151 5503 41157
rect 6362 41148 6368 41160
rect 6420 41148 6426 41200
rect 6914 41148 6920 41200
rect 6972 41188 6978 41200
rect 7558 41188 7564 41200
rect 6972 41160 7564 41188
rect 6972 41148 6978 41160
rect 7558 41148 7564 41160
rect 7616 41148 7622 41200
rect 3605 41123 3663 41129
rect 3605 41120 3617 41123
rect 2608 41092 3617 41120
rect 1673 41083 1731 41089
rect 3605 41089 3617 41092
rect 3651 41120 3663 41123
rect 3694 41120 3700 41132
rect 3651 41092 3700 41120
rect 3651 41089 3663 41092
rect 3605 41083 3663 41089
rect 1688 41052 1716 41083
rect 3694 41080 3700 41092
rect 3752 41080 3758 41132
rect 3970 41120 3976 41132
rect 3931 41092 3976 41120
rect 3970 41080 3976 41092
rect 4028 41080 4034 41132
rect 4157 41123 4215 41129
rect 4157 41089 4169 41123
rect 4203 41120 4215 41123
rect 4430 41120 4436 41132
rect 4203 41092 4436 41120
rect 4203 41089 4215 41092
rect 4157 41083 4215 41089
rect 4430 41080 4436 41092
rect 4488 41080 4494 41132
rect 4617 41123 4675 41129
rect 4617 41089 4629 41123
rect 4663 41120 4675 41123
rect 5810 41120 5816 41132
rect 4663 41092 5816 41120
rect 4663 41089 4675 41092
rect 4617 41083 4675 41089
rect 5810 41080 5816 41092
rect 5868 41120 5874 41132
rect 6638 41120 6644 41132
rect 5868 41092 6644 41120
rect 5868 41080 5874 41092
rect 6638 41080 6644 41092
rect 6696 41080 6702 41132
rect 6730 41080 6736 41132
rect 6788 41120 6794 41132
rect 7662 41123 7720 41129
rect 7662 41120 7674 41123
rect 6788 41092 7674 41120
rect 6788 41080 6794 41092
rect 7662 41089 7674 41092
rect 7708 41089 7720 41123
rect 7662 41083 7720 41089
rect 7834 41080 7840 41132
rect 7892 41120 7898 41132
rect 8665 41123 8723 41129
rect 8665 41120 8677 41123
rect 7892 41092 8677 41120
rect 7892 41080 7898 41092
rect 8665 41089 8677 41092
rect 8711 41089 8723 41123
rect 8665 41083 8723 41089
rect 14458 41080 14464 41132
rect 14516 41120 14522 41132
rect 15013 41123 15071 41129
rect 15013 41120 15025 41123
rect 14516 41092 15025 41120
rect 14516 41080 14522 41092
rect 15013 41089 15025 41092
rect 15059 41089 15071 41123
rect 15013 41083 15071 41089
rect 15105 41123 15163 41129
rect 15105 41089 15117 41123
rect 15151 41120 15163 41123
rect 15562 41120 15568 41132
rect 15151 41092 15568 41120
rect 15151 41089 15163 41092
rect 15105 41083 15163 41089
rect 15562 41080 15568 41092
rect 15620 41120 15626 41132
rect 15657 41123 15715 41129
rect 15657 41120 15669 41123
rect 15620 41092 15669 41120
rect 15620 41080 15626 41092
rect 15657 41089 15669 41092
rect 15703 41089 15715 41123
rect 15657 41083 15715 41089
rect 15841 41123 15899 41129
rect 15841 41089 15853 41123
rect 15887 41089 15899 41123
rect 15841 41083 15899 41089
rect 3234 41052 3240 41064
rect 1688 41024 3240 41052
rect 3234 41012 3240 41024
rect 3292 41012 3298 41064
rect 3789 41055 3847 41061
rect 3789 41021 3801 41055
rect 3835 41021 3847 41055
rect 3789 41015 3847 41021
rect 3881 41055 3939 41061
rect 3881 41021 3893 41055
rect 3927 41052 3939 41055
rect 4246 41052 4252 41064
rect 3927 41024 4252 41052
rect 3927 41021 3939 41024
rect 3881 41015 3939 41021
rect 2958 40984 2964 40996
rect 2919 40956 2964 40984
rect 2958 40944 2964 40956
rect 3016 40944 3022 40996
rect 3804 40984 3832 41015
rect 4246 41012 4252 41024
rect 4304 41012 4310 41064
rect 4706 41052 4712 41064
rect 4540 41024 4712 41052
rect 4154 40984 4160 40996
rect 3804 40956 4160 40984
rect 4154 40944 4160 40956
rect 4212 40984 4218 40996
rect 4540 40984 4568 41024
rect 4706 41012 4712 41024
rect 4764 41012 4770 41064
rect 5442 41012 5448 41064
rect 5500 41052 5506 41064
rect 6914 41052 6920 41064
rect 5500 41024 6920 41052
rect 5500 41012 5506 41024
rect 6914 41012 6920 41024
rect 6972 41012 6978 41064
rect 7926 41052 7932 41064
rect 7887 41024 7932 41052
rect 7926 41012 7932 41024
rect 7984 41012 7990 41064
rect 8389 41055 8447 41061
rect 8389 41021 8401 41055
rect 8435 41021 8447 41055
rect 12618 41052 12624 41064
rect 12579 41024 12624 41052
rect 8389 41015 8447 41021
rect 5350 40984 5356 40996
rect 4212 40956 4568 40984
rect 4632 40956 5356 40984
rect 4212 40944 4218 40956
rect 1486 40916 1492 40928
rect 1447 40888 1492 40916
rect 1486 40876 1492 40888
rect 1544 40876 1550 40928
rect 2593 40919 2651 40925
rect 2593 40885 2605 40919
rect 2639 40916 2651 40919
rect 4632 40916 4660 40956
rect 5350 40944 5356 40956
rect 5408 40984 5414 40996
rect 5408 40956 5488 40984
rect 5408 40944 5414 40956
rect 4798 40916 4804 40928
rect 2639 40888 4660 40916
rect 4759 40888 4804 40916
rect 2639 40885 2651 40888
rect 2593 40879 2651 40885
rect 4798 40876 4804 40888
rect 4856 40876 4862 40928
rect 5460 40925 5488 40956
rect 5718 40944 5724 40996
rect 5776 40984 5782 40996
rect 5813 40987 5871 40993
rect 5813 40984 5825 40987
rect 5776 40956 5825 40984
rect 5776 40944 5782 40956
rect 5813 40953 5825 40956
rect 5859 40984 5871 40987
rect 6270 40984 6276 40996
rect 5859 40956 6276 40984
rect 5859 40953 5871 40956
rect 5813 40947 5871 40953
rect 6270 40944 6276 40956
rect 6328 40984 6334 40996
rect 6822 40984 6828 40996
rect 6328 40956 6828 40984
rect 6328 40944 6334 40956
rect 6822 40944 6828 40956
rect 6880 40944 6886 40996
rect 5445 40919 5503 40925
rect 5445 40885 5457 40919
rect 5491 40885 5503 40919
rect 5445 40879 5503 40885
rect 7190 40876 7196 40928
rect 7248 40916 7254 40928
rect 8404 40916 8432 41015
rect 12618 41012 12624 41024
rect 12676 41012 12682 41064
rect 12805 41055 12863 41061
rect 12805 41021 12817 41055
rect 12851 41052 12863 41055
rect 12894 41052 12900 41064
rect 12851 41024 12900 41052
rect 12851 41021 12863 41024
rect 12805 41015 12863 41021
rect 12894 41012 12900 41024
rect 12952 41012 12958 41064
rect 13538 41052 13544 41064
rect 13499 41024 13544 41052
rect 13538 41012 13544 41024
rect 13596 41012 13602 41064
rect 13722 41061 13728 41064
rect 13679 41055 13728 41061
rect 13679 41021 13691 41055
rect 13725 41021 13728 41055
rect 13679 41015 13728 41021
rect 13722 41012 13728 41015
rect 13780 41012 13786 41064
rect 13817 41055 13875 41061
rect 13817 41021 13829 41055
rect 13863 41052 13875 41055
rect 13998 41052 14004 41064
rect 13863 41024 14004 41052
rect 13863 41021 13875 41024
rect 13817 41015 13875 41021
rect 13998 41012 14004 41024
rect 14056 41012 14062 41064
rect 13265 40987 13323 40993
rect 13265 40953 13277 40987
rect 13311 40953 13323 40987
rect 14918 40984 14924 40996
rect 13265 40947 13323 40953
rect 14200 40956 14924 40984
rect 7248 40888 8432 40916
rect 13280 40916 13308 40947
rect 14200 40916 14228 40956
rect 14918 40944 14924 40956
rect 14976 40984 14982 40996
rect 15856 40984 15884 41083
rect 16298 41080 16304 41132
rect 16356 41120 16362 41132
rect 16669 41123 16727 41129
rect 16669 41120 16681 41123
rect 16356 41092 16681 41120
rect 16356 41080 16362 41092
rect 16669 41089 16681 41092
rect 16715 41089 16727 41123
rect 17402 41120 17408 41132
rect 17363 41092 17408 41120
rect 16669 41083 16727 41089
rect 17402 41080 17408 41092
rect 17460 41080 17466 41132
rect 22002 41080 22008 41132
rect 22060 41120 22066 41132
rect 22097 41123 22155 41129
rect 22097 41120 22109 41123
rect 22060 41092 22109 41120
rect 22060 41080 22066 41092
rect 22097 41089 22109 41092
rect 22143 41089 22155 41123
rect 30098 41120 30104 41132
rect 30059 41092 30104 41120
rect 22097 41083 22155 41089
rect 30098 41080 30104 41092
rect 30156 41080 30162 41132
rect 22281 41055 22339 41061
rect 22281 41021 22293 41055
rect 22327 41052 22339 41055
rect 22327 41024 26234 41052
rect 22327 41021 22339 41024
rect 22281 41015 22339 41021
rect 14976 40956 15884 40984
rect 26206 40984 26234 41024
rect 29917 40987 29975 40993
rect 29917 40984 29929 40987
rect 26206 40956 29929 40984
rect 14976 40944 14982 40956
rect 29917 40953 29929 40956
rect 29963 40953 29975 40987
rect 29917 40947 29975 40953
rect 13280 40888 14228 40916
rect 14461 40919 14519 40925
rect 7248 40876 7254 40888
rect 14461 40885 14473 40919
rect 14507 40916 14519 40919
rect 14734 40916 14740 40928
rect 14507 40888 14740 40916
rect 14507 40885 14519 40888
rect 14461 40879 14519 40885
rect 14734 40876 14740 40888
rect 14792 40876 14798 40928
rect 16025 40919 16083 40925
rect 16025 40885 16037 40919
rect 16071 40916 16083 40919
rect 16482 40916 16488 40928
rect 16071 40888 16488 40916
rect 16071 40885 16083 40888
rect 16025 40879 16083 40885
rect 16482 40876 16488 40888
rect 16540 40876 16546 40928
rect 16666 40916 16672 40928
rect 16627 40888 16672 40916
rect 16666 40876 16672 40888
rect 16724 40876 16730 40928
rect 17034 40876 17040 40928
rect 17092 40916 17098 40928
rect 17405 40919 17463 40925
rect 17405 40916 17417 40919
rect 17092 40888 17417 40916
rect 17092 40876 17098 40888
rect 17405 40885 17417 40888
rect 17451 40885 17463 40919
rect 17405 40879 17463 40885
rect 1104 40826 30820 40848
rect 1104 40774 5915 40826
rect 5967 40774 5979 40826
rect 6031 40774 6043 40826
rect 6095 40774 6107 40826
rect 6159 40774 6171 40826
rect 6223 40774 15846 40826
rect 15898 40774 15910 40826
rect 15962 40774 15974 40826
rect 16026 40774 16038 40826
rect 16090 40774 16102 40826
rect 16154 40774 25776 40826
rect 25828 40774 25840 40826
rect 25892 40774 25904 40826
rect 25956 40774 25968 40826
rect 26020 40774 26032 40826
rect 26084 40774 30820 40826
rect 1104 40752 30820 40774
rect 3970 40672 3976 40724
rect 4028 40712 4034 40724
rect 6641 40715 6699 40721
rect 4028 40684 6592 40712
rect 4028 40672 4034 40684
rect 2222 40604 2228 40656
rect 2280 40644 2286 40656
rect 4985 40647 5043 40653
rect 4985 40644 4997 40647
rect 2280 40616 4997 40644
rect 2280 40604 2286 40616
rect 4985 40613 4997 40616
rect 5031 40613 5043 40647
rect 6454 40644 6460 40656
rect 4985 40607 5043 40613
rect 5920 40616 6460 40644
rect 4246 40576 4252 40588
rect 4207 40548 4252 40576
rect 4246 40536 4252 40548
rect 4304 40536 4310 40588
rect 1673 40511 1731 40517
rect 1673 40477 1685 40511
rect 1719 40508 1731 40511
rect 1946 40508 1952 40520
rect 1719 40480 1952 40508
rect 1719 40477 1731 40480
rect 1673 40471 1731 40477
rect 1946 40468 1952 40480
rect 2004 40468 2010 40520
rect 2593 40511 2651 40517
rect 2593 40477 2605 40511
rect 2639 40508 2651 40511
rect 2774 40508 2780 40520
rect 2639 40480 2780 40508
rect 2639 40477 2651 40480
rect 2593 40471 2651 40477
rect 2774 40468 2780 40480
rect 2832 40468 2838 40520
rect 3970 40508 3976 40520
rect 3931 40480 3976 40508
rect 3970 40468 3976 40480
rect 4028 40468 4034 40520
rect 4154 40508 4160 40520
rect 4115 40480 4160 40508
rect 4154 40468 4160 40480
rect 4212 40468 4218 40520
rect 4341 40511 4399 40517
rect 4341 40477 4353 40511
rect 4387 40477 4399 40511
rect 4341 40471 4399 40477
rect 4356 40440 4384 40471
rect 4430 40468 4436 40520
rect 4488 40508 4494 40520
rect 4525 40511 4583 40517
rect 4525 40508 4537 40511
rect 4488 40480 4537 40508
rect 4488 40468 4494 40480
rect 4525 40477 4537 40480
rect 4571 40508 4583 40511
rect 4614 40508 4620 40520
rect 4571 40480 4620 40508
rect 4571 40477 4583 40480
rect 4525 40471 4583 40477
rect 4614 40468 4620 40480
rect 4672 40468 4678 40520
rect 5074 40468 5080 40520
rect 5132 40508 5138 40520
rect 5920 40517 5948 40616
rect 6454 40604 6460 40616
rect 6512 40604 6518 40656
rect 6564 40644 6592 40684
rect 6641 40681 6653 40715
rect 6687 40712 6699 40715
rect 6730 40712 6736 40724
rect 6687 40684 6736 40712
rect 6687 40681 6699 40684
rect 6641 40675 6699 40681
rect 6730 40672 6736 40684
rect 6788 40672 6794 40724
rect 6822 40672 6828 40724
rect 6880 40712 6886 40724
rect 9585 40715 9643 40721
rect 9585 40712 9597 40715
rect 6880 40684 9597 40712
rect 6880 40672 6886 40684
rect 9585 40681 9597 40684
rect 9631 40681 9643 40715
rect 9585 40675 9643 40681
rect 12529 40715 12587 40721
rect 12529 40681 12541 40715
rect 12575 40712 12587 40715
rect 12986 40712 12992 40724
rect 12575 40684 12992 40712
rect 12575 40681 12587 40684
rect 12529 40675 12587 40681
rect 12986 40672 12992 40684
rect 13044 40672 13050 40724
rect 17310 40712 17316 40724
rect 16868 40684 17316 40712
rect 16868 40656 16896 40684
rect 17310 40672 17316 40684
rect 17368 40672 17374 40724
rect 7282 40644 7288 40656
rect 6564 40616 7288 40644
rect 7282 40604 7288 40616
rect 7340 40604 7346 40656
rect 16850 40644 16856 40656
rect 14568 40616 16856 40644
rect 6273 40579 6331 40585
rect 6273 40545 6285 40579
rect 6319 40576 6331 40579
rect 7377 40579 7435 40585
rect 6319 40548 6960 40576
rect 6319 40545 6331 40548
rect 6273 40539 6331 40545
rect 6932 40520 6960 40548
rect 7377 40545 7389 40579
rect 7423 40576 7435 40579
rect 7742 40576 7748 40588
rect 7423 40548 7748 40576
rect 7423 40545 7435 40548
rect 7377 40539 7435 40545
rect 7742 40536 7748 40548
rect 7800 40536 7806 40588
rect 13538 40576 13544 40588
rect 12360 40548 13544 40576
rect 5169 40511 5227 40517
rect 5169 40508 5181 40511
rect 5132 40480 5181 40508
rect 5132 40468 5138 40480
rect 5169 40477 5181 40480
rect 5215 40477 5227 40511
rect 5169 40471 5227 40477
rect 5905 40511 5963 40517
rect 5905 40477 5917 40511
rect 5951 40477 5963 40511
rect 5905 40471 5963 40477
rect 6089 40511 6147 40517
rect 6089 40477 6101 40511
rect 6135 40477 6147 40511
rect 6089 40471 6147 40477
rect 6181 40511 6239 40517
rect 6181 40477 6193 40511
rect 6227 40477 6239 40511
rect 6181 40471 6239 40477
rect 6457 40511 6515 40517
rect 6457 40477 6469 40511
rect 6503 40508 6515 40511
rect 6546 40508 6552 40520
rect 6503 40480 6552 40508
rect 6503 40477 6515 40480
rect 6457 40471 6515 40477
rect 5442 40440 5448 40452
rect 4356 40412 5448 40440
rect 5442 40400 5448 40412
rect 5500 40400 5506 40452
rect 1486 40372 1492 40384
rect 1447 40344 1492 40372
rect 1486 40332 1492 40344
rect 1544 40332 1550 40384
rect 2777 40375 2835 40381
rect 2777 40341 2789 40375
rect 2823 40372 2835 40375
rect 3050 40372 3056 40384
rect 2823 40344 3056 40372
rect 2823 40341 2835 40344
rect 2777 40335 2835 40341
rect 3050 40332 3056 40344
rect 3108 40332 3114 40384
rect 3786 40372 3792 40384
rect 3747 40344 3792 40372
rect 3786 40332 3792 40344
rect 3844 40332 3850 40384
rect 6104 40372 6132 40471
rect 6196 40440 6224 40471
rect 6546 40468 6552 40480
rect 6604 40468 6610 40520
rect 6914 40468 6920 40520
rect 6972 40508 6978 40520
rect 7101 40511 7159 40517
rect 7101 40508 7113 40511
rect 6972 40480 7113 40508
rect 6972 40468 6978 40480
rect 7101 40477 7113 40480
rect 7147 40477 7159 40511
rect 7101 40471 7159 40477
rect 8570 40468 8576 40520
rect 8628 40508 8634 40520
rect 8941 40511 8999 40517
rect 8941 40508 8953 40511
rect 8628 40480 8953 40508
rect 8628 40468 8634 40480
rect 8941 40477 8953 40480
rect 8987 40477 8999 40511
rect 9766 40508 9772 40520
rect 9727 40480 9772 40508
rect 8941 40471 8999 40477
rect 9766 40468 9772 40480
rect 9824 40468 9830 40520
rect 12360 40517 12388 40548
rect 13538 40536 13544 40548
rect 13596 40536 13602 40588
rect 14568 40585 14596 40616
rect 16850 40604 16856 40616
rect 16908 40604 16914 40656
rect 14553 40579 14611 40585
rect 14553 40545 14565 40579
rect 14599 40545 14611 40579
rect 14734 40576 14740 40588
rect 14695 40548 14740 40576
rect 14553 40539 14611 40545
rect 14734 40536 14740 40548
rect 14792 40536 14798 40588
rect 16117 40579 16175 40585
rect 16117 40545 16129 40579
rect 16163 40576 16175 40579
rect 16666 40576 16672 40588
rect 16163 40548 16672 40576
rect 16163 40545 16175 40548
rect 16117 40539 16175 40545
rect 16666 40536 16672 40548
rect 16724 40536 16730 40588
rect 16758 40536 16764 40588
rect 16816 40576 16822 40588
rect 17034 40576 17040 40588
rect 16816 40548 16861 40576
rect 16995 40548 17040 40576
rect 16816 40536 16822 40548
rect 17034 40536 17040 40548
rect 17092 40536 17098 40588
rect 17175 40579 17233 40585
rect 17175 40545 17187 40579
rect 17221 40576 17233 40579
rect 17494 40576 17500 40588
rect 17221 40548 17500 40576
rect 17221 40545 17233 40548
rect 17175 40539 17233 40545
rect 17494 40536 17500 40548
rect 17552 40536 17558 40588
rect 12345 40511 12403 40517
rect 12345 40477 12357 40511
rect 12391 40477 12403 40511
rect 12986 40508 12992 40520
rect 12947 40480 12992 40508
rect 12345 40471 12403 40477
rect 12986 40468 12992 40480
rect 13044 40468 13050 40520
rect 16298 40508 16304 40520
rect 16259 40480 16304 40508
rect 16298 40468 16304 40480
rect 16356 40468 16362 40520
rect 17310 40508 17316 40520
rect 17271 40480 17316 40508
rect 17310 40468 17316 40480
rect 17368 40468 17374 40520
rect 18598 40508 18604 40520
rect 18559 40480 18604 40508
rect 18598 40468 18604 40480
rect 18656 40468 18662 40520
rect 6730 40440 6736 40452
rect 6196 40412 6736 40440
rect 6730 40400 6736 40412
rect 6788 40400 6794 40452
rect 19794 40440 19800 40452
rect 17788 40412 19800 40440
rect 8938 40372 8944 40384
rect 6104 40344 8944 40372
rect 8938 40332 8944 40344
rect 8996 40332 9002 40384
rect 9122 40372 9128 40384
rect 9083 40344 9128 40372
rect 9122 40332 9128 40344
rect 9180 40332 9186 40384
rect 13173 40375 13231 40381
rect 13173 40341 13185 40375
rect 13219 40372 13231 40375
rect 13814 40372 13820 40384
rect 13219 40344 13820 40372
rect 13219 40341 13231 40344
rect 13173 40335 13231 40341
rect 13814 40332 13820 40344
rect 13872 40332 13878 40384
rect 14826 40332 14832 40384
rect 14884 40372 14890 40384
rect 15197 40375 15255 40381
rect 14884 40344 14929 40372
rect 14884 40332 14890 40344
rect 15197 40341 15209 40375
rect 15243 40372 15255 40375
rect 17788 40372 17816 40412
rect 19794 40400 19800 40412
rect 19852 40400 19858 40452
rect 17954 40372 17960 40384
rect 15243 40344 17816 40372
rect 17915 40344 17960 40372
rect 15243 40341 15255 40344
rect 15197 40335 15255 40341
rect 17954 40332 17960 40344
rect 18012 40332 18018 40384
rect 18414 40372 18420 40384
rect 18375 40344 18420 40372
rect 18414 40332 18420 40344
rect 18472 40332 18478 40384
rect 1104 40282 30820 40304
rect 1104 40230 10880 40282
rect 10932 40230 10944 40282
rect 10996 40230 11008 40282
rect 11060 40230 11072 40282
rect 11124 40230 11136 40282
rect 11188 40230 20811 40282
rect 20863 40230 20875 40282
rect 20927 40230 20939 40282
rect 20991 40230 21003 40282
rect 21055 40230 21067 40282
rect 21119 40230 30820 40282
rect 1104 40208 30820 40230
rect 2225 40171 2283 40177
rect 2225 40137 2237 40171
rect 2271 40168 2283 40171
rect 3970 40168 3976 40180
rect 2271 40140 3976 40168
rect 2271 40137 2283 40140
rect 2225 40131 2283 40137
rect 3970 40128 3976 40140
rect 4028 40168 4034 40180
rect 4249 40171 4307 40177
rect 4249 40168 4261 40171
rect 4028 40140 4261 40168
rect 4028 40128 4034 40140
rect 4249 40137 4261 40140
rect 4295 40137 4307 40171
rect 4249 40131 4307 40137
rect 4798 40128 4804 40180
rect 4856 40168 4862 40180
rect 7653 40171 7711 40177
rect 4856 40140 7420 40168
rect 4856 40128 4862 40140
rect 3136 40103 3194 40109
rect 3136 40069 3148 40103
rect 3182 40100 3194 40103
rect 3786 40100 3792 40112
rect 3182 40072 3792 40100
rect 3182 40069 3194 40072
rect 3136 40063 3194 40069
rect 3786 40060 3792 40072
rect 3844 40060 3850 40112
rect 5445 40103 5503 40109
rect 5445 40069 5457 40103
rect 5491 40100 5503 40103
rect 7282 40100 7288 40112
rect 5491 40072 7288 40100
rect 5491 40069 5503 40072
rect 5445 40063 5503 40069
rect 7282 40060 7288 40072
rect 7340 40060 7346 40112
rect 7392 40100 7420 40140
rect 7653 40137 7665 40171
rect 7699 40168 7711 40171
rect 7926 40168 7932 40180
rect 7699 40140 7932 40168
rect 7699 40137 7711 40140
rect 7653 40131 7711 40137
rect 7926 40128 7932 40140
rect 7984 40128 7990 40180
rect 8570 40168 8576 40180
rect 8531 40140 8576 40168
rect 8570 40128 8576 40140
rect 8628 40128 8634 40180
rect 9217 40171 9275 40177
rect 9217 40137 9229 40171
rect 9263 40137 9275 40171
rect 9217 40131 9275 40137
rect 14645 40171 14703 40177
rect 14645 40137 14657 40171
rect 14691 40168 14703 40171
rect 14826 40168 14832 40180
rect 14691 40140 14832 40168
rect 14691 40137 14703 40140
rect 14645 40131 14703 40137
rect 7392 40072 7512 40100
rect 1857 40035 1915 40041
rect 1857 40001 1869 40035
rect 1903 40032 1915 40035
rect 2958 40032 2964 40044
rect 1903 40004 2964 40032
rect 1903 40001 1915 40004
rect 1857 39995 1915 40001
rect 2958 39992 2964 40004
rect 3016 39992 3022 40044
rect 5718 39992 5724 40044
rect 5776 40032 5782 40044
rect 5813 40035 5871 40041
rect 5813 40032 5825 40035
rect 5776 40004 5825 40032
rect 5776 39992 5782 40004
rect 5813 40001 5825 40004
rect 5859 40001 5871 40035
rect 5813 39995 5871 40001
rect 6730 39992 6736 40044
rect 6788 40032 6794 40044
rect 6825 40035 6883 40041
rect 6825 40032 6837 40035
rect 6788 40004 6837 40032
rect 6788 39992 6794 40004
rect 6825 40001 6837 40004
rect 6871 40032 6883 40035
rect 7190 40032 7196 40044
rect 6871 40004 7196 40032
rect 6871 40001 6883 40004
rect 6825 39995 6883 40001
rect 7190 39992 7196 40004
rect 7248 40032 7254 40044
rect 7374 40032 7380 40044
rect 7248 40004 7380 40032
rect 7248 39992 7254 40004
rect 7374 39992 7380 40004
rect 7432 39992 7438 40044
rect 7484 40041 7512 40072
rect 8018 40060 8024 40112
rect 8076 40100 8082 40112
rect 9232 40100 9260 40131
rect 14826 40128 14832 40140
rect 14884 40128 14890 40180
rect 16574 40128 16580 40180
rect 16632 40168 16638 40180
rect 16853 40171 16911 40177
rect 16632 40140 16804 40168
rect 16632 40128 16638 40140
rect 15562 40100 15568 40112
rect 8076 40072 9076 40100
rect 9232 40072 9904 40100
rect 15523 40072 15568 40100
rect 8076 40060 8082 40072
rect 8404 40041 8432 40072
rect 9048 40041 9076 40072
rect 9876 40041 9904 40072
rect 15562 40060 15568 40072
rect 15620 40060 15626 40112
rect 16482 40060 16488 40112
rect 16540 40100 16546 40112
rect 16776 40100 16804 40140
rect 16853 40137 16865 40171
rect 16899 40168 16911 40171
rect 17402 40168 17408 40180
rect 16899 40140 17408 40168
rect 16899 40137 16911 40140
rect 16853 40131 16911 40137
rect 17402 40128 17408 40140
rect 17460 40128 17466 40180
rect 17497 40171 17555 40177
rect 17497 40137 17509 40171
rect 17543 40137 17555 40171
rect 17497 40131 17555 40137
rect 17865 40171 17923 40177
rect 17865 40137 17877 40171
rect 17911 40168 17923 40171
rect 18414 40168 18420 40180
rect 17911 40140 18420 40168
rect 17911 40137 17923 40140
rect 17865 40131 17923 40137
rect 17512 40100 17540 40131
rect 18414 40128 18420 40140
rect 18472 40128 18478 40180
rect 18892 40140 20024 40168
rect 17954 40100 17960 40112
rect 16540 40072 16712 40100
rect 16776 40072 17540 40100
rect 17915 40072 17960 40100
rect 16540 40060 16546 40072
rect 7469 40035 7527 40041
rect 7469 40001 7481 40035
rect 7515 40001 7527 40035
rect 7469 39995 7527 40001
rect 8389 40035 8447 40041
rect 8389 40001 8401 40035
rect 8435 40001 8447 40035
rect 8389 39995 8447 40001
rect 9033 40035 9091 40041
rect 9033 40001 9045 40035
rect 9079 40001 9091 40035
rect 9033 39995 9091 40001
rect 9861 40035 9919 40041
rect 9861 40001 9873 40035
rect 9907 40001 9919 40035
rect 9861 39995 9919 40001
rect 12618 39992 12624 40044
rect 12676 40032 12682 40044
rect 12805 40035 12863 40041
rect 12805 40032 12817 40035
rect 12676 40004 12817 40032
rect 12676 39992 12682 40004
rect 12805 40001 12817 40004
rect 12851 40001 12863 40035
rect 12805 39995 12863 40001
rect 12894 39992 12900 40044
rect 12952 40032 12958 40044
rect 12989 40035 13047 40041
rect 12989 40032 13001 40035
rect 12952 40004 13001 40032
rect 12952 39992 12958 40004
rect 12989 40001 13001 40004
rect 13035 40001 13047 40035
rect 12989 39995 13047 40001
rect 15654 39992 15660 40044
rect 15712 40032 15718 40044
rect 16684 40041 16712 40072
rect 17954 40060 17960 40072
rect 18012 40060 18018 40112
rect 18046 40060 18052 40112
rect 18104 40100 18110 40112
rect 18892 40109 18920 40140
rect 18877 40103 18935 40109
rect 18877 40100 18889 40103
rect 18104 40072 18889 40100
rect 18104 40060 18110 40072
rect 18877 40069 18889 40072
rect 18923 40069 18935 40103
rect 19794 40100 19800 40112
rect 19755 40072 19800 40100
rect 18877 40063 18935 40069
rect 19794 40060 19800 40072
rect 19852 40060 19858 40112
rect 19996 40109 20024 40140
rect 19981 40103 20039 40109
rect 19981 40069 19993 40103
rect 20027 40069 20039 40103
rect 19981 40063 20039 40069
rect 15749 40035 15807 40041
rect 15749 40032 15761 40035
rect 15712 40004 15761 40032
rect 15712 39992 15718 40004
rect 15749 40001 15761 40004
rect 15795 40001 15807 40035
rect 15749 39995 15807 40001
rect 16669 40035 16727 40041
rect 16669 40001 16681 40035
rect 16715 40001 16727 40035
rect 18690 40032 18696 40044
rect 18651 40004 18696 40032
rect 16669 39995 16727 40001
rect 18690 39992 18696 40004
rect 18748 39992 18754 40044
rect 2866 39964 2872 39976
rect 2827 39936 2872 39964
rect 2866 39924 2872 39936
rect 2924 39924 2930 39976
rect 13538 39924 13544 39976
rect 13596 39964 13602 39976
rect 13725 39967 13783 39973
rect 13725 39964 13737 39967
rect 13596 39936 13737 39964
rect 13596 39924 13602 39936
rect 13725 39933 13737 39936
rect 13771 39933 13783 39967
rect 13725 39927 13783 39933
rect 13814 39924 13820 39976
rect 13872 39973 13878 39976
rect 13872 39967 13900 39973
rect 13888 39933 13900 39967
rect 13872 39927 13900 39933
rect 13872 39924 13878 39927
rect 13998 39924 14004 39976
rect 14056 39964 14062 39976
rect 16206 39964 16212 39976
rect 14056 39936 16212 39964
rect 14056 39924 14062 39936
rect 16206 39924 16212 39936
rect 16264 39964 16270 39976
rect 16758 39964 16764 39976
rect 16264 39936 16764 39964
rect 16264 39924 16270 39936
rect 16758 39924 16764 39936
rect 16816 39964 16822 39976
rect 18049 39967 18107 39973
rect 18049 39964 18061 39967
rect 16816 39936 18061 39964
rect 16816 39924 16822 39936
rect 18049 39933 18061 39936
rect 18095 39964 18107 39967
rect 18874 39964 18880 39976
rect 18095 39936 18880 39964
rect 18095 39933 18107 39936
rect 18049 39927 18107 39933
rect 18874 39924 18880 39936
rect 18932 39924 18938 39976
rect 4522 39856 4528 39908
rect 4580 39896 4586 39908
rect 5261 39899 5319 39905
rect 5261 39896 5273 39899
rect 4580 39868 5273 39896
rect 4580 39856 4586 39868
rect 5261 39865 5273 39868
rect 5307 39865 5319 39899
rect 5261 39859 5319 39865
rect 13449 39899 13507 39905
rect 13449 39865 13461 39899
rect 13495 39865 13507 39899
rect 13449 39859 13507 39865
rect 2222 39828 2228 39840
rect 2183 39800 2228 39828
rect 2222 39788 2228 39800
rect 2280 39788 2286 39840
rect 2409 39831 2467 39837
rect 2409 39797 2421 39831
rect 2455 39828 2467 39831
rect 3510 39828 3516 39840
rect 2455 39800 3516 39828
rect 2455 39797 2467 39800
rect 2409 39791 2467 39797
rect 3510 39788 3516 39800
rect 3568 39788 3574 39840
rect 4338 39788 4344 39840
rect 4396 39828 4402 39840
rect 4890 39828 4896 39840
rect 4396 39800 4896 39828
rect 4396 39788 4402 39800
rect 4890 39788 4896 39800
rect 4948 39788 4954 39840
rect 5350 39788 5356 39840
rect 5408 39828 5414 39840
rect 5445 39831 5503 39837
rect 5445 39828 5457 39831
rect 5408 39800 5457 39828
rect 5408 39788 5414 39800
rect 5445 39797 5457 39800
rect 5491 39797 5503 39831
rect 6914 39828 6920 39840
rect 6875 39800 6920 39828
rect 5445 39791 5503 39797
rect 6914 39788 6920 39800
rect 6972 39788 6978 39840
rect 9674 39828 9680 39840
rect 9635 39800 9680 39828
rect 9674 39788 9680 39800
rect 9732 39788 9738 39840
rect 13464 39828 13492 39859
rect 15746 39856 15752 39908
rect 15804 39896 15810 39908
rect 15933 39899 15991 39905
rect 15933 39896 15945 39899
rect 15804 39868 15945 39896
rect 15804 39856 15810 39868
rect 15933 39865 15945 39868
rect 15979 39865 15991 39899
rect 15933 39859 15991 39865
rect 15654 39828 15660 39840
rect 13464 39800 15660 39828
rect 15654 39788 15660 39800
rect 15712 39788 15718 39840
rect 19061 39831 19119 39837
rect 19061 39797 19073 39831
rect 19107 39828 19119 39831
rect 19426 39828 19432 39840
rect 19107 39800 19432 39828
rect 19107 39797 19119 39800
rect 19061 39791 19119 39797
rect 19426 39788 19432 39800
rect 19484 39788 19490 39840
rect 20070 39788 20076 39840
rect 20128 39828 20134 39840
rect 20165 39831 20223 39837
rect 20165 39828 20177 39831
rect 20128 39800 20177 39828
rect 20128 39788 20134 39800
rect 20165 39797 20177 39800
rect 20211 39797 20223 39831
rect 20165 39791 20223 39797
rect 1104 39738 30820 39760
rect 1104 39686 5915 39738
rect 5967 39686 5979 39738
rect 6031 39686 6043 39738
rect 6095 39686 6107 39738
rect 6159 39686 6171 39738
rect 6223 39686 15846 39738
rect 15898 39686 15910 39738
rect 15962 39686 15974 39738
rect 16026 39686 16038 39738
rect 16090 39686 16102 39738
rect 16154 39686 25776 39738
rect 25828 39686 25840 39738
rect 25892 39686 25904 39738
rect 25956 39686 25968 39738
rect 26020 39686 26032 39738
rect 26084 39686 30820 39738
rect 1104 39664 30820 39686
rect 2866 39624 2872 39636
rect 2827 39596 2872 39624
rect 2866 39584 2872 39596
rect 2924 39584 2930 39636
rect 5810 39624 5816 39636
rect 5771 39596 5816 39624
rect 5810 39584 5816 39596
rect 5868 39584 5874 39636
rect 6638 39584 6644 39636
rect 6696 39624 6702 39636
rect 6696 39596 7144 39624
rect 6696 39584 6702 39596
rect 4522 39516 4528 39568
rect 4580 39556 4586 39568
rect 7006 39556 7012 39568
rect 4580 39528 7012 39556
rect 4580 39516 4586 39528
rect 7006 39516 7012 39528
rect 7064 39516 7070 39568
rect 7116 39556 7144 39596
rect 8018 39584 8024 39636
rect 8076 39624 8082 39636
rect 8205 39627 8263 39633
rect 8205 39624 8217 39627
rect 8076 39596 8217 39624
rect 8076 39584 8082 39596
rect 8205 39593 8217 39596
rect 8251 39593 8263 39627
rect 9674 39624 9680 39636
rect 8205 39587 8263 39593
rect 9416 39596 9680 39624
rect 8846 39556 8852 39568
rect 7116 39528 8852 39556
rect 8846 39516 8852 39528
rect 8904 39516 8910 39568
rect 4062 39488 4068 39500
rect 2424 39460 4068 39488
rect 1578 39380 1584 39432
rect 1636 39420 1642 39432
rect 2424 39429 2452 39460
rect 4062 39448 4068 39460
rect 4120 39448 4126 39500
rect 6362 39448 6368 39500
rect 6420 39488 6426 39500
rect 9416 39497 9444 39596
rect 9674 39584 9680 39596
rect 9732 39584 9738 39636
rect 12986 39624 12992 39636
rect 12947 39596 12992 39624
rect 12986 39584 12992 39596
rect 13044 39584 13050 39636
rect 15654 39624 15660 39636
rect 15304 39596 15660 39624
rect 15304 39565 15332 39596
rect 15654 39584 15660 39596
rect 15712 39584 15718 39636
rect 18509 39627 18567 39633
rect 18509 39593 18521 39627
rect 18555 39624 18567 39627
rect 18598 39624 18604 39636
rect 18555 39596 18604 39624
rect 18555 39593 18567 39596
rect 18509 39587 18567 39593
rect 18598 39584 18604 39596
rect 18656 39584 18662 39636
rect 15289 39559 15347 39565
rect 15289 39525 15301 39559
rect 15335 39525 15347 39559
rect 15289 39519 15347 39525
rect 20533 39559 20591 39565
rect 20533 39525 20545 39559
rect 20579 39556 20591 39559
rect 22278 39556 22284 39568
rect 20579 39528 22284 39556
rect 20579 39525 20591 39528
rect 20533 39519 20591 39525
rect 22278 39516 22284 39528
rect 22336 39516 22342 39568
rect 9401 39491 9459 39497
rect 6420 39460 7052 39488
rect 6420 39448 6426 39460
rect 1673 39423 1731 39429
rect 1673 39420 1685 39423
rect 1636 39392 1685 39420
rect 1636 39380 1642 39392
rect 1673 39389 1685 39392
rect 1719 39389 1731 39423
rect 1673 39383 1731 39389
rect 2409 39423 2467 39429
rect 2409 39389 2421 39423
rect 2455 39389 2467 39423
rect 3050 39420 3056 39432
rect 3011 39392 3056 39420
rect 2409 39383 2467 39389
rect 3050 39380 3056 39392
rect 3108 39380 3114 39432
rect 3786 39420 3792 39432
rect 3747 39392 3792 39420
rect 3786 39380 3792 39392
rect 3844 39380 3850 39432
rect 4525 39423 4583 39429
rect 4525 39389 4537 39423
rect 4571 39420 4583 39423
rect 5353 39423 5411 39429
rect 4571 39392 5212 39420
rect 4571 39389 4583 39392
rect 4525 39383 4583 39389
rect 1486 39284 1492 39296
rect 1447 39256 1492 39284
rect 1486 39244 1492 39256
rect 1544 39244 1550 39296
rect 2222 39284 2228 39296
rect 2183 39256 2228 39284
rect 2222 39244 2228 39256
rect 2280 39244 2286 39296
rect 3970 39284 3976 39296
rect 3931 39256 3976 39284
rect 3970 39244 3976 39256
rect 4028 39244 4034 39296
rect 4706 39284 4712 39296
rect 4667 39256 4712 39284
rect 4706 39244 4712 39256
rect 4764 39244 4770 39296
rect 5184 39293 5212 39392
rect 5353 39389 5365 39423
rect 5399 39420 5411 39423
rect 5810 39420 5816 39432
rect 5399 39392 5816 39420
rect 5399 39389 5411 39392
rect 5353 39383 5411 39389
rect 5810 39380 5816 39392
rect 5868 39380 5874 39432
rect 5997 39423 6055 39429
rect 5997 39389 6009 39423
rect 6043 39420 6055 39423
rect 6454 39420 6460 39432
rect 6043 39392 6316 39420
rect 6415 39392 6460 39420
rect 6043 39389 6055 39392
rect 5997 39383 6055 39389
rect 5169 39287 5227 39293
rect 5169 39253 5181 39287
rect 5215 39253 5227 39287
rect 6288 39284 6316 39392
rect 6454 39380 6460 39392
rect 6512 39380 6518 39432
rect 6638 39420 6644 39432
rect 6599 39392 6644 39420
rect 6638 39380 6644 39392
rect 6696 39380 6702 39432
rect 6730 39380 6736 39432
rect 6788 39420 6794 39432
rect 6914 39429 6920 39432
rect 6871 39423 6920 39429
rect 6788 39392 6833 39420
rect 6788 39380 6794 39392
rect 6871 39389 6883 39423
rect 6917 39389 6920 39423
rect 6871 39383 6920 39389
rect 6914 39380 6920 39383
rect 6972 39380 6978 39432
rect 7024 39429 7052 39460
rect 9401 39457 9413 39491
rect 9447 39457 9459 39491
rect 9401 39451 9459 39457
rect 14274 39448 14280 39500
rect 14332 39488 14338 39500
rect 14645 39491 14703 39497
rect 14645 39488 14657 39491
rect 14332 39460 14657 39488
rect 14332 39448 14338 39460
rect 14645 39457 14657 39460
rect 14691 39488 14703 39491
rect 15010 39488 15016 39500
rect 14691 39460 15016 39488
rect 14691 39457 14703 39460
rect 14645 39451 14703 39457
rect 15010 39448 15016 39460
rect 15068 39448 15074 39500
rect 15378 39448 15384 39500
rect 15436 39488 15442 39500
rect 15682 39491 15740 39497
rect 15682 39488 15694 39491
rect 15436 39460 15694 39488
rect 15436 39448 15442 39460
rect 15682 39457 15694 39460
rect 15728 39457 15740 39491
rect 15682 39451 15740 39457
rect 16850 39448 16856 39500
rect 16908 39488 16914 39500
rect 17037 39491 17095 39497
rect 17037 39488 17049 39491
rect 16908 39460 17049 39488
rect 16908 39448 16914 39460
rect 17037 39457 17049 39460
rect 17083 39457 17095 39491
rect 17037 39451 17095 39457
rect 7009 39423 7067 39429
rect 7009 39389 7021 39423
rect 7055 39389 7067 39423
rect 7009 39383 7067 39389
rect 8389 39423 8447 39429
rect 8389 39389 8401 39423
rect 8435 39389 8447 39423
rect 8389 39383 8447 39389
rect 12621 39423 12679 39429
rect 12621 39389 12633 39423
rect 12667 39420 12679 39423
rect 12894 39420 12900 39432
rect 12667 39392 12900 39420
rect 12667 39389 12679 39392
rect 12621 39383 12679 39389
rect 8404 39352 8432 39383
rect 12894 39380 12900 39392
rect 12952 39380 12958 39432
rect 14826 39420 14832 39432
rect 14787 39392 14832 39420
rect 14826 39380 14832 39392
rect 14884 39380 14890 39432
rect 15562 39380 15568 39432
rect 15620 39420 15626 39432
rect 15838 39420 15844 39432
rect 15620 39392 15665 39420
rect 15799 39392 15844 39420
rect 15620 39380 15626 39392
rect 15838 39380 15844 39392
rect 15896 39380 15902 39432
rect 17954 39380 17960 39432
rect 18012 39420 18018 39432
rect 18141 39423 18199 39429
rect 18141 39420 18153 39423
rect 18012 39392 18153 39420
rect 18012 39380 18018 39392
rect 18141 39389 18153 39392
rect 18187 39389 18199 39423
rect 19426 39420 19432 39432
rect 19387 39392 19432 39420
rect 18141 39383 18199 39389
rect 19426 39380 19432 39392
rect 19484 39380 19490 39432
rect 21729 39423 21787 39429
rect 21729 39389 21741 39423
rect 21775 39389 21787 39423
rect 21729 39383 21787 39389
rect 21913 39423 21971 39429
rect 21913 39389 21925 39423
rect 21959 39420 21971 39423
rect 30098 39420 30104 39432
rect 21959 39392 26234 39420
rect 30059 39392 30104 39420
rect 21959 39389 21971 39392
rect 21913 39383 21971 39389
rect 9674 39361 9680 39364
rect 6840 39324 8432 39352
rect 6840 39296 6868 39324
rect 9668 39315 9680 39361
rect 9732 39352 9738 39364
rect 12805 39355 12863 39361
rect 9732 39324 9768 39352
rect 9674 39312 9680 39315
rect 9732 39312 9738 39324
rect 12805 39321 12817 39355
rect 12851 39352 12863 39355
rect 14090 39352 14096 39364
rect 12851 39324 14096 39352
rect 12851 39321 12863 39324
rect 12805 39315 12863 39321
rect 14090 39312 14096 39324
rect 14148 39352 14154 39364
rect 14458 39352 14464 39364
rect 14148 39324 14464 39352
rect 14148 39312 14154 39324
rect 14458 39312 14464 39324
rect 14516 39312 14522 39364
rect 16485 39355 16543 39361
rect 16485 39321 16497 39355
rect 16531 39352 16543 39355
rect 17313 39355 17371 39361
rect 17313 39352 17325 39355
rect 16531 39324 17325 39352
rect 16531 39321 16543 39324
rect 16485 39315 16543 39321
rect 17313 39321 17325 39324
rect 17359 39321 17371 39355
rect 17313 39315 17371 39321
rect 18046 39312 18052 39364
rect 18104 39352 18110 39364
rect 18325 39355 18383 39361
rect 18325 39352 18337 39355
rect 18104 39324 18337 39352
rect 18104 39312 18110 39324
rect 18325 39321 18337 39324
rect 18371 39321 18383 39355
rect 18325 39315 18383 39321
rect 18874 39312 18880 39364
rect 18932 39352 18938 39364
rect 19981 39355 20039 39361
rect 19981 39352 19993 39355
rect 18932 39324 19993 39352
rect 18932 39312 18938 39324
rect 19981 39321 19993 39324
rect 20027 39321 20039 39355
rect 20254 39352 20260 39364
rect 20215 39324 20260 39352
rect 19981 39315 20039 39321
rect 20254 39312 20260 39324
rect 20312 39312 20318 39364
rect 21744 39352 21772 39383
rect 22002 39352 22008 39364
rect 21744 39324 22008 39352
rect 22002 39312 22008 39324
rect 22060 39312 22066 39364
rect 6822 39284 6828 39296
rect 6288 39256 6828 39284
rect 5169 39247 5227 39253
rect 6822 39244 6828 39256
rect 6880 39284 6886 39296
rect 7190 39284 7196 39296
rect 6880 39256 6973 39284
rect 7151 39256 7196 39284
rect 6880 39244 6886 39256
rect 7190 39244 7196 39256
rect 7248 39244 7254 39296
rect 10778 39284 10784 39296
rect 10739 39256 10784 39284
rect 10778 39244 10784 39256
rect 10836 39244 10842 39296
rect 15010 39244 15016 39296
rect 15068 39284 15074 39296
rect 15562 39284 15568 39296
rect 15068 39256 15568 39284
rect 15068 39244 15074 39256
rect 15562 39244 15568 39256
rect 15620 39244 15626 39296
rect 16114 39244 16120 39296
rect 16172 39284 16178 39296
rect 17221 39287 17279 39293
rect 17221 39284 17233 39287
rect 16172 39256 17233 39284
rect 16172 39244 16178 39256
rect 17221 39253 17233 39256
rect 17267 39253 17279 39287
rect 17221 39247 17279 39253
rect 17681 39287 17739 39293
rect 17681 39253 17693 39287
rect 17727 39284 17739 39287
rect 18690 39284 18696 39296
rect 17727 39256 18696 39284
rect 17727 39253 17739 39256
rect 17681 39247 17739 39253
rect 18690 39244 18696 39256
rect 18748 39244 18754 39296
rect 19150 39244 19156 39296
rect 19208 39284 19214 39296
rect 19245 39287 19303 39293
rect 19245 39284 19257 39287
rect 19208 39256 19257 39284
rect 19208 39244 19214 39256
rect 19245 39253 19257 39256
rect 19291 39253 19303 39287
rect 19245 39247 19303 39253
rect 19794 39244 19800 39296
rect 19852 39284 19858 39296
rect 20073 39287 20131 39293
rect 20073 39284 20085 39287
rect 19852 39256 20085 39284
rect 19852 39244 19858 39256
rect 20073 39253 20085 39256
rect 20119 39253 20131 39287
rect 21542 39284 21548 39296
rect 21503 39256 21548 39284
rect 20073 39247 20131 39253
rect 21542 39244 21548 39256
rect 21600 39244 21606 39296
rect 26206 39284 26234 39392
rect 30098 39380 30104 39392
rect 30156 39380 30162 39432
rect 29917 39287 29975 39293
rect 29917 39284 29929 39287
rect 26206 39256 29929 39284
rect 29917 39253 29929 39256
rect 29963 39253 29975 39287
rect 29917 39247 29975 39253
rect 1104 39194 30820 39216
rect 1104 39142 10880 39194
rect 10932 39142 10944 39194
rect 10996 39142 11008 39194
rect 11060 39142 11072 39194
rect 11124 39142 11136 39194
rect 11188 39142 20811 39194
rect 20863 39142 20875 39194
rect 20927 39142 20939 39194
rect 20991 39142 21003 39194
rect 21055 39142 21067 39194
rect 21119 39142 30820 39194
rect 1104 39120 30820 39142
rect 2409 39083 2467 39089
rect 2409 39049 2421 39083
rect 2455 39080 2467 39083
rect 2498 39080 2504 39092
rect 2455 39052 2504 39080
rect 2455 39049 2467 39052
rect 2409 39043 2467 39049
rect 2498 39040 2504 39052
rect 2556 39040 2562 39092
rect 6362 39040 6368 39092
rect 6420 39080 6426 39092
rect 8205 39083 8263 39089
rect 8205 39080 8217 39083
rect 6420 39052 8217 39080
rect 6420 39040 6426 39052
rect 8205 39049 8217 39052
rect 8251 39049 8263 39083
rect 13538 39080 13544 39092
rect 13499 39052 13544 39080
rect 8205 39043 8263 39049
rect 13538 39040 13544 39052
rect 13596 39080 13602 39092
rect 15286 39080 15292 39092
rect 13596 39052 15292 39080
rect 13596 39040 13602 39052
rect 15286 39040 15292 39052
rect 15344 39040 15350 39092
rect 16114 39080 16120 39092
rect 16075 39052 16120 39080
rect 16114 39040 16120 39052
rect 16172 39040 16178 39092
rect 19150 39080 19156 39092
rect 19111 39052 19156 39080
rect 19150 39040 19156 39052
rect 19208 39040 19214 39092
rect 20254 39080 20260 39092
rect 20215 39052 20260 39080
rect 20254 39040 20260 39052
rect 20312 39040 20318 39092
rect 2225 39015 2283 39021
rect 2225 38981 2237 39015
rect 2271 39012 2283 39015
rect 2271 38984 4108 39012
rect 2271 38981 2283 38984
rect 2225 38975 2283 38981
rect 2869 38947 2927 38953
rect 2869 38913 2881 38947
rect 2915 38944 2927 38947
rect 3142 38944 3148 38956
rect 2915 38916 3148 38944
rect 2915 38913 2927 38916
rect 2869 38907 2927 38913
rect 3142 38904 3148 38916
rect 3200 38904 3206 38956
rect 4080 38953 4108 38984
rect 4706 38972 4712 39024
rect 4764 39012 4770 39024
rect 7092 39015 7150 39021
rect 4764 38984 6868 39012
rect 4764 38972 4770 38984
rect 4065 38947 4123 38953
rect 4065 38913 4077 38947
rect 4111 38944 4123 38947
rect 4154 38944 4160 38956
rect 4111 38916 4160 38944
rect 4111 38913 4123 38916
rect 4065 38907 4123 38913
rect 4154 38904 4160 38916
rect 4212 38904 4218 38956
rect 4430 38944 4436 38956
rect 4391 38916 4436 38944
rect 4430 38904 4436 38916
rect 4488 38904 4494 38956
rect 4614 38944 4620 38956
rect 4575 38916 4620 38944
rect 4614 38904 4620 38916
rect 4672 38904 4678 38956
rect 5810 38944 5816 38956
rect 5771 38916 5816 38944
rect 5810 38904 5816 38916
rect 5868 38904 5874 38956
rect 6840 38953 6868 38984
rect 7092 38981 7104 39015
rect 7138 39012 7150 39015
rect 7190 39012 7196 39024
rect 7138 38984 7196 39012
rect 7138 38981 7150 38984
rect 7092 38975 7150 38981
rect 7190 38972 7196 38984
rect 7248 38972 7254 39024
rect 13814 39012 13820 39024
rect 13775 38984 13820 39012
rect 13814 38972 13820 38984
rect 13872 38972 13878 39024
rect 18690 38972 18696 39024
rect 18748 39012 18754 39024
rect 19061 39015 19119 39021
rect 19061 39012 19073 39015
rect 18748 38984 19073 39012
rect 18748 38972 18754 38984
rect 19061 38981 19073 38984
rect 19107 38981 19119 39015
rect 19061 38975 19119 38981
rect 6825 38947 6883 38953
rect 6825 38913 6837 38947
rect 6871 38913 6883 38947
rect 6825 38907 6883 38913
rect 9122 38904 9128 38956
rect 9180 38944 9186 38956
rect 9490 38953 9496 38956
rect 9217 38947 9275 38953
rect 9217 38944 9229 38947
rect 9180 38916 9229 38944
rect 9180 38904 9186 38916
rect 9217 38913 9229 38916
rect 9263 38913 9275 38947
rect 9217 38907 9275 38913
rect 9484 38907 9496 38953
rect 9548 38944 9554 38956
rect 9548 38916 9584 38944
rect 9490 38904 9496 38907
rect 9548 38904 9554 38916
rect 12618 38904 12624 38956
rect 12676 38944 12682 38956
rect 13265 38947 13323 38953
rect 13265 38944 13277 38947
rect 12676 38916 13277 38944
rect 12676 38904 12682 38916
rect 13265 38913 13277 38916
rect 13311 38913 13323 38947
rect 14274 38944 14280 38956
rect 14235 38916 14280 38944
rect 13265 38907 13323 38913
rect 14274 38904 14280 38916
rect 14332 38904 14338 38956
rect 15286 38904 15292 38956
rect 15344 38953 15350 38956
rect 15344 38947 15372 38953
rect 15360 38913 15372 38947
rect 20070 38944 20076 38956
rect 20031 38916 20076 38944
rect 15344 38907 15372 38913
rect 15344 38904 15350 38907
rect 20070 38904 20076 38916
rect 20128 38904 20134 38956
rect 1857 38879 1915 38885
rect 1857 38845 1869 38879
rect 1903 38876 1915 38879
rect 2958 38876 2964 38888
rect 1903 38848 2964 38876
rect 1903 38845 1915 38848
rect 1857 38839 1915 38845
rect 2958 38836 2964 38848
rect 3016 38836 3022 38888
rect 4246 38876 4252 38888
rect 4159 38848 4252 38876
rect 4246 38836 4252 38848
rect 4304 38836 4310 38888
rect 4338 38836 4344 38888
rect 4396 38876 4402 38888
rect 13173 38879 13231 38885
rect 4396 38848 4441 38876
rect 4396 38836 4402 38848
rect 13173 38845 13185 38879
rect 13219 38876 13231 38879
rect 13998 38876 14004 38888
rect 13219 38848 14004 38876
rect 13219 38845 13231 38848
rect 13173 38839 13231 38845
rect 13998 38836 14004 38848
rect 14056 38836 14062 38888
rect 14461 38879 14519 38885
rect 14461 38845 14473 38879
rect 14507 38876 14519 38879
rect 14826 38876 14832 38888
rect 14507 38848 14832 38876
rect 14507 38845 14519 38848
rect 14461 38839 14519 38845
rect 14826 38836 14832 38848
rect 14884 38836 14890 38888
rect 14921 38879 14979 38885
rect 14921 38845 14933 38879
rect 14967 38845 14979 38879
rect 15194 38876 15200 38888
rect 15155 38848 15200 38876
rect 14921 38839 14979 38845
rect 2866 38768 2872 38820
rect 2924 38808 2930 38820
rect 4264 38808 4292 38836
rect 4982 38808 4988 38820
rect 2924 38780 4988 38808
rect 2924 38768 2930 38780
rect 4982 38768 4988 38780
rect 5040 38768 5046 38820
rect 14936 38752 14964 38839
rect 15194 38836 15200 38848
rect 15252 38836 15258 38888
rect 15473 38879 15531 38885
rect 15473 38845 15485 38879
rect 15519 38876 15531 38879
rect 15838 38876 15844 38888
rect 15519 38848 15844 38876
rect 15519 38845 15531 38848
rect 15473 38839 15531 38845
rect 15838 38836 15844 38848
rect 15896 38876 15902 38888
rect 16206 38876 16212 38888
rect 15896 38848 16212 38876
rect 15896 38836 15902 38848
rect 16206 38836 16212 38848
rect 16264 38836 16270 38888
rect 18874 38876 18880 38888
rect 18835 38848 18880 38876
rect 18874 38836 18880 38848
rect 18932 38836 18938 38888
rect 1946 38700 1952 38752
rect 2004 38740 2010 38752
rect 2225 38743 2283 38749
rect 2225 38740 2237 38743
rect 2004 38712 2237 38740
rect 2004 38700 2010 38712
rect 2225 38709 2237 38712
rect 2271 38740 2283 38743
rect 2314 38740 2320 38752
rect 2271 38712 2320 38740
rect 2271 38709 2283 38712
rect 2225 38703 2283 38709
rect 2314 38700 2320 38712
rect 2372 38700 2378 38752
rect 3050 38740 3056 38752
rect 3011 38712 3056 38740
rect 3050 38700 3056 38712
rect 3108 38700 3114 38752
rect 3881 38743 3939 38749
rect 3881 38709 3893 38743
rect 3927 38740 3939 38743
rect 4246 38740 4252 38752
rect 3927 38712 4252 38740
rect 3927 38709 3939 38712
rect 3881 38703 3939 38709
rect 4246 38700 4252 38712
rect 4304 38700 4310 38752
rect 5718 38740 5724 38752
rect 5679 38712 5724 38740
rect 5718 38700 5724 38712
rect 5776 38700 5782 38752
rect 6454 38700 6460 38752
rect 6512 38740 6518 38752
rect 7006 38740 7012 38752
rect 6512 38712 7012 38740
rect 6512 38700 6518 38712
rect 7006 38700 7012 38712
rect 7064 38700 7070 38752
rect 9214 38700 9220 38752
rect 9272 38740 9278 38752
rect 10597 38743 10655 38749
rect 10597 38740 10609 38743
rect 9272 38712 10609 38740
rect 9272 38700 9278 38712
rect 10597 38709 10609 38712
rect 10643 38709 10655 38743
rect 10597 38703 10655 38709
rect 14918 38700 14924 38752
rect 14976 38700 14982 38752
rect 19521 38743 19579 38749
rect 19521 38709 19533 38743
rect 19567 38740 19579 38743
rect 20254 38740 20260 38752
rect 19567 38712 20260 38740
rect 19567 38709 19579 38712
rect 19521 38703 19579 38709
rect 20254 38700 20260 38712
rect 20312 38700 20318 38752
rect 1104 38650 30820 38672
rect 1104 38598 5915 38650
rect 5967 38598 5979 38650
rect 6031 38598 6043 38650
rect 6095 38598 6107 38650
rect 6159 38598 6171 38650
rect 6223 38598 15846 38650
rect 15898 38598 15910 38650
rect 15962 38598 15974 38650
rect 16026 38598 16038 38650
rect 16090 38598 16102 38650
rect 16154 38598 25776 38650
rect 25828 38598 25840 38650
rect 25892 38598 25904 38650
rect 25956 38598 25968 38650
rect 26020 38598 26032 38650
rect 26084 38598 30820 38650
rect 1104 38576 30820 38598
rect 1857 38539 1915 38545
rect 1857 38505 1869 38539
rect 1903 38536 1915 38539
rect 1946 38536 1952 38548
rect 1903 38508 1952 38536
rect 1903 38505 1915 38508
rect 1857 38499 1915 38505
rect 1946 38496 1952 38508
rect 2004 38496 2010 38548
rect 2041 38539 2099 38545
rect 2041 38505 2053 38539
rect 2087 38536 2099 38539
rect 2130 38536 2136 38548
rect 2087 38508 2136 38536
rect 2087 38505 2099 38508
rect 2041 38499 2099 38505
rect 2130 38496 2136 38508
rect 2188 38496 2194 38548
rect 4154 38496 4160 38548
rect 4212 38536 4218 38548
rect 5353 38539 5411 38545
rect 5353 38536 5365 38539
rect 4212 38508 5365 38536
rect 4212 38496 4218 38508
rect 5353 38505 5365 38508
rect 5399 38505 5411 38539
rect 9306 38536 9312 38548
rect 5353 38499 5411 38505
rect 6840 38508 9312 38536
rect 1489 38471 1547 38477
rect 1489 38437 1501 38471
rect 1535 38468 1547 38471
rect 2958 38468 2964 38480
rect 1535 38440 2964 38468
rect 1535 38437 1547 38440
rect 1489 38431 1547 38437
rect 2958 38428 2964 38440
rect 3016 38428 3022 38480
rect 2866 38400 2872 38412
rect 2827 38372 2872 38400
rect 2866 38360 2872 38372
rect 2924 38360 2930 38412
rect 3789 38403 3847 38409
rect 3789 38400 3801 38403
rect 2976 38372 3801 38400
rect 2682 38332 2688 38344
rect 2643 38304 2688 38332
rect 2682 38292 2688 38304
rect 2740 38292 2746 38344
rect 2976 38341 3004 38372
rect 3789 38369 3801 38372
rect 3835 38369 3847 38403
rect 3970 38400 3976 38412
rect 3931 38372 3976 38400
rect 3789 38363 3847 38369
rect 3970 38360 3976 38372
rect 4028 38360 4034 38412
rect 4982 38360 4988 38412
rect 5040 38400 5046 38412
rect 6089 38403 6147 38409
rect 6089 38400 6101 38403
rect 5040 38372 6101 38400
rect 5040 38360 5046 38372
rect 6089 38369 6101 38372
rect 6135 38369 6147 38403
rect 6089 38363 6147 38369
rect 2961 38335 3019 38341
rect 2961 38301 2973 38335
rect 3007 38301 3019 38335
rect 2961 38295 3019 38301
rect 3053 38335 3111 38341
rect 3053 38301 3065 38335
rect 3099 38332 3111 38335
rect 3142 38332 3148 38344
rect 3099 38304 3148 38332
rect 3099 38301 3111 38304
rect 3053 38295 3111 38301
rect 3142 38292 3148 38304
rect 3200 38292 3206 38344
rect 3237 38335 3295 38341
rect 3237 38301 3249 38335
rect 3283 38332 3295 38335
rect 4062 38332 4068 38344
rect 3283 38304 4068 38332
rect 3283 38301 3295 38304
rect 3237 38295 3295 38301
rect 4062 38292 4068 38304
rect 4120 38292 4126 38344
rect 4246 38341 4252 38344
rect 4240 38332 4252 38341
rect 4207 38304 4252 38332
rect 4240 38295 4252 38304
rect 4246 38292 4252 38295
rect 4304 38292 4310 38344
rect 5810 38332 5816 38344
rect 5723 38304 5816 38332
rect 5810 38292 5816 38304
rect 5868 38332 5874 38344
rect 6840 38332 6868 38508
rect 9306 38496 9312 38508
rect 9364 38496 9370 38548
rect 9398 38496 9404 38548
rect 9456 38536 9462 38548
rect 12529 38539 12587 38545
rect 9456 38508 12434 38536
rect 9456 38496 9462 38508
rect 7006 38428 7012 38480
rect 7064 38468 7070 38480
rect 10778 38468 10784 38480
rect 7064 38440 7788 38468
rect 7064 38428 7070 38440
rect 6914 38360 6920 38412
rect 6972 38400 6978 38412
rect 7469 38403 7527 38409
rect 7469 38400 7481 38403
rect 6972 38372 7481 38400
rect 6972 38360 6978 38372
rect 7469 38369 7481 38372
rect 7515 38369 7527 38403
rect 7760 38400 7788 38440
rect 7944 38440 10784 38468
rect 7760 38372 7880 38400
rect 7469 38363 7527 38369
rect 7282 38332 7288 38344
rect 5868 38304 6868 38332
rect 7243 38304 7288 38332
rect 5868 38292 5874 38304
rect 7282 38292 7288 38304
rect 7340 38292 7346 38344
rect 7374 38292 7380 38344
rect 7432 38332 7438 38344
rect 7561 38335 7619 38341
rect 7561 38332 7573 38335
rect 7432 38304 7573 38332
rect 7432 38292 7438 38304
rect 7561 38301 7573 38304
rect 7607 38301 7619 38335
rect 7561 38295 7619 38301
rect 7650 38292 7656 38344
rect 7708 38332 7714 38344
rect 7852 38341 7880 38372
rect 7837 38335 7895 38341
rect 7708 38304 7753 38332
rect 7708 38292 7714 38304
rect 7837 38301 7849 38335
rect 7883 38301 7895 38335
rect 7837 38295 7895 38301
rect 1857 38267 1915 38273
rect 1857 38233 1869 38267
rect 1903 38264 1915 38267
rect 1903 38236 7604 38264
rect 1903 38233 1915 38236
rect 1857 38227 1915 38233
rect 2498 38196 2504 38208
rect 2459 38168 2504 38196
rect 2498 38156 2504 38168
rect 2556 38156 2562 38208
rect 3789 38199 3847 38205
rect 3789 38165 3801 38199
rect 3835 38196 3847 38199
rect 4338 38196 4344 38208
rect 3835 38168 4344 38196
rect 3835 38165 3847 38168
rect 3789 38159 3847 38165
rect 4338 38156 4344 38168
rect 4396 38156 4402 38208
rect 7098 38196 7104 38208
rect 7059 38168 7104 38196
rect 7098 38156 7104 38168
rect 7156 38156 7162 38208
rect 7576 38196 7604 38236
rect 7944 38196 7972 38440
rect 8754 38360 8760 38412
rect 8812 38400 8818 38412
rect 9217 38403 9275 38409
rect 9217 38400 9229 38403
rect 8812 38372 9229 38400
rect 8812 38360 8818 38372
rect 9217 38369 9229 38372
rect 9263 38369 9275 38403
rect 9217 38363 9275 38369
rect 8941 38335 8999 38341
rect 8941 38301 8953 38335
rect 8987 38301 8999 38335
rect 8941 38295 8999 38301
rect 8662 38224 8668 38276
rect 8720 38264 8726 38276
rect 8956 38264 8984 38295
rect 9030 38292 9036 38344
rect 9088 38332 9094 38344
rect 9125 38335 9183 38341
rect 9125 38332 9137 38335
rect 9088 38304 9137 38332
rect 9088 38292 9094 38304
rect 9125 38301 9137 38304
rect 9171 38301 9183 38335
rect 9306 38332 9312 38344
rect 9267 38304 9312 38332
rect 9125 38295 9183 38301
rect 9306 38292 9312 38304
rect 9364 38292 9370 38344
rect 9508 38341 9536 38440
rect 10778 38428 10784 38440
rect 10836 38428 10842 38480
rect 12406 38468 12434 38508
rect 12529 38505 12541 38539
rect 12575 38536 12587 38539
rect 12894 38536 12900 38548
rect 12575 38508 12900 38536
rect 12575 38505 12587 38508
rect 12529 38499 12587 38505
rect 12894 38496 12900 38508
rect 12952 38496 12958 38548
rect 14277 38539 14335 38545
rect 14277 38505 14289 38539
rect 14323 38536 14335 38539
rect 14826 38536 14832 38548
rect 14323 38508 14832 38536
rect 14323 38505 14335 38508
rect 14277 38499 14335 38505
rect 14826 38496 14832 38508
rect 14884 38496 14890 38548
rect 17402 38536 17408 38548
rect 17315 38508 17408 38536
rect 17402 38496 17408 38508
rect 17460 38536 17466 38548
rect 19426 38536 19432 38548
rect 17460 38508 19432 38536
rect 17460 38496 17466 38508
rect 19426 38496 19432 38508
rect 19484 38496 19490 38548
rect 12406 38440 12848 38468
rect 9582 38360 9588 38412
rect 9640 38400 9646 38412
rect 9640 38372 11008 38400
rect 9640 38360 9646 38372
rect 9493 38335 9551 38341
rect 9493 38301 9505 38335
rect 9539 38301 9551 38335
rect 9674 38332 9680 38344
rect 9635 38304 9680 38332
rect 9493 38295 9551 38301
rect 9674 38292 9680 38304
rect 9732 38292 9738 38344
rect 10594 38292 10600 38344
rect 10652 38332 10658 38344
rect 10873 38335 10931 38341
rect 10873 38332 10885 38335
rect 10652 38304 10885 38332
rect 10652 38292 10658 38304
rect 10873 38301 10885 38304
rect 10919 38301 10931 38335
rect 10873 38295 10931 38301
rect 10980 38264 11008 38372
rect 12345 38335 12403 38341
rect 12345 38301 12357 38335
rect 12391 38332 12403 38335
rect 12710 38332 12716 38344
rect 12391 38304 12716 38332
rect 12391 38301 12403 38304
rect 12345 38295 12403 38301
rect 12710 38292 12716 38304
rect 12768 38292 12774 38344
rect 12820 38264 12848 38440
rect 12912 38400 12940 38496
rect 18601 38471 18659 38477
rect 18601 38437 18613 38471
rect 18647 38437 18659 38471
rect 18601 38431 18659 38437
rect 12989 38403 13047 38409
rect 12989 38400 13001 38403
rect 12912 38372 13001 38400
rect 12989 38369 13001 38372
rect 13035 38369 13047 38403
rect 12989 38363 13047 38369
rect 13170 38332 13176 38344
rect 13131 38304 13176 38332
rect 13170 38292 13176 38304
rect 13228 38292 13234 38344
rect 13357 38335 13415 38341
rect 13357 38301 13369 38335
rect 13403 38332 13415 38335
rect 14093 38335 14151 38341
rect 14093 38332 14105 38335
rect 13403 38304 14105 38332
rect 13403 38301 13415 38304
rect 13357 38295 13415 38301
rect 14093 38301 14105 38304
rect 14139 38301 14151 38335
rect 17586 38332 17592 38344
rect 17547 38304 17592 38332
rect 14093 38295 14151 38301
rect 17586 38292 17592 38304
rect 17644 38292 17650 38344
rect 18414 38332 18420 38344
rect 18375 38304 18420 38332
rect 18414 38292 18420 38304
rect 18472 38292 18478 38344
rect 18616 38332 18644 38431
rect 19429 38335 19487 38341
rect 19429 38332 19441 38335
rect 18616 38304 19441 38332
rect 19429 38301 19441 38304
rect 19475 38301 19487 38335
rect 30098 38332 30104 38344
rect 30059 38304 30104 38332
rect 19429 38295 19487 38301
rect 30098 38292 30104 38304
rect 30156 38292 30162 38344
rect 21542 38264 21548 38276
rect 8720 38236 10824 38264
rect 10980 38236 12756 38264
rect 12820 38236 21548 38264
rect 8720 38224 8726 38236
rect 7576 38168 7972 38196
rect 8846 38156 8852 38208
rect 8904 38196 8910 38208
rect 9582 38196 9588 38208
rect 8904 38168 9588 38196
rect 8904 38156 8910 38168
rect 9582 38156 9588 38168
rect 9640 38156 9646 38208
rect 9950 38156 9956 38208
rect 10008 38196 10014 38208
rect 10689 38199 10747 38205
rect 10689 38196 10701 38199
rect 10008 38168 10701 38196
rect 10008 38156 10014 38168
rect 10689 38165 10701 38168
rect 10735 38165 10747 38199
rect 10796 38196 10824 38236
rect 12526 38196 12532 38208
rect 10796 38168 12532 38196
rect 10689 38159 10747 38165
rect 12526 38156 12532 38168
rect 12584 38156 12590 38208
rect 12728 38196 12756 38236
rect 21542 38224 21548 38236
rect 21600 38224 21606 38276
rect 17310 38196 17316 38208
rect 12728 38168 17316 38196
rect 17310 38156 17316 38168
rect 17368 38156 17374 38208
rect 18966 38156 18972 38208
rect 19024 38196 19030 38208
rect 19245 38199 19303 38205
rect 19245 38196 19257 38199
rect 19024 38168 19257 38196
rect 19024 38156 19030 38168
rect 19245 38165 19257 38168
rect 19291 38165 19303 38199
rect 29914 38196 29920 38208
rect 29875 38168 29920 38196
rect 19245 38159 19303 38165
rect 29914 38156 29920 38168
rect 29972 38156 29978 38208
rect 1104 38106 30820 38128
rect 1104 38054 10880 38106
rect 10932 38054 10944 38106
rect 10996 38054 11008 38106
rect 11060 38054 11072 38106
rect 11124 38054 11136 38106
rect 11188 38054 20811 38106
rect 20863 38054 20875 38106
rect 20927 38054 20939 38106
rect 20991 38054 21003 38106
rect 21055 38054 21067 38106
rect 21119 38054 30820 38106
rect 1104 38032 30820 38054
rect 1854 37952 1860 38004
rect 1912 37992 1918 38004
rect 1949 37995 2007 38001
rect 1949 37992 1961 37995
rect 1912 37964 1961 37992
rect 1912 37952 1918 37964
rect 1949 37961 1961 37964
rect 1995 37961 2007 37995
rect 1949 37955 2007 37961
rect 2133 37995 2191 38001
rect 2133 37961 2145 37995
rect 2179 37992 2191 37995
rect 2682 37992 2688 38004
rect 2179 37964 2688 37992
rect 2179 37961 2191 37964
rect 2133 37955 2191 37961
rect 2682 37952 2688 37964
rect 2740 37992 2746 38004
rect 3053 37995 3111 38001
rect 3053 37992 3065 37995
rect 2740 37964 3065 37992
rect 2740 37952 2746 37964
rect 3053 37961 3065 37964
rect 3099 37961 3111 37995
rect 3053 37955 3111 37961
rect 3142 37952 3148 38004
rect 3200 37992 3206 38004
rect 3694 37992 3700 38004
rect 3200 37964 3700 37992
rect 3200 37952 3206 37964
rect 3694 37952 3700 37964
rect 3752 37992 3758 38004
rect 7466 37992 7472 38004
rect 3752 37964 7472 37992
rect 3752 37952 3758 37964
rect 7466 37952 7472 37964
rect 7524 37952 7530 38004
rect 9401 37995 9459 38001
rect 7576 37964 9352 37992
rect 2498 37884 2504 37936
rect 2556 37924 2562 37936
rect 4166 37927 4224 37933
rect 4166 37924 4178 37927
rect 2556 37896 4178 37924
rect 2556 37884 2562 37896
rect 4166 37893 4178 37896
rect 4212 37893 4224 37927
rect 4166 37887 4224 37893
rect 6362 37884 6368 37936
rect 6420 37924 6426 37936
rect 6546 37924 6552 37936
rect 6420 37896 6552 37924
rect 6420 37884 6426 37896
rect 6546 37884 6552 37896
rect 6604 37924 6610 37936
rect 7576 37924 7604 37964
rect 6604 37896 7604 37924
rect 9324 37924 9352 37964
rect 9401 37961 9413 37995
rect 9447 37992 9459 37995
rect 9490 37992 9496 38004
rect 9447 37964 9496 37992
rect 9447 37961 9459 37964
rect 9401 37955 9459 37961
rect 9490 37952 9496 37964
rect 9548 37952 9554 38004
rect 12710 37992 12716 38004
rect 12671 37964 12716 37992
rect 12710 37952 12716 37964
rect 12768 37952 12774 38004
rect 13817 37995 13875 38001
rect 13817 37961 13829 37995
rect 13863 37992 13875 37995
rect 15102 37992 15108 38004
rect 13863 37964 15108 37992
rect 13863 37961 13875 37964
rect 13817 37955 13875 37961
rect 15102 37952 15108 37964
rect 15160 37952 15166 38004
rect 17310 37952 17316 38004
rect 17368 37992 17374 38004
rect 21913 37995 21971 38001
rect 21913 37992 21925 37995
rect 17368 37964 21925 37992
rect 17368 37952 17374 37964
rect 21913 37961 21925 37964
rect 21959 37961 21971 37995
rect 21913 37955 21971 37961
rect 9324 37896 12434 37924
rect 6604 37884 6610 37896
rect 4338 37816 4344 37868
rect 4396 37856 4402 37868
rect 5537 37859 5595 37865
rect 5537 37856 5549 37859
rect 4396 37828 5549 37856
rect 4396 37816 4402 37828
rect 5537 37825 5549 37828
rect 5583 37825 5595 37859
rect 5537 37819 5595 37825
rect 5718 37816 5724 37868
rect 5776 37856 5782 37868
rect 5813 37859 5871 37865
rect 5813 37856 5825 37859
rect 5776 37828 5825 37856
rect 5776 37816 5782 37828
rect 5813 37825 5825 37828
rect 5859 37856 5871 37859
rect 8018 37856 8024 37868
rect 5859 37828 7696 37856
rect 7979 37828 8024 37856
rect 5859 37825 5871 37828
rect 5813 37819 5871 37825
rect 2501 37791 2559 37797
rect 2501 37757 2513 37791
rect 2547 37788 2559 37791
rect 2958 37788 2964 37800
rect 2547 37760 2964 37788
rect 2547 37757 2559 37760
rect 2501 37751 2559 37757
rect 2958 37748 2964 37760
rect 3016 37748 3022 37800
rect 4430 37788 4436 37800
rect 4391 37760 4436 37788
rect 4430 37748 4436 37760
rect 4488 37748 4494 37800
rect 6362 37788 6368 37800
rect 6323 37760 6368 37788
rect 6362 37748 6368 37760
rect 6420 37748 6426 37800
rect 6641 37791 6699 37797
rect 6641 37757 6653 37791
rect 6687 37757 6699 37791
rect 7668 37788 7696 37828
rect 8018 37816 8024 37828
rect 8076 37816 8082 37868
rect 8294 37816 8300 37868
rect 8352 37856 8358 37868
rect 8662 37856 8668 37868
rect 8352 37828 8668 37856
rect 8352 37816 8358 37828
rect 8662 37816 8668 37828
rect 8720 37816 8726 37868
rect 8846 37856 8852 37868
rect 8807 37828 8852 37856
rect 8846 37816 8852 37828
rect 8904 37816 8910 37868
rect 9214 37856 9220 37868
rect 9127 37828 9220 37856
rect 9214 37816 9220 37828
rect 9272 37856 9278 37868
rect 9950 37856 9956 37868
rect 9272 37828 9444 37856
rect 9911 37828 9956 37856
rect 9272 37816 9278 37828
rect 8478 37788 8484 37800
rect 7668 37760 8484 37788
rect 6641 37751 6699 37757
rect 4614 37680 4620 37732
rect 4672 37720 4678 37732
rect 6656 37720 6684 37751
rect 8478 37748 8484 37760
rect 8536 37788 8542 37800
rect 8754 37788 8760 37800
rect 8536 37760 8760 37788
rect 8536 37748 8542 37760
rect 8754 37748 8760 37760
rect 8812 37788 8818 37800
rect 8941 37791 8999 37797
rect 8941 37788 8953 37791
rect 8812 37760 8953 37788
rect 8812 37748 8818 37760
rect 8941 37757 8953 37760
rect 8987 37757 8999 37791
rect 8941 37751 8999 37757
rect 9033 37791 9091 37797
rect 9033 37757 9045 37791
rect 9079 37788 9091 37791
rect 9122 37788 9128 37800
rect 9079 37760 9128 37788
rect 9079 37757 9091 37760
rect 9033 37751 9091 37757
rect 9122 37748 9128 37760
rect 9180 37788 9186 37800
rect 9306 37788 9312 37800
rect 9180 37760 9312 37788
rect 9180 37748 9186 37760
rect 9306 37748 9312 37760
rect 9364 37748 9370 37800
rect 9416 37720 9444 37828
rect 9950 37816 9956 37828
rect 10008 37816 10014 37868
rect 10042 37816 10048 37868
rect 10100 37856 10106 37868
rect 10594 37856 10600 37868
rect 10100 37828 10600 37856
rect 10100 37816 10106 37828
rect 10594 37816 10600 37828
rect 10652 37816 10658 37868
rect 11701 37859 11759 37865
rect 11701 37856 11713 37859
rect 10796 37828 11713 37856
rect 10796 37729 10824 37828
rect 11701 37825 11713 37828
rect 11747 37825 11759 37859
rect 11701 37819 11759 37825
rect 4672 37692 6684 37720
rect 8137 37692 9444 37720
rect 10781 37723 10839 37729
rect 4672 37680 4678 37692
rect 1946 37612 1952 37664
rect 2004 37652 2010 37664
rect 2133 37655 2191 37661
rect 2133 37652 2145 37655
rect 2004 37624 2145 37652
rect 2004 37612 2010 37624
rect 2133 37621 2145 37624
rect 2179 37621 2191 37655
rect 2133 37615 2191 37621
rect 4154 37612 4160 37664
rect 4212 37652 4218 37664
rect 4632 37652 4660 37680
rect 4212 37624 4660 37652
rect 4212 37612 4218 37624
rect 5442 37612 5448 37664
rect 5500 37652 5506 37664
rect 8137 37652 8165 37692
rect 10781 37689 10793 37723
rect 10827 37689 10839 37723
rect 12406 37720 12434 37896
rect 12526 37884 12532 37936
rect 12584 37924 12590 37936
rect 17402 37924 17408 37936
rect 12584 37896 17408 37924
rect 12584 37884 12590 37896
rect 17402 37884 17408 37896
rect 17460 37884 17466 37936
rect 17681 37927 17739 37933
rect 17681 37893 17693 37927
rect 17727 37924 17739 37927
rect 18046 37924 18052 37936
rect 17727 37896 18052 37924
rect 17727 37893 17739 37896
rect 17681 37887 17739 37893
rect 18046 37884 18052 37896
rect 18104 37884 18110 37936
rect 18414 37924 18420 37936
rect 18327 37896 18420 37924
rect 12618 37816 12624 37868
rect 12676 37856 12682 37868
rect 12897 37859 12955 37865
rect 12897 37856 12909 37859
rect 12676 37828 12909 37856
rect 12676 37816 12682 37828
rect 12897 37825 12909 37828
rect 12943 37825 12955 37859
rect 13078 37856 13084 37868
rect 13039 37828 13084 37856
rect 12897 37819 12955 37825
rect 13078 37816 13084 37828
rect 13136 37816 13142 37868
rect 13998 37856 14004 37868
rect 13959 37828 14004 37856
rect 13998 37816 14004 37828
rect 14056 37816 14062 37868
rect 14918 37856 14924 37868
rect 14108 37828 14924 37856
rect 13725 37791 13783 37797
rect 13725 37757 13737 37791
rect 13771 37788 13783 37791
rect 14108 37788 14136 37828
rect 14918 37816 14924 37828
rect 14976 37816 14982 37868
rect 16853 37859 16911 37865
rect 16853 37825 16865 37859
rect 16899 37856 16911 37859
rect 17497 37859 17555 37865
rect 17497 37856 17509 37859
rect 16899 37828 17509 37856
rect 16899 37825 16911 37828
rect 16853 37819 16911 37825
rect 17497 37825 17509 37828
rect 17543 37825 17555 37859
rect 17862 37856 17868 37868
rect 17823 37828 17868 37856
rect 17497 37819 17555 37825
rect 17862 37816 17868 37828
rect 17920 37816 17926 37868
rect 18340 37865 18368 37896
rect 18414 37884 18420 37896
rect 18472 37924 18478 37936
rect 20714 37924 20720 37936
rect 18472 37896 20720 37924
rect 18472 37884 18478 37896
rect 20714 37884 20720 37896
rect 20772 37884 20778 37936
rect 18325 37859 18383 37865
rect 18325 37825 18337 37859
rect 18371 37825 18383 37859
rect 18966 37856 18972 37868
rect 18927 37828 18972 37856
rect 18325 37819 18383 37825
rect 18966 37816 18972 37828
rect 19024 37816 19030 37868
rect 19242 37865 19248 37868
rect 19236 37819 19248 37865
rect 19300 37856 19306 37868
rect 19300 37828 19336 37856
rect 19242 37816 19248 37819
rect 19300 37816 19306 37828
rect 22002 37816 22008 37868
rect 22060 37856 22066 37868
rect 22097 37859 22155 37865
rect 22097 37856 22109 37859
rect 22060 37828 22109 37856
rect 22060 37816 22066 37828
rect 22097 37825 22109 37828
rect 22143 37825 22155 37859
rect 22097 37819 22155 37825
rect 14274 37788 14280 37800
rect 13771 37760 14136 37788
rect 14235 37760 14280 37788
rect 13771 37757 13783 37760
rect 13725 37751 13783 37757
rect 14274 37748 14280 37760
rect 14332 37788 14338 37800
rect 14829 37791 14887 37797
rect 14829 37788 14841 37791
rect 14332 37760 14841 37788
rect 14332 37748 14338 37760
rect 14829 37757 14841 37760
rect 14875 37757 14887 37791
rect 14829 37751 14887 37757
rect 22281 37791 22339 37797
rect 22281 37757 22293 37791
rect 22327 37788 22339 37791
rect 29914 37788 29920 37800
rect 22327 37760 29920 37788
rect 22327 37757 22339 37760
rect 22281 37751 22339 37757
rect 29914 37748 29920 37760
rect 29972 37748 29978 37800
rect 17586 37720 17592 37732
rect 12406 37692 17592 37720
rect 10781 37683 10839 37689
rect 17586 37680 17592 37692
rect 17644 37680 17650 37732
rect 5500 37624 8165 37652
rect 8205 37655 8263 37661
rect 5500 37612 5506 37624
rect 8205 37621 8217 37655
rect 8251 37652 8263 37655
rect 9306 37652 9312 37664
rect 8251 37624 9312 37652
rect 8251 37621 8263 37624
rect 8205 37615 8263 37621
rect 9306 37612 9312 37624
rect 9364 37612 9370 37664
rect 10137 37655 10195 37661
rect 10137 37621 10149 37655
rect 10183 37652 10195 37655
rect 10870 37652 10876 37664
rect 10183 37624 10876 37652
rect 10183 37621 10195 37624
rect 10137 37615 10195 37621
rect 10870 37612 10876 37624
rect 10928 37612 10934 37664
rect 11514 37652 11520 37664
rect 11475 37624 11520 37652
rect 11514 37612 11520 37624
rect 11572 37612 11578 37664
rect 12710 37612 12716 37664
rect 12768 37652 12774 37664
rect 13081 37655 13139 37661
rect 13081 37652 13093 37655
rect 12768 37624 13093 37652
rect 12768 37612 12774 37624
rect 13081 37621 13093 37624
rect 13127 37652 13139 37655
rect 13725 37655 13783 37661
rect 13725 37652 13737 37655
rect 13127 37624 13737 37652
rect 13127 37621 13139 37624
rect 13081 37615 13139 37621
rect 13725 37621 13737 37624
rect 13771 37621 13783 37655
rect 14182 37652 14188 37664
rect 14143 37624 14188 37652
rect 13725 37615 13783 37621
rect 14182 37612 14188 37624
rect 14240 37612 14246 37664
rect 17037 37655 17095 37661
rect 17037 37621 17049 37655
rect 17083 37652 17095 37655
rect 17954 37652 17960 37664
rect 17083 37624 17960 37652
rect 17083 37621 17095 37624
rect 17037 37615 17095 37621
rect 17954 37612 17960 37624
rect 18012 37612 18018 37664
rect 18509 37655 18567 37661
rect 18509 37621 18521 37655
rect 18555 37652 18567 37655
rect 19334 37652 19340 37664
rect 18555 37624 19340 37652
rect 18555 37621 18567 37624
rect 18509 37615 18567 37621
rect 19334 37612 19340 37624
rect 19392 37612 19398 37664
rect 20346 37652 20352 37664
rect 20307 37624 20352 37652
rect 20346 37612 20352 37624
rect 20404 37612 20410 37664
rect 1104 37562 30820 37584
rect 1104 37510 5915 37562
rect 5967 37510 5979 37562
rect 6031 37510 6043 37562
rect 6095 37510 6107 37562
rect 6159 37510 6171 37562
rect 6223 37510 15846 37562
rect 15898 37510 15910 37562
rect 15962 37510 15974 37562
rect 16026 37510 16038 37562
rect 16090 37510 16102 37562
rect 16154 37510 25776 37562
rect 25828 37510 25840 37562
rect 25892 37510 25904 37562
rect 25956 37510 25968 37562
rect 26020 37510 26032 37562
rect 26084 37510 30820 37562
rect 1104 37488 30820 37510
rect 1946 37408 1952 37460
rect 2004 37448 2010 37460
rect 2225 37451 2283 37457
rect 2225 37448 2237 37451
rect 2004 37420 2237 37448
rect 2004 37408 2010 37420
rect 2225 37417 2237 37420
rect 2271 37417 2283 37451
rect 2225 37411 2283 37417
rect 6917 37451 6975 37457
rect 6917 37417 6929 37451
rect 6963 37448 6975 37451
rect 7282 37448 7288 37460
rect 6963 37420 7288 37448
rect 6963 37417 6975 37420
rect 6917 37411 6975 37417
rect 7282 37408 7288 37420
rect 7340 37408 7346 37460
rect 7469 37451 7527 37457
rect 7469 37417 7481 37451
rect 7515 37417 7527 37451
rect 7469 37411 7527 37417
rect 12897 37451 12955 37457
rect 12897 37417 12909 37451
rect 12943 37448 12955 37451
rect 13170 37448 13176 37460
rect 12943 37420 13176 37448
rect 12943 37417 12955 37420
rect 12897 37411 12955 37417
rect 7190 37340 7196 37392
rect 7248 37380 7254 37392
rect 7484 37380 7512 37411
rect 13170 37408 13176 37420
rect 13228 37408 13234 37460
rect 14093 37451 14151 37457
rect 14093 37417 14105 37451
rect 14139 37448 14151 37451
rect 14182 37448 14188 37460
rect 14139 37420 14188 37448
rect 14139 37417 14151 37420
rect 14093 37411 14151 37417
rect 14182 37408 14188 37420
rect 14240 37408 14246 37460
rect 15102 37408 15108 37460
rect 15160 37448 15166 37460
rect 16298 37448 16304 37460
rect 15160 37420 16304 37448
rect 15160 37408 15166 37420
rect 16298 37408 16304 37420
rect 16356 37408 16362 37460
rect 7248 37352 7512 37380
rect 12805 37383 12863 37389
rect 7248 37340 7254 37352
rect 12805 37349 12817 37383
rect 12851 37380 12863 37383
rect 13078 37380 13084 37392
rect 12851 37352 13084 37380
rect 12851 37349 12863 37352
rect 12805 37343 12863 37349
rect 13078 37340 13084 37352
rect 13136 37340 13142 37392
rect 15304 37352 15700 37380
rect 5442 37312 5448 37324
rect 2516 37284 5448 37312
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37244 1915 37247
rect 2314 37244 2320 37256
rect 1903 37216 2320 37244
rect 1903 37213 1915 37216
rect 1857 37207 1915 37213
rect 2314 37204 2320 37216
rect 2372 37204 2378 37256
rect 2225 37179 2283 37185
rect 2225 37145 2237 37179
rect 2271 37176 2283 37179
rect 2516 37176 2544 37284
rect 5442 37272 5448 37284
rect 5500 37272 5506 37324
rect 10870 37312 10876 37324
rect 10831 37284 10876 37312
rect 10870 37272 10876 37284
rect 10928 37272 10934 37324
rect 12618 37272 12624 37324
rect 12676 37312 12682 37324
rect 12989 37315 13047 37321
rect 12989 37312 13001 37315
rect 12676 37284 13001 37312
rect 12676 37272 12682 37284
rect 12989 37281 13001 37284
rect 13035 37281 13047 37315
rect 15194 37312 15200 37324
rect 12989 37275 13047 37281
rect 14936 37284 15200 37312
rect 2590 37204 2596 37256
rect 2648 37244 2654 37256
rect 2869 37247 2927 37253
rect 2869 37246 2881 37247
rect 2746 37244 2881 37246
rect 2648 37218 2881 37244
rect 2648 37216 2774 37218
rect 2648 37204 2654 37216
rect 2869 37213 2881 37218
rect 2915 37213 2927 37247
rect 2869 37207 2927 37213
rect 2958 37204 2964 37256
rect 3016 37244 3022 37256
rect 3970 37244 3976 37256
rect 3016 37216 3976 37244
rect 3016 37204 3022 37216
rect 3970 37204 3976 37216
rect 4028 37204 4034 37256
rect 4617 37247 4675 37253
rect 4617 37213 4629 37247
rect 4663 37213 4675 37247
rect 4617 37207 4675 37213
rect 4632 37176 4660 37207
rect 4982 37204 4988 37256
rect 5040 37244 5046 37256
rect 5537 37247 5595 37253
rect 5537 37244 5549 37247
rect 5040 37216 5549 37244
rect 5040 37204 5046 37216
rect 5537 37213 5549 37216
rect 5583 37213 5595 37247
rect 5537 37207 5595 37213
rect 5804 37247 5862 37253
rect 5804 37213 5816 37247
rect 5850 37244 5862 37247
rect 7098 37244 7104 37256
rect 5850 37216 7104 37244
rect 5850 37213 5862 37216
rect 5804 37207 5862 37213
rect 7098 37204 7104 37216
rect 7156 37204 7162 37256
rect 7377 37247 7435 37253
rect 7377 37213 7389 37247
rect 7423 37244 7435 37247
rect 9674 37244 9680 37256
rect 7423 37216 9680 37244
rect 7423 37213 7435 37216
rect 7377 37207 7435 37213
rect 9674 37204 9680 37216
rect 9732 37204 9738 37256
rect 9766 37204 9772 37256
rect 9824 37244 9830 37256
rect 10321 37247 10379 37253
rect 10321 37244 10333 37247
rect 9824 37216 10333 37244
rect 9824 37204 9830 37216
rect 10321 37213 10333 37216
rect 10367 37213 10379 37247
rect 12710 37244 12716 37256
rect 12671 37216 12716 37244
rect 10321 37207 10379 37213
rect 12710 37204 12716 37216
rect 12768 37204 12774 37256
rect 14090 37244 14096 37256
rect 14051 37216 14096 37244
rect 14090 37204 14096 37216
rect 14148 37204 14154 37256
rect 14936 37253 14964 37284
rect 15194 37272 15200 37284
rect 15252 37312 15258 37324
rect 15304 37312 15332 37352
rect 15562 37312 15568 37324
rect 15252 37284 15332 37312
rect 15523 37284 15568 37312
rect 15252 37272 15258 37284
rect 15562 37272 15568 37284
rect 15620 37272 15626 37324
rect 15672 37312 15700 37352
rect 15841 37315 15899 37321
rect 15841 37312 15853 37315
rect 15672 37284 15853 37312
rect 15841 37281 15853 37284
rect 15887 37281 15899 37315
rect 15841 37275 15899 37281
rect 15979 37315 16037 37321
rect 15979 37281 15991 37315
rect 16025 37312 16037 37315
rect 16298 37312 16304 37324
rect 16025 37284 16304 37312
rect 16025 37281 16037 37284
rect 15979 37275 16037 37281
rect 16298 37272 16304 37284
rect 16356 37272 16362 37324
rect 17681 37315 17739 37321
rect 17681 37281 17693 37315
rect 17727 37281 17739 37315
rect 17862 37312 17868 37324
rect 17823 37284 17868 37312
rect 17681 37275 17739 37281
rect 14277 37247 14335 37253
rect 14277 37213 14289 37247
rect 14323 37213 14335 37247
rect 14277 37207 14335 37213
rect 14921 37247 14979 37253
rect 14921 37213 14933 37247
rect 14967 37213 14979 37247
rect 15102 37244 15108 37256
rect 15063 37216 15108 37244
rect 14921 37207 14979 37213
rect 2271 37148 2544 37176
rect 2884 37148 4660 37176
rect 2271 37145 2283 37148
rect 2225 37139 2283 37145
rect 2884 37120 2912 37148
rect 9030 37136 9036 37188
rect 9088 37176 9094 37188
rect 10054 37179 10112 37185
rect 10054 37176 10066 37179
rect 9088 37148 10066 37176
rect 9088 37136 9094 37148
rect 10054 37145 10066 37148
rect 10100 37145 10112 37179
rect 10054 37139 10112 37145
rect 11140 37179 11198 37185
rect 11140 37145 11152 37179
rect 11186 37176 11198 37179
rect 11238 37176 11244 37188
rect 11186 37148 11244 37176
rect 11186 37145 11198 37148
rect 11140 37139 11198 37145
rect 11238 37136 11244 37148
rect 11296 37136 11302 37188
rect 13078 37136 13084 37188
rect 13136 37176 13142 37188
rect 14292 37176 14320 37207
rect 15102 37204 15108 37216
rect 15160 37204 15166 37256
rect 16114 37244 16120 37256
rect 16075 37216 16120 37244
rect 16114 37204 16120 37216
rect 16172 37204 16178 37256
rect 14550 37176 14556 37188
rect 13136 37148 14556 37176
rect 13136 37136 13142 37148
rect 14550 37136 14556 37148
rect 14608 37136 14614 37188
rect 17696 37176 17724 37275
rect 17862 37272 17868 37284
rect 17920 37272 17926 37324
rect 17954 37244 17960 37256
rect 17915 37216 17960 37244
rect 17954 37204 17960 37216
rect 18012 37204 18018 37256
rect 19334 37204 19340 37256
rect 19392 37244 19398 37256
rect 19429 37247 19487 37253
rect 19429 37244 19441 37247
rect 19392 37216 19441 37244
rect 19392 37204 19398 37216
rect 19429 37213 19441 37216
rect 19475 37213 19487 37247
rect 19429 37207 19487 37213
rect 19978 37204 19984 37256
rect 20036 37244 20042 37256
rect 20257 37247 20315 37253
rect 20257 37244 20269 37247
rect 20036 37216 20269 37244
rect 20036 37204 20042 37216
rect 20257 37213 20269 37216
rect 20303 37213 20315 37247
rect 20257 37207 20315 37213
rect 20346 37204 20352 37256
rect 20404 37244 20410 37256
rect 20441 37247 20499 37253
rect 20441 37244 20453 37247
rect 20404 37216 20453 37244
rect 20404 37204 20410 37216
rect 20441 37213 20453 37216
rect 20487 37213 20499 37247
rect 20441 37207 20499 37213
rect 16592 37148 17724 37176
rect 2406 37108 2412 37120
rect 2367 37080 2412 37108
rect 2406 37068 2412 37080
rect 2464 37068 2470 37120
rect 2866 37068 2872 37120
rect 2924 37068 2930 37120
rect 3050 37108 3056 37120
rect 3011 37080 3056 37108
rect 3050 37068 3056 37080
rect 3108 37068 3114 37120
rect 3786 37108 3792 37120
rect 3747 37080 3792 37108
rect 3786 37068 3792 37080
rect 3844 37068 3850 37120
rect 3878 37068 3884 37120
rect 3936 37108 3942 37120
rect 4433 37111 4491 37117
rect 4433 37108 4445 37111
rect 3936 37080 4445 37108
rect 3936 37068 3942 37080
rect 4433 37077 4445 37080
rect 4479 37077 4491 37111
rect 4433 37071 4491 37077
rect 7837 37111 7895 37117
rect 7837 37077 7849 37111
rect 7883 37108 7895 37111
rect 8570 37108 8576 37120
rect 7883 37080 8576 37108
rect 7883 37077 7895 37080
rect 7837 37071 7895 37077
rect 8570 37068 8576 37080
rect 8628 37068 8634 37120
rect 8754 37068 8760 37120
rect 8812 37108 8818 37120
rect 8941 37111 8999 37117
rect 8941 37108 8953 37111
rect 8812 37080 8953 37108
rect 8812 37068 8818 37080
rect 8941 37077 8953 37080
rect 8987 37077 8999 37111
rect 8941 37071 8999 37077
rect 11422 37068 11428 37120
rect 11480 37108 11486 37120
rect 12253 37111 12311 37117
rect 12253 37108 12265 37111
rect 11480 37080 12265 37108
rect 11480 37068 11486 37080
rect 12253 37077 12265 37080
rect 12299 37077 12311 37111
rect 14568 37108 14596 37136
rect 15286 37108 15292 37120
rect 14568 37080 15292 37108
rect 12253 37071 12311 37077
rect 15286 37068 15292 37080
rect 15344 37068 15350 37120
rect 16206 37068 16212 37120
rect 16264 37108 16270 37120
rect 16592 37108 16620 37148
rect 20070 37136 20076 37188
rect 20128 37176 20134 37188
rect 20364 37176 20392 37204
rect 20128 37148 20392 37176
rect 20128 37136 20134 37148
rect 16758 37108 16764 37120
rect 16264 37080 16620 37108
rect 16719 37080 16764 37108
rect 16264 37068 16270 37080
rect 16758 37068 16764 37080
rect 16816 37068 16822 37120
rect 18138 37068 18144 37120
rect 18196 37108 18202 37120
rect 18325 37111 18383 37117
rect 18325 37108 18337 37111
rect 18196 37080 18337 37108
rect 18196 37068 18202 37080
rect 18325 37077 18337 37080
rect 18371 37077 18383 37111
rect 18325 37071 18383 37077
rect 18414 37068 18420 37120
rect 18472 37108 18478 37120
rect 19245 37111 19303 37117
rect 19245 37108 19257 37111
rect 18472 37080 19257 37108
rect 18472 37068 18478 37080
rect 19245 37077 19257 37080
rect 19291 37077 19303 37111
rect 20346 37108 20352 37120
rect 20307 37080 20352 37108
rect 19245 37071 19303 37077
rect 20346 37068 20352 37080
rect 20404 37068 20410 37120
rect 1104 37018 30820 37040
rect 1104 36966 10880 37018
rect 10932 36966 10944 37018
rect 10996 36966 11008 37018
rect 11060 36966 11072 37018
rect 11124 36966 11136 37018
rect 11188 36966 20811 37018
rect 20863 36966 20875 37018
rect 20927 36966 20939 37018
rect 20991 36966 21003 37018
rect 21055 36966 21067 37018
rect 21119 36966 30820 37018
rect 1104 36944 30820 36966
rect 1394 36864 1400 36916
rect 1452 36904 1458 36916
rect 2590 36904 2596 36916
rect 1452 36876 2596 36904
rect 1452 36864 1458 36876
rect 2590 36864 2596 36876
rect 2648 36864 2654 36916
rect 3697 36907 3755 36913
rect 3697 36873 3709 36907
rect 3743 36904 3755 36907
rect 4430 36904 4436 36916
rect 3743 36876 4436 36904
rect 3743 36873 3755 36876
rect 3697 36867 3755 36873
rect 4430 36864 4436 36876
rect 4488 36864 4494 36916
rect 4982 36904 4988 36916
rect 4943 36876 4988 36904
rect 4982 36864 4988 36876
rect 5040 36864 5046 36916
rect 6822 36864 6828 36916
rect 6880 36904 6886 36916
rect 8941 36907 8999 36913
rect 6880 36876 8524 36904
rect 6880 36864 6886 36876
rect 6730 36836 6736 36848
rect 1688 36808 6736 36836
rect 1688 36777 1716 36808
rect 6730 36796 6736 36808
rect 6788 36796 6794 36848
rect 8496 36836 8524 36876
rect 8941 36873 8953 36907
rect 8987 36904 8999 36907
rect 9030 36904 9036 36916
rect 8987 36876 9036 36904
rect 8987 36873 8999 36876
rect 8941 36867 8999 36873
rect 9030 36864 9036 36876
rect 9088 36864 9094 36916
rect 9858 36864 9864 36916
rect 9916 36904 9922 36916
rect 10318 36904 10324 36916
rect 9916 36876 10324 36904
rect 9916 36864 9922 36876
rect 10318 36864 10324 36876
rect 10376 36864 10382 36916
rect 12897 36907 12955 36913
rect 12897 36904 12909 36907
rect 10796 36876 12909 36904
rect 8496 36808 9628 36836
rect 1673 36771 1731 36777
rect 1673 36737 1685 36771
rect 1719 36737 1731 36771
rect 1673 36731 1731 36737
rect 2038 36728 2044 36780
rect 2096 36768 2102 36780
rect 2133 36771 2191 36777
rect 2133 36768 2145 36771
rect 2096 36740 2145 36768
rect 2096 36728 2102 36740
rect 2133 36737 2145 36740
rect 2179 36737 2191 36771
rect 2133 36731 2191 36737
rect 2774 36728 2780 36780
rect 2832 36768 2838 36780
rect 2869 36771 2927 36777
rect 2869 36768 2881 36771
rect 2832 36740 2881 36768
rect 2832 36728 2838 36740
rect 2869 36737 2881 36740
rect 2915 36737 2927 36771
rect 3513 36771 3571 36777
rect 3513 36768 3525 36771
rect 2869 36731 2927 36737
rect 3068 36740 3525 36768
rect 2406 36592 2412 36644
rect 2464 36632 2470 36644
rect 3068 36641 3096 36740
rect 3513 36737 3525 36740
rect 3559 36737 3571 36771
rect 3513 36731 3571 36737
rect 4154 36728 4160 36780
rect 4212 36768 4218 36780
rect 4341 36771 4399 36777
rect 4341 36768 4353 36771
rect 4212 36740 4353 36768
rect 4212 36728 4218 36740
rect 4341 36737 4353 36740
rect 4387 36737 4399 36771
rect 4341 36731 4399 36737
rect 4801 36771 4859 36777
rect 4801 36737 4813 36771
rect 4847 36768 4859 36771
rect 5166 36768 5172 36780
rect 4847 36740 5172 36768
rect 4847 36737 4859 36740
rect 4801 36731 4859 36737
rect 4356 36700 4384 36731
rect 5166 36728 5172 36740
rect 5224 36728 5230 36780
rect 5626 36768 5632 36780
rect 5587 36740 5632 36768
rect 5626 36728 5632 36740
rect 5684 36728 5690 36780
rect 6825 36771 6883 36777
rect 6825 36768 6837 36771
rect 6288 36740 6837 36768
rect 4890 36700 4896 36712
rect 4356 36672 4896 36700
rect 4890 36660 4896 36672
rect 4948 36700 4954 36712
rect 6288 36700 6316 36740
rect 6825 36737 6837 36740
rect 6871 36768 6883 36771
rect 7190 36768 7196 36780
rect 6871 36740 7196 36768
rect 6871 36737 6883 36740
rect 6825 36731 6883 36737
rect 7190 36728 7196 36740
rect 7248 36728 7254 36780
rect 8205 36771 8263 36777
rect 8205 36737 8217 36771
rect 8251 36768 8263 36771
rect 8294 36768 8300 36780
rect 8251 36740 8300 36768
rect 8251 36737 8263 36740
rect 8205 36731 8263 36737
rect 8294 36728 8300 36740
rect 8352 36728 8358 36780
rect 8386 36728 8392 36780
rect 8444 36768 8450 36780
rect 8754 36768 8760 36780
rect 8444 36740 8489 36768
rect 8715 36740 8760 36768
rect 8444 36728 8450 36740
rect 8754 36728 8760 36740
rect 8812 36728 8818 36780
rect 9600 36777 9628 36808
rect 9674 36796 9680 36848
rect 9732 36836 9738 36848
rect 10796 36836 10824 36876
rect 12897 36873 12909 36876
rect 12943 36873 12955 36907
rect 12897 36867 12955 36873
rect 13449 36907 13507 36913
rect 13449 36873 13461 36907
rect 13495 36904 13507 36907
rect 13495 36876 14780 36904
rect 13495 36873 13507 36876
rect 13449 36867 13507 36873
rect 9732 36808 10824 36836
rect 9732 36796 9738 36808
rect 9585 36771 9643 36777
rect 9585 36737 9597 36771
rect 9631 36737 9643 36771
rect 9585 36731 9643 36737
rect 10229 36771 10287 36777
rect 10229 36737 10241 36771
rect 10275 36737 10287 36771
rect 10410 36768 10416 36780
rect 10371 36740 10416 36768
rect 10229 36731 10287 36737
rect 4948 36672 6316 36700
rect 6549 36703 6607 36709
rect 4948 36660 4954 36672
rect 6549 36669 6561 36703
rect 6595 36700 6607 36703
rect 8478 36700 8484 36712
rect 6595 36672 6684 36700
rect 8439 36672 8484 36700
rect 6595 36669 6607 36672
rect 6549 36663 6607 36669
rect 3053 36635 3111 36641
rect 2464 36604 2774 36632
rect 2464 36592 2470 36604
rect 1394 36524 1400 36576
rect 1452 36564 1458 36576
rect 1489 36567 1547 36573
rect 1489 36564 1501 36567
rect 1452 36536 1501 36564
rect 1452 36524 1458 36536
rect 1489 36533 1501 36536
rect 1535 36533 1547 36567
rect 2314 36564 2320 36576
rect 2275 36536 2320 36564
rect 1489 36527 1547 36533
rect 2314 36524 2320 36536
rect 2372 36524 2378 36576
rect 2746 36564 2774 36604
rect 3053 36601 3065 36635
rect 3099 36601 3111 36635
rect 3053 36595 3111 36601
rect 3970 36592 3976 36644
rect 4028 36632 4034 36644
rect 5445 36635 5503 36641
rect 5445 36632 5457 36635
rect 4028 36604 5457 36632
rect 4028 36592 4034 36604
rect 5445 36601 5457 36604
rect 5491 36601 5503 36635
rect 5445 36595 5503 36601
rect 6656 36576 6684 36672
rect 8478 36660 8484 36672
rect 8536 36660 8542 36712
rect 8573 36703 8631 36709
rect 8573 36669 8585 36703
rect 8619 36700 8631 36703
rect 9030 36700 9036 36712
rect 8619 36672 9036 36700
rect 8619 36669 8631 36672
rect 8573 36663 8631 36669
rect 9030 36660 9036 36672
rect 9088 36660 9094 36712
rect 10244 36700 10272 36731
rect 10410 36728 10416 36740
rect 10468 36728 10474 36780
rect 10502 36728 10508 36780
rect 10560 36768 10566 36780
rect 10796 36777 10824 36808
rect 10965 36839 11023 36845
rect 10965 36805 10977 36839
rect 11011 36836 11023 36839
rect 11762 36839 11820 36845
rect 11762 36836 11774 36839
rect 11011 36808 11774 36836
rect 11011 36805 11023 36808
rect 10965 36799 11023 36805
rect 11762 36805 11774 36808
rect 11808 36805 11820 36839
rect 11762 36799 11820 36805
rect 13078 36796 13084 36848
rect 13136 36836 13142 36848
rect 13136 36808 13400 36836
rect 13136 36796 13142 36808
rect 10781 36771 10839 36777
rect 10560 36740 10605 36768
rect 10560 36728 10566 36740
rect 10781 36737 10793 36771
rect 10827 36737 10839 36771
rect 11514 36768 11520 36780
rect 11475 36740 11520 36768
rect 10781 36731 10839 36737
rect 11514 36728 11520 36740
rect 11572 36728 11578 36780
rect 13262 36768 13268 36780
rect 11624 36740 13268 36768
rect 10318 36700 10324 36712
rect 10244 36672 10324 36700
rect 10318 36660 10324 36672
rect 10376 36660 10382 36712
rect 10597 36703 10655 36709
rect 10597 36669 10609 36703
rect 10643 36700 10655 36703
rect 10686 36700 10692 36712
rect 10643 36672 10692 36700
rect 10643 36669 10655 36672
rect 10597 36663 10655 36669
rect 10686 36660 10692 36672
rect 10744 36660 10750 36712
rect 11624 36700 11652 36740
rect 13262 36728 13268 36740
rect 13320 36728 13326 36780
rect 13372 36777 13400 36808
rect 13357 36771 13415 36777
rect 13357 36737 13369 36771
rect 13403 36737 13415 36771
rect 13357 36731 13415 36737
rect 11532 36672 11652 36700
rect 7650 36592 7656 36644
rect 7708 36632 7714 36644
rect 8386 36632 8392 36644
rect 7708 36604 8392 36632
rect 7708 36592 7714 36604
rect 8386 36592 8392 36604
rect 8444 36632 8450 36644
rect 11532 36632 11560 36672
rect 8444 36604 11560 36632
rect 8444 36592 8450 36604
rect 4157 36567 4215 36573
rect 4157 36564 4169 36567
rect 2746 36536 4169 36564
rect 4157 36533 4169 36536
rect 4203 36533 4215 36567
rect 6638 36564 6644 36576
rect 6551 36536 6644 36564
rect 4157 36527 4215 36533
rect 6638 36524 6644 36536
rect 6696 36564 6702 36576
rect 9214 36564 9220 36576
rect 6696 36536 9220 36564
rect 6696 36524 6702 36536
rect 9214 36524 9220 36536
rect 9272 36564 9278 36576
rect 9582 36564 9588 36576
rect 9272 36536 9588 36564
rect 9272 36524 9278 36536
rect 9582 36524 9588 36536
rect 9640 36524 9646 36576
rect 9769 36567 9827 36573
rect 9769 36533 9781 36567
rect 9815 36564 9827 36567
rect 9950 36564 9956 36576
rect 9815 36536 9956 36564
rect 9815 36533 9827 36536
rect 9769 36527 9827 36533
rect 9950 36524 9956 36536
rect 10008 36524 10014 36576
rect 11882 36524 11888 36576
rect 11940 36564 11946 36576
rect 13464 36564 13492 36867
rect 14752 36836 14780 36876
rect 15102 36864 15108 36916
rect 15160 36904 15166 36916
rect 15749 36907 15807 36913
rect 15749 36904 15761 36907
rect 15160 36876 15761 36904
rect 15160 36864 15166 36876
rect 15749 36873 15761 36876
rect 15795 36873 15807 36907
rect 15749 36867 15807 36873
rect 16758 36864 16764 36916
rect 16816 36904 16822 36916
rect 17129 36907 17187 36913
rect 17129 36904 17141 36907
rect 16816 36876 17141 36904
rect 16816 36864 16822 36876
rect 17129 36873 17141 36876
rect 17175 36873 17187 36907
rect 17129 36867 17187 36873
rect 17497 36907 17555 36913
rect 17497 36873 17509 36907
rect 17543 36904 17555 36907
rect 17862 36904 17868 36916
rect 17543 36876 17868 36904
rect 17543 36873 17555 36876
rect 17497 36867 17555 36873
rect 17862 36864 17868 36876
rect 17920 36864 17926 36916
rect 14752 36808 15516 36836
rect 14182 36768 14188 36780
rect 14143 36740 14188 36768
rect 14182 36728 14188 36740
rect 14240 36728 14246 36780
rect 14550 36768 14556 36780
rect 14511 36740 14556 36768
rect 14550 36728 14556 36740
rect 14608 36728 14614 36780
rect 14826 36728 14832 36780
rect 14884 36768 14890 36780
rect 15488 36777 15516 36808
rect 19058 36796 19064 36848
rect 19116 36836 19122 36848
rect 20438 36836 20444 36848
rect 19116 36808 20444 36836
rect 19116 36796 19122 36808
rect 20438 36796 20444 36808
rect 20496 36836 20502 36848
rect 20496 36808 20668 36836
rect 20496 36796 20502 36808
rect 15197 36774 15255 36777
rect 15028 36771 15255 36774
rect 15028 36768 15209 36771
rect 14884 36746 15209 36768
rect 14884 36740 15056 36746
rect 14884 36728 14890 36740
rect 15197 36737 15209 36746
rect 15243 36737 15255 36771
rect 15197 36731 15255 36737
rect 15473 36771 15531 36777
rect 15473 36737 15485 36771
rect 15519 36737 15531 36771
rect 15473 36731 15531 36737
rect 15565 36771 15623 36777
rect 15565 36737 15577 36771
rect 15611 36737 15623 36771
rect 15565 36731 15623 36737
rect 18325 36771 18383 36777
rect 18325 36737 18337 36771
rect 18371 36768 18383 36771
rect 18414 36768 18420 36780
rect 18371 36740 18420 36768
rect 18371 36737 18383 36740
rect 18325 36731 18383 36737
rect 14090 36660 14096 36712
rect 14148 36700 14154 36712
rect 14642 36700 14648 36712
rect 14148 36672 14648 36700
rect 14148 36660 14154 36672
rect 14642 36660 14648 36672
rect 14700 36700 14706 36712
rect 14737 36703 14795 36709
rect 14737 36700 14749 36703
rect 14700 36672 14749 36700
rect 14700 36660 14706 36672
rect 14737 36669 14749 36672
rect 14783 36669 14795 36703
rect 15286 36700 15292 36712
rect 15247 36672 15292 36700
rect 14737 36663 14795 36669
rect 15286 36660 15292 36672
rect 15344 36660 15350 36712
rect 15580 36700 15608 36731
rect 18414 36728 18420 36740
rect 18472 36728 18478 36780
rect 18598 36777 18604 36780
rect 18592 36731 18604 36777
rect 18656 36768 18662 36780
rect 20530 36768 20536 36780
rect 18656 36740 18692 36768
rect 20491 36740 20536 36768
rect 18598 36728 18604 36731
rect 18656 36728 18662 36740
rect 20530 36728 20536 36740
rect 20588 36728 20594 36780
rect 20640 36768 20668 36808
rect 20640 36740 20760 36768
rect 15488 36672 15608 36700
rect 14277 36635 14335 36641
rect 14277 36601 14289 36635
rect 14323 36601 14335 36635
rect 14277 36595 14335 36601
rect 11940 36536 13492 36564
rect 14292 36564 14320 36595
rect 14366 36592 14372 36644
rect 14424 36632 14430 36644
rect 14424 36604 15332 36632
rect 14424 36592 14430 36604
rect 15194 36564 15200 36576
rect 14292 36536 15200 36564
rect 11940 36524 11946 36536
rect 15194 36524 15200 36536
rect 15252 36524 15258 36576
rect 15304 36564 15332 36604
rect 15488 36564 15516 36672
rect 16758 36660 16764 36712
rect 16816 36700 16822 36712
rect 16853 36703 16911 36709
rect 16853 36700 16865 36703
rect 16816 36672 16865 36700
rect 16816 36660 16822 36672
rect 16853 36669 16865 36672
rect 16899 36669 16911 36703
rect 17034 36700 17040 36712
rect 16995 36672 17040 36700
rect 16853 36663 16911 36669
rect 17034 36660 17040 36672
rect 17092 36660 17098 36712
rect 20622 36700 20628 36712
rect 20583 36672 20628 36700
rect 20622 36660 20628 36672
rect 20680 36660 20686 36712
rect 20732 36709 20760 36740
rect 21358 36728 21364 36780
rect 21416 36768 21422 36780
rect 22002 36768 22008 36780
rect 21416 36740 22008 36768
rect 21416 36728 21422 36740
rect 22002 36728 22008 36740
rect 22060 36768 22066 36780
rect 22097 36771 22155 36777
rect 22097 36768 22109 36771
rect 22060 36740 22109 36768
rect 22060 36728 22066 36740
rect 22097 36737 22109 36740
rect 22143 36737 22155 36771
rect 30098 36768 30104 36780
rect 30059 36740 30104 36768
rect 22097 36731 22155 36737
rect 30098 36728 30104 36740
rect 30156 36728 30162 36780
rect 20717 36703 20775 36709
rect 20717 36669 20729 36703
rect 20763 36669 20775 36703
rect 20717 36663 20775 36669
rect 22281 36703 22339 36709
rect 22281 36669 22293 36703
rect 22327 36700 22339 36703
rect 22327 36672 26234 36700
rect 22327 36669 22339 36672
rect 22281 36663 22339 36669
rect 19705 36635 19763 36641
rect 19705 36601 19717 36635
rect 19751 36632 19763 36635
rect 19978 36632 19984 36644
rect 19751 36604 19984 36632
rect 19751 36601 19763 36604
rect 19705 36595 19763 36601
rect 19978 36592 19984 36604
rect 20036 36592 20042 36644
rect 26206 36632 26234 36672
rect 29917 36635 29975 36641
rect 29917 36632 29929 36635
rect 26206 36604 29929 36632
rect 29917 36601 29929 36604
rect 29963 36601 29975 36635
rect 29917 36595 29975 36601
rect 15304 36536 15516 36564
rect 19794 36524 19800 36576
rect 19852 36564 19858 36576
rect 20165 36567 20223 36573
rect 20165 36564 20177 36567
rect 19852 36536 20177 36564
rect 19852 36524 19858 36536
rect 20165 36533 20177 36536
rect 20211 36533 20223 36567
rect 20165 36527 20223 36533
rect 20806 36524 20812 36576
rect 20864 36564 20870 36576
rect 21913 36567 21971 36573
rect 21913 36564 21925 36567
rect 20864 36536 21925 36564
rect 20864 36524 20870 36536
rect 21913 36533 21925 36536
rect 21959 36533 21971 36567
rect 21913 36527 21971 36533
rect 1104 36474 30820 36496
rect 1104 36422 5915 36474
rect 5967 36422 5979 36474
rect 6031 36422 6043 36474
rect 6095 36422 6107 36474
rect 6159 36422 6171 36474
rect 6223 36422 15846 36474
rect 15898 36422 15910 36474
rect 15962 36422 15974 36474
rect 16026 36422 16038 36474
rect 16090 36422 16102 36474
rect 16154 36422 25776 36474
rect 25828 36422 25840 36474
rect 25892 36422 25904 36474
rect 25956 36422 25968 36474
rect 26020 36422 26032 36474
rect 26084 36422 30820 36474
rect 1104 36400 30820 36422
rect 5166 36360 5172 36372
rect 5127 36332 5172 36360
rect 5166 36320 5172 36332
rect 5224 36320 5230 36372
rect 7190 36360 7196 36372
rect 7151 36332 7196 36360
rect 7190 36320 7196 36332
rect 7248 36320 7254 36372
rect 9766 36360 9772 36372
rect 9727 36332 9772 36360
rect 9766 36320 9772 36332
rect 9824 36320 9830 36372
rect 10410 36320 10416 36372
rect 10468 36360 10474 36372
rect 10468 36332 10536 36360
rect 10468 36320 10474 36332
rect 3789 36295 3847 36301
rect 3789 36261 3801 36295
rect 3835 36261 3847 36295
rect 3789 36255 3847 36261
rect 4709 36295 4767 36301
rect 4709 36261 4721 36295
rect 4755 36292 4767 36295
rect 9674 36292 9680 36304
rect 4755 36264 9680 36292
rect 4755 36261 4767 36264
rect 4709 36255 4767 36261
rect 1670 36156 1676 36168
rect 1631 36128 1676 36156
rect 1670 36116 1676 36128
rect 1728 36116 1734 36168
rect 2317 36159 2375 36165
rect 2317 36125 2329 36159
rect 2363 36125 2375 36159
rect 2317 36119 2375 36125
rect 2777 36159 2835 36165
rect 2777 36125 2789 36159
rect 2823 36156 2835 36159
rect 3804 36156 3832 36255
rect 9674 36252 9680 36264
rect 9732 36252 9738 36304
rect 4264 36196 5396 36224
rect 4264 36168 4292 36196
rect 2823 36128 3832 36156
rect 3973 36159 4031 36165
rect 2823 36125 2835 36128
rect 2777 36119 2835 36125
rect 3973 36125 3985 36159
rect 4019 36156 4031 36159
rect 4246 36156 4252 36168
rect 4019 36128 4252 36156
rect 4019 36125 4031 36128
rect 3973 36119 4031 36125
rect 2332 36088 2360 36119
rect 4246 36116 4252 36128
rect 4304 36116 4310 36168
rect 5368 36165 5396 36196
rect 5534 36184 5540 36236
rect 5592 36224 5598 36236
rect 6365 36227 6423 36233
rect 6365 36224 6377 36227
rect 5592 36196 6377 36224
rect 5592 36184 5598 36196
rect 6365 36193 6377 36196
rect 6411 36224 6423 36227
rect 6454 36224 6460 36236
rect 6411 36196 6460 36224
rect 6411 36193 6423 36196
rect 6365 36187 6423 36193
rect 6454 36184 6460 36196
rect 6512 36184 6518 36236
rect 6638 36224 6644 36236
rect 6599 36196 6644 36224
rect 6638 36184 6644 36196
rect 6696 36184 6702 36236
rect 6730 36184 6736 36236
rect 6788 36224 6794 36236
rect 10042 36224 10048 36236
rect 6788 36196 10048 36224
rect 6788 36184 6794 36196
rect 10042 36184 10048 36196
rect 10100 36184 10106 36236
rect 4525 36159 4583 36165
rect 4525 36125 4537 36159
rect 4571 36125 4583 36159
rect 4525 36119 4583 36125
rect 5353 36159 5411 36165
rect 5353 36125 5365 36159
rect 5399 36125 5411 36159
rect 5353 36119 5411 36125
rect 7101 36159 7159 36165
rect 7101 36125 7113 36159
rect 7147 36125 7159 36159
rect 8018 36156 8024 36168
rect 7979 36128 8024 36156
rect 7101 36119 7159 36125
rect 3510 36088 3516 36100
rect 2332 36060 3516 36088
rect 3510 36048 3516 36060
rect 3568 36048 3574 36100
rect 4540 36088 4568 36119
rect 5442 36088 5448 36100
rect 4540 36060 5448 36088
rect 5442 36048 5448 36060
rect 5500 36048 5506 36100
rect 7116 36088 7144 36119
rect 8018 36116 8024 36128
rect 8076 36116 8082 36168
rect 9122 36156 9128 36168
rect 9083 36128 9128 36156
rect 9122 36116 9128 36128
rect 9180 36116 9186 36168
rect 9306 36116 9312 36168
rect 9364 36156 9370 36168
rect 9585 36159 9643 36165
rect 9585 36156 9597 36159
rect 9364 36128 9597 36156
rect 9364 36116 9370 36128
rect 9585 36125 9597 36128
rect 9631 36125 9643 36159
rect 10318 36156 10324 36168
rect 10279 36128 10324 36156
rect 9585 36119 9643 36125
rect 10318 36116 10324 36128
rect 10376 36116 10382 36168
rect 10508 36165 10536 36332
rect 10594 36320 10600 36372
rect 10652 36320 10658 36372
rect 10686 36320 10692 36372
rect 10744 36320 10750 36372
rect 11057 36363 11115 36369
rect 11057 36329 11069 36363
rect 11103 36360 11115 36363
rect 11238 36360 11244 36372
rect 11103 36332 11244 36360
rect 11103 36329 11115 36332
rect 11057 36323 11115 36329
rect 11238 36320 11244 36332
rect 11296 36320 11302 36372
rect 11330 36320 11336 36372
rect 11388 36360 11394 36372
rect 11388 36332 12434 36360
rect 11388 36320 11394 36332
rect 10612 36233 10640 36320
rect 10704 36233 10732 36320
rect 11514 36292 11520 36304
rect 11475 36264 11520 36292
rect 11514 36252 11520 36264
rect 11572 36252 11578 36304
rect 12406 36292 12434 36332
rect 13998 36320 14004 36372
rect 14056 36360 14062 36372
rect 14185 36363 14243 36369
rect 14185 36360 14197 36363
rect 14056 36332 14197 36360
rect 14056 36320 14062 36332
rect 14185 36329 14197 36332
rect 14231 36329 14243 36363
rect 16761 36363 16819 36369
rect 14185 36323 14243 36329
rect 14844 36332 16712 36360
rect 14844 36292 14872 36332
rect 15194 36292 15200 36304
rect 12406 36264 14872 36292
rect 14936 36264 15200 36292
rect 14936 36233 14964 36264
rect 15194 36252 15200 36264
rect 15252 36292 15258 36304
rect 16684 36292 16712 36332
rect 16761 36329 16773 36363
rect 16807 36360 16819 36363
rect 17034 36360 17040 36372
rect 16807 36332 17040 36360
rect 16807 36329 16819 36332
rect 16761 36323 16819 36329
rect 17034 36320 17040 36332
rect 17092 36320 17098 36372
rect 18598 36360 18604 36372
rect 18559 36332 18604 36360
rect 18598 36320 18604 36332
rect 18656 36320 18662 36372
rect 20533 36363 20591 36369
rect 20533 36329 20545 36363
rect 20579 36360 20591 36363
rect 20622 36360 20628 36372
rect 20579 36332 20628 36360
rect 20579 36329 20591 36332
rect 20533 36323 20591 36329
rect 20622 36320 20628 36332
rect 20680 36320 20686 36372
rect 19610 36292 19616 36304
rect 15252 36264 15700 36292
rect 16684 36264 19616 36292
rect 15252 36252 15258 36264
rect 10597 36227 10655 36233
rect 10597 36193 10609 36227
rect 10643 36193 10655 36227
rect 10597 36187 10655 36193
rect 10689 36227 10747 36233
rect 10689 36193 10701 36227
rect 10735 36193 10747 36227
rect 10689 36187 10747 36193
rect 14921 36227 14979 36233
rect 14921 36193 14933 36227
rect 14967 36193 14979 36227
rect 15102 36224 15108 36236
rect 15063 36196 15108 36224
rect 14921 36187 14979 36193
rect 15102 36184 15108 36196
rect 15160 36184 15166 36236
rect 15565 36227 15623 36233
rect 15565 36224 15577 36227
rect 15212 36196 15577 36224
rect 10505 36159 10563 36165
rect 10505 36125 10517 36159
rect 10551 36125 10563 36159
rect 10505 36119 10563 36125
rect 10873 36159 10931 36165
rect 10873 36125 10885 36159
rect 10919 36156 10931 36159
rect 11422 36156 11428 36168
rect 10919 36128 11428 36156
rect 10919 36125 10931 36128
rect 10873 36119 10931 36125
rect 10888 36088 10916 36119
rect 11422 36116 11428 36128
rect 11480 36116 11486 36168
rect 11698 36156 11704 36168
rect 11659 36128 11704 36156
rect 11698 36116 11704 36128
rect 11756 36116 11762 36168
rect 14093 36159 14151 36165
rect 14093 36125 14105 36159
rect 14139 36156 14151 36159
rect 14182 36156 14188 36168
rect 14139 36128 14188 36156
rect 14139 36125 14151 36128
rect 14093 36119 14151 36125
rect 14182 36116 14188 36128
rect 14240 36116 14246 36168
rect 14274 36116 14280 36168
rect 14332 36156 14338 36168
rect 14332 36128 14377 36156
rect 14332 36116 14338 36128
rect 15010 36116 15016 36168
rect 15068 36156 15074 36168
rect 15212 36156 15240 36196
rect 15565 36193 15577 36196
rect 15611 36193 15623 36227
rect 15672 36224 15700 36264
rect 19610 36252 19616 36264
rect 19668 36252 19674 36304
rect 15841 36227 15899 36233
rect 15841 36224 15853 36227
rect 15672 36196 15853 36224
rect 15565 36187 15623 36193
rect 15841 36193 15853 36196
rect 15887 36193 15899 36227
rect 15841 36187 15899 36193
rect 15979 36227 16037 36233
rect 15979 36193 15991 36227
rect 16025 36224 16037 36227
rect 16298 36224 16304 36236
rect 16025 36196 16304 36224
rect 16025 36193 16037 36196
rect 15979 36187 16037 36193
rect 16298 36184 16304 36196
rect 16356 36184 16362 36236
rect 20806 36224 20812 36236
rect 16684 36196 20812 36224
rect 16114 36156 16120 36168
rect 15068 36128 15240 36156
rect 16075 36128 16120 36156
rect 15068 36116 15074 36128
rect 16114 36116 16120 36128
rect 16172 36116 16178 36168
rect 7116 36060 10916 36088
rect 1486 36020 1492 36032
rect 1447 35992 1492 36020
rect 1486 35980 1492 35992
rect 1544 35980 1550 36032
rect 2133 36023 2191 36029
rect 2133 35989 2145 36023
rect 2179 36020 2191 36023
rect 2222 36020 2228 36032
rect 2179 35992 2228 36020
rect 2179 35989 2191 35992
rect 2133 35983 2191 35989
rect 2222 35980 2228 35992
rect 2280 35980 2286 36032
rect 2958 36020 2964 36032
rect 2919 35992 2964 36020
rect 2958 35980 2964 35992
rect 3016 35980 3022 36032
rect 3528 36020 3556 36048
rect 5074 36020 5080 36032
rect 3528 35992 5080 36020
rect 5074 35980 5080 35992
rect 5132 35980 5138 36032
rect 7466 35980 7472 36032
rect 7524 36020 7530 36032
rect 7561 36023 7619 36029
rect 7561 36020 7573 36023
rect 7524 35992 7573 36020
rect 7524 35980 7530 35992
rect 7561 35989 7573 35992
rect 7607 35989 7619 36023
rect 7561 35983 7619 35989
rect 8205 36023 8263 36029
rect 8205 35989 8217 36023
rect 8251 36020 8263 36023
rect 8386 36020 8392 36032
rect 8251 35992 8392 36020
rect 8251 35989 8263 35992
rect 8205 35983 8263 35989
rect 8386 35980 8392 35992
rect 8444 35980 8450 36032
rect 8938 36020 8944 36032
rect 8899 35992 8944 36020
rect 8938 35980 8944 35992
rect 8996 35980 9002 36032
rect 9030 35980 9036 36032
rect 9088 36020 9094 36032
rect 11330 36020 11336 36032
rect 9088 35992 11336 36020
rect 9088 35980 9094 35992
rect 11330 35980 11336 35992
rect 11388 35980 11394 36032
rect 13262 35980 13268 36032
rect 13320 36020 13326 36032
rect 16684 36020 16712 36196
rect 20806 36184 20812 36196
rect 20864 36184 20870 36236
rect 21358 36224 21364 36236
rect 21319 36196 21364 36224
rect 21358 36184 21364 36196
rect 21416 36184 21422 36236
rect 17497 36159 17555 36165
rect 17497 36125 17509 36159
rect 17543 36156 17555 36159
rect 18230 36156 18236 36168
rect 17543 36128 18236 36156
rect 17543 36125 17555 36128
rect 17497 36119 17555 36125
rect 18230 36116 18236 36128
rect 18288 36116 18294 36168
rect 18417 36159 18475 36165
rect 18417 36125 18429 36159
rect 18463 36125 18475 36159
rect 18598 36156 18604 36168
rect 18559 36128 18604 36156
rect 18417 36119 18475 36125
rect 18046 36048 18052 36100
rect 18104 36088 18110 36100
rect 18432 36088 18460 36119
rect 18598 36116 18604 36128
rect 18656 36116 18662 36168
rect 19886 36116 19892 36168
rect 19944 36156 19950 36168
rect 20070 36156 20076 36168
rect 19944 36128 20076 36156
rect 19944 36116 19950 36128
rect 20070 36116 20076 36128
rect 20128 36116 20134 36168
rect 20346 36156 20352 36168
rect 20307 36128 20352 36156
rect 20346 36116 20352 36128
rect 20404 36116 20410 36168
rect 21085 36159 21143 36165
rect 21085 36125 21097 36159
rect 21131 36156 21143 36159
rect 21542 36156 21548 36168
rect 21131 36128 21548 36156
rect 21131 36125 21143 36128
rect 21085 36119 21143 36125
rect 21542 36116 21548 36128
rect 21600 36116 21606 36168
rect 18104 36060 18460 36088
rect 18104 36048 18110 36060
rect 13320 35992 16712 36020
rect 13320 35980 13326 35992
rect 17218 35980 17224 36032
rect 17276 36020 17282 36032
rect 17313 36023 17371 36029
rect 17313 36020 17325 36023
rect 17276 35992 17325 36020
rect 17276 35980 17282 35992
rect 17313 35989 17325 35992
rect 17359 35989 17371 36023
rect 17313 35983 17371 35989
rect 19978 35980 19984 36032
rect 20036 36020 20042 36032
rect 20165 36023 20223 36029
rect 20165 36020 20177 36023
rect 20036 35992 20177 36020
rect 20036 35980 20042 35992
rect 20165 35989 20177 35992
rect 20211 35989 20223 36023
rect 20165 35983 20223 35989
rect 1104 35930 30820 35952
rect 1104 35878 10880 35930
rect 10932 35878 10944 35930
rect 10996 35878 11008 35930
rect 11060 35878 11072 35930
rect 11124 35878 11136 35930
rect 11188 35878 20811 35930
rect 20863 35878 20875 35930
rect 20927 35878 20939 35930
rect 20991 35878 21003 35930
rect 21055 35878 21067 35930
rect 21119 35878 30820 35930
rect 1104 35856 30820 35878
rect 2409 35819 2467 35825
rect 2409 35785 2421 35819
rect 2455 35816 2467 35819
rect 7009 35819 7067 35825
rect 2455 35788 6960 35816
rect 2455 35785 2467 35788
rect 2409 35779 2467 35785
rect 2225 35751 2283 35757
rect 2225 35717 2237 35751
rect 2271 35748 2283 35751
rect 6932 35748 6960 35788
rect 7009 35785 7021 35819
rect 7055 35816 7067 35819
rect 8018 35816 8024 35828
rect 7055 35788 8024 35816
rect 7055 35785 7067 35788
rect 7009 35779 7067 35785
rect 8018 35776 8024 35788
rect 8076 35776 8082 35828
rect 8205 35819 8263 35825
rect 8205 35785 8217 35819
rect 8251 35816 8263 35819
rect 9122 35816 9128 35828
rect 8251 35788 9128 35816
rect 8251 35785 8263 35788
rect 8205 35779 8263 35785
rect 9122 35776 9128 35788
rect 9180 35776 9186 35828
rect 11698 35816 11704 35828
rect 9232 35788 11704 35816
rect 9232 35748 9260 35788
rect 11698 35776 11704 35788
rect 11756 35776 11762 35828
rect 18230 35816 18236 35828
rect 18191 35788 18236 35816
rect 18230 35776 18236 35788
rect 18288 35776 18294 35828
rect 18598 35776 18604 35828
rect 18656 35816 18662 35828
rect 18969 35819 19027 35825
rect 18969 35816 18981 35819
rect 18656 35788 18981 35816
rect 18656 35776 18662 35788
rect 18969 35785 18981 35788
rect 19015 35785 19027 35819
rect 19150 35816 19156 35828
rect 19111 35788 19156 35816
rect 18969 35779 19027 35785
rect 19150 35776 19156 35788
rect 19208 35776 19214 35828
rect 20438 35776 20444 35828
rect 20496 35816 20502 35828
rect 20901 35819 20959 35825
rect 20901 35816 20913 35819
rect 20496 35788 20913 35816
rect 20496 35776 20502 35788
rect 20901 35785 20913 35788
rect 20947 35785 20959 35819
rect 20901 35779 20959 35785
rect 2271 35720 5764 35748
rect 6932 35720 9260 35748
rect 2271 35717 2283 35720
rect 2225 35711 2283 35717
rect 1854 35680 1860 35692
rect 1767 35652 1860 35680
rect 1854 35640 1860 35652
rect 1912 35680 1918 35692
rect 2406 35680 2412 35692
rect 1912 35652 2412 35680
rect 1912 35640 1918 35652
rect 2406 35640 2412 35652
rect 2464 35640 2470 35692
rect 2958 35640 2964 35692
rect 3016 35680 3022 35692
rect 3418 35689 3424 35692
rect 3145 35683 3203 35689
rect 3145 35680 3157 35683
rect 3016 35652 3157 35680
rect 3016 35640 3022 35652
rect 3145 35649 3157 35652
rect 3191 35649 3203 35683
rect 3145 35643 3203 35649
rect 3412 35643 3424 35689
rect 3476 35680 3482 35692
rect 3476 35652 3512 35680
rect 3418 35640 3424 35643
rect 3476 35640 3482 35652
rect 4430 35640 4436 35692
rect 4488 35680 4494 35692
rect 5169 35683 5227 35689
rect 5169 35680 5181 35683
rect 4488 35652 5181 35680
rect 4488 35640 4494 35652
rect 5169 35649 5181 35652
rect 5215 35649 5227 35683
rect 5169 35643 5227 35649
rect 5736 35612 5764 35720
rect 9674 35708 9680 35760
rect 9732 35708 9738 35760
rect 10410 35748 10416 35760
rect 9784 35720 10416 35748
rect 5813 35683 5871 35689
rect 5813 35649 5825 35683
rect 5859 35680 5871 35683
rect 6270 35680 6276 35692
rect 5859 35652 6276 35680
rect 5859 35649 5871 35652
rect 5813 35643 5871 35649
rect 6270 35640 6276 35652
rect 6328 35680 6334 35692
rect 6730 35680 6736 35692
rect 6328 35652 6736 35680
rect 6328 35640 6334 35652
rect 6730 35640 6736 35652
rect 6788 35640 6794 35692
rect 6825 35683 6883 35689
rect 6825 35649 6837 35683
rect 6871 35680 6883 35683
rect 7558 35680 7564 35692
rect 6871 35652 7564 35680
rect 6871 35649 6883 35652
rect 6825 35643 6883 35649
rect 7558 35640 7564 35652
rect 7616 35680 7622 35692
rect 8021 35683 8079 35689
rect 8021 35680 8033 35683
rect 7616 35652 8033 35680
rect 7616 35640 7622 35652
rect 8021 35649 8033 35652
rect 8067 35649 8079 35683
rect 8021 35643 8079 35649
rect 9401 35683 9459 35689
rect 9401 35649 9413 35683
rect 9447 35680 9459 35683
rect 9692 35680 9720 35708
rect 9784 35689 9812 35720
rect 10410 35708 10416 35720
rect 10468 35708 10474 35760
rect 20530 35748 20536 35760
rect 18984 35720 20536 35748
rect 18984 35692 19012 35720
rect 20530 35708 20536 35720
rect 20588 35708 20594 35760
rect 9447 35652 9720 35680
rect 9769 35683 9827 35689
rect 9447 35649 9459 35652
rect 9401 35643 9459 35649
rect 9769 35649 9781 35683
rect 9815 35649 9827 35683
rect 9769 35643 9827 35649
rect 9953 35683 10011 35689
rect 9953 35649 9965 35683
rect 9999 35680 10011 35683
rect 10042 35680 10048 35692
rect 9999 35652 10048 35680
rect 9999 35649 10011 35652
rect 9953 35643 10011 35649
rect 10042 35640 10048 35652
rect 10100 35640 10106 35692
rect 10778 35680 10784 35692
rect 10739 35652 10784 35680
rect 10778 35640 10784 35652
rect 10836 35640 10842 35692
rect 11514 35680 11520 35692
rect 11475 35652 11520 35680
rect 11514 35640 11520 35652
rect 11572 35640 11578 35692
rect 16390 35640 16396 35692
rect 16448 35680 16454 35692
rect 17037 35683 17095 35689
rect 17037 35680 17049 35683
rect 16448 35652 17049 35680
rect 16448 35640 16454 35652
rect 17037 35649 17049 35652
rect 17083 35649 17095 35683
rect 17865 35683 17923 35689
rect 17865 35680 17877 35683
rect 17037 35643 17095 35649
rect 17420 35652 17877 35680
rect 8754 35612 8760 35624
rect 5736 35584 8760 35612
rect 8754 35572 8760 35584
rect 8812 35572 8818 35624
rect 9585 35615 9643 35621
rect 9585 35581 9597 35615
rect 9631 35581 9643 35615
rect 9585 35575 9643 35581
rect 9677 35615 9735 35621
rect 9677 35581 9689 35615
rect 9723 35612 9735 35615
rect 10226 35612 10232 35624
rect 9723 35584 10232 35612
rect 9723 35581 9735 35584
rect 9677 35575 9735 35581
rect 9600 35544 9628 35575
rect 10226 35572 10232 35584
rect 10284 35572 10290 35624
rect 10318 35572 10324 35624
rect 10376 35612 10382 35624
rect 10376 35584 12434 35612
rect 10376 35572 10382 35584
rect 10686 35544 10692 35556
rect 9600 35516 10692 35544
rect 10686 35504 10692 35516
rect 10744 35504 10750 35556
rect 12406 35544 12434 35584
rect 14458 35572 14464 35624
rect 14516 35612 14522 35624
rect 16758 35612 16764 35624
rect 14516 35584 16764 35612
rect 14516 35572 14522 35584
rect 16758 35572 16764 35584
rect 16816 35572 16822 35624
rect 16850 35572 16856 35624
rect 16908 35612 16914 35624
rect 16945 35615 17003 35621
rect 16945 35612 16957 35615
rect 16908 35584 16957 35612
rect 16908 35572 16914 35584
rect 16945 35581 16957 35584
rect 16991 35581 17003 35615
rect 16945 35575 17003 35581
rect 17126 35544 17132 35556
rect 12406 35516 17132 35544
rect 17126 35504 17132 35516
rect 17184 35504 17190 35556
rect 17420 35488 17448 35652
rect 17865 35649 17877 35652
rect 17911 35649 17923 35683
rect 17865 35643 17923 35649
rect 17954 35640 17960 35692
rect 18012 35680 18018 35692
rect 18049 35683 18107 35689
rect 18049 35680 18061 35683
rect 18012 35652 18061 35680
rect 18012 35640 18018 35652
rect 18049 35649 18061 35652
rect 18095 35680 18107 35683
rect 18966 35680 18972 35692
rect 18095 35652 18972 35680
rect 18095 35649 18107 35652
rect 18049 35643 18107 35649
rect 18966 35640 18972 35652
rect 19024 35640 19030 35692
rect 19150 35683 19208 35689
rect 19150 35649 19162 35683
rect 19196 35680 19208 35683
rect 19794 35680 19800 35692
rect 19196 35652 19800 35680
rect 19196 35649 19208 35652
rect 19150 35643 19208 35649
rect 19794 35640 19800 35652
rect 19852 35640 19858 35692
rect 20073 35683 20131 35689
rect 20073 35649 20085 35683
rect 20119 35680 20131 35683
rect 20162 35680 20168 35692
rect 20119 35652 20168 35680
rect 20119 35649 20131 35652
rect 20073 35643 20131 35649
rect 20162 35640 20168 35652
rect 20220 35640 20226 35692
rect 20257 35683 20315 35689
rect 20257 35649 20269 35683
rect 20303 35680 20315 35683
rect 20346 35680 20352 35692
rect 20303 35652 20352 35680
rect 20303 35649 20315 35652
rect 20257 35643 20315 35649
rect 20346 35640 20352 35652
rect 20404 35640 20410 35692
rect 20809 35683 20867 35689
rect 20809 35649 20821 35683
rect 20855 35680 20867 35683
rect 21542 35680 21548 35692
rect 20855 35652 21548 35680
rect 20855 35649 20867 35652
rect 20809 35643 20867 35649
rect 21542 35640 21548 35652
rect 21600 35640 21606 35692
rect 19518 35572 19524 35624
rect 19576 35612 19582 35624
rect 19613 35615 19671 35621
rect 19613 35612 19625 35615
rect 19576 35584 19625 35612
rect 19576 35572 19582 35584
rect 19613 35581 19625 35584
rect 19659 35581 19671 35615
rect 19613 35575 19671 35581
rect 2222 35476 2228 35488
rect 2183 35448 2228 35476
rect 2222 35436 2228 35448
rect 2280 35436 2286 35488
rect 3786 35436 3792 35488
rect 3844 35476 3850 35488
rect 4525 35479 4583 35485
rect 4525 35476 4537 35479
rect 3844 35448 4537 35476
rect 3844 35436 3850 35448
rect 4525 35445 4537 35448
rect 4571 35445 4583 35479
rect 4525 35439 4583 35445
rect 4890 35436 4896 35488
rect 4948 35476 4954 35488
rect 4985 35479 5043 35485
rect 4985 35476 4997 35479
rect 4948 35448 4997 35476
rect 4948 35436 4954 35448
rect 4985 35445 4997 35448
rect 5031 35445 5043 35479
rect 4985 35439 5043 35445
rect 5534 35436 5540 35488
rect 5592 35476 5598 35488
rect 5629 35479 5687 35485
rect 5629 35476 5641 35479
rect 5592 35448 5641 35476
rect 5592 35436 5598 35448
rect 5629 35445 5641 35448
rect 5675 35445 5687 35479
rect 9214 35476 9220 35488
rect 9175 35448 9220 35476
rect 5629 35439 5687 35445
rect 9214 35436 9220 35448
rect 9272 35436 9278 35488
rect 10594 35476 10600 35488
rect 10555 35448 10600 35476
rect 10594 35436 10600 35448
rect 10652 35436 10658 35488
rect 11701 35479 11759 35485
rect 11701 35445 11713 35479
rect 11747 35476 11759 35479
rect 17310 35476 17316 35488
rect 11747 35448 17316 35476
rect 11747 35445 11759 35448
rect 11701 35439 11759 35445
rect 17310 35436 17316 35448
rect 17368 35436 17374 35488
rect 17402 35436 17408 35488
rect 17460 35476 17466 35488
rect 17460 35448 17505 35476
rect 17460 35436 17466 35448
rect 19426 35436 19432 35488
rect 19484 35476 19490 35488
rect 19521 35479 19579 35485
rect 19521 35476 19533 35479
rect 19484 35448 19533 35476
rect 19484 35436 19490 35448
rect 19521 35445 19533 35448
rect 19567 35445 19579 35479
rect 19521 35439 19579 35445
rect 20165 35479 20223 35485
rect 20165 35445 20177 35479
rect 20211 35476 20223 35479
rect 20622 35476 20628 35488
rect 20211 35448 20628 35476
rect 20211 35445 20223 35448
rect 20165 35439 20223 35445
rect 20622 35436 20628 35448
rect 20680 35436 20686 35488
rect 1104 35386 30820 35408
rect 1104 35334 5915 35386
rect 5967 35334 5979 35386
rect 6031 35334 6043 35386
rect 6095 35334 6107 35386
rect 6159 35334 6171 35386
rect 6223 35334 15846 35386
rect 15898 35334 15910 35386
rect 15962 35334 15974 35386
rect 16026 35334 16038 35386
rect 16090 35334 16102 35386
rect 16154 35334 25776 35386
rect 25828 35334 25840 35386
rect 25892 35334 25904 35386
rect 25956 35334 25968 35386
rect 26020 35334 26032 35386
rect 26084 35334 30820 35386
rect 1104 35312 30820 35334
rect 2222 35272 2228 35284
rect 2183 35244 2228 35272
rect 2222 35232 2228 35244
rect 2280 35232 2286 35284
rect 4430 35272 4436 35284
rect 4391 35244 4436 35272
rect 4430 35232 4436 35244
rect 4488 35232 4494 35284
rect 4908 35244 8432 35272
rect 1854 35204 1860 35216
rect 1815 35176 1860 35204
rect 1854 35164 1860 35176
rect 1912 35164 1918 35216
rect 2409 35207 2467 35213
rect 2409 35173 2421 35207
rect 2455 35204 2467 35207
rect 4908 35204 4936 35244
rect 2455 35176 4936 35204
rect 8404 35204 8432 35244
rect 8662 35232 8668 35284
rect 8720 35272 8726 35284
rect 10042 35272 10048 35284
rect 8720 35244 10048 35272
rect 8720 35232 8726 35244
rect 10042 35232 10048 35244
rect 10100 35232 10106 35284
rect 10778 35272 10784 35284
rect 10739 35244 10784 35272
rect 10778 35232 10784 35244
rect 10836 35232 10842 35284
rect 12434 35272 12440 35284
rect 11716 35244 12440 35272
rect 8846 35204 8852 35216
rect 8404 35176 8852 35204
rect 2455 35173 2467 35176
rect 2409 35167 2467 35173
rect 8846 35164 8852 35176
rect 8904 35164 8910 35216
rect 4890 35136 4896 35148
rect 3160 35108 4752 35136
rect 4851 35108 4896 35136
rect 3160 35077 3188 35108
rect 3145 35071 3203 35077
rect 3145 35037 3157 35071
rect 3191 35037 3203 35071
rect 4246 35068 4252 35080
rect 4207 35040 4252 35068
rect 3145 35031 3203 35037
rect 4246 35028 4252 35040
rect 4304 35028 4310 35080
rect 4724 35068 4752 35108
rect 4890 35096 4896 35108
rect 4948 35096 4954 35148
rect 8386 35136 8392 35148
rect 8347 35108 8392 35136
rect 8386 35096 8392 35108
rect 8444 35096 8450 35148
rect 8938 35136 8944 35148
rect 8899 35108 8944 35136
rect 8938 35096 8944 35108
rect 8996 35096 9002 35148
rect 11716 35145 11744 35244
rect 12434 35232 12440 35244
rect 12492 35232 12498 35284
rect 13078 35272 13084 35284
rect 13039 35244 13084 35272
rect 13078 35232 13084 35244
rect 13136 35232 13142 35284
rect 15562 35272 15568 35284
rect 15212 35244 15568 35272
rect 11701 35139 11759 35145
rect 11701 35105 11713 35139
rect 11747 35105 11759 35139
rect 13096 35136 13124 35232
rect 15212 35213 15240 35244
rect 15562 35232 15568 35244
rect 15620 35232 15626 35284
rect 16390 35272 16396 35284
rect 16351 35244 16396 35272
rect 16390 35232 16396 35244
rect 16448 35232 16454 35284
rect 20346 35232 20352 35284
rect 20404 35272 20410 35284
rect 20993 35275 21051 35281
rect 20993 35272 21005 35275
rect 20404 35244 21005 35272
rect 20404 35232 20410 35244
rect 20993 35241 21005 35244
rect 21039 35241 21051 35275
rect 20993 35235 21051 35241
rect 15197 35207 15255 35213
rect 15197 35173 15209 35207
rect 15243 35173 15255 35207
rect 15197 35167 15255 35173
rect 18693 35207 18751 35213
rect 18693 35173 18705 35207
rect 18739 35204 18751 35207
rect 20162 35204 20168 35216
rect 18739 35176 20168 35204
rect 18739 35173 18751 35176
rect 18693 35167 18751 35173
rect 20162 35164 20168 35176
rect 20220 35164 20226 35216
rect 13722 35136 13728 35148
rect 13096 35108 13728 35136
rect 11701 35099 11759 35105
rect 13722 35096 13728 35108
rect 13780 35136 13786 35148
rect 14737 35139 14795 35145
rect 14737 35136 14749 35139
rect 13780 35108 14749 35136
rect 13780 35096 13786 35108
rect 14737 35105 14749 35108
rect 14783 35105 14795 35139
rect 14737 35099 14795 35105
rect 15286 35096 15292 35148
rect 15344 35136 15350 35148
rect 15590 35139 15648 35145
rect 15590 35136 15602 35139
rect 15344 35108 15602 35136
rect 15344 35096 15350 35108
rect 15590 35105 15602 35108
rect 15636 35105 15648 35139
rect 17310 35136 17316 35148
rect 17271 35108 17316 35136
rect 15590 35099 15648 35105
rect 17310 35096 17316 35108
rect 17368 35096 17374 35148
rect 20349 35139 20407 35145
rect 20349 35105 20361 35139
rect 20395 35136 20407 35139
rect 20438 35136 20444 35148
rect 20395 35108 20444 35136
rect 20395 35105 20407 35108
rect 20349 35099 20407 35105
rect 20438 35096 20444 35108
rect 20496 35096 20502 35148
rect 20622 35096 20628 35148
rect 20680 35136 20686 35148
rect 20680 35108 21220 35136
rect 20680 35096 20686 35108
rect 6362 35068 6368 35080
rect 4724 35040 6368 35068
rect 6362 35028 6368 35040
rect 6420 35028 6426 35080
rect 9214 35077 9220 35080
rect 9208 35068 9220 35077
rect 9175 35040 9220 35068
rect 9208 35031 9220 35040
rect 9214 35028 9220 35031
rect 9272 35028 9278 35080
rect 9950 35028 9956 35080
rect 10008 35068 10014 35080
rect 10965 35071 11023 35077
rect 10965 35068 10977 35071
rect 10008 35040 10977 35068
rect 10008 35028 10014 35040
rect 10965 35037 10977 35040
rect 11011 35068 11023 35071
rect 14366 35068 14372 35080
rect 11011 35040 14372 35068
rect 11011 35037 11023 35040
rect 10965 35031 11023 35037
rect 14366 35028 14372 35040
rect 14424 35028 14430 35080
rect 14553 35071 14611 35077
rect 14553 35037 14565 35071
rect 14599 35068 14611 35071
rect 14642 35068 14648 35080
rect 14599 35040 14648 35068
rect 14599 35037 14611 35040
rect 14553 35031 14611 35037
rect 14642 35028 14648 35040
rect 14700 35028 14706 35080
rect 15470 35028 15476 35080
rect 15528 35068 15534 35080
rect 15746 35068 15752 35080
rect 15528 35040 15573 35068
rect 15707 35040 15752 35068
rect 15528 35028 15534 35040
rect 15746 35028 15752 35040
rect 15804 35028 15810 35080
rect 20162 35028 20168 35080
rect 20220 35068 20226 35080
rect 21192 35077 21220 35108
rect 20901 35071 20959 35077
rect 20901 35068 20913 35071
rect 20220 35040 20913 35068
rect 20220 35028 20226 35040
rect 20901 35037 20913 35040
rect 20947 35037 20959 35071
rect 20901 35031 20959 35037
rect 21177 35071 21235 35077
rect 21177 35037 21189 35071
rect 21223 35037 21235 35071
rect 21177 35031 21235 35037
rect 2225 35003 2283 35009
rect 2225 34969 2237 35003
rect 2271 35000 2283 35003
rect 3786 35000 3792 35012
rect 2271 34972 3792 35000
rect 2271 34969 2283 34972
rect 2225 34963 2283 34969
rect 3786 34960 3792 34972
rect 3844 34960 3850 35012
rect 4706 34960 4712 35012
rect 4764 35000 4770 35012
rect 5138 35003 5196 35009
rect 5138 35000 5150 35003
rect 4764 34972 5150 35000
rect 4764 34960 4770 34972
rect 5138 34969 5150 34972
rect 5184 34969 5196 35003
rect 5138 34963 5196 34969
rect 7650 34960 7656 35012
rect 7708 35000 7714 35012
rect 8122 35003 8180 35009
rect 8122 35000 8134 35003
rect 7708 34972 8134 35000
rect 7708 34960 7714 34972
rect 8122 34969 8134 34972
rect 8168 34969 8180 35003
rect 8122 34963 8180 34969
rect 11968 35003 12026 35009
rect 11968 34969 11980 35003
rect 12014 35000 12026 35003
rect 12066 35000 12072 35012
rect 12014 34972 12072 35000
rect 12014 34969 12026 34972
rect 11968 34963 12026 34969
rect 12066 34960 12072 34972
rect 12124 34960 12130 35012
rect 2958 34932 2964 34944
rect 2919 34904 2964 34932
rect 2958 34892 2964 34904
rect 3016 34892 3022 34944
rect 4890 34892 4896 34944
rect 4948 34932 4954 34944
rect 6273 34935 6331 34941
rect 6273 34932 6285 34935
rect 4948 34904 6285 34932
rect 4948 34892 4954 34904
rect 6273 34901 6285 34904
rect 6319 34901 6331 34935
rect 7006 34932 7012 34944
rect 6967 34904 7012 34932
rect 6273 34895 6331 34901
rect 7006 34892 7012 34904
rect 7064 34892 7070 34944
rect 9674 34892 9680 34944
rect 9732 34932 9738 34944
rect 10321 34935 10379 34941
rect 10321 34932 10333 34935
rect 9732 34904 10333 34932
rect 9732 34892 9738 34904
rect 10321 34901 10333 34904
rect 10367 34932 10379 34935
rect 10502 34932 10508 34944
rect 10367 34904 10508 34932
rect 10367 34901 10379 34904
rect 10321 34895 10379 34901
rect 10502 34892 10508 34904
rect 10560 34892 10566 34944
rect 14660 34932 14688 35028
rect 17580 35003 17638 35009
rect 17580 34969 17592 35003
rect 17626 35000 17638 35003
rect 18230 35000 18236 35012
rect 17626 34972 18236 35000
rect 17626 34969 17638 34972
rect 17580 34963 17638 34969
rect 18230 34960 18236 34972
rect 18288 34960 18294 35012
rect 15470 34932 15476 34944
rect 14660 34904 15476 34932
rect 15470 34892 15476 34904
rect 15528 34892 15534 34944
rect 19702 34932 19708 34944
rect 19663 34904 19708 34932
rect 19702 34892 19708 34904
rect 19760 34892 19766 34944
rect 20070 34932 20076 34944
rect 20031 34904 20076 34932
rect 20070 34892 20076 34904
rect 20128 34892 20134 34944
rect 20165 34935 20223 34941
rect 20165 34901 20177 34935
rect 20211 34932 20223 34935
rect 21361 34935 21419 34941
rect 21361 34932 21373 34935
rect 20211 34904 21373 34932
rect 20211 34901 20223 34904
rect 20165 34895 20223 34901
rect 21361 34901 21373 34904
rect 21407 34901 21419 34935
rect 21361 34895 21419 34901
rect 1104 34842 30820 34864
rect 1104 34790 10880 34842
rect 10932 34790 10944 34842
rect 10996 34790 11008 34842
rect 11060 34790 11072 34842
rect 11124 34790 11136 34842
rect 11188 34790 20811 34842
rect 20863 34790 20875 34842
rect 20927 34790 20939 34842
rect 20991 34790 21003 34842
rect 21055 34790 21067 34842
rect 21119 34790 30820 34842
rect 1104 34768 30820 34790
rect 1762 34688 1768 34740
rect 1820 34728 1826 34740
rect 1857 34731 1915 34737
rect 1857 34728 1869 34731
rect 1820 34700 1869 34728
rect 1820 34688 1826 34700
rect 1857 34697 1869 34700
rect 1903 34697 1915 34731
rect 1857 34691 1915 34697
rect 3418 34688 3424 34740
rect 3476 34728 3482 34740
rect 3513 34731 3571 34737
rect 3513 34728 3525 34731
rect 3476 34700 3525 34728
rect 3476 34688 3482 34700
rect 3513 34697 3525 34700
rect 3559 34697 3571 34731
rect 4706 34728 4712 34740
rect 4667 34700 4712 34728
rect 3513 34691 3571 34697
rect 4706 34688 4712 34700
rect 4764 34688 4770 34740
rect 7561 34731 7619 34737
rect 7561 34697 7573 34731
rect 7607 34728 7619 34731
rect 7650 34728 7656 34740
rect 7607 34700 7656 34728
rect 7607 34697 7619 34700
rect 7561 34691 7619 34697
rect 7650 34688 7656 34700
rect 7708 34688 7714 34740
rect 10318 34688 10324 34740
rect 10376 34728 10382 34740
rect 11609 34731 11667 34737
rect 11609 34728 11621 34731
rect 10376 34700 11621 34728
rect 10376 34688 10382 34700
rect 11609 34697 11621 34700
rect 11655 34697 11667 34731
rect 11609 34691 11667 34697
rect 16117 34731 16175 34737
rect 16117 34697 16129 34731
rect 16163 34728 16175 34731
rect 16850 34728 16856 34740
rect 16163 34700 16856 34728
rect 16163 34697 16175 34700
rect 16117 34691 16175 34697
rect 16850 34688 16856 34700
rect 16908 34688 16914 34740
rect 16945 34731 17003 34737
rect 16945 34697 16957 34731
rect 16991 34728 17003 34731
rect 17034 34728 17040 34740
rect 16991 34700 17040 34728
rect 16991 34697 17003 34700
rect 16945 34691 17003 34697
rect 17034 34688 17040 34700
rect 17092 34688 17098 34740
rect 17218 34688 17224 34740
rect 17276 34728 17282 34740
rect 17313 34731 17371 34737
rect 17313 34728 17325 34731
rect 17276 34700 17325 34728
rect 17276 34688 17282 34700
rect 17313 34697 17325 34700
rect 17359 34697 17371 34731
rect 17313 34691 17371 34697
rect 17402 34688 17408 34740
rect 17460 34728 17466 34740
rect 18230 34728 18236 34740
rect 17460 34700 17505 34728
rect 18191 34700 18236 34728
rect 17460 34688 17466 34700
rect 18230 34688 18236 34700
rect 18288 34688 18294 34740
rect 18877 34731 18935 34737
rect 18877 34697 18889 34731
rect 18923 34697 18935 34731
rect 18877 34691 18935 34697
rect 19061 34731 19119 34737
rect 19061 34697 19073 34731
rect 19107 34728 19119 34731
rect 19150 34728 19156 34740
rect 19107 34700 19156 34728
rect 19107 34697 19119 34700
rect 19061 34691 19119 34697
rect 2041 34663 2099 34669
rect 2041 34629 2053 34663
rect 2087 34660 2099 34663
rect 6914 34660 6920 34672
rect 2087 34632 4936 34660
rect 2087 34629 2099 34632
rect 2041 34623 2099 34629
rect 4908 34604 4936 34632
rect 5736 34632 6920 34660
rect 5736 34604 5764 34632
rect 6914 34620 6920 34632
rect 6972 34620 6978 34672
rect 9766 34660 9772 34672
rect 9232 34632 9772 34660
rect 2406 34592 2412 34604
rect 2367 34564 2412 34592
rect 2406 34552 2412 34564
rect 2464 34552 2470 34604
rect 2866 34592 2872 34604
rect 2827 34564 2872 34592
rect 2866 34552 2872 34564
rect 2924 34552 2930 34604
rect 3697 34595 3755 34601
rect 3697 34561 3709 34595
rect 3743 34592 3755 34595
rect 3786 34592 3792 34604
rect 3743 34564 3792 34592
rect 3743 34561 3755 34564
rect 3697 34555 3755 34561
rect 3786 34552 3792 34564
rect 3844 34552 3850 34604
rect 4062 34592 4068 34604
rect 4023 34564 4068 34592
rect 4062 34552 4068 34564
rect 4120 34552 4126 34604
rect 4249 34595 4307 34601
rect 4249 34561 4261 34595
rect 4295 34592 4307 34595
rect 4338 34592 4344 34604
rect 4295 34564 4344 34592
rect 4295 34561 4307 34564
rect 4249 34555 4307 34561
rect 4338 34552 4344 34564
rect 4396 34552 4402 34604
rect 4890 34592 4896 34604
rect 4851 34564 4896 34592
rect 4890 34552 4896 34564
rect 4948 34552 4954 34604
rect 5074 34592 5080 34604
rect 5035 34564 5080 34592
rect 5074 34552 5080 34564
rect 5132 34552 5138 34604
rect 5258 34592 5264 34604
rect 5219 34564 5264 34592
rect 5258 34552 5264 34564
rect 5316 34552 5322 34604
rect 5445 34595 5503 34601
rect 5445 34561 5457 34595
rect 5491 34592 5503 34595
rect 5718 34592 5724 34604
rect 5491 34564 5724 34592
rect 5491 34561 5503 34564
rect 5445 34555 5503 34561
rect 5718 34552 5724 34564
rect 5776 34552 5782 34604
rect 6365 34595 6423 34601
rect 6365 34561 6377 34595
rect 6411 34592 6423 34595
rect 7006 34592 7012 34604
rect 6411 34564 7012 34592
rect 6411 34561 6423 34564
rect 6365 34555 6423 34561
rect 7006 34552 7012 34564
rect 7064 34592 7070 34604
rect 7745 34595 7803 34601
rect 7745 34592 7757 34595
rect 7064 34564 7757 34592
rect 7064 34552 7070 34564
rect 7745 34561 7757 34564
rect 7791 34561 7803 34595
rect 7745 34555 7803 34561
rect 8113 34595 8171 34601
rect 8113 34561 8125 34595
rect 8159 34592 8171 34595
rect 8202 34592 8208 34604
rect 8159 34564 8208 34592
rect 8159 34561 8171 34564
rect 8113 34555 8171 34561
rect 8202 34552 8208 34564
rect 8260 34552 8266 34604
rect 8297 34595 8355 34601
rect 8297 34561 8309 34595
rect 8343 34592 8355 34595
rect 8662 34592 8668 34604
rect 8343 34564 8668 34592
rect 8343 34561 8355 34564
rect 8297 34555 8355 34561
rect 8662 34552 8668 34564
rect 8720 34552 8726 34604
rect 9232 34601 9260 34632
rect 9766 34620 9772 34632
rect 9824 34660 9830 34672
rect 12434 34660 12440 34672
rect 9824 34632 10640 34660
rect 9824 34620 9830 34632
rect 9217 34595 9275 34601
rect 9217 34561 9229 34595
rect 9263 34561 9275 34595
rect 10226 34592 10232 34604
rect 10187 34564 10232 34592
rect 9217 34555 9275 34561
rect 10226 34552 10232 34564
rect 10284 34552 10290 34604
rect 10410 34592 10416 34604
rect 10371 34564 10416 34592
rect 10410 34552 10416 34564
rect 10468 34552 10474 34604
rect 10612 34601 10640 34632
rect 12360 34632 12440 34660
rect 10597 34595 10655 34601
rect 10597 34561 10609 34595
rect 10643 34592 10655 34595
rect 10686 34592 10692 34604
rect 10643 34564 10692 34592
rect 10643 34561 10655 34564
rect 10597 34555 10655 34561
rect 10686 34552 10692 34564
rect 10744 34552 10750 34604
rect 10781 34595 10839 34601
rect 10781 34561 10793 34595
rect 10827 34592 10839 34595
rect 11238 34592 11244 34604
rect 10827 34564 11244 34592
rect 10827 34561 10839 34564
rect 10781 34555 10839 34561
rect 11238 34552 11244 34564
rect 11296 34552 11302 34604
rect 11514 34552 11520 34604
rect 11572 34592 11578 34604
rect 12360 34601 12388 34632
rect 12434 34620 12440 34632
rect 12492 34620 12498 34672
rect 13722 34620 13728 34672
rect 13780 34660 13786 34672
rect 13780 34632 14504 34660
rect 13780 34620 13786 34632
rect 11793 34595 11851 34601
rect 11793 34592 11805 34595
rect 11572 34564 11805 34592
rect 11572 34552 11578 34564
rect 11793 34561 11805 34564
rect 11839 34561 11851 34595
rect 11793 34555 11851 34561
rect 12345 34595 12403 34601
rect 12345 34561 12357 34595
rect 12391 34561 12403 34595
rect 12345 34555 12403 34561
rect 12612 34595 12670 34601
rect 12612 34561 12624 34595
rect 12658 34592 12670 34595
rect 14090 34592 14096 34604
rect 12658 34564 14096 34592
rect 12658 34561 12670 34564
rect 12612 34555 12670 34561
rect 14090 34552 14096 34564
rect 14148 34552 14154 34604
rect 14476 34601 14504 34632
rect 14461 34595 14519 34601
rect 14461 34561 14473 34595
rect 14507 34561 14519 34595
rect 14461 34555 14519 34561
rect 15286 34552 15292 34604
rect 15344 34601 15350 34604
rect 15344 34595 15372 34601
rect 15360 34561 15372 34595
rect 15344 34555 15372 34561
rect 15344 34552 15350 34555
rect 18046 34552 18052 34604
rect 18104 34592 18110 34604
rect 18141 34595 18199 34601
rect 18141 34592 18153 34595
rect 18104 34564 18153 34592
rect 18104 34552 18110 34564
rect 18141 34561 18153 34564
rect 18187 34561 18199 34595
rect 18141 34555 18199 34561
rect 18325 34595 18383 34601
rect 18325 34561 18337 34595
rect 18371 34592 18383 34595
rect 18892 34592 18920 34691
rect 19150 34688 19156 34700
rect 19208 34688 19214 34740
rect 19518 34620 19524 34672
rect 19576 34660 19582 34672
rect 20257 34663 20315 34669
rect 20257 34660 20269 34663
rect 19576 34632 20269 34660
rect 19576 34620 19582 34632
rect 20257 34629 20269 34632
rect 20303 34629 20315 34663
rect 20257 34623 20315 34629
rect 18371 34564 18920 34592
rect 19058 34595 19116 34601
rect 18371 34561 18383 34564
rect 18325 34555 18383 34561
rect 19058 34561 19070 34595
rect 19104 34592 19116 34595
rect 19702 34592 19708 34604
rect 19104 34564 19708 34592
rect 19104 34561 19116 34564
rect 19058 34555 19116 34561
rect 19702 34552 19708 34564
rect 19760 34552 19766 34604
rect 19794 34552 19800 34604
rect 19852 34592 19858 34604
rect 19978 34592 19984 34604
rect 19852 34564 19984 34592
rect 19852 34552 19858 34564
rect 19978 34552 19984 34564
rect 20036 34592 20042 34604
rect 20165 34595 20223 34601
rect 20165 34592 20177 34595
rect 20036 34564 20177 34592
rect 20036 34552 20042 34564
rect 20165 34561 20177 34564
rect 20211 34561 20223 34595
rect 30098 34592 30104 34604
rect 30059 34564 30104 34592
rect 20165 34555 20223 34561
rect 30098 34552 30104 34564
rect 30156 34552 30162 34604
rect 3881 34527 3939 34533
rect 3881 34493 3893 34527
rect 3927 34493 3939 34527
rect 3881 34487 3939 34493
rect 3973 34527 4031 34533
rect 3973 34493 3985 34527
rect 4019 34524 4031 34527
rect 5169 34527 5227 34533
rect 5169 34524 5181 34527
rect 4019 34496 5181 34524
rect 4019 34493 4031 34496
rect 3973 34487 4031 34493
rect 3896 34456 3924 34487
rect 4080 34468 4108 34496
rect 5169 34493 5181 34496
rect 5215 34493 5227 34527
rect 5169 34487 5227 34493
rect 6825 34527 6883 34533
rect 6825 34493 6837 34527
rect 6871 34524 6883 34527
rect 7282 34524 7288 34536
rect 6871 34496 7288 34524
rect 6871 34493 6883 34496
rect 6825 34487 6883 34493
rect 7282 34484 7288 34496
rect 7340 34484 7346 34536
rect 7929 34527 7987 34533
rect 7929 34493 7941 34527
rect 7975 34493 7987 34527
rect 7929 34487 7987 34493
rect 3896 34428 4016 34456
rect 3988 34400 4016 34428
rect 4062 34416 4068 34468
rect 4120 34416 4126 34468
rect 7944 34456 7972 34487
rect 8018 34484 8024 34536
rect 8076 34524 8082 34536
rect 8938 34524 8944 34536
rect 8076 34496 8121 34524
rect 8899 34496 8944 34524
rect 8076 34484 8082 34496
rect 8938 34484 8944 34496
rect 8996 34484 9002 34536
rect 9674 34484 9680 34536
rect 9732 34524 9738 34536
rect 10505 34527 10563 34533
rect 10505 34524 10517 34527
rect 9732 34496 10517 34524
rect 9732 34484 9738 34496
rect 10505 34493 10517 34496
rect 10551 34493 10563 34527
rect 10505 34487 10563 34493
rect 14277 34527 14335 34533
rect 14277 34493 14289 34527
rect 14323 34524 14335 34527
rect 14642 34524 14648 34536
rect 14323 34496 14648 34524
rect 14323 34493 14335 34496
rect 14277 34487 14335 34493
rect 14642 34484 14648 34496
rect 14700 34524 14706 34536
rect 15197 34527 15255 34533
rect 15197 34524 15209 34527
rect 14700 34496 15209 34524
rect 14700 34484 14706 34496
rect 15197 34493 15209 34496
rect 15243 34493 15255 34527
rect 15197 34487 15255 34493
rect 15473 34527 15531 34533
rect 15473 34493 15485 34527
rect 15519 34524 15531 34527
rect 15654 34524 15660 34536
rect 15519 34496 15660 34524
rect 15519 34493 15531 34496
rect 15473 34487 15531 34493
rect 15654 34484 15660 34496
rect 15712 34524 15718 34536
rect 17586 34524 17592 34536
rect 15712 34496 17592 34524
rect 15712 34484 15718 34496
rect 17586 34484 17592 34496
rect 17644 34484 17650 34536
rect 19426 34524 19432 34536
rect 19387 34496 19432 34524
rect 19426 34484 19432 34496
rect 19484 34484 19490 34536
rect 19521 34527 19579 34533
rect 19521 34493 19533 34527
rect 19567 34524 19579 34527
rect 20254 34524 20260 34536
rect 19567 34496 20260 34524
rect 19567 34493 19579 34496
rect 19521 34487 19579 34493
rect 20254 34484 20260 34496
rect 20312 34484 20318 34536
rect 29822 34524 29828 34536
rect 29783 34496 29828 34524
rect 29822 34484 29828 34496
rect 29880 34484 29886 34536
rect 8956 34456 8984 34484
rect 14921 34459 14979 34465
rect 7944 34428 8984 34456
rect 9048 34428 11100 34456
rect 2041 34391 2099 34397
rect 2041 34357 2053 34391
rect 2087 34388 2099 34391
rect 2222 34388 2228 34400
rect 2087 34360 2228 34388
rect 2087 34357 2099 34360
rect 2041 34351 2099 34357
rect 2222 34348 2228 34360
rect 2280 34348 2286 34400
rect 3050 34388 3056 34400
rect 3011 34360 3056 34388
rect 3050 34348 3056 34360
rect 3108 34348 3114 34400
rect 3970 34388 3976 34400
rect 3883 34360 3976 34388
rect 3970 34348 3976 34360
rect 4028 34388 4034 34400
rect 5074 34388 5080 34400
rect 4028 34360 5080 34388
rect 4028 34348 4034 34360
rect 5074 34348 5080 34360
rect 5132 34348 5138 34400
rect 6454 34388 6460 34400
rect 6415 34360 6460 34388
rect 6454 34348 6460 34360
rect 6512 34348 6518 34400
rect 7374 34348 7380 34400
rect 7432 34388 7438 34400
rect 9048 34388 9076 34428
rect 7432 34360 9076 34388
rect 7432 34348 7438 34360
rect 10870 34348 10876 34400
rect 10928 34388 10934 34400
rect 10965 34391 11023 34397
rect 10965 34388 10977 34391
rect 10928 34360 10977 34388
rect 10928 34348 10934 34360
rect 10965 34357 10977 34360
rect 11011 34357 11023 34391
rect 11072 34388 11100 34428
rect 13648 34428 14872 34456
rect 13648 34388 13676 34428
rect 11072 34360 13676 34388
rect 13725 34391 13783 34397
rect 10965 34351 11023 34357
rect 13725 34357 13737 34391
rect 13771 34388 13783 34391
rect 14458 34388 14464 34400
rect 13771 34360 14464 34388
rect 13771 34357 13783 34360
rect 13725 34351 13783 34357
rect 14458 34348 14464 34360
rect 14516 34348 14522 34400
rect 14844 34388 14872 34428
rect 14921 34425 14933 34459
rect 14967 34456 14979 34459
rect 15010 34456 15016 34468
rect 14967 34428 15016 34456
rect 14967 34425 14979 34428
rect 14921 34419 14979 34425
rect 15010 34416 15016 34428
rect 15068 34416 15074 34468
rect 19334 34416 19340 34468
rect 19392 34456 19398 34468
rect 19978 34456 19984 34468
rect 19392 34428 19984 34456
rect 19392 34416 19398 34428
rect 19978 34416 19984 34428
rect 20036 34416 20042 34468
rect 20438 34388 20444 34400
rect 14844 34360 20444 34388
rect 20438 34348 20444 34360
rect 20496 34348 20502 34400
rect 1104 34298 30820 34320
rect 1104 34246 5915 34298
rect 5967 34246 5979 34298
rect 6031 34246 6043 34298
rect 6095 34246 6107 34298
rect 6159 34246 6171 34298
rect 6223 34246 15846 34298
rect 15898 34246 15910 34298
rect 15962 34246 15974 34298
rect 16026 34246 16038 34298
rect 16090 34246 16102 34298
rect 16154 34246 25776 34298
rect 25828 34246 25840 34298
rect 25892 34246 25904 34298
rect 25956 34246 25968 34298
rect 26020 34246 26032 34298
rect 26084 34246 30820 34298
rect 1104 34224 30820 34246
rect 2222 34184 2228 34196
rect 2183 34156 2228 34184
rect 2222 34144 2228 34156
rect 2280 34144 2286 34196
rect 6089 34187 6147 34193
rect 6089 34153 6101 34187
rect 6135 34184 6147 34187
rect 6270 34184 6276 34196
rect 6135 34156 6276 34184
rect 6135 34153 6147 34156
rect 6089 34147 6147 34153
rect 6270 34144 6276 34156
rect 6328 34144 6334 34196
rect 7558 34184 7564 34196
rect 7519 34156 7564 34184
rect 7558 34144 7564 34156
rect 7616 34144 7622 34196
rect 7650 34144 7656 34196
rect 7708 34184 7714 34196
rect 20714 34184 20720 34196
rect 7708 34156 20720 34184
rect 7708 34144 7714 34156
rect 20714 34144 20720 34156
rect 20772 34184 20778 34196
rect 20772 34156 21772 34184
rect 20772 34144 20778 34156
rect 1857 34119 1915 34125
rect 1857 34085 1869 34119
rect 1903 34116 1915 34119
rect 2406 34116 2412 34128
rect 1903 34088 2412 34116
rect 1903 34085 1915 34088
rect 1857 34079 1915 34085
rect 2406 34076 2412 34088
rect 2464 34076 2470 34128
rect 4798 34076 4804 34128
rect 4856 34116 4862 34128
rect 5350 34116 5356 34128
rect 4856 34088 5356 34116
rect 4856 34076 4862 34088
rect 5350 34076 5356 34088
rect 5408 34116 5414 34128
rect 9674 34116 9680 34128
rect 5408 34088 9680 34116
rect 5408 34076 5414 34088
rect 9674 34076 9680 34088
rect 9732 34076 9738 34128
rect 10134 34076 10140 34128
rect 10192 34076 10198 34128
rect 12526 34076 12532 34128
rect 12584 34116 12590 34128
rect 14090 34116 14096 34128
rect 12584 34088 13584 34116
rect 14051 34088 14096 34116
rect 12584 34076 12590 34088
rect 3050 34008 3056 34060
rect 3108 34048 3114 34060
rect 3789 34051 3847 34057
rect 3789 34048 3801 34051
rect 3108 34020 3801 34048
rect 3108 34008 3114 34020
rect 3789 34017 3801 34020
rect 3835 34017 3847 34051
rect 8294 34048 8300 34060
rect 3789 34011 3847 34017
rect 6932 34020 8300 34048
rect 3145 33983 3203 33989
rect 3145 33949 3157 33983
rect 3191 33980 3203 33983
rect 3878 33980 3884 33992
rect 3191 33952 3884 33980
rect 3191 33949 3203 33952
rect 3145 33943 3203 33949
rect 3878 33940 3884 33952
rect 3936 33940 3942 33992
rect 6932 33989 6960 34020
rect 8294 34008 8300 34020
rect 8352 34008 8358 34060
rect 9766 34048 9772 34060
rect 9727 34020 9772 34048
rect 9766 34008 9772 34020
rect 9824 34008 9830 34060
rect 9861 34051 9919 34057
rect 9861 34017 9873 34051
rect 9907 34048 9919 34051
rect 10152 34048 10180 34076
rect 10594 34048 10600 34060
rect 9907 34020 10180 34048
rect 10555 34020 10600 34048
rect 9907 34017 9919 34020
rect 9861 34011 9919 34017
rect 10594 34008 10600 34020
rect 10652 34008 10658 34060
rect 13446 34048 13452 34060
rect 12452 34020 13452 34048
rect 6273 33983 6331 33989
rect 6273 33949 6285 33983
rect 6319 33949 6331 33983
rect 6273 33943 6331 33949
rect 6917 33983 6975 33989
rect 6917 33949 6929 33983
rect 6963 33949 6975 33983
rect 6917 33943 6975 33949
rect 7377 33983 7435 33989
rect 7377 33949 7389 33983
rect 7423 33980 7435 33983
rect 7650 33980 7656 33992
rect 7423 33952 7656 33980
rect 7423 33949 7435 33952
rect 7377 33943 7435 33949
rect 2225 33915 2283 33921
rect 2225 33881 2237 33915
rect 2271 33912 2283 33915
rect 2271 33884 3556 33912
rect 2271 33881 2283 33884
rect 2225 33875 2283 33881
rect 2409 33847 2467 33853
rect 2409 33813 2421 33847
rect 2455 33844 2467 33847
rect 2774 33844 2780 33856
rect 2455 33816 2780 33844
rect 2455 33813 2467 33816
rect 2409 33807 2467 33813
rect 2774 33804 2780 33816
rect 2832 33804 2838 33856
rect 2958 33844 2964 33856
rect 2919 33816 2964 33844
rect 2958 33804 2964 33816
rect 3016 33804 3022 33856
rect 3528 33844 3556 33884
rect 3602 33872 3608 33924
rect 3660 33912 3666 33924
rect 4034 33915 4092 33921
rect 4034 33912 4046 33915
rect 3660 33884 4046 33912
rect 3660 33872 3666 33884
rect 4034 33881 4046 33884
rect 4080 33881 4092 33915
rect 6288 33912 6316 33943
rect 7650 33940 7656 33952
rect 7708 33940 7714 33992
rect 8202 33980 8208 33992
rect 8163 33952 8208 33980
rect 8202 33940 8208 33952
rect 8260 33940 8266 33992
rect 9585 33983 9643 33989
rect 9585 33949 9597 33983
rect 9631 33980 9643 33983
rect 9674 33980 9680 33992
rect 9631 33952 9680 33980
rect 9631 33949 9643 33952
rect 9585 33943 9643 33949
rect 9674 33940 9680 33952
rect 9732 33940 9738 33992
rect 9953 33983 10011 33989
rect 9953 33949 9965 33983
rect 9999 33949 10011 33983
rect 9953 33943 10011 33949
rect 10137 33983 10195 33989
rect 10137 33949 10149 33983
rect 10183 33980 10195 33983
rect 10686 33980 10692 33992
rect 10183 33952 10692 33980
rect 10183 33949 10195 33952
rect 10137 33943 10195 33949
rect 8386 33912 8392 33924
rect 6288 33884 8392 33912
rect 4034 33875 4092 33881
rect 8386 33872 8392 33884
rect 8444 33872 8450 33924
rect 9968 33912 9996 33943
rect 10686 33940 10692 33952
rect 10744 33940 10750 33992
rect 10870 33989 10876 33992
rect 10864 33980 10876 33989
rect 10831 33952 10876 33980
rect 10864 33943 10876 33952
rect 10870 33940 10876 33943
rect 10928 33940 10934 33992
rect 12452 33989 12480 34020
rect 13446 34008 13452 34020
rect 13504 34008 13510 34060
rect 13556 34048 13584 34088
rect 14090 34076 14096 34088
rect 14148 34076 14154 34128
rect 14366 34076 14372 34128
rect 14424 34116 14430 34128
rect 15010 34116 15016 34128
rect 14424 34088 15016 34116
rect 14424 34076 14430 34088
rect 15010 34076 15016 34088
rect 15068 34116 15074 34128
rect 15657 34119 15715 34125
rect 15068 34088 15516 34116
rect 15068 34076 15074 34088
rect 13556 34020 14381 34048
rect 12437 33983 12495 33989
rect 12437 33949 12449 33983
rect 12483 33949 12495 33983
rect 12437 33943 12495 33949
rect 12526 33940 12532 33992
rect 12584 33980 12590 33992
rect 12986 33989 12992 33992
rect 12941 33983 12992 33989
rect 12584 33952 12629 33980
rect 12584 33940 12590 33952
rect 12941 33949 12953 33983
rect 12987 33949 12992 33983
rect 12941 33943 12992 33949
rect 12986 33940 12992 33943
rect 13044 33982 13050 33992
rect 14231 33983 14289 33989
rect 13044 33980 13135 33982
rect 14231 33980 14243 33983
rect 13044 33954 14243 33980
rect 13044 33940 13050 33954
rect 13096 33952 14243 33954
rect 14231 33949 14243 33952
rect 14277 33949 14289 33983
rect 14353 33980 14381 34020
rect 15488 33989 15516 34088
rect 15657 34085 15669 34119
rect 15703 34085 15715 34119
rect 15657 34079 15715 34085
rect 18601 34119 18659 34125
rect 18601 34085 18613 34119
rect 18647 34116 18659 34119
rect 19426 34116 19432 34128
rect 18647 34088 19432 34116
rect 18647 34085 18659 34088
rect 18601 34079 18659 34085
rect 14589 33983 14647 33989
rect 14589 33980 14601 33983
rect 14353 33952 14601 33980
rect 14231 33943 14289 33949
rect 14589 33949 14601 33952
rect 14635 33949 14647 33983
rect 14589 33943 14647 33949
rect 14737 33983 14795 33989
rect 14737 33949 14749 33983
rect 14783 33949 14795 33983
rect 14737 33943 14795 33949
rect 15473 33983 15531 33989
rect 15473 33949 15485 33983
rect 15519 33949 15531 33983
rect 15672 33980 15700 34079
rect 19426 34076 19432 34088
rect 19484 34076 19490 34128
rect 20438 34116 20444 34128
rect 20399 34088 20444 34116
rect 20438 34076 20444 34088
rect 20496 34076 20502 34128
rect 18064 34020 19932 34048
rect 16117 33983 16175 33989
rect 16117 33980 16129 33983
rect 15672 33952 16129 33980
rect 15473 33943 15531 33949
rect 16117 33949 16129 33952
rect 16163 33949 16175 33983
rect 16117 33943 16175 33949
rect 10410 33912 10416 33924
rect 9968 33884 10416 33912
rect 10410 33872 10416 33884
rect 10468 33872 10474 33924
rect 12710 33912 12716 33924
rect 12671 33884 12716 33912
rect 12710 33872 12716 33884
rect 12768 33872 12774 33924
rect 12802 33872 12808 33924
rect 12860 33912 12866 33924
rect 14366 33912 14372 33924
rect 12860 33884 12905 33912
rect 14327 33884 14372 33912
rect 12860 33872 12866 33884
rect 14366 33872 14372 33884
rect 14424 33872 14430 33924
rect 14458 33872 14464 33924
rect 14516 33912 14522 33924
rect 14516 33884 14561 33912
rect 14516 33872 14522 33884
rect 3786 33844 3792 33856
rect 3528 33816 3792 33844
rect 3786 33804 3792 33816
rect 3844 33844 3850 33856
rect 5169 33847 5227 33853
rect 5169 33844 5181 33847
rect 3844 33816 5181 33844
rect 3844 33804 3850 33816
rect 5169 33813 5181 33816
rect 5215 33813 5227 33847
rect 5169 33807 5227 33813
rect 6546 33804 6552 33856
rect 6604 33844 6610 33856
rect 6825 33847 6883 33853
rect 6825 33844 6837 33847
rect 6604 33816 6837 33844
rect 6604 33804 6610 33816
rect 6825 33813 6837 33816
rect 6871 33813 6883 33847
rect 6825 33807 6883 33813
rect 8297 33847 8355 33853
rect 8297 33813 8309 33847
rect 8343 33844 8355 33847
rect 8478 33844 8484 33856
rect 8343 33816 8484 33844
rect 8343 33813 8355 33816
rect 8297 33807 8355 33813
rect 8478 33804 8484 33816
rect 8536 33844 8542 33856
rect 8938 33844 8944 33856
rect 8536 33816 8944 33844
rect 8536 33804 8542 33816
rect 8938 33804 8944 33816
rect 8996 33804 9002 33856
rect 9398 33844 9404 33856
rect 9359 33816 9404 33844
rect 9398 33804 9404 33816
rect 9456 33804 9462 33856
rect 11238 33804 11244 33856
rect 11296 33844 11302 33856
rect 11977 33847 12035 33853
rect 11977 33844 11989 33847
rect 11296 33816 11989 33844
rect 11296 33804 11302 33816
rect 11977 33813 11989 33816
rect 12023 33813 12035 33847
rect 11977 33807 12035 33813
rect 13081 33847 13139 33853
rect 13081 33813 13093 33847
rect 13127 33844 13139 33847
rect 13170 33844 13176 33856
rect 13127 33816 13176 33844
rect 13127 33813 13139 33816
rect 13081 33807 13139 33813
rect 13170 33804 13176 33816
rect 13228 33804 13234 33856
rect 13446 33804 13452 33856
rect 13504 33844 13510 33856
rect 14752 33844 14780 33943
rect 17402 33940 17408 33992
rect 17460 33980 17466 33992
rect 18064 33989 18092 34020
rect 19904 33992 19932 34020
rect 17865 33983 17923 33989
rect 17865 33980 17877 33983
rect 17460 33952 17877 33980
rect 17460 33940 17466 33952
rect 17865 33949 17877 33952
rect 17911 33949 17923 33983
rect 17865 33943 17923 33949
rect 18049 33983 18107 33989
rect 18049 33949 18061 33983
rect 18095 33949 18107 33983
rect 18506 33980 18512 33992
rect 18467 33952 18512 33980
rect 18049 33943 18107 33949
rect 18506 33940 18512 33952
rect 18564 33940 18570 33992
rect 19886 33940 19892 33992
rect 19944 33980 19950 33992
rect 19981 33983 20039 33989
rect 19981 33980 19993 33983
rect 19944 33952 19993 33980
rect 19944 33940 19950 33952
rect 19981 33949 19993 33952
rect 20027 33949 20039 33983
rect 20622 33980 20628 33992
rect 20583 33952 20628 33980
rect 19981 33943 20039 33949
rect 20622 33940 20628 33952
rect 20680 33940 20686 33992
rect 21634 33980 21640 33992
rect 20916 33952 21640 33980
rect 17957 33915 18015 33921
rect 17957 33881 17969 33915
rect 18003 33912 18015 33915
rect 18874 33912 18880 33924
rect 18003 33884 18880 33912
rect 18003 33881 18015 33884
rect 17957 33875 18015 33881
rect 18874 33872 18880 33884
rect 18932 33872 18938 33924
rect 20916 33912 20944 33952
rect 21634 33940 21640 33952
rect 21692 33940 21698 33992
rect 21744 33989 21772 34156
rect 21729 33983 21787 33989
rect 21729 33949 21741 33983
rect 21775 33949 21787 33983
rect 21729 33943 21787 33949
rect 19904 33884 20944 33912
rect 20993 33915 21051 33921
rect 13504 33816 14780 33844
rect 16301 33847 16359 33853
rect 13504 33804 13510 33816
rect 16301 33813 16313 33847
rect 16347 33844 16359 33847
rect 16942 33844 16948 33856
rect 16347 33816 16948 33844
rect 16347 33813 16359 33816
rect 16301 33807 16359 33813
rect 16942 33804 16948 33816
rect 17000 33804 17006 33856
rect 19334 33804 19340 33856
rect 19392 33844 19398 33856
rect 19904 33853 19932 33884
rect 20993 33881 21005 33915
rect 21039 33912 21051 33915
rect 21174 33912 21180 33924
rect 21039 33884 21180 33912
rect 21039 33881 21051 33884
rect 20993 33875 21051 33881
rect 21174 33872 21180 33884
rect 21232 33872 21238 33924
rect 19889 33847 19947 33853
rect 19889 33844 19901 33847
rect 19392 33816 19901 33844
rect 19392 33804 19398 33816
rect 19889 33813 19901 33816
rect 19935 33813 19947 33847
rect 20714 33844 20720 33856
rect 20675 33816 20720 33844
rect 19889 33807 19947 33813
rect 20714 33804 20720 33816
rect 20772 33804 20778 33856
rect 20809 33847 20867 33853
rect 20809 33813 20821 33847
rect 20855 33844 20867 33847
rect 21266 33844 21272 33856
rect 20855 33816 21272 33844
rect 20855 33813 20867 33816
rect 20809 33807 20867 33813
rect 21266 33804 21272 33816
rect 21324 33804 21330 33856
rect 21913 33847 21971 33853
rect 21913 33813 21925 33847
rect 21959 33844 21971 33847
rect 22646 33844 22652 33856
rect 21959 33816 22652 33844
rect 21959 33813 21971 33816
rect 21913 33807 21971 33813
rect 22646 33804 22652 33816
rect 22704 33804 22710 33856
rect 1104 33754 30820 33776
rect 1104 33702 10880 33754
rect 10932 33702 10944 33754
rect 10996 33702 11008 33754
rect 11060 33702 11072 33754
rect 11124 33702 11136 33754
rect 11188 33702 20811 33754
rect 20863 33702 20875 33754
rect 20927 33702 20939 33754
rect 20991 33702 21003 33754
rect 21055 33702 21067 33754
rect 21119 33702 30820 33754
rect 1104 33680 30820 33702
rect 2866 33600 2872 33652
rect 2924 33640 2930 33652
rect 2961 33643 3019 33649
rect 2961 33640 2973 33643
rect 2924 33612 2973 33640
rect 2924 33600 2930 33612
rect 2961 33609 2973 33612
rect 3007 33609 3019 33643
rect 3602 33640 3608 33652
rect 3563 33612 3608 33640
rect 2961 33603 3019 33609
rect 3602 33600 3608 33612
rect 3660 33600 3666 33652
rect 5626 33600 5632 33652
rect 5684 33640 5690 33652
rect 6365 33643 6423 33649
rect 6365 33640 6377 33643
rect 5684 33612 6377 33640
rect 5684 33600 5690 33612
rect 6365 33609 6377 33612
rect 6411 33640 6423 33643
rect 7650 33640 7656 33652
rect 6411 33612 7656 33640
rect 6411 33609 6423 33612
rect 6365 33603 6423 33609
rect 7650 33600 7656 33612
rect 7708 33600 7714 33652
rect 7834 33600 7840 33652
rect 7892 33640 7898 33652
rect 8754 33640 8760 33652
rect 7892 33612 8760 33640
rect 7892 33600 7898 33612
rect 8754 33600 8760 33612
rect 8812 33600 8818 33652
rect 10686 33640 10692 33652
rect 8864 33612 10692 33640
rect 4798 33572 4804 33584
rect 4172 33544 4804 33572
rect 1673 33507 1731 33513
rect 1673 33473 1685 33507
rect 1719 33504 1731 33507
rect 2038 33504 2044 33516
rect 1719 33476 2044 33504
rect 1719 33473 1731 33476
rect 1673 33467 1731 33473
rect 2038 33464 2044 33476
rect 2096 33464 2102 33516
rect 2317 33507 2375 33513
rect 2317 33473 2329 33507
rect 2363 33473 2375 33507
rect 3142 33504 3148 33516
rect 3103 33476 3148 33504
rect 2317 33467 2375 33473
rect 2332 33368 2360 33467
rect 3142 33464 3148 33476
rect 3200 33464 3206 33516
rect 3786 33504 3792 33516
rect 3747 33476 3792 33504
rect 3786 33464 3792 33476
rect 3844 33464 3850 33516
rect 4062 33504 4068 33516
rect 4023 33476 4068 33504
rect 4062 33464 4068 33476
rect 4120 33464 4126 33516
rect 4172 33513 4200 33544
rect 4798 33532 4804 33544
rect 4856 33532 4862 33584
rect 7558 33532 7564 33584
rect 7616 33572 7622 33584
rect 7616 33544 8800 33572
rect 7616 33532 7622 33544
rect 4157 33507 4215 33513
rect 4157 33473 4169 33507
rect 4203 33473 4215 33507
rect 4338 33504 4344 33516
rect 4299 33476 4344 33504
rect 4157 33467 4215 33473
rect 4338 33464 4344 33476
rect 4396 33464 4402 33516
rect 5537 33507 5595 33513
rect 5537 33473 5549 33507
rect 5583 33504 5595 33507
rect 6270 33504 6276 33516
rect 5583 33476 6276 33504
rect 5583 33473 5595 33476
rect 5537 33467 5595 33473
rect 6270 33464 6276 33476
rect 6328 33464 6334 33516
rect 6546 33504 6552 33516
rect 6507 33476 6552 33504
rect 6546 33464 6552 33476
rect 6604 33464 6610 33516
rect 7742 33504 7748 33516
rect 7703 33476 7748 33504
rect 7742 33464 7748 33476
rect 7800 33464 7806 33516
rect 7834 33464 7840 33516
rect 7892 33504 7898 33516
rect 8021 33507 8079 33513
rect 8021 33504 8033 33507
rect 7892 33476 8033 33504
rect 7892 33464 7898 33476
rect 8021 33473 8033 33476
rect 8067 33473 8079 33507
rect 8021 33467 8079 33473
rect 8113 33507 8171 33513
rect 8113 33473 8125 33507
rect 8159 33473 8171 33507
rect 8113 33467 8171 33473
rect 8297 33507 8355 33513
rect 8297 33473 8309 33507
rect 8343 33504 8355 33507
rect 8662 33504 8668 33516
rect 8343 33476 8668 33504
rect 8343 33473 8355 33476
rect 8297 33467 8355 33473
rect 3970 33436 3976 33448
rect 3931 33408 3976 33436
rect 3970 33396 3976 33408
rect 4028 33396 4034 33448
rect 7929 33439 7987 33445
rect 7929 33405 7941 33439
rect 7975 33405 7987 33439
rect 8128 33436 8156 33467
rect 8662 33464 8668 33476
rect 8720 33464 8726 33516
rect 8772 33513 8800 33544
rect 8757 33507 8815 33513
rect 8757 33473 8769 33507
rect 8803 33473 8815 33507
rect 8757 33467 8815 33473
rect 8202 33436 8208 33448
rect 8115 33408 8208 33436
rect 7929 33399 7987 33405
rect 2332 33340 2774 33368
rect 1486 33300 1492 33312
rect 1447 33272 1492 33300
rect 1486 33260 1492 33272
rect 1544 33260 1550 33312
rect 2130 33300 2136 33312
rect 2091 33272 2136 33300
rect 2130 33260 2136 33272
rect 2188 33260 2194 33312
rect 2746 33300 2774 33340
rect 3142 33328 3148 33380
rect 3200 33368 3206 33380
rect 4246 33368 4252 33380
rect 3200 33340 4252 33368
rect 3200 33328 3206 33340
rect 4246 33328 4252 33340
rect 4304 33368 4310 33380
rect 5353 33371 5411 33377
rect 5353 33368 5365 33371
rect 4304 33340 5365 33368
rect 4304 33328 4310 33340
rect 5353 33337 5365 33340
rect 5399 33337 5411 33371
rect 7944 33368 7972 33399
rect 8202 33396 8208 33408
rect 8260 33436 8266 33448
rect 8680 33436 8708 33464
rect 8864 33436 8892 33612
rect 10686 33600 10692 33612
rect 10744 33600 10750 33652
rect 12710 33600 12716 33652
rect 12768 33640 12774 33652
rect 14277 33643 14335 33649
rect 14277 33640 14289 33643
rect 12768 33612 14289 33640
rect 12768 33600 12774 33612
rect 14277 33609 14289 33612
rect 14323 33640 14335 33643
rect 14918 33640 14924 33652
rect 14323 33612 14924 33640
rect 14323 33609 14335 33612
rect 14277 33603 14335 33609
rect 14918 33600 14924 33612
rect 14976 33600 14982 33652
rect 19521 33643 19579 33649
rect 17328 33612 18552 33640
rect 17328 33584 17356 33612
rect 9490 33532 9496 33584
rect 9548 33572 9554 33584
rect 14366 33572 14372 33584
rect 9548 33544 14372 33572
rect 9548 33532 9554 33544
rect 14366 33532 14372 33544
rect 14424 33532 14430 33584
rect 15381 33575 15439 33581
rect 15381 33541 15393 33575
rect 15427 33572 15439 33575
rect 15562 33572 15568 33584
rect 15427 33544 15568 33572
rect 15427 33541 15439 33544
rect 15381 33535 15439 33541
rect 15562 33532 15568 33544
rect 15620 33572 15626 33584
rect 16390 33572 16396 33584
rect 15620 33544 16396 33572
rect 15620 33532 15626 33544
rect 16390 33532 16396 33544
rect 16448 33532 16454 33584
rect 17310 33572 17316 33584
rect 17223 33544 17316 33572
rect 17310 33532 17316 33544
rect 17368 33532 17374 33584
rect 18322 33572 18328 33584
rect 18283 33544 18328 33572
rect 18322 33532 18328 33544
rect 18380 33532 18386 33584
rect 18524 33581 18552 33612
rect 19521 33609 19533 33643
rect 19567 33640 19579 33643
rect 19886 33640 19892 33652
rect 19567 33612 19892 33640
rect 19567 33609 19579 33612
rect 19521 33603 19579 33609
rect 19886 33600 19892 33612
rect 19944 33600 19950 33652
rect 19981 33643 20039 33649
rect 19981 33609 19993 33643
rect 20027 33640 20039 33643
rect 20027 33612 20668 33640
rect 20027 33609 20039 33612
rect 19981 33603 20039 33609
rect 20640 33581 20668 33612
rect 20714 33600 20720 33652
rect 20772 33640 20778 33652
rect 21266 33640 21272 33652
rect 20772 33612 20865 33640
rect 20916 33612 21272 33640
rect 20772 33600 20778 33612
rect 18509 33575 18567 33581
rect 18509 33541 18521 33575
rect 18555 33572 18567 33575
rect 20625 33575 20683 33581
rect 18555 33544 20300 33572
rect 18555 33541 18567 33544
rect 18509 33535 18567 33541
rect 9585 33507 9643 33513
rect 9585 33504 9597 33507
rect 8260 33408 8616 33436
rect 8680 33408 8892 33436
rect 8956 33476 9597 33504
rect 8260 33396 8266 33408
rect 8478 33368 8484 33380
rect 7944 33340 8484 33368
rect 5353 33331 5411 33337
rect 8478 33328 8484 33340
rect 8536 33328 8542 33380
rect 4154 33300 4160 33312
rect 2746 33272 4160 33300
rect 4154 33260 4160 33272
rect 4212 33260 4218 33312
rect 7098 33260 7104 33312
rect 7156 33300 7162 33312
rect 7561 33303 7619 33309
rect 7561 33300 7573 33303
rect 7156 33272 7573 33300
rect 7156 33260 7162 33272
rect 7561 33269 7573 33272
rect 7607 33269 7619 33303
rect 8588 33300 8616 33408
rect 8956 33377 8984 33476
rect 9585 33473 9597 33476
rect 9631 33473 9643 33507
rect 9585 33467 9643 33473
rect 10321 33507 10379 33513
rect 10321 33473 10333 33507
rect 10367 33504 10379 33507
rect 10410 33504 10416 33516
rect 10367 33476 10416 33504
rect 10367 33473 10379 33476
rect 10321 33467 10379 33473
rect 10410 33464 10416 33476
rect 10468 33464 10474 33516
rect 10686 33464 10692 33516
rect 10744 33504 10750 33516
rect 11793 33507 11851 33513
rect 11793 33504 11805 33507
rect 10744 33476 11805 33504
rect 10744 33464 10750 33476
rect 11793 33473 11805 33476
rect 11839 33473 11851 33507
rect 11793 33467 11851 33473
rect 12342 33464 12348 33516
rect 12400 33504 12406 33516
rect 12802 33504 12808 33516
rect 12400 33476 12808 33504
rect 12400 33464 12406 33476
rect 12802 33464 12808 33476
rect 12860 33464 12866 33516
rect 13170 33513 13176 33516
rect 13164 33504 13176 33513
rect 13131 33476 13176 33504
rect 13164 33467 13176 33476
rect 13170 33464 13176 33467
rect 13228 33464 13234 33516
rect 13446 33464 13452 33516
rect 13504 33504 13510 33516
rect 15013 33507 15071 33513
rect 15013 33504 15025 33507
rect 13504 33476 15025 33504
rect 13504 33464 13510 33476
rect 15013 33473 15025 33476
rect 15059 33473 15071 33507
rect 15013 33467 15071 33473
rect 15106 33507 15164 33513
rect 15106 33473 15118 33507
rect 15152 33473 15164 33507
rect 15286 33504 15292 33516
rect 15247 33476 15292 33504
rect 15106 33467 15164 33473
rect 10045 33439 10103 33445
rect 10045 33405 10057 33439
rect 10091 33405 10103 33439
rect 11514 33436 11520 33448
rect 11475 33408 11520 33436
rect 10045 33399 10103 33405
rect 8941 33371 8999 33377
rect 8941 33337 8953 33371
rect 8987 33337 8999 33371
rect 10060 33368 10088 33399
rect 11514 33396 11520 33408
rect 11572 33396 11578 33448
rect 12434 33396 12440 33448
rect 12492 33436 12498 33448
rect 12894 33436 12900 33448
rect 12492 33408 12900 33436
rect 12492 33396 12498 33408
rect 12894 33396 12900 33408
rect 12952 33396 12958 33448
rect 15120 33436 15148 33467
rect 15286 33464 15292 33476
rect 15344 33464 15350 33516
rect 15470 33464 15476 33516
rect 15528 33513 15534 33516
rect 15528 33504 15536 33513
rect 17497 33507 17555 33513
rect 15528 33476 15573 33504
rect 15528 33467 15536 33476
rect 17497 33473 17509 33507
rect 17543 33504 17555 33507
rect 17954 33504 17960 33516
rect 17543 33476 17960 33504
rect 17543 33473 17555 33476
rect 17497 33467 17555 33473
rect 15528 33464 15534 33467
rect 17954 33464 17960 33476
rect 18012 33464 18018 33516
rect 19334 33464 19340 33516
rect 19392 33504 19398 33516
rect 19613 33507 19671 33513
rect 19613 33504 19625 33507
rect 19392 33476 19625 33504
rect 19392 33464 19398 33476
rect 19613 33473 19625 33476
rect 19659 33473 19671 33507
rect 19613 33467 19671 33473
rect 19705 33507 19763 33513
rect 19705 33473 19717 33507
rect 19751 33504 19763 33507
rect 20162 33504 20168 33516
rect 19751 33476 20168 33504
rect 19751 33473 19763 33476
rect 19705 33467 19763 33473
rect 20162 33464 20168 33476
rect 20220 33464 20226 33516
rect 17129 33439 17187 33445
rect 17129 33436 17141 33439
rect 15120 33408 17141 33436
rect 17129 33405 17141 33408
rect 17175 33405 17187 33439
rect 17129 33399 17187 33405
rect 18233 33439 18291 33445
rect 18233 33405 18245 33439
rect 18279 33436 18291 33439
rect 19521 33439 19579 33445
rect 19521 33436 19533 33439
rect 18279 33408 19533 33436
rect 18279 33405 18291 33408
rect 18233 33399 18291 33405
rect 19521 33405 19533 33408
rect 19567 33405 19579 33439
rect 20272 33436 20300 33544
rect 20625 33541 20637 33575
rect 20671 33541 20683 33575
rect 20625 33535 20683 33541
rect 20732 33504 20760 33600
rect 20806 33532 20812 33584
rect 20864 33581 20870 33584
rect 20864 33575 20885 33581
rect 20873 33572 20885 33575
rect 20916 33572 20944 33612
rect 21266 33600 21272 33612
rect 21324 33600 21330 33652
rect 20873 33544 20944 33572
rect 20993 33575 21051 33581
rect 20873 33541 20885 33544
rect 20864 33535 20885 33541
rect 20993 33541 21005 33575
rect 21039 33572 21051 33575
rect 21174 33572 21180 33584
rect 21039 33544 21180 33572
rect 21039 33541 21051 33544
rect 20993 33535 21051 33541
rect 20864 33532 20870 33535
rect 21174 33532 21180 33544
rect 21232 33572 21238 33584
rect 21913 33575 21971 33581
rect 21913 33572 21925 33575
rect 21232 33544 21925 33572
rect 21232 33532 21238 33544
rect 21913 33541 21925 33544
rect 21959 33541 21971 33575
rect 21913 33535 21971 33541
rect 21450 33504 21456 33516
rect 20732 33476 21456 33504
rect 21450 33464 21456 33476
rect 21508 33464 21514 33516
rect 21818 33504 21824 33516
rect 21779 33476 21824 33504
rect 21818 33464 21824 33476
rect 21876 33464 21882 33516
rect 22646 33504 22652 33516
rect 22607 33476 22652 33504
rect 22646 33464 22652 33476
rect 22704 33464 22710 33516
rect 29825 33507 29883 33513
rect 29825 33473 29837 33507
rect 29871 33504 29883 33507
rect 30098 33504 30104 33516
rect 29871 33476 30104 33504
rect 29871 33473 29883 33476
rect 29825 33467 29883 33473
rect 30098 33464 30104 33476
rect 30156 33464 30162 33516
rect 20272 33408 22094 33436
rect 19521 33399 19579 33405
rect 20441 33371 20499 33377
rect 20441 33368 20453 33371
rect 8941 33331 8999 33337
rect 9048 33340 10088 33368
rect 9048 33300 9076 33340
rect 8588 33272 9076 33300
rect 7561 33263 7619 33269
rect 9306 33260 9312 33312
rect 9364 33300 9370 33312
rect 9401 33303 9459 33309
rect 9401 33300 9413 33303
rect 9364 33272 9413 33300
rect 9364 33260 9370 33272
rect 9401 33269 9413 33272
rect 9447 33269 9459 33303
rect 10060 33300 10088 33340
rect 14200 33340 20453 33368
rect 14200 33300 14228 33340
rect 20441 33337 20453 33340
rect 20487 33337 20499 33371
rect 22066 33368 22094 33408
rect 29822 33368 29828 33380
rect 22066 33340 29828 33368
rect 20441 33331 20499 33337
rect 29822 33328 29828 33340
rect 29880 33328 29886 33380
rect 15654 33300 15660 33312
rect 10060 33272 14228 33300
rect 15615 33272 15660 33300
rect 9401 33263 9459 33269
rect 15654 33260 15660 33272
rect 15712 33260 15718 33312
rect 18690 33260 18696 33312
rect 18748 33300 18754 33312
rect 18785 33303 18843 33309
rect 18785 33300 18797 33303
rect 18748 33272 18797 33300
rect 18748 33260 18754 33272
rect 18785 33269 18797 33272
rect 18831 33269 18843 33303
rect 19794 33300 19800 33312
rect 19755 33272 19800 33300
rect 18785 33263 18843 33269
rect 19794 33260 19800 33272
rect 19852 33260 19858 33312
rect 22370 33260 22376 33312
rect 22428 33300 22434 33312
rect 22465 33303 22523 33309
rect 22465 33300 22477 33303
rect 22428 33272 22477 33300
rect 22428 33260 22434 33272
rect 22465 33269 22477 33272
rect 22511 33269 22523 33303
rect 30006 33300 30012 33312
rect 29967 33272 30012 33300
rect 22465 33263 22523 33269
rect 30006 33260 30012 33272
rect 30064 33260 30070 33312
rect 1104 33210 30820 33232
rect 1104 33158 5915 33210
rect 5967 33158 5979 33210
rect 6031 33158 6043 33210
rect 6095 33158 6107 33210
rect 6159 33158 6171 33210
rect 6223 33158 15846 33210
rect 15898 33158 15910 33210
rect 15962 33158 15974 33210
rect 16026 33158 16038 33210
rect 16090 33158 16102 33210
rect 16154 33158 25776 33210
rect 25828 33158 25840 33210
rect 25892 33158 25904 33210
rect 25956 33158 25968 33210
rect 26020 33158 26032 33210
rect 26084 33158 30820 33210
rect 1104 33136 30820 33158
rect 2222 33096 2228 33108
rect 2183 33068 2228 33096
rect 2222 33056 2228 33068
rect 2280 33056 2286 33108
rect 5718 33096 5724 33108
rect 5679 33068 5724 33096
rect 5718 33056 5724 33068
rect 5776 33056 5782 33108
rect 7926 33056 7932 33108
rect 7984 33096 7990 33108
rect 9214 33096 9220 33108
rect 7984 33068 9220 33096
rect 7984 33056 7990 33068
rect 9214 33056 9220 33068
rect 9272 33056 9278 33108
rect 9674 33056 9680 33108
rect 9732 33096 9738 33108
rect 10318 33096 10324 33108
rect 9732 33068 10324 33096
rect 9732 33056 9738 33068
rect 10318 33056 10324 33068
rect 10376 33096 10382 33108
rect 10689 33099 10747 33105
rect 10689 33096 10701 33099
rect 10376 33068 10701 33096
rect 10376 33056 10382 33068
rect 10689 33065 10701 33068
rect 10735 33065 10747 33099
rect 12066 33096 12072 33108
rect 12027 33068 12072 33096
rect 10689 33059 10747 33065
rect 12066 33056 12072 33068
rect 12124 33056 12130 33108
rect 19058 33096 19064 33108
rect 12406 33068 19064 33096
rect 1857 33031 1915 33037
rect 1857 32997 1869 33031
rect 1903 33028 1915 33031
rect 2130 33028 2136 33040
rect 1903 33000 2136 33028
rect 1903 32997 1915 33000
rect 1857 32991 1915 32997
rect 2130 32988 2136 33000
rect 2188 32988 2194 33040
rect 10410 32988 10416 33040
rect 10468 33028 10474 33040
rect 12406 33028 12434 33068
rect 19058 33056 19064 33068
rect 19116 33056 19122 33108
rect 19150 33056 19156 33108
rect 19208 33096 19214 33108
rect 19245 33099 19303 33105
rect 19245 33096 19257 33099
rect 19208 33068 19257 33096
rect 19208 33056 19214 33068
rect 19245 33065 19257 33068
rect 19291 33065 19303 33099
rect 19794 33096 19800 33108
rect 19707 33068 19800 33096
rect 19245 33059 19303 33065
rect 19794 33056 19800 33068
rect 19852 33096 19858 33108
rect 20438 33096 20444 33108
rect 19852 33068 20444 33096
rect 19852 33056 19858 33068
rect 20438 33056 20444 33068
rect 20496 33056 20502 33108
rect 20530 33056 20536 33108
rect 20588 33096 20594 33108
rect 21545 33099 21603 33105
rect 20588 33068 20944 33096
rect 20588 33056 20594 33068
rect 16390 33028 16396 33040
rect 10468 33000 12434 33028
rect 16351 33000 16396 33028
rect 10468 32988 10474 33000
rect 16390 32988 16396 33000
rect 16448 32988 16454 33040
rect 7926 32960 7932 32972
rect 7887 32932 7932 32960
rect 7926 32920 7932 32932
rect 7984 32920 7990 32972
rect 8021 32963 8079 32969
rect 8021 32929 8033 32963
rect 8067 32960 8079 32963
rect 8478 32960 8484 32972
rect 8067 32932 8484 32960
rect 8067 32929 8079 32932
rect 8021 32923 8079 32929
rect 8478 32920 8484 32932
rect 8536 32920 8542 32972
rect 9306 32960 9312 32972
rect 9267 32932 9312 32960
rect 9306 32920 9312 32932
rect 9364 32920 9370 32972
rect 10778 32920 10784 32972
rect 10836 32960 10842 32972
rect 11609 32963 11667 32969
rect 11609 32960 11621 32963
rect 10836 32932 11621 32960
rect 10836 32920 10842 32932
rect 11609 32929 11621 32932
rect 11655 32929 11667 32963
rect 12986 32960 12992 32972
rect 11609 32923 11667 32929
rect 11808 32932 12992 32960
rect 11808 32904 11836 32932
rect 12986 32920 12992 32932
rect 13044 32920 13050 32972
rect 15010 32960 15016 32972
rect 14971 32932 15016 32960
rect 15010 32920 15016 32932
rect 15068 32920 15074 32972
rect 16942 32960 16948 32972
rect 16903 32932 16948 32960
rect 16942 32920 16948 32932
rect 17000 32920 17006 32972
rect 19705 32963 19763 32969
rect 19705 32929 19717 32963
rect 19751 32960 19763 32963
rect 19886 32960 19892 32972
rect 19751 32932 19892 32960
rect 19751 32929 19763 32932
rect 19705 32923 19763 32929
rect 19886 32920 19892 32932
rect 19944 32960 19950 32972
rect 20916 32969 20944 33068
rect 21545 33065 21557 33099
rect 21591 33096 21603 33099
rect 21818 33096 21824 33108
rect 21591 33068 21824 33096
rect 21591 33065 21603 33068
rect 21545 33059 21603 33065
rect 21818 33056 21824 33068
rect 21876 33056 21882 33108
rect 22189 33099 22247 33105
rect 22189 33065 22201 33099
rect 22235 33065 22247 33099
rect 22189 33059 22247 33065
rect 22204 33028 22232 33059
rect 22066 33000 22232 33028
rect 20901 32963 20959 32969
rect 19944 32932 20852 32960
rect 19944 32920 19950 32932
rect 2869 32895 2927 32901
rect 2869 32861 2881 32895
rect 2915 32892 2927 32895
rect 3142 32892 3148 32904
rect 2915 32864 3148 32892
rect 2915 32861 2927 32864
rect 2869 32855 2927 32861
rect 3142 32852 3148 32864
rect 3200 32852 3206 32904
rect 3326 32852 3332 32904
rect 3384 32892 3390 32904
rect 3789 32895 3847 32901
rect 3789 32892 3801 32895
rect 3384 32864 3801 32892
rect 3384 32852 3390 32864
rect 3789 32861 3801 32864
rect 3835 32861 3847 32895
rect 3789 32855 3847 32861
rect 7009 32895 7067 32901
rect 7009 32861 7021 32895
rect 7055 32892 7067 32895
rect 7558 32892 7564 32904
rect 7055 32864 7564 32892
rect 7055 32861 7067 32864
rect 7009 32855 7067 32861
rect 7558 32852 7564 32864
rect 7616 32852 7622 32904
rect 7653 32895 7711 32901
rect 7653 32861 7665 32895
rect 7699 32861 7711 32895
rect 7653 32855 7711 32861
rect 7837 32895 7895 32901
rect 7837 32861 7849 32895
rect 7883 32892 7895 32895
rect 8110 32892 8116 32904
rect 7883 32864 8116 32892
rect 7883 32861 7895 32864
rect 7837 32855 7895 32861
rect 2225 32827 2283 32833
rect 2225 32793 2237 32827
rect 2271 32824 2283 32827
rect 2271 32796 3832 32824
rect 2271 32793 2283 32796
rect 2225 32787 2283 32793
rect 2406 32756 2412 32768
rect 2367 32728 2412 32756
rect 2406 32716 2412 32728
rect 2464 32716 2470 32768
rect 3053 32759 3111 32765
rect 3053 32725 3065 32759
rect 3099 32756 3111 32759
rect 3142 32756 3148 32768
rect 3099 32728 3148 32756
rect 3099 32725 3111 32728
rect 3053 32719 3111 32725
rect 3142 32716 3148 32728
rect 3200 32716 3206 32768
rect 3804 32756 3832 32796
rect 3878 32784 3884 32836
rect 3936 32824 3942 32836
rect 4034 32827 4092 32833
rect 4034 32824 4046 32827
rect 3936 32796 4046 32824
rect 3936 32784 3942 32796
rect 4034 32793 4046 32796
rect 4080 32793 4092 32827
rect 4034 32787 4092 32793
rect 5626 32784 5632 32836
rect 5684 32824 5690 32836
rect 5813 32827 5871 32833
rect 5813 32824 5825 32827
rect 5684 32796 5825 32824
rect 5684 32784 5690 32796
rect 5813 32793 5825 32796
rect 5859 32793 5871 32827
rect 7668 32824 7696 32855
rect 8110 32852 8116 32864
rect 8168 32852 8174 32904
rect 8205 32895 8263 32901
rect 8205 32861 8217 32895
rect 8251 32892 8263 32895
rect 9214 32892 9220 32904
rect 8251 32864 9220 32892
rect 8251 32861 8263 32864
rect 8205 32855 8263 32861
rect 9214 32852 9220 32864
rect 9272 32852 9278 32904
rect 9398 32852 9404 32904
rect 9456 32892 9462 32904
rect 9565 32895 9623 32901
rect 9565 32892 9577 32895
rect 9456 32864 9577 32892
rect 9456 32852 9462 32864
rect 9565 32861 9577 32864
rect 9611 32861 9623 32895
rect 9565 32855 9623 32861
rect 11517 32895 11575 32901
rect 11517 32861 11529 32895
rect 11563 32861 11575 32895
rect 11790 32892 11796 32904
rect 11703 32864 11796 32892
rect 11517 32855 11575 32861
rect 8662 32824 8668 32836
rect 7668 32796 8668 32824
rect 5813 32787 5871 32793
rect 8662 32784 8668 32796
rect 8720 32784 8726 32836
rect 11532 32824 11560 32855
rect 11790 32852 11796 32864
rect 11848 32852 11854 32904
rect 11882 32852 11888 32904
rect 11940 32892 11946 32904
rect 11940 32864 11985 32892
rect 11940 32852 11946 32864
rect 12066 32852 12072 32904
rect 12124 32892 12130 32904
rect 15280 32895 15338 32901
rect 12124 32864 12169 32892
rect 12124 32852 12130 32864
rect 15280 32861 15292 32895
rect 15326 32892 15338 32895
rect 15654 32892 15660 32904
rect 15326 32864 15660 32892
rect 15326 32861 15338 32864
rect 15280 32855 15338 32861
rect 15654 32852 15660 32864
rect 15712 32852 15718 32904
rect 19426 32852 19432 32904
rect 19484 32892 19490 32904
rect 19521 32895 19579 32901
rect 19521 32892 19533 32895
rect 19484 32864 19533 32892
rect 19484 32852 19490 32864
rect 19521 32861 19533 32864
rect 19567 32861 19579 32895
rect 19521 32855 19579 32861
rect 19610 32852 19616 32904
rect 19668 32892 19674 32904
rect 19981 32895 20039 32901
rect 19668 32864 19713 32892
rect 19668 32852 19674 32864
rect 19981 32861 19993 32895
rect 20027 32892 20039 32895
rect 20162 32892 20168 32904
rect 20027 32864 20168 32892
rect 20027 32861 20039 32864
rect 19981 32855 20039 32861
rect 20162 32852 20168 32864
rect 20220 32852 20226 32904
rect 20824 32892 20852 32932
rect 20901 32929 20913 32963
rect 20947 32929 20959 32963
rect 20901 32923 20959 32929
rect 22066 32892 22094 33000
rect 20824 32864 22094 32892
rect 12526 32824 12532 32836
rect 11532 32796 12532 32824
rect 12526 32784 12532 32796
rect 12584 32824 12590 32836
rect 12986 32824 12992 32836
rect 12584 32796 12992 32824
rect 12584 32784 12590 32796
rect 12986 32784 12992 32796
rect 13044 32784 13050 32836
rect 17212 32827 17270 32833
rect 17212 32793 17224 32827
rect 17258 32824 17270 32827
rect 17862 32824 17868 32836
rect 17258 32796 17868 32824
rect 17258 32793 17270 32796
rect 17212 32787 17270 32793
rect 17862 32784 17868 32796
rect 17920 32784 17926 32836
rect 20622 32784 20628 32836
rect 20680 32824 20686 32836
rect 21177 32827 21235 32833
rect 21177 32824 21189 32827
rect 20680 32796 21189 32824
rect 20680 32784 20686 32796
rect 21177 32793 21189 32796
rect 21223 32793 21235 32827
rect 21177 32787 21235 32793
rect 21910 32784 21916 32836
rect 21968 32824 21974 32836
rect 22373 32827 22431 32833
rect 22373 32824 22385 32827
rect 21968 32796 22385 32824
rect 21968 32784 21974 32796
rect 22373 32793 22385 32796
rect 22419 32793 22431 32827
rect 22373 32787 22431 32793
rect 5166 32756 5172 32768
rect 3804 32728 5172 32756
rect 5166 32716 5172 32728
rect 5224 32716 5230 32768
rect 6822 32756 6828 32768
rect 6783 32728 6828 32756
rect 6822 32716 6828 32728
rect 6880 32716 6886 32768
rect 8389 32759 8447 32765
rect 8389 32725 8401 32759
rect 8435 32756 8447 32759
rect 8754 32756 8760 32768
rect 8435 32728 8760 32756
rect 8435 32725 8447 32728
rect 8389 32719 8447 32725
rect 8754 32716 8760 32728
rect 8812 32716 8818 32768
rect 18322 32756 18328 32768
rect 18283 32728 18328 32756
rect 18322 32716 18328 32728
rect 18380 32716 18386 32768
rect 18414 32716 18420 32768
rect 18472 32756 18478 32768
rect 20530 32756 20536 32768
rect 18472 32728 20536 32756
rect 18472 32716 18478 32728
rect 20530 32716 20536 32728
rect 20588 32716 20594 32768
rect 20714 32716 20720 32768
rect 20772 32756 20778 32768
rect 21085 32759 21143 32765
rect 21085 32756 21097 32759
rect 20772 32728 21097 32756
rect 20772 32716 20778 32728
rect 21085 32725 21097 32728
rect 21131 32725 21143 32759
rect 21085 32719 21143 32725
rect 21358 32716 21364 32768
rect 21416 32756 21422 32768
rect 22186 32765 22192 32768
rect 22005 32759 22063 32765
rect 22005 32756 22017 32759
rect 21416 32728 22017 32756
rect 21416 32716 21422 32728
rect 22005 32725 22017 32728
rect 22051 32725 22063 32759
rect 22005 32719 22063 32725
rect 22173 32759 22192 32765
rect 22173 32725 22185 32759
rect 22173 32719 22192 32725
rect 22186 32716 22192 32719
rect 22244 32716 22250 32768
rect 1104 32666 30820 32688
rect 1104 32614 10880 32666
rect 10932 32614 10944 32666
rect 10996 32614 11008 32666
rect 11060 32614 11072 32666
rect 11124 32614 11136 32666
rect 11188 32614 20811 32666
rect 20863 32614 20875 32666
rect 20927 32614 20939 32666
rect 20991 32614 21003 32666
rect 21055 32614 21067 32666
rect 21119 32614 30820 32666
rect 1104 32592 30820 32614
rect 3326 32552 3332 32564
rect 3287 32524 3332 32552
rect 3326 32512 3332 32524
rect 3384 32512 3390 32564
rect 3789 32555 3847 32561
rect 3789 32521 3801 32555
rect 3835 32552 3847 32555
rect 3878 32552 3884 32564
rect 3835 32524 3884 32552
rect 3835 32521 3847 32524
rect 3789 32515 3847 32521
rect 3878 32512 3884 32524
rect 3936 32512 3942 32564
rect 7742 32512 7748 32564
rect 7800 32552 7806 32564
rect 8110 32552 8116 32564
rect 7800 32524 8116 32552
rect 7800 32512 7806 32524
rect 8110 32512 8116 32524
rect 8168 32552 8174 32564
rect 8205 32555 8263 32561
rect 8205 32552 8217 32555
rect 8168 32524 8217 32552
rect 8168 32512 8174 32524
rect 8205 32521 8217 32524
rect 8251 32521 8263 32555
rect 8205 32515 8263 32521
rect 9214 32512 9220 32564
rect 9272 32552 9278 32564
rect 10045 32555 10103 32561
rect 10045 32552 10057 32555
rect 9272 32524 10057 32552
rect 9272 32512 9278 32524
rect 10045 32521 10057 32524
rect 10091 32521 10103 32555
rect 15470 32552 15476 32564
rect 10045 32515 10103 32521
rect 10612 32524 13952 32552
rect 15431 32524 15476 32552
rect 5166 32484 5172 32496
rect 3988 32456 5172 32484
rect 1673 32419 1731 32425
rect 1673 32385 1685 32419
rect 1719 32385 1731 32419
rect 1673 32379 1731 32385
rect 2409 32419 2467 32425
rect 2409 32385 2421 32419
rect 2455 32416 2467 32419
rect 2774 32416 2780 32428
rect 2455 32388 2780 32416
rect 2455 32385 2467 32388
rect 2409 32379 2467 32385
rect 1688 32348 1716 32379
rect 2774 32376 2780 32388
rect 2832 32376 2838 32428
rect 3142 32416 3148 32428
rect 3103 32388 3148 32416
rect 3142 32376 3148 32388
rect 3200 32376 3206 32428
rect 3988 32425 4016 32456
rect 5166 32444 5172 32456
rect 5224 32444 5230 32496
rect 7098 32493 7104 32496
rect 7092 32484 7104 32493
rect 7059 32456 7104 32484
rect 7092 32447 7104 32456
rect 7098 32444 7104 32447
rect 7156 32444 7162 32496
rect 9950 32484 9956 32496
rect 7208 32456 9956 32484
rect 3973 32419 4031 32425
rect 3973 32385 3985 32419
rect 4019 32385 4031 32419
rect 4246 32416 4252 32428
rect 4207 32388 4252 32416
rect 3973 32379 4031 32385
rect 4246 32376 4252 32388
rect 4304 32376 4310 32428
rect 4341 32419 4399 32425
rect 4341 32385 4353 32419
rect 4387 32385 4399 32419
rect 4341 32379 4399 32385
rect 2958 32348 2964 32360
rect 1688 32320 2964 32348
rect 2958 32308 2964 32320
rect 3016 32308 3022 32360
rect 4062 32308 4068 32360
rect 4120 32348 4126 32360
rect 4157 32351 4215 32357
rect 4157 32348 4169 32351
rect 4120 32320 4169 32348
rect 4120 32308 4126 32320
rect 4157 32317 4169 32320
rect 4203 32317 4215 32351
rect 4157 32311 4215 32317
rect 4356 32280 4384 32379
rect 4430 32376 4436 32428
rect 4488 32416 4494 32428
rect 4525 32419 4583 32425
rect 4525 32416 4537 32419
rect 4488 32388 4537 32416
rect 4488 32376 4494 32388
rect 4525 32385 4537 32388
rect 4571 32385 4583 32419
rect 4525 32379 4583 32385
rect 5353 32419 5411 32425
rect 5353 32385 5365 32419
rect 5399 32416 5411 32419
rect 5626 32416 5632 32428
rect 5399 32388 5632 32416
rect 5399 32385 5411 32388
rect 5353 32379 5411 32385
rect 5626 32376 5632 32388
rect 5684 32416 5690 32428
rect 7208 32416 7236 32456
rect 9950 32444 9956 32456
rect 10008 32444 10014 32496
rect 5684 32388 7236 32416
rect 5684 32376 5690 32388
rect 8754 32376 8760 32428
rect 8812 32416 8818 32428
rect 8921 32419 8979 32425
rect 8921 32416 8933 32419
rect 8812 32388 8933 32416
rect 8812 32376 8818 32388
rect 8921 32385 8933 32388
rect 8967 32385 8979 32419
rect 8921 32379 8979 32385
rect 5537 32351 5595 32357
rect 5537 32317 5549 32351
rect 5583 32317 5595 32351
rect 5537 32311 5595 32317
rect 4522 32280 4528 32292
rect 4356 32252 4528 32280
rect 4522 32240 4528 32252
rect 4580 32240 4586 32292
rect 5552 32280 5580 32311
rect 6362 32308 6368 32360
rect 6420 32348 6426 32360
rect 6825 32351 6883 32357
rect 6825 32348 6837 32351
rect 6420 32320 6837 32348
rect 6420 32308 6426 32320
rect 6825 32317 6837 32320
rect 6871 32317 6883 32351
rect 8662 32348 8668 32360
rect 8623 32320 8668 32348
rect 6825 32311 6883 32317
rect 8662 32308 8668 32320
rect 8720 32308 8726 32360
rect 6638 32280 6644 32292
rect 5552 32252 6644 32280
rect 6638 32240 6644 32252
rect 6696 32240 6702 32292
rect 10410 32280 10416 32292
rect 9646 32252 10416 32280
rect 1486 32212 1492 32224
rect 1447 32184 1492 32212
rect 1486 32172 1492 32184
rect 1544 32172 1550 32224
rect 2222 32212 2228 32224
rect 2183 32184 2228 32212
rect 2222 32172 2228 32184
rect 2280 32172 2286 32224
rect 6730 32172 6736 32224
rect 6788 32212 6794 32224
rect 9646 32212 9674 32252
rect 10410 32240 10416 32252
rect 10468 32240 10474 32292
rect 6788 32184 9674 32212
rect 6788 32172 6794 32184
rect 9766 32172 9772 32224
rect 9824 32212 9830 32224
rect 10612 32221 10640 32524
rect 13924 32496 13952 32524
rect 15470 32512 15476 32524
rect 15528 32512 15534 32564
rect 17862 32552 17868 32564
rect 17823 32524 17868 32552
rect 17862 32512 17868 32524
rect 17920 32512 17926 32564
rect 19242 32552 19248 32564
rect 19203 32524 19248 32552
rect 19242 32512 19248 32524
rect 19300 32512 19306 32564
rect 19702 32512 19708 32564
rect 19760 32552 19766 32564
rect 19760 32524 20116 32552
rect 19760 32512 19766 32524
rect 11514 32484 11520 32496
rect 10888 32456 11520 32484
rect 10888 32428 10916 32456
rect 11514 32444 11520 32456
rect 11572 32484 11578 32496
rect 12066 32484 12072 32496
rect 11572 32456 12072 32484
rect 11572 32444 11578 32456
rect 12066 32444 12072 32456
rect 12124 32444 12130 32496
rect 12526 32444 12532 32496
rect 12584 32484 12590 32496
rect 13694 32487 13752 32493
rect 13694 32484 13706 32487
rect 12584 32456 13706 32484
rect 12584 32444 12590 32456
rect 13694 32453 13706 32456
rect 13740 32453 13752 32487
rect 13694 32447 13752 32453
rect 13906 32444 13912 32496
rect 13964 32484 13970 32496
rect 13964 32456 18552 32484
rect 13964 32444 13970 32456
rect 10870 32416 10876 32428
rect 10831 32388 10876 32416
rect 10870 32376 10876 32388
rect 10928 32376 10934 32428
rect 11784 32419 11842 32425
rect 11784 32385 11796 32419
rect 11830 32416 11842 32419
rect 12250 32416 12256 32428
rect 11830 32388 12256 32416
rect 11830 32385 11842 32388
rect 11784 32379 11842 32385
rect 12250 32376 12256 32388
rect 12308 32376 12314 32428
rect 12894 32376 12900 32428
rect 12952 32416 12958 32428
rect 13449 32419 13507 32425
rect 13449 32416 13461 32419
rect 12952 32388 13461 32416
rect 12952 32376 12958 32388
rect 13449 32385 13461 32388
rect 13495 32385 13507 32419
rect 13449 32379 13507 32385
rect 15286 32376 15292 32428
rect 15344 32416 15350 32428
rect 15381 32419 15439 32425
rect 15381 32416 15393 32419
rect 15344 32388 15393 32416
rect 15344 32376 15350 32388
rect 15381 32385 15393 32388
rect 15427 32385 15439 32419
rect 17126 32416 17132 32428
rect 17087 32388 17132 32416
rect 15381 32379 15439 32385
rect 17126 32376 17132 32388
rect 17184 32376 17190 32428
rect 17310 32416 17316 32428
rect 17271 32388 17316 32416
rect 17310 32376 17316 32388
rect 17368 32376 17374 32428
rect 17681 32419 17739 32425
rect 17681 32385 17693 32419
rect 17727 32416 17739 32419
rect 18322 32416 18328 32428
rect 17727 32388 18328 32416
rect 17727 32385 17739 32388
rect 17681 32379 17739 32385
rect 18322 32376 18328 32388
rect 18380 32376 18386 32428
rect 18524 32425 18552 32456
rect 18598 32444 18604 32496
rect 18656 32484 18662 32496
rect 18656 32456 19104 32484
rect 18656 32444 18662 32456
rect 18509 32419 18567 32425
rect 18509 32385 18521 32419
rect 18555 32385 18567 32419
rect 18693 32419 18751 32425
rect 18693 32416 18705 32419
rect 18509 32379 18567 32385
rect 18616 32388 18705 32416
rect 11330 32308 11336 32360
rect 11388 32348 11394 32360
rect 11517 32351 11575 32357
rect 11517 32348 11529 32351
rect 11388 32320 11529 32348
rect 11388 32308 11394 32320
rect 11517 32317 11529 32320
rect 11563 32317 11575 32351
rect 11517 32311 11575 32317
rect 17144 32280 17172 32376
rect 17402 32348 17408 32360
rect 17363 32320 17408 32348
rect 17402 32308 17408 32320
rect 17460 32308 17466 32360
rect 17497 32351 17555 32357
rect 17497 32317 17509 32351
rect 17543 32348 17555 32351
rect 18414 32348 18420 32360
rect 17543 32320 18420 32348
rect 17543 32317 17555 32320
rect 17497 32311 17555 32317
rect 18414 32308 18420 32320
rect 18472 32308 18478 32360
rect 17770 32280 17776 32292
rect 17144 32252 17776 32280
rect 17770 32240 17776 32252
rect 17828 32240 17834 32292
rect 10597 32215 10655 32221
rect 10597 32212 10609 32215
rect 9824 32184 10609 32212
rect 9824 32172 9830 32184
rect 10597 32181 10609 32184
rect 10643 32181 10655 32215
rect 10597 32175 10655 32181
rect 12158 32172 12164 32224
rect 12216 32212 12222 32224
rect 12897 32215 12955 32221
rect 12897 32212 12909 32215
rect 12216 32184 12909 32212
rect 12216 32172 12222 32184
rect 12897 32181 12909 32184
rect 12943 32212 12955 32215
rect 14642 32212 14648 32224
rect 12943 32184 14648 32212
rect 12943 32181 12955 32184
rect 12897 32175 12955 32181
rect 14642 32172 14648 32184
rect 14700 32172 14706 32224
rect 14734 32172 14740 32224
rect 14792 32212 14798 32224
rect 14829 32215 14887 32221
rect 14829 32212 14841 32215
rect 14792 32184 14841 32212
rect 14792 32172 14798 32184
rect 14829 32181 14841 32184
rect 14875 32181 14887 32215
rect 18616 32212 18644 32388
rect 18693 32385 18705 32388
rect 18739 32385 18751 32419
rect 18874 32416 18880 32428
rect 18835 32388 18880 32416
rect 18693 32379 18751 32385
rect 18874 32376 18880 32388
rect 18932 32376 18938 32428
rect 19076 32425 19104 32456
rect 19794 32444 19800 32496
rect 19852 32484 19858 32496
rect 19981 32487 20039 32493
rect 19981 32484 19993 32487
rect 19852 32456 19993 32484
rect 19852 32444 19858 32456
rect 19981 32453 19993 32456
rect 20027 32453 20039 32487
rect 20088 32484 20116 32524
rect 20254 32512 20260 32564
rect 20312 32552 20318 32564
rect 20312 32524 21496 32552
rect 20312 32512 20318 32524
rect 20622 32484 20628 32496
rect 20088 32456 20628 32484
rect 19981 32447 20039 32453
rect 20622 32444 20628 32456
rect 20680 32444 20686 32496
rect 21358 32484 21364 32496
rect 20916 32456 21364 32484
rect 19061 32419 19119 32425
rect 19061 32385 19073 32419
rect 19107 32385 19119 32419
rect 19061 32379 19119 32385
rect 19610 32376 19616 32428
rect 19668 32416 19674 32428
rect 20438 32416 20444 32428
rect 19668 32388 20444 32416
rect 19668 32376 19674 32388
rect 20438 32376 20444 32388
rect 20496 32416 20502 32428
rect 20916 32425 20944 32456
rect 21358 32444 21364 32456
rect 21416 32444 21422 32496
rect 21468 32484 21496 32524
rect 21634 32512 21640 32564
rect 21692 32552 21698 32564
rect 21979 32555 22037 32561
rect 21979 32552 21991 32555
rect 21692 32524 21991 32552
rect 21692 32512 21698 32524
rect 21979 32521 21991 32524
rect 22025 32521 22037 32555
rect 21979 32515 22037 32521
rect 22186 32484 22192 32496
rect 21468 32456 22192 32484
rect 22186 32444 22192 32456
rect 22244 32444 22250 32496
rect 20533 32419 20591 32425
rect 20533 32416 20545 32419
rect 20496 32388 20545 32416
rect 20496 32376 20502 32388
rect 20533 32385 20545 32388
rect 20579 32385 20591 32419
rect 20533 32379 20591 32385
rect 20901 32419 20959 32425
rect 20901 32385 20913 32419
rect 20947 32385 20959 32419
rect 21266 32416 21272 32428
rect 21227 32388 21272 32416
rect 20901 32379 20959 32385
rect 21266 32376 21272 32388
rect 21324 32376 21330 32428
rect 18785 32351 18843 32357
rect 18785 32317 18797 32351
rect 18831 32348 18843 32351
rect 19150 32348 19156 32360
rect 18831 32320 19156 32348
rect 18831 32317 18843 32320
rect 18785 32311 18843 32317
rect 19150 32308 19156 32320
rect 19208 32308 19214 32360
rect 20625 32351 20683 32357
rect 20625 32348 20637 32351
rect 20088 32320 20637 32348
rect 18690 32240 18696 32292
rect 18748 32280 18754 32292
rect 20088 32280 20116 32320
rect 20625 32317 20637 32320
rect 20671 32348 20683 32351
rect 20714 32348 20720 32360
rect 20671 32320 20720 32348
rect 20671 32317 20683 32320
rect 20625 32311 20683 32317
rect 20714 32308 20720 32320
rect 20772 32308 20778 32360
rect 21085 32351 21143 32357
rect 21085 32317 21097 32351
rect 21131 32348 21143 32351
rect 21174 32348 21180 32360
rect 21131 32320 21180 32348
rect 21131 32317 21143 32320
rect 21085 32311 21143 32317
rect 21174 32308 21180 32320
rect 21232 32308 21238 32360
rect 18748 32252 20116 32280
rect 18748 32240 18754 32252
rect 20530 32240 20536 32292
rect 20588 32280 20594 32292
rect 20588 32252 21956 32280
rect 20588 32240 20594 32252
rect 21928 32224 21956 32252
rect 19886 32212 19892 32224
rect 18616 32184 19892 32212
rect 14829 32175 14887 32181
rect 19886 32172 19892 32184
rect 19944 32172 19950 32224
rect 20898 32172 20904 32224
rect 20956 32212 20962 32224
rect 21821 32215 21879 32221
rect 21821 32212 21833 32215
rect 20956 32184 21833 32212
rect 20956 32172 20962 32184
rect 21821 32181 21833 32184
rect 21867 32181 21879 32215
rect 21821 32175 21879 32181
rect 21910 32172 21916 32224
rect 21968 32212 21974 32224
rect 22005 32215 22063 32221
rect 22005 32212 22017 32215
rect 21968 32184 22017 32212
rect 21968 32172 21974 32184
rect 22005 32181 22017 32184
rect 22051 32181 22063 32215
rect 22005 32175 22063 32181
rect 1104 32122 30820 32144
rect 1104 32070 5915 32122
rect 5967 32070 5979 32122
rect 6031 32070 6043 32122
rect 6095 32070 6107 32122
rect 6159 32070 6171 32122
rect 6223 32070 15846 32122
rect 15898 32070 15910 32122
rect 15962 32070 15974 32122
rect 16026 32070 16038 32122
rect 16090 32070 16102 32122
rect 16154 32070 25776 32122
rect 25828 32070 25840 32122
rect 25892 32070 25904 32122
rect 25956 32070 25968 32122
rect 26020 32070 26032 32122
rect 26084 32070 30820 32122
rect 1104 32048 30820 32070
rect 2314 32008 2320 32020
rect 2275 31980 2320 32008
rect 2314 31968 2320 31980
rect 2372 31968 2378 32020
rect 2958 32008 2964 32020
rect 2919 31980 2964 32008
rect 2958 31968 2964 31980
rect 3016 31968 3022 32020
rect 6362 32008 6368 32020
rect 6323 31980 6368 32008
rect 6362 31968 6368 31980
rect 6420 31968 6426 32020
rect 7009 32011 7067 32017
rect 7009 31977 7021 32011
rect 7055 32008 7067 32011
rect 8662 32008 8668 32020
rect 7055 31980 8668 32008
rect 7055 31977 7067 31980
rect 7009 31971 7067 31977
rect 8662 31968 8668 31980
rect 8720 31968 8726 32020
rect 9674 32008 9680 32020
rect 9635 31980 9680 32008
rect 9674 31968 9680 31980
rect 9732 31968 9738 32020
rect 10134 31968 10140 32020
rect 10192 32008 10198 32020
rect 10870 32008 10876 32020
rect 10192 31980 10876 32008
rect 10192 31968 10198 31980
rect 10870 31968 10876 31980
rect 10928 31968 10934 32020
rect 18506 32008 18512 32020
rect 18467 31980 18512 32008
rect 18506 31968 18512 31980
rect 18564 31968 18570 32020
rect 19058 31968 19064 32020
rect 19116 32008 19122 32020
rect 20533 32011 20591 32017
rect 20533 32008 20545 32011
rect 19116 31980 20545 32008
rect 19116 31968 19122 31980
rect 20533 31977 20545 31980
rect 20579 31977 20591 32011
rect 20533 31971 20591 31977
rect 1949 31943 2007 31949
rect 1949 31909 1961 31943
rect 1995 31940 2007 31943
rect 2130 31940 2136 31952
rect 1995 31912 2136 31940
rect 1995 31909 2007 31912
rect 1949 31903 2007 31909
rect 2130 31900 2136 31912
rect 2188 31900 2194 31952
rect 2501 31943 2559 31949
rect 2501 31909 2513 31943
rect 2547 31909 2559 31943
rect 2501 31903 2559 31909
rect 2516 31872 2544 31903
rect 3786 31900 3792 31952
rect 3844 31940 3850 31952
rect 4062 31940 4068 31952
rect 3844 31912 4068 31940
rect 3844 31900 3850 31912
rect 4062 31900 4068 31912
rect 4120 31900 4126 31952
rect 7469 31943 7527 31949
rect 7469 31909 7481 31943
rect 7515 31909 7527 31943
rect 7469 31903 7527 31909
rect 8113 31943 8171 31949
rect 8113 31909 8125 31943
rect 8159 31909 8171 31943
rect 8113 31903 8171 31909
rect 2958 31872 2964 31884
rect 2516 31844 2964 31872
rect 2958 31832 2964 31844
rect 3016 31832 3022 31884
rect 5626 31872 5632 31884
rect 5587 31844 5632 31872
rect 5626 31832 5632 31844
rect 5684 31832 5690 31884
rect 7484 31872 7512 31903
rect 8128 31872 8156 31903
rect 9858 31900 9864 31952
rect 9916 31940 9922 31952
rect 10597 31943 10655 31949
rect 10597 31940 10609 31943
rect 9916 31912 10609 31940
rect 9916 31900 9922 31912
rect 10597 31909 10609 31912
rect 10643 31940 10655 31943
rect 11146 31940 11152 31952
rect 10643 31912 11152 31940
rect 10643 31909 10655 31912
rect 10597 31903 10655 31909
rect 11146 31900 11152 31912
rect 11204 31900 11210 31952
rect 11238 31900 11244 31952
rect 11296 31900 11302 31952
rect 12618 31940 12624 31952
rect 12579 31912 12624 31940
rect 12618 31900 12624 31912
rect 12676 31900 12682 31952
rect 12894 31900 12900 31952
rect 12952 31940 12958 31952
rect 13081 31943 13139 31949
rect 13081 31940 13093 31943
rect 12952 31912 13093 31940
rect 12952 31900 12958 31912
rect 13081 31909 13093 31912
rect 13127 31909 13139 31943
rect 13081 31903 13139 31909
rect 17402 31900 17408 31952
rect 17460 31940 17466 31952
rect 19613 31943 19671 31949
rect 19613 31940 19625 31943
rect 17460 31912 19625 31940
rect 17460 31900 17466 31912
rect 19613 31909 19625 31912
rect 19659 31909 19671 31943
rect 19613 31903 19671 31909
rect 6196 31844 7512 31872
rect 7760 31844 8156 31872
rect 3142 31804 3148 31816
rect 3103 31776 3148 31804
rect 3142 31764 3148 31776
rect 3200 31764 3206 31816
rect 4522 31764 4528 31816
rect 4580 31804 4586 31816
rect 5166 31804 5172 31816
rect 4580 31776 5172 31804
rect 4580 31764 4586 31776
rect 5166 31764 5172 31776
rect 5224 31804 5230 31816
rect 6196 31813 6224 31844
rect 5353 31807 5411 31813
rect 5353 31804 5365 31807
rect 5224 31776 5365 31804
rect 5224 31764 5230 31776
rect 5353 31773 5365 31776
rect 5399 31773 5411 31807
rect 5353 31767 5411 31773
rect 6181 31807 6239 31813
rect 6181 31773 6193 31807
rect 6227 31773 6239 31807
rect 6181 31767 6239 31773
rect 6454 31764 6460 31816
rect 6512 31804 6518 31816
rect 6822 31804 6828 31816
rect 6512 31776 6684 31804
rect 6783 31776 6828 31804
rect 6512 31764 6518 31776
rect 4249 31739 4307 31745
rect 4249 31705 4261 31739
rect 4295 31736 4307 31739
rect 4798 31736 4804 31748
rect 4295 31708 4804 31736
rect 4295 31705 4307 31708
rect 4249 31699 4307 31705
rect 4798 31696 4804 31708
rect 4856 31696 4862 31748
rect 6656 31736 6684 31776
rect 6822 31764 6828 31776
rect 6880 31764 6886 31816
rect 6932 31776 7512 31804
rect 6932 31736 6960 31776
rect 6656 31708 6960 31736
rect 7484 31736 7512 31776
rect 7558 31764 7564 31816
rect 7616 31804 7622 31816
rect 7653 31807 7711 31813
rect 7653 31804 7665 31807
rect 7616 31776 7665 31804
rect 7616 31764 7622 31776
rect 7653 31773 7665 31776
rect 7699 31773 7711 31807
rect 7653 31767 7711 31773
rect 7760 31736 7788 31844
rect 9122 31832 9128 31884
rect 9180 31872 9186 31884
rect 9493 31875 9551 31881
rect 9493 31872 9505 31875
rect 9180 31844 9505 31872
rect 9180 31832 9186 31844
rect 9493 31841 9505 31844
rect 9539 31841 9551 31875
rect 11256 31872 11284 31900
rect 9493 31835 9551 31841
rect 9968 31844 11284 31872
rect 8297 31807 8355 31813
rect 8297 31773 8309 31807
rect 8343 31804 8355 31807
rect 8846 31804 8852 31816
rect 8343 31776 8852 31804
rect 8343 31773 8355 31776
rect 8297 31767 8355 31773
rect 8846 31764 8852 31776
rect 8904 31764 8910 31816
rect 9968 31813 9996 31844
rect 9953 31807 10011 31813
rect 9953 31773 9965 31807
rect 9999 31773 10011 31807
rect 9953 31767 10011 31773
rect 10042 31764 10048 31816
rect 10100 31804 10106 31816
rect 10413 31807 10471 31813
rect 10413 31804 10425 31807
rect 10100 31776 10425 31804
rect 10100 31764 10106 31776
rect 10413 31773 10425 31776
rect 10459 31773 10471 31807
rect 10413 31767 10471 31773
rect 11241 31807 11299 31813
rect 11241 31773 11253 31807
rect 11287 31804 11299 31807
rect 11330 31804 11336 31816
rect 11287 31776 11336 31804
rect 11287 31773 11299 31776
rect 11241 31767 11299 31773
rect 11330 31764 11336 31776
rect 11388 31804 11394 31816
rect 12912 31804 12940 31900
rect 18414 31872 18420 31884
rect 13280 31844 14228 31872
rect 18375 31844 18420 31872
rect 13280 31813 13308 31844
rect 13265 31807 13323 31813
rect 11388 31776 13216 31804
rect 11388 31764 11394 31776
rect 7484 31708 7788 31736
rect 11508 31739 11566 31745
rect 11508 31705 11520 31739
rect 11554 31736 11566 31739
rect 11882 31736 11888 31748
rect 11554 31708 11888 31736
rect 11554 31705 11566 31708
rect 11508 31699 11566 31705
rect 11882 31696 11888 31708
rect 11940 31696 11946 31748
rect 13188 31736 13216 31776
rect 13265 31773 13277 31807
rect 13311 31773 13323 31807
rect 14093 31807 14151 31813
rect 14093 31804 14105 31807
rect 13265 31767 13323 31773
rect 13372 31776 14105 31804
rect 13372 31736 13400 31776
rect 14093 31773 14105 31776
rect 14139 31773 14151 31807
rect 14200 31804 14228 31844
rect 18414 31832 18420 31844
rect 18472 31832 18478 31884
rect 18601 31875 18659 31881
rect 18601 31841 18613 31875
rect 18647 31872 18659 31875
rect 19978 31872 19984 31884
rect 18647 31844 19984 31872
rect 18647 31841 18659 31844
rect 18601 31835 18659 31841
rect 19978 31832 19984 31844
rect 20036 31872 20042 31884
rect 20714 31872 20720 31884
rect 20036 31844 20720 31872
rect 20036 31832 20042 31844
rect 20714 31832 20720 31844
rect 20772 31832 20778 31884
rect 20898 31872 20904 31884
rect 20859 31844 20904 31872
rect 20898 31832 20904 31844
rect 20956 31832 20962 31884
rect 21266 31832 21272 31884
rect 21324 31832 21330 31884
rect 15470 31804 15476 31816
rect 14200 31776 15476 31804
rect 14093 31767 14151 31773
rect 15470 31764 15476 31776
rect 15528 31764 15534 31816
rect 18690 31804 18696 31816
rect 18651 31776 18696 31804
rect 18690 31764 18696 31776
rect 18748 31764 18754 31816
rect 20622 31804 20628 31816
rect 20583 31776 20628 31804
rect 20622 31764 20628 31776
rect 20680 31764 20686 31816
rect 20732 31804 20760 31832
rect 20809 31807 20867 31813
rect 20809 31804 20821 31807
rect 20732 31776 20821 31804
rect 20809 31773 20821 31776
rect 20855 31773 20867 31807
rect 20994 31807 21052 31813
rect 20994 31804 21006 31807
rect 20809 31767 20867 31773
rect 20916 31776 21006 31804
rect 13188 31708 13400 31736
rect 13814 31696 13820 31748
rect 13872 31736 13878 31748
rect 14338 31739 14396 31745
rect 14338 31736 14350 31739
rect 13872 31708 14350 31736
rect 13872 31696 13878 31708
rect 14338 31705 14350 31708
rect 14384 31705 14396 31739
rect 14338 31699 14396 31705
rect 19797 31739 19855 31745
rect 19797 31705 19809 31739
rect 19843 31736 19855 31739
rect 20438 31736 20444 31748
rect 19843 31708 20444 31736
rect 19843 31705 19855 31708
rect 19797 31699 19855 31705
rect 20438 31696 20444 31708
rect 20496 31696 20502 31748
rect 20916 31736 20944 31776
rect 20994 31773 21006 31776
rect 21040 31773 21052 31807
rect 20994 31767 21052 31773
rect 21177 31807 21235 31813
rect 21177 31773 21189 31807
rect 21223 31804 21235 31807
rect 21284 31804 21312 31832
rect 21910 31804 21916 31816
rect 21223 31776 21916 31804
rect 21223 31773 21235 31776
rect 21177 31767 21235 31773
rect 21910 31764 21916 31776
rect 21968 31764 21974 31816
rect 29822 31804 29828 31816
rect 29783 31776 29828 31804
rect 29822 31764 29828 31776
rect 29880 31764 29886 31816
rect 21082 31736 21088 31748
rect 20916 31708 21088 31736
rect 21082 31696 21088 31708
rect 21140 31696 21146 31748
rect 2317 31671 2375 31677
rect 2317 31637 2329 31671
rect 2363 31668 2375 31671
rect 4154 31668 4160 31680
rect 2363 31640 4160 31668
rect 2363 31637 2375 31640
rect 2317 31631 2375 31637
rect 4154 31628 4160 31640
rect 4212 31628 4218 31680
rect 7098 31628 7104 31680
rect 7156 31668 7162 31680
rect 9766 31668 9772 31680
rect 7156 31640 9772 31668
rect 7156 31628 7162 31640
rect 9766 31628 9772 31640
rect 9824 31628 9830 31680
rect 15378 31628 15384 31680
rect 15436 31668 15442 31680
rect 15473 31671 15531 31677
rect 15473 31668 15485 31671
rect 15436 31640 15485 31668
rect 15436 31628 15442 31640
rect 15473 31637 15485 31640
rect 15519 31637 15531 31671
rect 30006 31668 30012 31680
rect 29967 31640 30012 31668
rect 15473 31631 15531 31637
rect 30006 31628 30012 31640
rect 30064 31628 30070 31680
rect 1104 31578 30820 31600
rect 1104 31526 10880 31578
rect 10932 31526 10944 31578
rect 10996 31526 11008 31578
rect 11060 31526 11072 31578
rect 11124 31526 11136 31578
rect 11188 31526 20811 31578
rect 20863 31526 20875 31578
rect 20927 31526 20939 31578
rect 20991 31526 21003 31578
rect 21055 31526 21067 31578
rect 21119 31526 30820 31578
rect 1104 31504 30820 31526
rect 2501 31467 2559 31473
rect 2501 31433 2513 31467
rect 2547 31464 2559 31467
rect 3142 31464 3148 31476
rect 2547 31436 3148 31464
rect 2547 31433 2559 31436
rect 2501 31427 2559 31433
rect 3142 31424 3148 31436
rect 3200 31424 3206 31476
rect 8297 31467 8355 31473
rect 8297 31433 8309 31467
rect 8343 31464 8355 31467
rect 8386 31464 8392 31476
rect 8343 31436 8392 31464
rect 8343 31433 8355 31436
rect 8297 31427 8355 31433
rect 8386 31424 8392 31436
rect 8444 31424 8450 31476
rect 11793 31467 11851 31473
rect 11793 31433 11805 31467
rect 11839 31464 11851 31467
rect 12526 31464 12532 31476
rect 11839 31436 12532 31464
rect 11839 31433 11851 31436
rect 11793 31427 11851 31433
rect 12526 31424 12532 31436
rect 12584 31424 12590 31476
rect 12894 31424 12900 31476
rect 12952 31464 12958 31476
rect 13446 31464 13452 31476
rect 12952 31436 13452 31464
rect 12952 31424 12958 31436
rect 13446 31424 13452 31436
rect 13504 31424 13510 31476
rect 13541 31467 13599 31473
rect 13541 31433 13553 31467
rect 13587 31464 13599 31467
rect 13814 31464 13820 31476
rect 13587 31436 13820 31464
rect 13587 31433 13599 31436
rect 13541 31427 13599 31433
rect 13814 31424 13820 31436
rect 13872 31424 13878 31476
rect 15286 31424 15292 31476
rect 15344 31464 15350 31476
rect 15381 31467 15439 31473
rect 15381 31464 15393 31467
rect 15344 31436 15393 31464
rect 15344 31424 15350 31436
rect 15381 31433 15393 31436
rect 15427 31433 15439 31467
rect 15381 31427 15439 31433
rect 17034 31424 17040 31476
rect 17092 31464 17098 31476
rect 17221 31467 17279 31473
rect 17221 31464 17233 31467
rect 17092 31436 17233 31464
rect 17092 31424 17098 31436
rect 17221 31433 17233 31436
rect 17267 31433 17279 31467
rect 17221 31427 17279 31433
rect 18322 31424 18328 31476
rect 18380 31464 18386 31476
rect 18693 31467 18751 31473
rect 18693 31464 18705 31467
rect 18380 31436 18705 31464
rect 18380 31424 18386 31436
rect 18693 31433 18705 31436
rect 18739 31433 18751 31467
rect 18693 31427 18751 31433
rect 19061 31467 19119 31473
rect 19061 31433 19073 31467
rect 19107 31433 19119 31467
rect 21910 31464 21916 31476
rect 21871 31436 21916 31464
rect 19061 31427 19119 31433
rect 2317 31399 2375 31405
rect 2317 31365 2329 31399
rect 2363 31365 2375 31399
rect 2317 31359 2375 31365
rect 1949 31331 2007 31337
rect 1949 31297 1961 31331
rect 1995 31328 2007 31331
rect 2130 31328 2136 31340
rect 1995 31300 2136 31328
rect 1995 31297 2007 31300
rect 1949 31291 2007 31297
rect 2130 31288 2136 31300
rect 2188 31288 2194 31340
rect 2332 31192 2360 31359
rect 3694 31356 3700 31408
rect 3752 31396 3758 31408
rect 4246 31396 4252 31408
rect 3752 31368 4016 31396
rect 3752 31356 3758 31368
rect 3605 31331 3663 31337
rect 3605 31297 3617 31331
rect 3651 31297 3663 31331
rect 3786 31328 3792 31340
rect 3747 31300 3792 31328
rect 3605 31291 3663 31297
rect 3510 31192 3516 31204
rect 2332 31164 3516 31192
rect 3510 31152 3516 31164
rect 3568 31152 3574 31204
rect 3620 31192 3648 31291
rect 3786 31288 3792 31300
rect 3844 31288 3850 31340
rect 3988 31337 4016 31368
rect 4080 31368 4252 31396
rect 3973 31331 4031 31337
rect 3973 31297 3985 31331
rect 4019 31297 4031 31331
rect 3973 31291 4031 31297
rect 3881 31263 3939 31269
rect 3881 31229 3893 31263
rect 3927 31260 3939 31263
rect 4080 31260 4108 31368
rect 4246 31356 4252 31368
rect 4304 31396 4310 31408
rect 7834 31396 7840 31408
rect 4304 31368 4568 31396
rect 4304 31356 4310 31368
rect 4157 31331 4215 31337
rect 4157 31297 4169 31331
rect 4203 31328 4215 31331
rect 4430 31328 4436 31340
rect 4203 31300 4436 31328
rect 4203 31297 4215 31300
rect 4157 31291 4215 31297
rect 4430 31288 4436 31300
rect 4488 31288 4494 31340
rect 4540 31328 4568 31368
rect 6932 31368 7840 31396
rect 5077 31331 5135 31337
rect 5077 31328 5089 31331
rect 4540 31300 5089 31328
rect 5077 31297 5089 31300
rect 5123 31297 5135 31331
rect 6546 31328 6552 31340
rect 6507 31300 6552 31328
rect 5077 31291 5135 31297
rect 6546 31288 6552 31300
rect 6604 31288 6610 31340
rect 6730 31328 6736 31340
rect 6691 31300 6736 31328
rect 6730 31288 6736 31300
rect 6788 31288 6794 31340
rect 6932 31337 6960 31368
rect 7834 31356 7840 31368
rect 7892 31356 7898 31408
rect 12710 31396 12716 31408
rect 11987 31368 12716 31396
rect 6917 31331 6975 31337
rect 6917 31297 6929 31331
rect 6963 31297 6975 31331
rect 7098 31328 7104 31340
rect 7059 31300 7104 31328
rect 6917 31291 6975 31297
rect 7098 31288 7104 31300
rect 7156 31288 7162 31340
rect 7282 31288 7288 31340
rect 7340 31328 7346 31340
rect 7745 31331 7803 31337
rect 7745 31328 7757 31331
rect 7340 31300 7757 31328
rect 7340 31288 7346 31300
rect 7745 31297 7757 31300
rect 7791 31297 7803 31331
rect 7745 31291 7803 31297
rect 8294 31288 8300 31340
rect 8352 31328 8358 31340
rect 8389 31331 8447 31337
rect 8389 31328 8401 31331
rect 8352 31300 8401 31328
rect 8352 31288 8358 31300
rect 8389 31297 8401 31300
rect 8435 31297 8447 31331
rect 9030 31328 9036 31340
rect 8991 31300 9036 31328
rect 8389 31291 8447 31297
rect 3927 31232 4108 31260
rect 4801 31263 4859 31269
rect 3927 31229 3939 31232
rect 3881 31223 3939 31229
rect 4801 31229 4813 31263
rect 4847 31260 4859 31263
rect 4847 31232 5120 31260
rect 4847 31229 4859 31232
rect 4801 31223 4859 31229
rect 5092 31204 5120 31232
rect 6822 31220 6828 31272
rect 6880 31260 6886 31272
rect 6880 31232 6925 31260
rect 6880 31220 6886 31232
rect 3620 31164 4292 31192
rect 4264 31136 4292 31164
rect 5074 31152 5080 31204
rect 5132 31152 5138 31204
rect 6914 31152 6920 31204
rect 6972 31192 6978 31204
rect 8404 31192 8432 31291
rect 9030 31288 9036 31300
rect 9088 31288 9094 31340
rect 9493 31331 9551 31337
rect 9493 31297 9505 31331
rect 9539 31328 9551 31331
rect 10318 31328 10324 31340
rect 9539 31300 10324 31328
rect 9539 31297 9551 31300
rect 9493 31291 9551 31297
rect 10318 31288 10324 31300
rect 10376 31288 10382 31340
rect 10413 31331 10471 31337
rect 10413 31297 10425 31331
rect 10459 31328 10471 31331
rect 10502 31328 10508 31340
rect 10459 31300 10508 31328
rect 10459 31297 10471 31300
rect 10413 31291 10471 31297
rect 10502 31288 10508 31300
rect 10560 31288 10566 31340
rect 11987 31337 12015 31368
rect 12710 31356 12716 31368
rect 12768 31396 12774 31408
rect 12768 31368 13446 31396
rect 12768 31356 12774 31368
rect 11972 31331 12030 31337
rect 11972 31297 11984 31331
rect 12018 31297 12030 31331
rect 11972 31291 12030 31297
rect 12069 31331 12127 31337
rect 12069 31297 12081 31331
rect 12115 31297 12127 31331
rect 12069 31291 12127 31297
rect 12161 31331 12219 31337
rect 12161 31297 12173 31331
rect 12207 31297 12219 31331
rect 12161 31291 12219 31297
rect 12344 31331 12402 31337
rect 12344 31297 12356 31331
rect 12390 31297 12402 31331
rect 12344 31291 12402 31297
rect 10226 31220 10232 31272
rect 10284 31260 10290 31272
rect 12084 31260 12112 31291
rect 10284 31232 12112 31260
rect 10284 31220 10290 31232
rect 12176 31192 12204 31291
rect 12360 31260 12388 31291
rect 12434 31288 12440 31340
rect 12492 31328 12498 31340
rect 12894 31328 12900 31340
rect 12492 31300 12537 31328
rect 12855 31300 12900 31328
rect 12492 31288 12498 31300
rect 12894 31288 12900 31300
rect 12952 31288 12958 31340
rect 12986 31288 12992 31340
rect 13044 31328 13050 31340
rect 13173 31331 13231 31337
rect 13044 31300 13089 31328
rect 13044 31288 13050 31300
rect 13173 31297 13185 31331
rect 13219 31297 13231 31331
rect 13173 31291 13231 31297
rect 13078 31260 13084 31272
rect 12360 31232 13084 31260
rect 13078 31220 13084 31232
rect 13136 31220 13142 31272
rect 13188 31260 13216 31291
rect 13262 31288 13268 31340
rect 13320 31328 13326 31340
rect 13418 31337 13446 31368
rect 15856 31368 17448 31396
rect 13401 31331 13459 31337
rect 13320 31300 13365 31328
rect 13320 31288 13326 31300
rect 13401 31297 13413 31331
rect 13447 31297 13459 31331
rect 13401 31291 13459 31297
rect 15562 31288 15568 31340
rect 15620 31328 15626 31340
rect 15749 31331 15807 31337
rect 15749 31328 15761 31331
rect 15620 31300 15761 31328
rect 15620 31288 15626 31300
rect 15749 31297 15761 31300
rect 15795 31297 15807 31331
rect 15749 31291 15807 31297
rect 15010 31260 15016 31272
rect 13188 31232 15016 31260
rect 15010 31220 15016 31232
rect 15068 31260 15074 31272
rect 15378 31260 15384 31272
rect 15068 31232 15384 31260
rect 15068 31220 15074 31232
rect 15378 31220 15384 31232
rect 15436 31220 15442 31272
rect 15856 31269 15884 31368
rect 17218 31288 17224 31340
rect 17276 31328 17282 31340
rect 17313 31331 17371 31337
rect 17313 31328 17325 31331
rect 17276 31300 17325 31328
rect 17276 31288 17282 31300
rect 17313 31297 17325 31300
rect 17359 31297 17371 31331
rect 17420 31328 17448 31368
rect 18414 31356 18420 31408
rect 18472 31396 18478 31408
rect 19076 31396 19104 31427
rect 21910 31424 21916 31436
rect 21968 31424 21974 31476
rect 18472 31368 19104 31396
rect 18472 31356 18478 31368
rect 19978 31356 19984 31408
rect 20036 31396 20042 31408
rect 20073 31399 20131 31405
rect 20073 31396 20085 31399
rect 20036 31368 20085 31396
rect 20036 31356 20042 31368
rect 20073 31365 20085 31368
rect 20119 31365 20131 31399
rect 20073 31359 20131 31365
rect 18601 31331 18659 31337
rect 18601 31328 18613 31331
rect 17420 31300 18613 31328
rect 17313 31291 17371 31297
rect 18601 31297 18613 31300
rect 18647 31297 18659 31331
rect 18601 31291 18659 31297
rect 20162 31288 20168 31340
rect 20220 31328 20226 31340
rect 20901 31331 20959 31337
rect 20901 31328 20913 31331
rect 20220 31300 20913 31328
rect 20220 31288 20226 31300
rect 20901 31297 20913 31300
rect 20947 31297 20959 31331
rect 20901 31291 20959 31297
rect 21634 31288 21640 31340
rect 21692 31328 21698 31340
rect 21821 31331 21879 31337
rect 21821 31328 21833 31331
rect 21692 31300 21833 31328
rect 21692 31288 21698 31300
rect 21821 31297 21833 31300
rect 21867 31297 21879 31331
rect 21821 31291 21879 31297
rect 15841 31263 15899 31269
rect 15841 31229 15853 31263
rect 15887 31229 15899 31263
rect 15841 31223 15899 31229
rect 16025 31263 16083 31269
rect 16025 31229 16037 31263
rect 16071 31229 16083 31263
rect 17126 31260 17132 31272
rect 17087 31232 17132 31260
rect 16025 31223 16083 31229
rect 14734 31192 14740 31204
rect 6972 31164 8432 31192
rect 9692 31164 10548 31192
rect 12176 31164 14740 31192
rect 6972 31152 6978 31164
rect 9692 31136 9720 31164
rect 2314 31124 2320 31136
rect 2275 31096 2320 31124
rect 2314 31084 2320 31096
rect 2372 31084 2378 31136
rect 3418 31124 3424 31136
rect 3379 31096 3424 31124
rect 3418 31084 3424 31096
rect 3476 31084 3482 31136
rect 4246 31084 4252 31136
rect 4304 31084 4310 31136
rect 6362 31124 6368 31136
rect 6323 31096 6368 31124
rect 6362 31084 6368 31096
rect 6420 31084 6426 31136
rect 7558 31124 7564 31136
rect 7519 31096 7564 31124
rect 7558 31084 7564 31096
rect 7616 31084 7622 31136
rect 8846 31124 8852 31136
rect 8807 31096 8852 31124
rect 8846 31084 8852 31096
rect 8904 31124 8910 31136
rect 9585 31127 9643 31133
rect 9585 31124 9597 31127
rect 8904 31096 9597 31124
rect 8904 31084 8910 31096
rect 9585 31093 9597 31096
rect 9631 31124 9643 31127
rect 9674 31124 9680 31136
rect 9631 31096 9680 31124
rect 9631 31093 9643 31096
rect 9585 31087 9643 31093
rect 9674 31084 9680 31096
rect 9732 31084 9738 31136
rect 9953 31127 10011 31133
rect 9953 31093 9965 31127
rect 9999 31124 10011 31127
rect 10042 31124 10048 31136
rect 9999 31096 10048 31124
rect 9999 31093 10011 31096
rect 9953 31087 10011 31093
rect 10042 31084 10048 31096
rect 10100 31084 10106 31136
rect 10520 31133 10548 31164
rect 14734 31152 14740 31164
rect 14792 31152 14798 31204
rect 15856 31192 15884 31223
rect 15396 31164 15884 31192
rect 16040 31192 16068 31223
rect 17126 31220 17132 31232
rect 17184 31220 17190 31272
rect 18417 31263 18475 31269
rect 18417 31229 18429 31263
rect 18463 31229 18475 31263
rect 18417 31223 18475 31229
rect 18432 31192 18460 31223
rect 19702 31192 19708 31204
rect 16040 31164 19708 31192
rect 15396 31136 15424 31164
rect 19702 31152 19708 31164
rect 19760 31152 19766 31204
rect 20257 31195 20315 31201
rect 20257 31161 20269 31195
rect 20303 31192 20315 31195
rect 20438 31192 20444 31204
rect 20303 31164 20444 31192
rect 20303 31161 20315 31164
rect 20257 31155 20315 31161
rect 20438 31152 20444 31164
rect 20496 31152 20502 31204
rect 10505 31127 10563 31133
rect 10505 31093 10517 31127
rect 10551 31093 10563 31127
rect 10505 31087 10563 31093
rect 10686 31084 10692 31136
rect 10744 31124 10750 31136
rect 10873 31127 10931 31133
rect 10873 31124 10885 31127
rect 10744 31096 10885 31124
rect 10744 31084 10750 31096
rect 10873 31093 10885 31096
rect 10919 31093 10931 31127
rect 10873 31087 10931 31093
rect 15378 31084 15384 31136
rect 15436 31084 15442 31136
rect 17681 31127 17739 31133
rect 17681 31093 17693 31127
rect 17727 31124 17739 31127
rect 17862 31124 17868 31136
rect 17727 31096 17868 31124
rect 17727 31093 17739 31096
rect 17681 31087 17739 31093
rect 17862 31084 17868 31096
rect 17920 31084 17926 31136
rect 20530 31084 20536 31136
rect 20588 31124 20594 31136
rect 20809 31127 20867 31133
rect 20809 31124 20821 31127
rect 20588 31096 20821 31124
rect 20588 31084 20594 31096
rect 20809 31093 20821 31096
rect 20855 31093 20867 31127
rect 20809 31087 20867 31093
rect 1104 31034 30820 31056
rect 1104 30982 5915 31034
rect 5967 30982 5979 31034
rect 6031 30982 6043 31034
rect 6095 30982 6107 31034
rect 6159 30982 6171 31034
rect 6223 30982 15846 31034
rect 15898 30982 15910 31034
rect 15962 30982 15974 31034
rect 16026 30982 16038 31034
rect 16090 30982 16102 31034
rect 16154 30982 25776 31034
rect 25828 30982 25840 31034
rect 25892 30982 25904 31034
rect 25956 30982 25968 31034
rect 26020 30982 26032 31034
rect 26084 30982 30820 31034
rect 1104 30960 30820 30982
rect 2314 30920 2320 30932
rect 2227 30892 2320 30920
rect 2314 30880 2320 30892
rect 2372 30920 2378 30932
rect 2682 30920 2688 30932
rect 2372 30892 2688 30920
rect 2372 30880 2378 30892
rect 2682 30880 2688 30892
rect 2740 30880 2746 30932
rect 8297 30923 8355 30929
rect 8297 30889 8309 30923
rect 8343 30920 8355 30923
rect 8846 30920 8852 30932
rect 8343 30892 8852 30920
rect 8343 30889 8355 30892
rect 8297 30883 8355 30889
rect 8846 30880 8852 30892
rect 8904 30920 8910 30932
rect 9125 30923 9183 30929
rect 9125 30920 9137 30923
rect 8904 30892 9137 30920
rect 8904 30880 8910 30892
rect 9125 30889 9137 30892
rect 9171 30889 9183 30923
rect 11882 30920 11888 30932
rect 11843 30892 11888 30920
rect 9125 30883 9183 30889
rect 11882 30880 11888 30892
rect 11940 30880 11946 30932
rect 29822 30880 29828 30932
rect 29880 30920 29886 30932
rect 29917 30923 29975 30929
rect 29917 30920 29929 30923
rect 29880 30892 29929 30920
rect 29880 30880 29886 30892
rect 29917 30889 29929 30892
rect 29963 30889 29975 30923
rect 29917 30883 29975 30889
rect 1949 30855 2007 30861
rect 1949 30821 1961 30855
rect 1995 30852 2007 30855
rect 2130 30852 2136 30864
rect 1995 30824 2136 30852
rect 1995 30821 2007 30824
rect 1949 30815 2007 30821
rect 2130 30812 2136 30824
rect 2188 30812 2194 30864
rect 3973 30855 4031 30861
rect 3973 30821 3985 30855
rect 4019 30852 4031 30855
rect 4019 30824 5672 30852
rect 4019 30821 4031 30824
rect 3973 30815 4031 30821
rect 3510 30744 3516 30796
rect 3568 30784 3574 30796
rect 4893 30787 4951 30793
rect 3568 30756 4660 30784
rect 3568 30744 3574 30756
rect 2961 30719 3019 30725
rect 2961 30685 2973 30719
rect 3007 30716 3019 30719
rect 3050 30716 3056 30728
rect 3007 30688 3056 30716
rect 3007 30685 3019 30688
rect 2961 30679 3019 30685
rect 3050 30676 3056 30688
rect 3108 30676 3114 30728
rect 3789 30719 3847 30725
rect 3789 30685 3801 30719
rect 3835 30716 3847 30719
rect 4522 30716 4528 30728
rect 3835 30688 4528 30716
rect 3835 30685 3847 30688
rect 3789 30679 3847 30685
rect 4522 30676 4528 30688
rect 4580 30676 4586 30728
rect 4632 30725 4660 30756
rect 4893 30753 4905 30787
rect 4939 30784 4951 30787
rect 5074 30784 5080 30796
rect 4939 30756 5080 30784
rect 4939 30753 4951 30756
rect 4893 30747 4951 30753
rect 5074 30744 5080 30756
rect 5132 30744 5138 30796
rect 5644 30793 5672 30824
rect 10318 30812 10324 30864
rect 10376 30852 10382 30864
rect 13262 30852 13268 30864
rect 10376 30824 13268 30852
rect 10376 30812 10382 30824
rect 13262 30812 13268 30824
rect 13320 30812 13326 30864
rect 20714 30812 20720 30864
rect 20772 30852 20778 30864
rect 20993 30855 21051 30861
rect 20993 30852 21005 30855
rect 20772 30824 21005 30852
rect 20772 30812 20778 30824
rect 20993 30821 21005 30824
rect 21039 30821 21051 30855
rect 20993 30815 21051 30821
rect 5629 30787 5687 30793
rect 5629 30753 5641 30787
rect 5675 30753 5687 30787
rect 5629 30747 5687 30753
rect 10594 30744 10600 30796
rect 10652 30784 10658 30796
rect 11517 30787 11575 30793
rect 10652 30756 11376 30784
rect 10652 30744 10658 30756
rect 4617 30719 4675 30725
rect 4617 30685 4629 30719
rect 4663 30716 4675 30719
rect 4706 30716 4712 30728
rect 4663 30688 4712 30716
rect 4663 30685 4675 30688
rect 4617 30679 4675 30685
rect 4706 30676 4712 30688
rect 4764 30676 4770 30728
rect 4798 30676 4804 30728
rect 4856 30716 4862 30728
rect 4985 30719 5043 30725
rect 4856 30688 4901 30716
rect 4856 30676 4862 30688
rect 4985 30685 4997 30719
rect 5031 30685 5043 30719
rect 5166 30716 5172 30728
rect 5127 30688 5172 30716
rect 4985 30679 5043 30685
rect 2317 30651 2375 30657
rect 2317 30617 2329 30651
rect 2363 30648 2375 30651
rect 5000 30648 5028 30679
rect 5166 30676 5172 30688
rect 5224 30676 5230 30728
rect 5896 30719 5954 30725
rect 5896 30685 5908 30719
rect 5942 30716 5954 30719
rect 6362 30716 6368 30728
rect 5942 30688 6368 30716
rect 5942 30685 5954 30688
rect 5896 30679 5954 30685
rect 6362 30676 6368 30688
rect 6420 30676 6426 30728
rect 7926 30676 7932 30728
rect 7984 30676 7990 30728
rect 8110 30676 8116 30728
rect 8168 30716 8174 30728
rect 8389 30719 8447 30725
rect 8389 30716 8401 30719
rect 8168 30688 8401 30716
rect 8168 30676 8174 30688
rect 8389 30685 8401 30688
rect 8435 30685 8447 30719
rect 8389 30679 8447 30685
rect 9214 30676 9220 30728
rect 9272 30716 9278 30728
rect 9401 30719 9459 30725
rect 9401 30716 9413 30719
rect 9272 30688 9413 30716
rect 9272 30676 9278 30688
rect 9401 30685 9413 30688
rect 9447 30685 9459 30719
rect 10042 30716 10048 30728
rect 10003 30688 10048 30716
rect 9401 30679 9459 30685
rect 10042 30676 10048 30688
rect 10100 30676 10106 30728
rect 10686 30716 10692 30728
rect 10647 30688 10692 30716
rect 10686 30676 10692 30688
rect 10744 30676 10750 30728
rect 11348 30725 11376 30756
rect 11517 30753 11529 30787
rect 11563 30784 11575 30787
rect 11882 30784 11888 30796
rect 11563 30756 11888 30784
rect 11563 30753 11575 30756
rect 11517 30747 11575 30753
rect 11882 30744 11888 30756
rect 11940 30744 11946 30796
rect 12802 30744 12808 30796
rect 12860 30784 12866 30796
rect 13173 30787 13231 30793
rect 13173 30784 13185 30787
rect 12860 30756 13185 30784
rect 12860 30744 12866 30756
rect 13173 30753 13185 30756
rect 13219 30753 13231 30787
rect 13173 30747 13231 30753
rect 16853 30787 16911 30793
rect 16853 30753 16865 30787
rect 16899 30784 16911 30787
rect 17126 30784 17132 30796
rect 16899 30756 17132 30784
rect 16899 30753 16911 30756
rect 16853 30747 16911 30753
rect 17126 30744 17132 30756
rect 17184 30784 17190 30796
rect 17494 30784 17500 30796
rect 17184 30756 17500 30784
rect 17184 30744 17190 30756
rect 17494 30744 17500 30756
rect 17552 30744 17558 30796
rect 17954 30784 17960 30796
rect 17915 30756 17960 30784
rect 17954 30744 17960 30756
rect 18012 30744 18018 30796
rect 19242 30784 19248 30796
rect 18156 30756 19248 30784
rect 11149 30719 11207 30725
rect 11149 30685 11161 30719
rect 11195 30685 11207 30719
rect 11149 30679 11207 30685
rect 11333 30719 11391 30725
rect 11333 30685 11345 30719
rect 11379 30685 11391 30719
rect 11333 30679 11391 30685
rect 7944 30648 7972 30676
rect 2363 30620 4936 30648
rect 5000 30620 7972 30648
rect 11164 30648 11192 30679
rect 11422 30676 11428 30728
rect 11480 30716 11486 30728
rect 11701 30719 11759 30725
rect 11480 30688 11525 30716
rect 11480 30676 11486 30688
rect 11701 30685 11713 30719
rect 11747 30716 11759 30719
rect 12618 30716 12624 30728
rect 11747 30688 12624 30716
rect 11747 30685 11759 30688
rect 11701 30679 11759 30685
rect 12618 30676 12624 30688
rect 12676 30676 12682 30728
rect 12897 30719 12955 30725
rect 12897 30685 12909 30719
rect 12943 30716 12955 30719
rect 12986 30716 12992 30728
rect 12943 30688 12992 30716
rect 12943 30685 12955 30688
rect 12897 30679 12955 30685
rect 12986 30676 12992 30688
rect 13044 30676 13050 30728
rect 14182 30676 14188 30728
rect 14240 30716 14246 30728
rect 14277 30719 14335 30725
rect 14277 30716 14289 30719
rect 14240 30688 14289 30716
rect 14240 30676 14246 30688
rect 14277 30685 14289 30688
rect 14323 30685 14335 30719
rect 14277 30679 14335 30685
rect 16945 30719 17003 30725
rect 16945 30685 16957 30719
rect 16991 30716 17003 30719
rect 17034 30716 17040 30728
rect 16991 30688 17040 30716
rect 16991 30685 17003 30688
rect 16945 30679 17003 30685
rect 17034 30676 17040 30688
rect 17092 30676 17098 30728
rect 17862 30716 17868 30728
rect 17823 30688 17868 30716
rect 17862 30676 17868 30688
rect 17920 30676 17926 30728
rect 18156 30725 18184 30756
rect 19242 30744 19248 30756
rect 19300 30744 19306 30796
rect 20254 30784 20260 30796
rect 20215 30756 20260 30784
rect 20254 30744 20260 30756
rect 20312 30744 20318 30796
rect 20530 30784 20536 30796
rect 20491 30756 20536 30784
rect 20530 30744 20536 30756
rect 20588 30744 20594 30796
rect 18141 30719 18199 30725
rect 18141 30685 18153 30719
rect 18187 30685 18199 30719
rect 18141 30679 18199 30685
rect 18233 30719 18291 30725
rect 18233 30685 18245 30719
rect 18279 30685 18291 30719
rect 18233 30679 18291 30685
rect 14544 30651 14602 30657
rect 11164 30620 11560 30648
rect 2363 30617 2375 30620
rect 2317 30611 2375 30617
rect 2498 30580 2504 30592
rect 2459 30552 2504 30580
rect 2498 30540 2504 30552
rect 2556 30540 2562 30592
rect 3142 30580 3148 30592
rect 3103 30552 3148 30580
rect 3142 30540 3148 30552
rect 3200 30540 3206 30592
rect 4154 30540 4160 30592
rect 4212 30580 4218 30592
rect 4433 30583 4491 30589
rect 4433 30580 4445 30583
rect 4212 30552 4445 30580
rect 4212 30540 4218 30552
rect 4433 30549 4445 30552
rect 4479 30549 4491 30583
rect 4908 30580 4936 30620
rect 11532 30592 11560 30620
rect 14544 30617 14556 30651
rect 14590 30648 14602 30651
rect 14734 30648 14740 30660
rect 14590 30620 14740 30648
rect 14590 30617 14602 30620
rect 14544 30611 14602 30617
rect 14734 30608 14740 30620
rect 14792 30608 14798 30660
rect 18248 30648 18276 30679
rect 29546 30676 29552 30728
rect 29604 30716 29610 30728
rect 29917 30719 29975 30725
rect 29917 30716 29929 30719
rect 29604 30688 29929 30716
rect 29604 30676 29610 30688
rect 29917 30685 29929 30688
rect 29963 30685 29975 30719
rect 30098 30716 30104 30728
rect 30059 30688 30104 30716
rect 29917 30679 29975 30685
rect 30098 30676 30104 30688
rect 30156 30676 30162 30728
rect 21174 30648 21180 30660
rect 17420 30620 18276 30648
rect 21135 30620 21180 30648
rect 6546 30580 6552 30592
rect 4908 30552 6552 30580
rect 4433 30543 4491 30549
rect 6546 30540 6552 30552
rect 6604 30580 6610 30592
rect 7009 30583 7067 30589
rect 7009 30580 7021 30583
rect 6604 30552 7021 30580
rect 6604 30540 6610 30552
rect 7009 30549 7021 30552
rect 7055 30549 7067 30583
rect 7926 30580 7932 30592
rect 7887 30552 7932 30580
rect 7009 30543 7067 30549
rect 7926 30540 7932 30552
rect 7984 30540 7990 30592
rect 8570 30540 8576 30592
rect 8628 30580 8634 30592
rect 8941 30583 8999 30589
rect 8941 30580 8953 30583
rect 8628 30552 8953 30580
rect 8628 30540 8634 30552
rect 8941 30549 8953 30552
rect 8987 30549 8999 30583
rect 8941 30543 8999 30549
rect 9214 30540 9220 30592
rect 9272 30580 9278 30592
rect 9861 30583 9919 30589
rect 9861 30580 9873 30583
rect 9272 30552 9873 30580
rect 9272 30540 9278 30552
rect 9861 30549 9873 30552
rect 9907 30549 9919 30583
rect 10502 30580 10508 30592
rect 10463 30552 10508 30580
rect 9861 30543 9919 30549
rect 10502 30540 10508 30552
rect 10560 30540 10566 30592
rect 11514 30540 11520 30592
rect 11572 30540 11578 30592
rect 15654 30580 15660 30592
rect 15615 30552 15660 30580
rect 15654 30540 15660 30552
rect 15712 30540 15718 30592
rect 17037 30583 17095 30589
rect 17037 30549 17049 30583
rect 17083 30580 17095 30583
rect 17218 30580 17224 30592
rect 17083 30552 17224 30580
rect 17083 30549 17095 30552
rect 17037 30543 17095 30549
rect 17218 30540 17224 30552
rect 17276 30540 17282 30592
rect 17420 30589 17448 30620
rect 21174 30608 21180 30620
rect 21232 30608 21238 30660
rect 21361 30651 21419 30657
rect 21361 30617 21373 30651
rect 21407 30648 21419 30651
rect 21634 30648 21640 30660
rect 21407 30620 21640 30648
rect 21407 30617 21419 30620
rect 21361 30611 21419 30617
rect 21634 30608 21640 30620
rect 21692 30608 21698 30660
rect 17405 30583 17463 30589
rect 17405 30549 17417 30583
rect 17451 30549 17463 30583
rect 17405 30543 17463 30549
rect 18417 30583 18475 30589
rect 18417 30549 18429 30583
rect 18463 30580 18475 30583
rect 19426 30580 19432 30592
rect 18463 30552 19432 30580
rect 18463 30549 18475 30552
rect 18417 30543 18475 30549
rect 19426 30540 19432 30552
rect 19484 30540 19490 30592
rect 1104 30490 30820 30512
rect 1104 30438 10880 30490
rect 10932 30438 10944 30490
rect 10996 30438 11008 30490
rect 11060 30438 11072 30490
rect 11124 30438 11136 30490
rect 11188 30438 20811 30490
rect 20863 30438 20875 30490
rect 20927 30438 20939 30490
rect 20991 30438 21003 30490
rect 21055 30438 21067 30490
rect 21119 30438 30820 30490
rect 1104 30416 30820 30438
rect 2225 30379 2283 30385
rect 2225 30345 2237 30379
rect 2271 30376 2283 30379
rect 4246 30376 4252 30388
rect 2271 30348 4108 30376
rect 4207 30348 4252 30376
rect 2271 30345 2283 30348
rect 2225 30339 2283 30345
rect 3136 30311 3194 30317
rect 3136 30277 3148 30311
rect 3182 30308 3194 30311
rect 3418 30308 3424 30320
rect 3182 30280 3424 30308
rect 3182 30277 3194 30280
rect 3136 30271 3194 30277
rect 3418 30268 3424 30280
rect 3476 30268 3482 30320
rect 4080 30308 4108 30348
rect 4246 30336 4252 30348
rect 4304 30336 4310 30388
rect 4522 30336 4528 30388
rect 4580 30376 4586 30388
rect 4709 30379 4767 30385
rect 4709 30376 4721 30379
rect 4580 30348 4721 30376
rect 4580 30336 4586 30348
rect 4709 30345 4721 30348
rect 4755 30345 4767 30379
rect 12986 30376 12992 30388
rect 4709 30339 4767 30345
rect 4816 30348 5580 30376
rect 4816 30320 4844 30348
rect 4798 30308 4804 30320
rect 4080 30280 4804 30308
rect 4798 30268 4804 30280
rect 4856 30268 4862 30320
rect 5442 30308 5448 30320
rect 4908 30280 5448 30308
rect 1857 30243 1915 30249
rect 1857 30209 1869 30243
rect 1903 30240 1915 30243
rect 2130 30240 2136 30252
rect 1903 30212 2136 30240
rect 1903 30209 1915 30212
rect 1857 30203 1915 30209
rect 2130 30200 2136 30212
rect 2188 30200 2194 30252
rect 4614 30200 4620 30252
rect 4672 30240 4678 30252
rect 4908 30249 4936 30280
rect 5442 30268 5448 30280
rect 5500 30268 5506 30320
rect 4893 30243 4951 30249
rect 4893 30240 4905 30243
rect 4672 30212 4905 30240
rect 4672 30200 4678 30212
rect 4893 30209 4905 30212
rect 4939 30209 4951 30243
rect 5350 30240 5356 30252
rect 5311 30212 5356 30240
rect 4893 30203 4951 30209
rect 5350 30200 5356 30212
rect 5408 30200 5414 30252
rect 5552 30240 5580 30348
rect 11716 30348 12992 30376
rect 8018 30308 8024 30320
rect 6932 30280 8024 30308
rect 6549 30243 6607 30249
rect 6549 30240 6561 30243
rect 5552 30212 6561 30240
rect 6549 30209 6561 30212
rect 6595 30209 6607 30243
rect 6822 30240 6828 30252
rect 6549 30203 6607 30209
rect 6656 30212 6828 30240
rect 2866 30172 2872 30184
rect 2827 30144 2872 30172
rect 2866 30132 2872 30144
rect 2924 30132 2930 30184
rect 5074 30132 5080 30184
rect 5132 30172 5138 30184
rect 5445 30175 5503 30181
rect 5445 30172 5457 30175
rect 5132 30144 5457 30172
rect 5132 30132 5138 30144
rect 5445 30141 5457 30144
rect 5491 30172 5503 30175
rect 6656 30172 6684 30212
rect 6822 30200 6828 30212
rect 6880 30200 6886 30252
rect 6932 30249 6960 30280
rect 8018 30268 8024 30280
rect 8076 30268 8082 30320
rect 10870 30268 10876 30320
rect 10928 30308 10934 30320
rect 10965 30311 11023 30317
rect 10965 30308 10977 30311
rect 10928 30280 10977 30308
rect 10928 30268 10934 30280
rect 10965 30277 10977 30280
rect 11011 30277 11023 30311
rect 10965 30271 11023 30277
rect 6917 30243 6975 30249
rect 6917 30209 6929 30243
rect 6963 30209 6975 30243
rect 7098 30240 7104 30252
rect 7059 30212 7104 30240
rect 6917 30203 6975 30209
rect 7098 30200 7104 30212
rect 7156 30200 7162 30252
rect 7926 30240 7932 30252
rect 7887 30212 7932 30240
rect 7926 30200 7932 30212
rect 7984 30200 7990 30252
rect 8570 30240 8576 30252
rect 8531 30212 8576 30240
rect 8570 30200 8576 30212
rect 8628 30200 8634 30252
rect 9122 30240 9128 30252
rect 9083 30212 9128 30240
rect 9122 30200 9128 30212
rect 9180 30200 9186 30252
rect 10410 30200 10416 30252
rect 10468 30240 10474 30252
rect 10781 30243 10839 30249
rect 10781 30240 10793 30243
rect 10468 30212 10793 30240
rect 10468 30200 10474 30212
rect 10781 30209 10793 30212
rect 10827 30209 10839 30243
rect 11514 30240 11520 30252
rect 11475 30212 11520 30240
rect 10781 30203 10839 30209
rect 11514 30200 11520 30212
rect 11572 30200 11578 30252
rect 11716 30249 11744 30348
rect 12986 30336 12992 30348
rect 13044 30336 13050 30388
rect 14734 30376 14740 30388
rect 14695 30348 14740 30376
rect 14734 30336 14740 30348
rect 14792 30336 14798 30388
rect 18969 30379 19027 30385
rect 18969 30345 18981 30379
rect 19015 30376 19027 30379
rect 19518 30376 19524 30388
rect 19015 30348 19524 30376
rect 19015 30345 19027 30348
rect 18969 30339 19027 30345
rect 19518 30336 19524 30348
rect 19576 30376 19582 30388
rect 19797 30379 19855 30385
rect 19797 30376 19809 30379
rect 19576 30348 19809 30376
rect 19576 30336 19582 30348
rect 19797 30345 19809 30348
rect 19843 30376 19855 30379
rect 20070 30376 20076 30388
rect 19843 30348 20076 30376
rect 19843 30345 19855 30348
rect 19797 30339 19855 30345
rect 20070 30336 20076 30348
rect 20128 30336 20134 30388
rect 12250 30308 12256 30320
rect 12211 30280 12256 30308
rect 12250 30268 12256 30280
rect 12308 30268 12314 30320
rect 12434 30268 12440 30320
rect 12492 30308 12498 30320
rect 12492 30280 13216 30308
rect 12492 30268 12498 30280
rect 11701 30243 11759 30249
rect 11701 30209 11713 30243
rect 11747 30209 11759 30243
rect 11701 30203 11759 30209
rect 12069 30243 12127 30249
rect 12069 30209 12081 30243
rect 12115 30240 12127 30243
rect 12158 30240 12164 30252
rect 12115 30212 12164 30240
rect 12115 30209 12127 30212
rect 12069 30203 12127 30209
rect 12158 30200 12164 30212
rect 12216 30200 12222 30252
rect 13078 30240 13084 30252
rect 13039 30212 13084 30240
rect 13078 30200 13084 30212
rect 13136 30200 13142 30252
rect 13188 30240 13216 30280
rect 13354 30268 13360 30320
rect 13412 30308 13418 30320
rect 15289 30311 15347 30317
rect 15289 30308 15301 30311
rect 13412 30280 15301 30308
rect 13412 30268 13418 30280
rect 15289 30277 15301 30280
rect 15335 30277 15347 30311
rect 15470 30308 15476 30320
rect 15431 30280 15476 30308
rect 15289 30271 15347 30277
rect 15470 30268 15476 30280
rect 15528 30268 15534 30320
rect 18887 30311 18945 30317
rect 18887 30277 18899 30311
rect 18933 30308 18945 30311
rect 19334 30308 19340 30320
rect 18933 30280 19340 30308
rect 18933 30277 18945 30280
rect 18887 30271 18945 30277
rect 19334 30268 19340 30280
rect 19392 30308 19398 30320
rect 19878 30311 19936 30317
rect 19878 30308 19890 30311
rect 19392 30280 19890 30308
rect 19392 30268 19398 30280
rect 19878 30277 19890 30280
rect 19924 30277 19936 30311
rect 19878 30271 19936 30277
rect 19981 30311 20039 30317
rect 19981 30277 19993 30311
rect 20027 30308 20039 30311
rect 20530 30308 20536 30320
rect 20027 30280 20536 30308
rect 20027 30277 20039 30280
rect 19981 30271 20039 30277
rect 20530 30268 20536 30280
rect 20588 30268 20594 30320
rect 30098 30308 30104 30320
rect 29196 30280 30104 30308
rect 14090 30240 14096 30252
rect 13188 30212 14096 30240
rect 14090 30200 14096 30212
rect 14148 30200 14154 30252
rect 14186 30243 14244 30249
rect 14186 30209 14198 30243
rect 14232 30209 14244 30243
rect 14186 30203 14244 30209
rect 14369 30243 14427 30249
rect 14369 30209 14381 30243
rect 14415 30209 14427 30243
rect 14369 30203 14427 30209
rect 5491 30144 6684 30172
rect 5491 30141 5503 30144
rect 5445 30135 5503 30141
rect 6730 30132 6736 30184
rect 6788 30172 6794 30184
rect 10505 30175 10563 30181
rect 6788 30144 6833 30172
rect 6788 30132 6794 30144
rect 10505 30141 10517 30175
rect 10551 30172 10563 30175
rect 10594 30172 10600 30184
rect 10551 30144 10600 30172
rect 10551 30141 10563 30144
rect 10505 30135 10563 30141
rect 10594 30132 10600 30144
rect 10652 30132 10658 30184
rect 10686 30132 10692 30184
rect 10744 30172 10750 30184
rect 11793 30175 11851 30181
rect 11793 30172 11805 30175
rect 10744 30144 11805 30172
rect 10744 30132 10750 30144
rect 11793 30141 11805 30144
rect 11839 30141 11851 30175
rect 11793 30135 11851 30141
rect 11882 30132 11888 30184
rect 11940 30172 11946 30184
rect 12802 30172 12808 30184
rect 11940 30144 11985 30172
rect 12763 30144 12808 30172
rect 11940 30132 11946 30144
rect 12802 30132 12808 30144
rect 12860 30132 12866 30184
rect 13096 30172 13124 30200
rect 13446 30172 13452 30184
rect 13096 30144 13452 30172
rect 13446 30132 13452 30144
rect 13504 30172 13510 30184
rect 14200 30172 14228 30203
rect 13504 30144 14228 30172
rect 13504 30132 13510 30144
rect 2682 30104 2688 30116
rect 2240 30076 2688 30104
rect 2240 30045 2268 30076
rect 2682 30064 2688 30076
rect 2740 30064 2746 30116
rect 4890 30064 4896 30116
rect 4948 30104 4954 30116
rect 5350 30104 5356 30116
rect 4948 30076 5356 30104
rect 4948 30064 4954 30076
rect 5350 30064 5356 30076
rect 5408 30104 5414 30116
rect 6748 30104 6776 30132
rect 5408 30076 6776 30104
rect 14384 30104 14412 30203
rect 14458 30200 14464 30252
rect 14516 30240 14522 30252
rect 14642 30249 14648 30252
rect 14599 30243 14648 30249
rect 14516 30212 14561 30240
rect 14516 30200 14522 30212
rect 14599 30209 14611 30243
rect 14645 30209 14648 30243
rect 14599 30203 14648 30209
rect 14642 30200 14648 30203
rect 14700 30200 14706 30252
rect 15933 30243 15991 30249
rect 15933 30209 15945 30243
rect 15979 30209 15991 30243
rect 15933 30203 15991 30209
rect 15654 30104 15660 30116
rect 14384 30076 15660 30104
rect 5408 30064 5414 30076
rect 15654 30064 15660 30076
rect 15712 30104 15718 30116
rect 15948 30104 15976 30203
rect 16850 30200 16856 30252
rect 16908 30240 16914 30252
rect 17037 30243 17095 30249
rect 17037 30240 17049 30243
rect 16908 30212 17049 30240
rect 16908 30200 16914 30212
rect 17037 30209 17049 30212
rect 17083 30209 17095 30243
rect 17862 30240 17868 30252
rect 17823 30212 17868 30240
rect 17037 30203 17095 30209
rect 17862 30200 17868 30212
rect 17920 30200 17926 30252
rect 18785 30243 18843 30249
rect 18785 30209 18797 30243
rect 18831 30209 18843 30243
rect 19150 30240 19156 30252
rect 19111 30212 19156 30240
rect 18785 30203 18843 30209
rect 17126 30172 17132 30184
rect 17087 30144 17132 30172
rect 17126 30132 17132 30144
rect 17184 30132 17190 30184
rect 17313 30175 17371 30181
rect 17313 30141 17325 30175
rect 17359 30172 17371 30175
rect 17494 30172 17500 30184
rect 17359 30144 17500 30172
rect 17359 30141 17371 30144
rect 17313 30135 17371 30141
rect 17494 30132 17500 30144
rect 17552 30132 17558 30184
rect 18800 30172 18828 30203
rect 19150 30200 19156 30212
rect 19208 30200 19214 30252
rect 19613 30243 19671 30249
rect 19613 30209 19625 30243
rect 19659 30240 19671 30243
rect 20714 30240 20720 30252
rect 19659 30212 20720 30240
rect 19659 30209 19671 30212
rect 19613 30203 19671 30209
rect 20714 30200 20720 30212
rect 20772 30240 20778 30252
rect 20901 30243 20959 30249
rect 20901 30240 20913 30243
rect 20772 30212 20913 30240
rect 20772 30200 20778 30212
rect 20901 30209 20913 30212
rect 20947 30209 20959 30243
rect 22922 30240 22928 30252
rect 22883 30212 22928 30240
rect 20901 30203 20959 30209
rect 22922 30200 22928 30212
rect 22980 30200 22986 30252
rect 29196 30249 29224 30280
rect 30098 30268 30104 30280
rect 30156 30268 30162 30320
rect 29181 30243 29239 30249
rect 29181 30209 29193 30243
rect 29227 30209 29239 30243
rect 29825 30243 29883 30249
rect 29825 30240 29837 30243
rect 29181 30203 29239 30209
rect 29380 30212 29837 30240
rect 20254 30172 20260 30184
rect 18800 30144 20260 30172
rect 20254 30132 20260 30144
rect 20312 30132 20318 30184
rect 15712 30076 15976 30104
rect 16025 30107 16083 30113
rect 15712 30064 15718 30076
rect 16025 30073 16037 30107
rect 16071 30104 16083 30107
rect 17034 30104 17040 30116
rect 16071 30076 17040 30104
rect 16071 30073 16083 30076
rect 16025 30067 16083 30073
rect 17034 30064 17040 30076
rect 17092 30064 17098 30116
rect 18230 30064 18236 30116
rect 18288 30104 18294 30116
rect 18601 30107 18659 30113
rect 18601 30104 18613 30107
rect 18288 30076 18613 30104
rect 18288 30064 18294 30076
rect 18601 30073 18613 30076
rect 18647 30073 18659 30107
rect 20162 30104 20168 30116
rect 20123 30076 20168 30104
rect 18601 30067 18659 30073
rect 20162 30064 20168 30076
rect 20220 30064 20226 30116
rect 29380 30113 29408 30212
rect 29825 30209 29837 30212
rect 29871 30209 29883 30243
rect 29825 30203 29883 30209
rect 29365 30107 29423 30113
rect 29365 30073 29377 30107
rect 29411 30073 29423 30107
rect 30006 30104 30012 30116
rect 29967 30076 30012 30104
rect 29365 30067 29423 30073
rect 30006 30064 30012 30076
rect 30064 30064 30070 30116
rect 2225 30039 2283 30045
rect 2225 30005 2237 30039
rect 2271 30005 2283 30039
rect 2225 29999 2283 30005
rect 2314 29996 2320 30048
rect 2372 30036 2378 30048
rect 2409 30039 2467 30045
rect 2409 30036 2421 30039
rect 2372 30008 2421 30036
rect 2372 29996 2378 30008
rect 2409 30005 2421 30008
rect 2455 30005 2467 30039
rect 6362 30036 6368 30048
rect 6323 30008 6368 30036
rect 2409 29999 2467 30005
rect 6362 29996 6368 30008
rect 6420 29996 6426 30048
rect 7282 29996 7288 30048
rect 7340 30036 7346 30048
rect 7745 30039 7803 30045
rect 7745 30036 7757 30039
rect 7340 30008 7757 30036
rect 7340 29996 7346 30008
rect 7745 30005 7757 30008
rect 7791 30005 7803 30039
rect 7745 29999 7803 30005
rect 7834 29996 7840 30048
rect 7892 30036 7898 30048
rect 8389 30039 8447 30045
rect 8389 30036 8401 30039
rect 7892 30008 8401 30036
rect 7892 29996 7898 30008
rect 8389 30005 8401 30008
rect 8435 30005 8447 30039
rect 9306 30036 9312 30048
rect 9267 30008 9312 30036
rect 8389 29999 8447 30005
rect 9306 29996 9312 30008
rect 9364 29996 9370 30048
rect 9674 29996 9680 30048
rect 9732 30036 9738 30048
rect 10226 30036 10232 30048
rect 9732 30008 10232 30036
rect 9732 29996 9738 30008
rect 10226 29996 10232 30008
rect 10284 30036 10290 30048
rect 10597 30039 10655 30045
rect 10597 30036 10609 30039
rect 10284 30008 10609 30036
rect 10284 29996 10290 30008
rect 10597 30005 10609 30008
rect 10643 30005 10655 30039
rect 10597 29999 10655 30005
rect 15194 29996 15200 30048
rect 15252 30036 15258 30048
rect 16669 30039 16727 30045
rect 16669 30036 16681 30039
rect 15252 30008 16681 30036
rect 15252 29996 15258 30008
rect 16669 30005 16681 30008
rect 16715 30005 16727 30039
rect 18046 30036 18052 30048
rect 18007 30008 18052 30036
rect 16669 29999 16727 30005
rect 18046 29996 18052 30008
rect 18104 29996 18110 30048
rect 20993 30039 21051 30045
rect 20993 30005 21005 30039
rect 21039 30036 21051 30039
rect 21266 30036 21272 30048
rect 21039 30008 21272 30036
rect 21039 30005 21051 30008
rect 20993 29999 21051 30005
rect 21266 29996 21272 30008
rect 21324 29996 21330 30048
rect 22646 29996 22652 30048
rect 22704 30036 22710 30048
rect 22741 30039 22799 30045
rect 22741 30036 22753 30039
rect 22704 30008 22753 30036
rect 22704 29996 22710 30008
rect 22741 30005 22753 30008
rect 22787 30005 22799 30039
rect 22741 29999 22799 30005
rect 1104 29946 30820 29968
rect 1104 29894 5915 29946
rect 5967 29894 5979 29946
rect 6031 29894 6043 29946
rect 6095 29894 6107 29946
rect 6159 29894 6171 29946
rect 6223 29894 15846 29946
rect 15898 29894 15910 29946
rect 15962 29894 15974 29946
rect 16026 29894 16038 29946
rect 16090 29894 16102 29946
rect 16154 29894 25776 29946
rect 25828 29894 25840 29946
rect 25892 29894 25904 29946
rect 25956 29894 25968 29946
rect 26020 29894 26032 29946
rect 26084 29894 30820 29946
rect 1104 29872 30820 29894
rect 1486 29832 1492 29844
rect 1447 29804 1492 29832
rect 1486 29792 1492 29804
rect 1544 29792 1550 29844
rect 2866 29792 2872 29844
rect 2924 29832 2930 29844
rect 2961 29835 3019 29841
rect 2961 29832 2973 29835
rect 2924 29804 2973 29832
rect 2924 29792 2930 29804
rect 2961 29801 2973 29804
rect 3007 29801 3019 29835
rect 2961 29795 3019 29801
rect 4798 29792 4804 29844
rect 4856 29832 4862 29844
rect 5077 29835 5135 29841
rect 5077 29832 5089 29835
rect 4856 29804 5089 29832
rect 4856 29792 4862 29804
rect 5077 29801 5089 29804
rect 5123 29801 5135 29835
rect 5077 29795 5135 29801
rect 11057 29835 11115 29841
rect 11057 29801 11069 29835
rect 11103 29832 11115 29835
rect 11698 29832 11704 29844
rect 11103 29804 11704 29832
rect 11103 29801 11115 29804
rect 11057 29795 11115 29801
rect 11698 29792 11704 29804
rect 11756 29832 11762 29844
rect 12342 29832 12348 29844
rect 11756 29804 12348 29832
rect 11756 29792 11762 29804
rect 12342 29792 12348 29804
rect 12400 29792 12406 29844
rect 13630 29792 13636 29844
rect 13688 29832 13694 29844
rect 15565 29835 15623 29841
rect 15565 29832 15577 29835
rect 13688 29804 15577 29832
rect 13688 29792 13694 29804
rect 15565 29801 15577 29804
rect 15611 29832 15623 29835
rect 17126 29832 17132 29844
rect 15611 29804 17132 29832
rect 15611 29801 15623 29804
rect 15565 29795 15623 29801
rect 17126 29792 17132 29804
rect 17184 29792 17190 29844
rect 17218 29792 17224 29844
rect 17276 29832 17282 29844
rect 19613 29835 19671 29841
rect 19613 29832 19625 29835
rect 17276 29804 19625 29832
rect 17276 29792 17282 29804
rect 19613 29801 19625 29804
rect 19659 29801 19671 29835
rect 19613 29795 19671 29801
rect 20070 29792 20076 29844
rect 20128 29832 20134 29844
rect 20165 29835 20223 29841
rect 20165 29832 20177 29835
rect 20128 29804 20177 29832
rect 20128 29792 20134 29804
rect 20165 29801 20177 29804
rect 20211 29801 20223 29835
rect 20165 29795 20223 29801
rect 2133 29767 2191 29773
rect 2133 29733 2145 29767
rect 2179 29733 2191 29767
rect 2133 29727 2191 29733
rect 3789 29767 3847 29773
rect 3789 29733 3801 29767
rect 3835 29733 3847 29767
rect 11790 29764 11796 29776
rect 11751 29736 11796 29764
rect 3789 29727 3847 29733
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29628 1731 29631
rect 2148 29628 2176 29727
rect 2314 29628 2320 29640
rect 1719 29600 2176 29628
rect 2275 29600 2320 29628
rect 1719 29597 1731 29600
rect 1673 29591 1731 29597
rect 2314 29588 2320 29600
rect 2372 29588 2378 29640
rect 3145 29631 3203 29637
rect 3145 29597 3157 29631
rect 3191 29628 3203 29631
rect 3804 29628 3832 29727
rect 11790 29724 11796 29736
rect 11848 29764 11854 29776
rect 12158 29764 12164 29776
rect 11848 29736 12164 29764
rect 11848 29724 11854 29736
rect 12158 29724 12164 29736
rect 12216 29724 12222 29776
rect 19150 29764 19156 29776
rect 18064 29736 19156 29764
rect 18064 29708 18092 29736
rect 19150 29724 19156 29736
rect 19208 29724 19214 29776
rect 21910 29764 21916 29776
rect 19720 29736 21916 29764
rect 12529 29699 12587 29705
rect 12529 29665 12541 29699
rect 12575 29696 12587 29699
rect 12710 29696 12716 29708
rect 12575 29668 12716 29696
rect 12575 29665 12587 29668
rect 12529 29659 12587 29665
rect 12710 29656 12716 29668
rect 12768 29656 12774 29708
rect 16853 29699 16911 29705
rect 16853 29665 16865 29699
rect 16899 29696 16911 29699
rect 17402 29696 17408 29708
rect 16899 29668 17408 29696
rect 16899 29665 16911 29668
rect 16853 29659 16911 29665
rect 17402 29656 17408 29668
rect 17460 29656 17466 29708
rect 17494 29656 17500 29708
rect 17552 29696 17558 29708
rect 18046 29696 18052 29708
rect 17552 29668 18052 29696
rect 17552 29656 17558 29668
rect 18046 29656 18052 29668
rect 18104 29656 18110 29708
rect 18138 29656 18144 29708
rect 18196 29696 18202 29708
rect 18233 29699 18291 29705
rect 18233 29696 18245 29699
rect 18196 29668 18245 29696
rect 18196 29656 18202 29668
rect 18233 29665 18245 29668
rect 18279 29665 18291 29699
rect 19426 29696 19432 29708
rect 19387 29668 19432 29696
rect 18233 29659 18291 29665
rect 19426 29656 19432 29668
rect 19484 29656 19490 29708
rect 3191 29600 3832 29628
rect 3973 29631 4031 29637
rect 3191 29597 3203 29600
rect 3145 29591 3203 29597
rect 3973 29597 3985 29631
rect 4019 29628 4031 29631
rect 4614 29628 4620 29640
rect 4019 29600 4620 29628
rect 4019 29597 4031 29600
rect 3973 29591 4031 29597
rect 4614 29588 4620 29600
rect 4672 29588 4678 29640
rect 5810 29588 5816 29640
rect 5868 29628 5874 29640
rect 6457 29631 6515 29637
rect 6457 29628 6469 29631
rect 5868 29600 6469 29628
rect 5868 29588 5874 29600
rect 6457 29597 6469 29600
rect 6503 29597 6515 29631
rect 6457 29591 6515 29597
rect 7466 29588 7472 29640
rect 7524 29628 7530 29640
rect 7837 29631 7895 29637
rect 7837 29628 7849 29631
rect 7524 29600 7849 29628
rect 7524 29588 7530 29600
rect 7837 29597 7849 29600
rect 7883 29597 7895 29631
rect 7837 29591 7895 29597
rect 9677 29631 9735 29637
rect 9677 29597 9689 29631
rect 9723 29628 9735 29631
rect 11330 29628 11336 29640
rect 9723 29600 11336 29628
rect 9723 29597 9735 29600
rect 9677 29591 9735 29597
rect 11330 29588 11336 29600
rect 11388 29588 11394 29640
rect 11606 29628 11612 29640
rect 11519 29600 11612 29628
rect 11606 29588 11612 29600
rect 11664 29628 11670 29640
rect 12253 29631 12311 29637
rect 12253 29628 12265 29631
rect 11664 29600 12265 29628
rect 11664 29588 11670 29600
rect 12253 29597 12265 29600
rect 12299 29597 12311 29631
rect 14182 29628 14188 29640
rect 14143 29600 14188 29628
rect 12253 29591 12311 29597
rect 14182 29588 14188 29600
rect 14240 29588 14246 29640
rect 15286 29588 15292 29640
rect 15344 29628 15350 29640
rect 16577 29631 16635 29637
rect 16577 29628 16589 29631
rect 15344 29600 16589 29628
rect 15344 29588 15350 29600
rect 16577 29597 16589 29600
rect 16623 29597 16635 29631
rect 16758 29628 16764 29640
rect 16719 29600 16764 29628
rect 16577 29591 16635 29597
rect 16758 29588 16764 29600
rect 16816 29588 16822 29640
rect 16942 29588 16948 29640
rect 17000 29628 17006 29640
rect 17126 29628 17132 29640
rect 17000 29600 17045 29628
rect 17087 29600 17132 29628
rect 17000 29588 17006 29600
rect 17126 29588 17132 29600
rect 17184 29588 17190 29640
rect 18325 29631 18383 29637
rect 18325 29597 18337 29631
rect 18371 29628 18383 29631
rect 18506 29628 18512 29640
rect 18371 29600 18512 29628
rect 18371 29597 18383 29600
rect 18325 29591 18383 29597
rect 18506 29588 18512 29600
rect 18564 29588 18570 29640
rect 19720 29637 19748 29736
rect 21910 29724 21916 29736
rect 21968 29724 21974 29776
rect 20165 29699 20223 29705
rect 20165 29665 20177 29699
rect 20211 29696 20223 29699
rect 20533 29699 20591 29705
rect 20533 29696 20545 29699
rect 20211 29668 20545 29696
rect 20211 29665 20223 29668
rect 20165 29659 20223 29665
rect 20533 29665 20545 29668
rect 20579 29665 20591 29699
rect 20533 29659 20591 29665
rect 20625 29699 20683 29705
rect 20625 29665 20637 29699
rect 20671 29696 20683 29699
rect 21542 29696 21548 29708
rect 20671 29668 21548 29696
rect 20671 29665 20683 29668
rect 20625 29659 20683 29665
rect 21542 29656 21548 29668
rect 21600 29656 21606 29708
rect 22370 29696 22376 29708
rect 22331 29668 22376 29696
rect 22370 29656 22376 29668
rect 22428 29656 22434 29708
rect 19337 29631 19395 29637
rect 19337 29597 19349 29631
rect 19383 29597 19395 29631
rect 19337 29591 19395 29597
rect 19705 29631 19763 29637
rect 19705 29597 19717 29631
rect 19751 29597 19763 29631
rect 19705 29591 19763 29597
rect 6212 29563 6270 29569
rect 6212 29529 6224 29563
rect 6258 29560 6270 29563
rect 6362 29560 6368 29572
rect 6258 29532 6368 29560
rect 6258 29529 6270 29532
rect 6212 29523 6270 29529
rect 6362 29520 6368 29532
rect 6420 29520 6426 29572
rect 6546 29520 6552 29572
rect 6604 29560 6610 29572
rect 7009 29563 7067 29569
rect 7009 29560 7021 29563
rect 6604 29532 7021 29560
rect 6604 29520 6610 29532
rect 7009 29529 7021 29532
rect 7055 29529 7067 29563
rect 7009 29523 7067 29529
rect 9766 29520 9772 29572
rect 9824 29560 9830 29572
rect 9922 29563 9980 29569
rect 9922 29560 9934 29563
rect 9824 29532 9934 29560
rect 9824 29520 9830 29532
rect 9922 29529 9934 29532
rect 9968 29529 9980 29563
rect 9922 29523 9980 29529
rect 13998 29520 14004 29572
rect 14056 29560 14062 29572
rect 14430 29563 14488 29569
rect 14430 29560 14442 29563
rect 14056 29532 14442 29560
rect 14056 29520 14062 29532
rect 14430 29529 14442 29532
rect 14476 29529 14488 29563
rect 14430 29523 14488 29529
rect 16393 29563 16451 29569
rect 16393 29529 16405 29563
rect 16439 29560 16451 29563
rect 19352 29560 19380 29591
rect 16439 29532 19380 29560
rect 16439 29529 16451 29532
rect 16393 29523 16451 29529
rect 19426 29520 19432 29572
rect 19484 29560 19490 29572
rect 19720 29560 19748 29591
rect 19978 29588 19984 29640
rect 20036 29628 20042 29640
rect 20349 29631 20407 29637
rect 20349 29628 20361 29631
rect 20036 29600 20361 29628
rect 20036 29588 20042 29600
rect 20349 29597 20361 29600
rect 20395 29597 20407 29631
rect 20349 29591 20407 29597
rect 20441 29631 20499 29637
rect 20441 29597 20453 29631
rect 20487 29597 20499 29631
rect 20441 29591 20499 29597
rect 19484 29532 19748 29560
rect 19484 29520 19490 29532
rect 20254 29520 20260 29572
rect 20312 29560 20318 29572
rect 20456 29560 20484 29591
rect 21450 29588 21456 29640
rect 21508 29628 21514 29640
rect 22646 29637 22652 29640
rect 21729 29631 21787 29637
rect 21729 29628 21741 29631
rect 21508 29600 21741 29628
rect 21508 29588 21514 29600
rect 21729 29597 21741 29600
rect 21775 29597 21787 29631
rect 22640 29628 22652 29637
rect 22607 29600 22652 29628
rect 21729 29591 21787 29597
rect 22640 29591 22652 29600
rect 22646 29588 22652 29591
rect 22704 29588 22710 29640
rect 20312 29532 20484 29560
rect 21545 29563 21603 29569
rect 20312 29520 20318 29532
rect 21545 29529 21557 29563
rect 21591 29560 21603 29563
rect 21634 29560 21640 29572
rect 21591 29532 21640 29560
rect 21591 29529 21603 29532
rect 21545 29523 21603 29529
rect 21634 29520 21640 29532
rect 21692 29520 21698 29572
rect 4430 29492 4436 29504
rect 4391 29464 4436 29492
rect 4430 29452 4436 29464
rect 4488 29452 4494 29504
rect 6914 29452 6920 29504
rect 6972 29492 6978 29504
rect 7101 29495 7159 29501
rect 7101 29492 7113 29495
rect 6972 29464 7113 29492
rect 6972 29452 6978 29464
rect 7101 29461 7113 29464
rect 7147 29461 7159 29495
rect 7650 29492 7656 29504
rect 7611 29464 7656 29492
rect 7101 29455 7159 29461
rect 7650 29452 7656 29464
rect 7708 29452 7714 29504
rect 18414 29452 18420 29504
rect 18472 29492 18478 29504
rect 18693 29495 18751 29501
rect 18693 29492 18705 29495
rect 18472 29464 18705 29492
rect 18472 29452 18478 29464
rect 18693 29461 18705 29464
rect 18739 29461 18751 29495
rect 19334 29492 19340 29504
rect 19295 29464 19340 29492
rect 18693 29455 18751 29461
rect 19334 29452 19340 29464
rect 19392 29452 19398 29504
rect 20809 29495 20867 29501
rect 20809 29461 20821 29495
rect 20855 29492 20867 29495
rect 21818 29492 21824 29504
rect 20855 29464 21824 29492
rect 20855 29461 20867 29464
rect 20809 29455 20867 29461
rect 21818 29452 21824 29464
rect 21876 29452 21882 29504
rect 23753 29495 23811 29501
rect 23753 29461 23765 29495
rect 23799 29492 23811 29495
rect 29730 29492 29736 29504
rect 23799 29464 29736 29492
rect 23799 29461 23811 29464
rect 23753 29455 23811 29461
rect 29730 29452 29736 29464
rect 29788 29452 29794 29504
rect 1104 29402 30820 29424
rect 1104 29350 10880 29402
rect 10932 29350 10944 29402
rect 10996 29350 11008 29402
rect 11060 29350 11072 29402
rect 11124 29350 11136 29402
rect 11188 29350 20811 29402
rect 20863 29350 20875 29402
rect 20927 29350 20939 29402
rect 20991 29350 21003 29402
rect 21055 29350 21067 29402
rect 21119 29350 30820 29402
rect 1104 29328 30820 29350
rect 2774 29248 2780 29300
rect 2832 29288 2838 29300
rect 2832 29260 2877 29288
rect 2832 29248 2838 29260
rect 4706 29248 4712 29300
rect 4764 29288 4770 29300
rect 5169 29291 5227 29297
rect 5169 29288 5181 29291
rect 4764 29260 5181 29288
rect 4764 29248 4770 29260
rect 5169 29257 5181 29260
rect 5215 29257 5227 29291
rect 5810 29288 5816 29300
rect 5771 29260 5816 29288
rect 5169 29251 5227 29257
rect 5810 29248 5816 29260
rect 5868 29248 5874 29300
rect 7285 29291 7343 29297
rect 7285 29257 7297 29291
rect 7331 29288 7343 29291
rect 8113 29291 8171 29297
rect 8113 29288 8125 29291
rect 7331 29260 8125 29288
rect 7331 29257 7343 29260
rect 7285 29251 7343 29257
rect 8113 29257 8125 29260
rect 8159 29257 8171 29291
rect 8113 29251 8171 29257
rect 9493 29291 9551 29297
rect 9493 29257 9505 29291
rect 9539 29288 9551 29291
rect 10502 29288 10508 29300
rect 9539 29260 10508 29288
rect 9539 29257 9551 29260
rect 9493 29251 9551 29257
rect 10502 29248 10508 29260
rect 10560 29248 10566 29300
rect 10873 29291 10931 29297
rect 10873 29257 10885 29291
rect 10919 29288 10931 29291
rect 11606 29288 11612 29300
rect 10919 29260 11612 29288
rect 10919 29257 10931 29260
rect 10873 29251 10931 29257
rect 11072 29232 11100 29260
rect 11606 29248 11612 29260
rect 11664 29248 11670 29300
rect 12802 29288 12808 29300
rect 12406 29260 12808 29288
rect 4056 29223 4114 29229
rect 4056 29189 4068 29223
rect 4102 29220 4114 29223
rect 4154 29220 4160 29232
rect 4102 29192 4160 29220
rect 4102 29189 4114 29192
rect 4056 29183 4114 29189
rect 4154 29180 4160 29192
rect 4212 29180 4218 29232
rect 9585 29223 9643 29229
rect 9585 29189 9597 29223
rect 9631 29220 9643 29223
rect 9674 29220 9680 29232
rect 9631 29192 9680 29220
rect 9631 29189 9643 29192
rect 9585 29183 9643 29189
rect 9674 29180 9680 29192
rect 9732 29180 9738 29232
rect 11054 29180 11060 29232
rect 11112 29180 11118 29232
rect 1670 29152 1676 29164
rect 1631 29124 1676 29152
rect 1670 29112 1676 29124
rect 1728 29112 1734 29164
rect 2133 29155 2191 29161
rect 2133 29121 2145 29155
rect 2179 29152 2191 29155
rect 2498 29152 2504 29164
rect 2179 29124 2504 29152
rect 2179 29121 2191 29124
rect 2133 29115 2191 29121
rect 2498 29112 2504 29124
rect 2556 29112 2562 29164
rect 2958 29152 2964 29164
rect 2919 29124 2964 29152
rect 2958 29112 2964 29124
rect 3016 29112 3022 29164
rect 5626 29152 5632 29164
rect 5587 29124 5632 29152
rect 5626 29112 5632 29124
rect 5684 29112 5690 29164
rect 8297 29155 8355 29161
rect 8297 29121 8309 29155
rect 8343 29152 8355 29155
rect 8478 29152 8484 29164
rect 8343 29124 8484 29152
rect 8343 29121 8355 29124
rect 8297 29115 8355 29121
rect 8478 29112 8484 29124
rect 8536 29112 8542 29164
rect 10965 29155 11023 29161
rect 10965 29121 10977 29155
rect 11011 29152 11023 29155
rect 11790 29152 11796 29164
rect 11011 29124 11796 29152
rect 11011 29121 11023 29124
rect 10965 29115 11023 29121
rect 11790 29112 11796 29124
rect 11848 29152 11854 29164
rect 12406 29152 12434 29260
rect 12802 29248 12808 29260
rect 12860 29248 12866 29300
rect 13998 29288 14004 29300
rect 13372 29260 13768 29288
rect 13959 29260 14004 29288
rect 12621 29223 12679 29229
rect 12621 29189 12633 29223
rect 12667 29220 12679 29223
rect 12710 29220 12716 29232
rect 12667 29192 12716 29220
rect 12667 29189 12679 29192
rect 12621 29183 12679 29189
rect 12710 29180 12716 29192
rect 12768 29180 12774 29232
rect 11848 29124 12434 29152
rect 11848 29112 11854 29124
rect 3786 29084 3792 29096
rect 3747 29056 3792 29084
rect 3786 29044 3792 29056
rect 3844 29044 3850 29096
rect 7374 29084 7380 29096
rect 7335 29056 7380 29084
rect 7374 29044 7380 29056
rect 7432 29044 7438 29096
rect 7561 29087 7619 29093
rect 7561 29053 7573 29087
rect 7607 29084 7619 29087
rect 7742 29084 7748 29096
rect 7607 29056 7748 29084
rect 7607 29053 7619 29056
rect 7561 29047 7619 29053
rect 7742 29044 7748 29056
rect 7800 29084 7806 29096
rect 9677 29087 9735 29093
rect 9677 29084 9689 29087
rect 7800 29056 9689 29084
rect 7800 29044 7806 29056
rect 9677 29053 9689 29056
rect 9723 29053 9735 29087
rect 12728 29084 12756 29180
rect 13372 29161 13400 29260
rect 13630 29220 13636 29232
rect 13591 29192 13636 29220
rect 13630 29180 13636 29192
rect 13688 29180 13694 29232
rect 13740 29220 13768 29260
rect 13998 29248 14004 29260
rect 14056 29248 14062 29300
rect 16025 29291 16083 29297
rect 16025 29257 16037 29291
rect 16071 29257 16083 29291
rect 16025 29251 16083 29257
rect 16669 29291 16727 29297
rect 16669 29257 16681 29291
rect 16715 29288 16727 29291
rect 16942 29288 16948 29300
rect 16715 29260 16948 29288
rect 16715 29257 16727 29260
rect 16669 29251 16727 29257
rect 14090 29220 14096 29232
rect 13740 29192 14096 29220
rect 14090 29180 14096 29192
rect 14148 29180 14154 29232
rect 15013 29223 15071 29229
rect 15013 29189 15025 29223
rect 15059 29220 15071 29223
rect 15562 29220 15568 29232
rect 15059 29192 15568 29220
rect 15059 29189 15071 29192
rect 15013 29183 15071 29189
rect 15562 29180 15568 29192
rect 15620 29180 15626 29232
rect 16040 29220 16068 29251
rect 16942 29248 16948 29260
rect 17000 29248 17006 29300
rect 17034 29248 17040 29300
rect 17092 29288 17098 29300
rect 17129 29291 17187 29297
rect 17129 29288 17141 29291
rect 17092 29260 17141 29288
rect 17092 29248 17098 29260
rect 17129 29257 17141 29260
rect 17175 29257 17187 29291
rect 17129 29251 17187 29257
rect 18230 29248 18236 29300
rect 18288 29288 18294 29300
rect 18690 29288 18696 29300
rect 18288 29260 18696 29288
rect 18288 29248 18294 29260
rect 18690 29248 18696 29260
rect 18748 29248 18754 29300
rect 20993 29291 21051 29297
rect 20993 29257 21005 29291
rect 21039 29288 21051 29291
rect 21542 29288 21548 29300
rect 21039 29260 21548 29288
rect 21039 29257 21051 29260
rect 20993 29251 21051 29257
rect 21542 29248 21548 29260
rect 21600 29288 21606 29300
rect 21726 29288 21732 29300
rect 21600 29260 21732 29288
rect 21600 29248 21606 29260
rect 21726 29248 21732 29260
rect 21784 29248 21790 29300
rect 23201 29291 23259 29297
rect 23201 29288 23213 29291
rect 21836 29260 23213 29288
rect 19978 29220 19984 29232
rect 16040 29192 19984 29220
rect 19978 29180 19984 29192
rect 20036 29220 20042 29232
rect 20036 29192 21404 29220
rect 20036 29180 20042 29192
rect 13357 29155 13415 29161
rect 13357 29121 13369 29155
rect 13403 29121 13415 29155
rect 13357 29115 13415 29121
rect 13446 29112 13452 29164
rect 13504 29152 13510 29164
rect 13722 29152 13728 29164
rect 13504 29124 13549 29152
rect 13683 29124 13728 29152
rect 13504 29112 13510 29124
rect 13722 29112 13728 29124
rect 13780 29112 13786 29164
rect 13822 29155 13880 29161
rect 13822 29121 13834 29155
rect 13868 29152 13880 29155
rect 14642 29152 14648 29164
rect 13868 29124 14648 29152
rect 13868 29121 13880 29124
rect 13822 29115 13880 29121
rect 13837 29084 13865 29115
rect 14642 29112 14648 29124
rect 14700 29112 14706 29164
rect 15197 29155 15255 29161
rect 15197 29121 15209 29155
rect 15243 29121 15255 29155
rect 15197 29115 15255 29121
rect 15381 29155 15439 29161
rect 15381 29121 15393 29155
rect 15427 29152 15439 29155
rect 15841 29155 15899 29161
rect 15841 29152 15853 29155
rect 15427 29124 15853 29152
rect 15427 29121 15439 29124
rect 15381 29115 15439 29121
rect 15841 29121 15853 29124
rect 15887 29121 15899 29155
rect 17034 29152 17040 29164
rect 16995 29124 17040 29152
rect 15841 29115 15899 29121
rect 12728 29056 13865 29084
rect 9677 29047 9735 29053
rect 14826 29044 14832 29096
rect 14884 29084 14890 29096
rect 15212 29084 15240 29115
rect 17034 29112 17040 29124
rect 17092 29112 17098 29164
rect 18138 29112 18144 29164
rect 18196 29152 18202 29164
rect 18417 29155 18475 29161
rect 18417 29152 18429 29155
rect 18196 29124 18429 29152
rect 18196 29112 18202 29124
rect 18417 29121 18429 29124
rect 18463 29121 18475 29155
rect 18417 29115 18475 29121
rect 18509 29155 18567 29161
rect 18509 29121 18521 29155
rect 18555 29121 18567 29155
rect 18782 29152 18788 29164
rect 18743 29124 18788 29152
rect 18509 29115 18567 29121
rect 14884 29056 15240 29084
rect 17313 29087 17371 29093
rect 14884 29044 14890 29056
rect 17313 29053 17325 29087
rect 17359 29084 17371 29087
rect 18230 29084 18236 29096
rect 17359 29056 18236 29084
rect 17359 29053 17371 29056
rect 17313 29047 17371 29053
rect 18230 29044 18236 29056
rect 18288 29044 18294 29096
rect 18524 29084 18552 29115
rect 18782 29112 18788 29124
rect 18840 29112 18846 29164
rect 19426 29152 19432 29164
rect 19387 29124 19432 29152
rect 19426 29112 19432 29124
rect 19484 29112 19490 29164
rect 19705 29155 19763 29161
rect 19705 29121 19717 29155
rect 19751 29152 19763 29155
rect 19794 29152 19800 29164
rect 19751 29124 19800 29152
rect 19751 29121 19763 29124
rect 19705 29115 19763 29121
rect 19794 29112 19800 29124
rect 19852 29112 19858 29164
rect 20901 29155 20959 29161
rect 20901 29121 20913 29155
rect 20947 29152 20959 29155
rect 21266 29152 21272 29164
rect 20947 29124 21272 29152
rect 20947 29121 20959 29124
rect 20901 29115 20959 29121
rect 21266 29112 21272 29124
rect 21324 29112 21330 29164
rect 21376 29152 21404 29192
rect 21450 29180 21456 29232
rect 21508 29220 21514 29232
rect 21836 29220 21864 29260
rect 23201 29257 23213 29260
rect 23247 29257 23259 29291
rect 23201 29251 23259 29257
rect 21508 29192 21864 29220
rect 21508 29180 21514 29192
rect 29362 29152 29368 29164
rect 21376 29124 29368 29152
rect 29362 29112 29368 29124
rect 29420 29112 29426 29164
rect 20438 29084 20444 29096
rect 18524 29056 20444 29084
rect 20438 29044 20444 29056
rect 20496 29044 20502 29096
rect 21821 29087 21879 29093
rect 21821 29053 21833 29087
rect 21867 29053 21879 29087
rect 21821 29047 21879 29053
rect 1486 29016 1492 29028
rect 1447 28988 1492 29016
rect 1486 28976 1492 28988
rect 1544 28976 1550 29028
rect 2317 29019 2375 29025
rect 2317 28985 2329 29019
rect 2363 29016 2375 29019
rect 3050 29016 3056 29028
rect 2363 28988 3056 29016
rect 2363 28985 2375 28988
rect 2317 28979 2375 28985
rect 3050 28976 3056 28988
rect 3108 28976 3114 29028
rect 6822 28976 6828 29028
rect 6880 29016 6886 29028
rect 9125 29019 9183 29025
rect 9125 29016 9137 29019
rect 6880 28988 9137 29016
rect 6880 28976 6886 28988
rect 9125 28985 9137 28988
rect 9171 28985 9183 29019
rect 9125 28979 9183 28985
rect 12342 28976 12348 29028
rect 12400 29016 12406 29028
rect 12437 29019 12495 29025
rect 12437 29016 12449 29019
rect 12400 28988 12449 29016
rect 12400 28976 12406 28988
rect 12437 28985 12449 28988
rect 12483 28985 12495 29019
rect 12437 28979 12495 28985
rect 14182 28976 14188 29028
rect 14240 29016 14246 29028
rect 15654 29016 15660 29028
rect 14240 28988 15660 29016
rect 14240 28976 14246 28988
rect 15654 28976 15660 28988
rect 15712 29016 15718 29028
rect 21836 29016 21864 29047
rect 22002 29044 22008 29096
rect 22060 29084 22066 29096
rect 22097 29087 22155 29093
rect 22097 29084 22109 29087
rect 22060 29056 22109 29084
rect 22060 29044 22066 29056
rect 22097 29053 22109 29056
rect 22143 29053 22155 29087
rect 22097 29047 22155 29053
rect 15712 28988 21864 29016
rect 15712 28976 15718 28988
rect 6917 28951 6975 28957
rect 6917 28917 6929 28951
rect 6963 28948 6975 28951
rect 7006 28948 7012 28960
rect 6963 28920 7012 28948
rect 6963 28917 6975 28920
rect 6917 28911 6975 28917
rect 7006 28908 7012 28920
rect 7064 28908 7070 28960
rect 18233 28951 18291 28957
rect 18233 28917 18245 28951
rect 18279 28948 18291 28951
rect 18322 28948 18328 28960
rect 18279 28920 18328 28948
rect 18279 28917 18291 28920
rect 18233 28911 18291 28917
rect 18322 28908 18328 28920
rect 18380 28908 18386 28960
rect 18693 28951 18751 28957
rect 18693 28917 18705 28951
rect 18739 28948 18751 28951
rect 19610 28948 19616 28960
rect 18739 28920 19616 28948
rect 18739 28917 18751 28920
rect 18693 28911 18751 28917
rect 19610 28908 19616 28920
rect 19668 28908 19674 28960
rect 1104 28858 30820 28880
rect 1104 28806 5915 28858
rect 5967 28806 5979 28858
rect 6031 28806 6043 28858
rect 6095 28806 6107 28858
rect 6159 28806 6171 28858
rect 6223 28806 15846 28858
rect 15898 28806 15910 28858
rect 15962 28806 15974 28858
rect 16026 28806 16038 28858
rect 16090 28806 16102 28858
rect 16154 28806 25776 28858
rect 25828 28806 25840 28858
rect 25892 28806 25904 28858
rect 25956 28806 25968 28858
rect 26020 28806 26032 28858
rect 26084 28806 30820 28858
rect 1104 28784 30820 28806
rect 1670 28704 1676 28756
rect 1728 28744 1734 28756
rect 2409 28747 2467 28753
rect 2409 28744 2421 28747
rect 1728 28716 2421 28744
rect 1728 28704 1734 28716
rect 2409 28713 2421 28716
rect 2455 28713 2467 28747
rect 3786 28744 3792 28756
rect 3747 28716 3792 28744
rect 2409 28707 2467 28713
rect 3786 28704 3792 28716
rect 3844 28704 3850 28756
rect 4801 28747 4859 28753
rect 4801 28713 4813 28747
rect 4847 28744 4859 28747
rect 5626 28744 5632 28756
rect 4847 28716 5632 28744
rect 4847 28713 4859 28716
rect 4801 28707 4859 28713
rect 5626 28704 5632 28716
rect 5684 28704 5690 28756
rect 6181 28747 6239 28753
rect 6181 28713 6193 28747
rect 6227 28744 6239 28747
rect 7374 28744 7380 28756
rect 6227 28716 7380 28744
rect 6227 28713 6239 28716
rect 6181 28707 6239 28713
rect 7374 28704 7380 28716
rect 7432 28704 7438 28756
rect 11422 28704 11428 28756
rect 11480 28744 11486 28756
rect 11885 28747 11943 28753
rect 11885 28744 11897 28747
rect 11480 28716 11897 28744
rect 11480 28704 11486 28716
rect 11885 28713 11897 28716
rect 11931 28744 11943 28747
rect 12250 28744 12256 28756
rect 11931 28716 12256 28744
rect 11931 28713 11943 28716
rect 11885 28707 11943 28713
rect 12250 28704 12256 28716
rect 12308 28704 12314 28756
rect 14185 28747 14243 28753
rect 14185 28713 14197 28747
rect 14231 28744 14243 28747
rect 15286 28744 15292 28756
rect 14231 28716 15292 28744
rect 14231 28713 14243 28716
rect 14185 28707 14243 28713
rect 15286 28704 15292 28716
rect 15344 28704 15350 28756
rect 15654 28744 15660 28756
rect 15615 28716 15660 28744
rect 15654 28704 15660 28716
rect 15712 28704 15718 28756
rect 16853 28747 16911 28753
rect 16853 28713 16865 28747
rect 16899 28744 16911 28747
rect 17218 28744 17224 28756
rect 16899 28716 17224 28744
rect 16899 28713 16911 28716
rect 16853 28707 16911 28713
rect 17218 28704 17224 28716
rect 17276 28704 17282 28756
rect 21174 28744 21180 28756
rect 20456 28716 21180 28744
rect 6641 28679 6699 28685
rect 6641 28645 6653 28679
rect 6687 28645 6699 28679
rect 6641 28639 6699 28645
rect 3145 28611 3203 28617
rect 3145 28608 3157 28611
rect 1688 28580 3157 28608
rect 1688 28549 1716 28580
rect 3145 28577 3157 28580
rect 3191 28577 3203 28611
rect 6656 28608 6684 28639
rect 12894 28636 12900 28688
rect 12952 28676 12958 28688
rect 18141 28679 18199 28685
rect 12952 28648 13584 28676
rect 12952 28636 12958 28648
rect 3145 28571 3203 28577
rect 3252 28580 6684 28608
rect 7285 28611 7343 28617
rect 3252 28549 3280 28580
rect 7285 28577 7297 28611
rect 7331 28608 7343 28611
rect 7742 28608 7748 28620
rect 7331 28580 7748 28608
rect 7331 28577 7343 28580
rect 7285 28571 7343 28577
rect 7742 28568 7748 28580
rect 7800 28608 7806 28620
rect 9493 28611 9551 28617
rect 9493 28608 9505 28611
rect 7800 28580 9505 28608
rect 7800 28568 7806 28580
rect 9493 28577 9505 28580
rect 9539 28577 9551 28611
rect 9493 28571 9551 28577
rect 11241 28611 11299 28617
rect 11241 28577 11253 28611
rect 11287 28608 11299 28611
rect 11882 28608 11888 28620
rect 11287 28580 11888 28608
rect 11287 28577 11299 28580
rect 11241 28571 11299 28577
rect 11882 28568 11888 28580
rect 11940 28568 11946 28620
rect 12526 28568 12532 28620
rect 12584 28608 12590 28620
rect 13446 28608 13452 28620
rect 12584 28580 13452 28608
rect 12584 28568 12590 28580
rect 1673 28543 1731 28549
rect 1673 28509 1685 28543
rect 1719 28509 1731 28543
rect 1673 28503 1731 28509
rect 2409 28543 2467 28549
rect 2409 28509 2421 28543
rect 2455 28509 2467 28543
rect 2409 28503 2467 28509
rect 2593 28543 2651 28549
rect 2593 28509 2605 28543
rect 2639 28540 2651 28543
rect 3053 28543 3111 28549
rect 3053 28540 3065 28543
rect 2639 28512 3065 28540
rect 2639 28509 2651 28512
rect 2593 28503 2651 28509
rect 3053 28509 3065 28512
rect 3099 28509 3111 28543
rect 3053 28503 3111 28509
rect 3237 28543 3295 28549
rect 3237 28509 3249 28543
rect 3283 28509 3295 28543
rect 3237 28503 3295 28509
rect 3973 28543 4031 28549
rect 3973 28509 3985 28543
rect 4019 28540 4031 28543
rect 4430 28540 4436 28552
rect 4019 28512 4436 28540
rect 4019 28509 4031 28512
rect 3973 28503 4031 28509
rect 2424 28472 2452 28503
rect 3068 28472 3096 28503
rect 4430 28500 4436 28512
rect 4488 28500 4494 28552
rect 4614 28540 4620 28552
rect 4575 28512 4620 28540
rect 4614 28500 4620 28512
rect 4672 28500 4678 28552
rect 5997 28543 6055 28549
rect 5997 28509 6009 28543
rect 6043 28540 6055 28543
rect 6454 28540 6460 28552
rect 6043 28512 6460 28540
rect 6043 28509 6055 28512
rect 5997 28503 6055 28509
rect 6454 28500 6460 28512
rect 6512 28500 6518 28552
rect 7009 28543 7067 28549
rect 7009 28509 7021 28543
rect 7055 28540 7067 28543
rect 7650 28540 7656 28552
rect 7055 28512 7656 28540
rect 7055 28509 7067 28512
rect 7009 28503 7067 28509
rect 7650 28500 7656 28512
rect 7708 28500 7714 28552
rect 8389 28543 8447 28549
rect 8389 28509 8401 28543
rect 8435 28509 8447 28543
rect 9306 28540 9312 28552
rect 9267 28512 9312 28540
rect 8389 28503 8447 28509
rect 3142 28472 3148 28484
rect 2424 28444 2774 28472
rect 3068 28444 3148 28472
rect 1486 28404 1492 28416
rect 1447 28376 1492 28404
rect 1486 28364 1492 28376
rect 1544 28364 1550 28416
rect 2746 28404 2774 28444
rect 3142 28432 3148 28444
rect 3200 28432 3206 28484
rect 8404 28472 8432 28503
rect 9306 28500 9312 28512
rect 9364 28500 9370 28552
rect 10318 28540 10324 28552
rect 10279 28512 10324 28540
rect 10318 28500 10324 28512
rect 10376 28540 10382 28552
rect 10778 28540 10784 28552
rect 10376 28512 10784 28540
rect 10376 28500 10382 28512
rect 10778 28500 10784 28512
rect 10836 28500 10842 28552
rect 11054 28540 11060 28552
rect 11015 28512 11060 28540
rect 11054 28500 11060 28512
rect 11112 28500 11118 28552
rect 11790 28540 11796 28552
rect 11751 28512 11796 28540
rect 11790 28500 11796 28512
rect 11848 28500 11854 28552
rect 11974 28500 11980 28552
rect 12032 28540 12038 28552
rect 13188 28549 13216 28580
rect 13446 28568 13452 28580
rect 13504 28568 13510 28620
rect 13556 28552 13584 28648
rect 18141 28645 18153 28679
rect 18187 28676 18199 28679
rect 19426 28676 19432 28688
rect 18187 28648 19432 28676
rect 18187 28645 18199 28648
rect 18141 28639 18199 28645
rect 19426 28636 19432 28648
rect 19484 28636 19490 28688
rect 14090 28568 14096 28620
rect 14148 28608 14154 28620
rect 15013 28611 15071 28617
rect 15013 28608 15025 28611
rect 14148 28580 15025 28608
rect 14148 28568 14154 28580
rect 15013 28577 15025 28580
rect 15059 28608 15071 28611
rect 17862 28608 17868 28620
rect 15059 28580 17868 28608
rect 15059 28577 15071 28580
rect 15013 28571 15071 28577
rect 17862 28568 17868 28580
rect 17920 28608 17926 28620
rect 17920 28580 20208 28608
rect 17920 28568 17926 28580
rect 12759 28543 12817 28549
rect 12759 28540 12771 28543
rect 12032 28512 12771 28540
rect 12032 28500 12038 28512
rect 12759 28509 12771 28512
rect 12805 28509 12817 28543
rect 12759 28503 12817 28509
rect 13172 28543 13230 28549
rect 13172 28509 13184 28543
rect 13218 28509 13230 28543
rect 13172 28503 13230 28509
rect 13265 28543 13323 28549
rect 13265 28509 13277 28543
rect 13311 28540 13323 28543
rect 13538 28540 13544 28552
rect 13311 28512 13544 28540
rect 13311 28509 13323 28512
rect 13265 28503 13323 28509
rect 13538 28500 13544 28512
rect 13596 28500 13602 28552
rect 14277 28543 14335 28549
rect 14277 28509 14289 28543
rect 14323 28540 14335 28543
rect 15194 28540 15200 28552
rect 14323 28512 15200 28540
rect 14323 28509 14335 28512
rect 14277 28503 14335 28509
rect 15194 28500 15200 28512
rect 15252 28500 15258 28552
rect 15470 28500 15476 28552
rect 15528 28540 15534 28552
rect 15565 28543 15623 28549
rect 15565 28540 15577 28543
rect 15528 28512 15577 28540
rect 15528 28500 15534 28512
rect 15565 28509 15577 28512
rect 15611 28509 15623 28543
rect 16942 28540 16948 28552
rect 16903 28512 16948 28540
rect 15565 28503 15623 28509
rect 16942 28500 16948 28512
rect 17000 28500 17006 28552
rect 17494 28500 17500 28552
rect 17552 28540 17558 28552
rect 18046 28540 18052 28552
rect 17552 28512 18052 28540
rect 17552 28500 17558 28512
rect 18046 28500 18052 28512
rect 18104 28500 18110 28552
rect 18233 28543 18291 28549
rect 18233 28509 18245 28543
rect 18279 28509 18291 28543
rect 18233 28503 18291 28509
rect 9490 28472 9496 28484
rect 8404 28444 9496 28472
rect 9490 28432 9496 28444
rect 9548 28432 9554 28484
rect 12158 28432 12164 28484
rect 12216 28472 12222 28484
rect 12897 28475 12955 28481
rect 12897 28472 12909 28475
rect 12216 28444 12909 28472
rect 12216 28432 12222 28444
rect 12897 28441 12909 28444
rect 12943 28441 12955 28475
rect 12897 28435 12955 28441
rect 12989 28475 13047 28481
rect 12989 28441 13001 28475
rect 13035 28472 13047 28475
rect 14090 28472 14096 28484
rect 13035 28444 14096 28472
rect 13035 28441 13047 28444
rect 12989 28435 13047 28441
rect 14090 28432 14096 28444
rect 14148 28432 14154 28484
rect 14826 28472 14832 28484
rect 14787 28444 14832 28472
rect 14826 28432 14832 28444
rect 14884 28432 14890 28484
rect 18248 28472 18276 28503
rect 18322 28500 18328 28552
rect 18380 28540 18386 28552
rect 18509 28543 18567 28549
rect 18380 28512 18425 28540
rect 18380 28500 18386 28512
rect 18509 28509 18521 28543
rect 18555 28540 18567 28543
rect 18598 28540 18604 28552
rect 18555 28512 18604 28540
rect 18555 28509 18567 28512
rect 18509 28503 18567 28509
rect 18598 28500 18604 28512
rect 18656 28500 18662 28552
rect 20180 28549 20208 28580
rect 20456 28549 20484 28716
rect 21174 28704 21180 28716
rect 21232 28744 21238 28756
rect 21542 28744 21548 28756
rect 21232 28716 21548 28744
rect 21232 28704 21238 28716
rect 21542 28704 21548 28716
rect 21600 28704 21606 28756
rect 22465 28747 22523 28753
rect 22465 28713 22477 28747
rect 22511 28744 22523 28747
rect 22922 28744 22928 28756
rect 22511 28716 22928 28744
rect 22511 28713 22523 28716
rect 22465 28707 22523 28713
rect 22922 28704 22928 28716
rect 22980 28704 22986 28756
rect 22002 28676 22008 28688
rect 20732 28648 22008 28676
rect 20732 28617 20760 28648
rect 22002 28636 22008 28648
rect 22060 28636 22066 28688
rect 20717 28611 20775 28617
rect 20717 28577 20729 28611
rect 20763 28577 20775 28611
rect 21818 28608 21824 28620
rect 21779 28580 21824 28608
rect 20717 28571 20775 28577
rect 21818 28568 21824 28580
rect 21876 28568 21882 28620
rect 21910 28568 21916 28620
rect 21968 28608 21974 28620
rect 22306 28611 22364 28617
rect 22306 28608 22318 28611
rect 21968 28580 22318 28608
rect 21968 28568 21974 28580
rect 22306 28577 22318 28580
rect 22352 28577 22364 28611
rect 22306 28571 22364 28577
rect 20165 28543 20223 28549
rect 20165 28509 20177 28543
rect 20211 28509 20223 28543
rect 20165 28503 20223 28509
rect 20257 28543 20315 28549
rect 20257 28509 20269 28543
rect 20303 28540 20315 28543
rect 20441 28543 20499 28549
rect 20303 28512 20392 28540
rect 20303 28509 20315 28512
rect 20257 28503 20315 28509
rect 18248 28444 18552 28472
rect 18524 28416 18552 28444
rect 7006 28404 7012 28416
rect 2746 28376 7012 28404
rect 7006 28364 7012 28376
rect 7064 28364 7070 28416
rect 7098 28364 7104 28416
rect 7156 28404 7162 28416
rect 8297 28407 8355 28413
rect 7156 28376 7201 28404
rect 7156 28364 7162 28376
rect 8297 28373 8309 28407
rect 8343 28404 8355 28407
rect 8662 28404 8668 28416
rect 8343 28376 8668 28404
rect 8343 28373 8355 28376
rect 8297 28367 8355 28373
rect 8662 28364 8668 28376
rect 8720 28364 8726 28416
rect 8938 28404 8944 28416
rect 8899 28376 8944 28404
rect 8938 28364 8944 28376
rect 8996 28364 9002 28416
rect 9398 28404 9404 28416
rect 9359 28376 9404 28404
rect 9398 28364 9404 28376
rect 9456 28364 9462 28416
rect 10226 28404 10232 28416
rect 10187 28376 10232 28404
rect 10226 28364 10232 28376
rect 10284 28364 10290 28416
rect 12621 28407 12679 28413
rect 12621 28373 12633 28407
rect 12667 28404 12679 28407
rect 13170 28404 13176 28416
rect 12667 28376 13176 28404
rect 12667 28373 12679 28376
rect 12621 28367 12679 28373
rect 13170 28364 13176 28376
rect 13228 28364 13234 28416
rect 17865 28407 17923 28413
rect 17865 28373 17877 28407
rect 17911 28404 17923 28407
rect 18230 28404 18236 28416
rect 17911 28376 18236 28404
rect 17911 28373 17923 28376
rect 17865 28367 17923 28373
rect 18230 28364 18236 28376
rect 18288 28364 18294 28416
rect 18506 28364 18512 28416
rect 18564 28364 18570 28416
rect 20364 28404 20392 28512
rect 20441 28509 20453 28543
rect 20487 28509 20499 28543
rect 20622 28540 20628 28552
rect 20583 28512 20628 28540
rect 20441 28503 20499 28509
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 22097 28543 22155 28549
rect 22097 28509 22109 28543
rect 22143 28540 22155 28543
rect 22554 28540 22560 28552
rect 22143 28512 22560 28540
rect 22143 28509 22155 28512
rect 22097 28503 22155 28509
rect 22554 28500 22560 28512
rect 22612 28500 22618 28552
rect 29822 28540 29828 28552
rect 29783 28512 29828 28540
rect 29822 28500 29828 28512
rect 29880 28500 29886 28552
rect 20533 28475 20591 28481
rect 20533 28441 20545 28475
rect 20579 28472 20591 28475
rect 20714 28472 20720 28484
rect 20579 28444 20720 28472
rect 20579 28441 20591 28444
rect 20533 28435 20591 28441
rect 20714 28432 20720 28444
rect 20772 28472 20778 28484
rect 21910 28472 21916 28484
rect 20772 28444 21916 28472
rect 20772 28432 20778 28444
rect 21910 28432 21916 28444
rect 21968 28432 21974 28484
rect 21818 28404 21824 28416
rect 20364 28376 21824 28404
rect 21818 28364 21824 28376
rect 21876 28364 21882 28416
rect 22186 28364 22192 28416
rect 22244 28404 22250 28416
rect 30006 28404 30012 28416
rect 22244 28376 22289 28404
rect 29967 28376 30012 28404
rect 22244 28364 22250 28376
rect 30006 28364 30012 28376
rect 30064 28364 30070 28416
rect 1104 28314 30820 28336
rect 1104 28262 10880 28314
rect 10932 28262 10944 28314
rect 10996 28262 11008 28314
rect 11060 28262 11072 28314
rect 11124 28262 11136 28314
rect 11188 28262 20811 28314
rect 20863 28262 20875 28314
rect 20927 28262 20939 28314
rect 20991 28262 21003 28314
rect 21055 28262 21067 28314
rect 21119 28262 30820 28314
rect 1104 28240 30820 28262
rect 2038 28160 2044 28212
rect 2096 28200 2102 28212
rect 2133 28203 2191 28209
rect 2133 28200 2145 28203
rect 2096 28172 2145 28200
rect 2096 28160 2102 28172
rect 2133 28169 2145 28172
rect 2179 28169 2191 28203
rect 2133 28163 2191 28169
rect 6733 28203 6791 28209
rect 6733 28169 6745 28203
rect 6779 28200 6791 28203
rect 7098 28200 7104 28212
rect 6779 28172 7104 28200
rect 6779 28169 6791 28172
rect 6733 28163 6791 28169
rect 7098 28160 7104 28172
rect 7156 28160 7162 28212
rect 8481 28203 8539 28209
rect 8481 28169 8493 28203
rect 8527 28200 8539 28203
rect 9398 28200 9404 28212
rect 8527 28172 9404 28200
rect 8527 28169 8539 28172
rect 8481 28163 8539 28169
rect 9398 28160 9404 28172
rect 9456 28160 9462 28212
rect 10042 28200 10048 28212
rect 9508 28172 10048 28200
rect 3697 28135 3755 28141
rect 3697 28132 3709 28135
rect 1688 28104 3709 28132
rect 1688 28073 1716 28104
rect 3697 28101 3709 28104
rect 3743 28101 3755 28135
rect 8938 28132 8944 28144
rect 3697 28095 3755 28101
rect 3804 28104 8944 28132
rect 1673 28067 1731 28073
rect 1673 28033 1685 28067
rect 1719 28033 1731 28067
rect 1673 28027 1731 28033
rect 2317 28067 2375 28073
rect 2317 28033 2329 28067
rect 2363 28064 2375 28067
rect 2406 28064 2412 28076
rect 2363 28036 2412 28064
rect 2363 28033 2375 28036
rect 2317 28027 2375 28033
rect 2406 28024 2412 28036
rect 2464 28024 2470 28076
rect 2869 28067 2927 28073
rect 2869 28033 2881 28067
rect 2915 28064 2927 28067
rect 3326 28064 3332 28076
rect 2915 28036 3332 28064
rect 2915 28033 2927 28036
rect 2869 28027 2927 28033
rect 3326 28024 3332 28036
rect 3384 28024 3390 28076
rect 3804 28073 3832 28104
rect 8938 28092 8944 28104
rect 8996 28092 9002 28144
rect 9508 28132 9536 28172
rect 10042 28160 10048 28172
rect 10100 28160 10106 28212
rect 14090 28160 14096 28212
rect 14148 28200 14154 28212
rect 14277 28203 14335 28209
rect 14277 28200 14289 28203
rect 14148 28172 14289 28200
rect 14148 28160 14154 28172
rect 14277 28169 14289 28172
rect 14323 28169 14335 28203
rect 14277 28163 14335 28169
rect 17037 28203 17095 28209
rect 17037 28169 17049 28203
rect 17083 28200 17095 28203
rect 17126 28200 17132 28212
rect 17083 28172 17132 28200
rect 17083 28169 17095 28172
rect 17037 28163 17095 28169
rect 17126 28160 17132 28172
rect 17184 28160 17190 28212
rect 18598 28200 18604 28212
rect 18559 28172 18604 28200
rect 18598 28160 18604 28172
rect 18656 28160 18662 28212
rect 18782 28160 18788 28212
rect 18840 28200 18846 28212
rect 19061 28203 19119 28209
rect 19061 28200 19073 28203
rect 18840 28172 19073 28200
rect 18840 28160 18846 28172
rect 19061 28169 19073 28172
rect 19107 28169 19119 28203
rect 19061 28163 19119 28169
rect 20622 28160 20628 28212
rect 20680 28200 20686 28212
rect 20901 28203 20959 28209
rect 20901 28200 20913 28203
rect 20680 28172 20913 28200
rect 20680 28160 20686 28172
rect 20901 28169 20913 28172
rect 20947 28169 20959 28203
rect 21910 28200 21916 28212
rect 21871 28172 21916 28200
rect 20901 28163 20959 28169
rect 21910 28160 21916 28172
rect 21968 28160 21974 28212
rect 22186 28160 22192 28212
rect 22244 28200 22250 28212
rect 29454 28200 29460 28212
rect 22244 28172 29460 28200
rect 22244 28160 22250 28172
rect 29454 28160 29460 28172
rect 29512 28160 29518 28212
rect 29822 28160 29828 28212
rect 29880 28200 29886 28212
rect 30009 28203 30067 28209
rect 30009 28200 30021 28203
rect 29880 28172 30021 28200
rect 29880 28160 29886 28172
rect 30009 28169 30021 28172
rect 30055 28169 30067 28203
rect 30009 28163 30067 28169
rect 11330 28132 11336 28144
rect 9048 28104 9536 28132
rect 9600 28104 11336 28132
rect 3605 28067 3663 28073
rect 3605 28033 3617 28067
rect 3651 28033 3663 28067
rect 3605 28027 3663 28033
rect 3789 28067 3847 28073
rect 3789 28033 3801 28067
rect 3835 28033 3847 28067
rect 3789 28027 3847 28033
rect 6549 28067 6607 28073
rect 6549 28033 6561 28067
rect 6595 28064 6607 28067
rect 7653 28067 7711 28073
rect 6595 28036 7236 28064
rect 6595 28033 6607 28036
rect 6549 28027 6607 28033
rect 3142 27956 3148 28008
rect 3200 27996 3206 28008
rect 3620 27996 3648 28027
rect 7208 28005 7236 28036
rect 7653 28033 7665 28067
rect 7699 28033 7711 28067
rect 8662 28064 8668 28076
rect 8623 28036 8668 28064
rect 7653 28027 7711 28033
rect 3200 27968 3648 27996
rect 7193 27999 7251 28005
rect 3200 27956 3206 27968
rect 7193 27965 7205 27999
rect 7239 27965 7251 27999
rect 7193 27959 7251 27965
rect 7668 27928 7696 28027
rect 8662 28024 8668 28036
rect 8720 28024 8726 28076
rect 8754 28024 8760 28076
rect 8812 28064 8818 28076
rect 9048 28073 9076 28104
rect 9600 28073 9628 28104
rect 11330 28092 11336 28104
rect 11388 28092 11394 28144
rect 12345 28135 12403 28141
rect 12345 28101 12357 28135
rect 12391 28132 12403 28135
rect 12526 28132 12532 28144
rect 12391 28104 12532 28132
rect 12391 28101 12403 28104
rect 12345 28095 12403 28101
rect 12526 28092 12532 28104
rect 12584 28092 12590 28144
rect 14182 28132 14188 28144
rect 12912 28104 14188 28132
rect 9858 28073 9864 28076
rect 9033 28067 9091 28073
rect 8812 28036 8857 28064
rect 8812 28024 8818 28036
rect 9033 28033 9045 28067
rect 9079 28033 9091 28067
rect 9033 28027 9091 28033
rect 9585 28067 9643 28073
rect 9585 28033 9597 28067
rect 9631 28033 9643 28067
rect 9585 28027 9643 28033
rect 9852 28027 9864 28073
rect 9916 28064 9922 28076
rect 9916 28036 9952 28064
rect 9858 28024 9864 28027
rect 9916 28024 9922 28036
rect 10318 28024 10324 28076
rect 10376 28064 10382 28076
rect 11609 28067 11667 28073
rect 11609 28064 11621 28067
rect 10376 28036 11621 28064
rect 10376 28024 10382 28036
rect 11609 28033 11621 28036
rect 11655 28033 11667 28067
rect 11609 28027 11667 28033
rect 11698 28024 11704 28076
rect 11756 28064 11762 28076
rect 11756 28036 11801 28064
rect 11756 28024 11762 28036
rect 12618 28024 12624 28076
rect 12676 28064 12682 28076
rect 12912 28073 12940 28104
rect 14182 28092 14188 28104
rect 14240 28092 14246 28144
rect 14737 28135 14795 28141
rect 14737 28132 14749 28135
rect 14292 28104 14749 28132
rect 13170 28073 13176 28076
rect 12897 28067 12955 28073
rect 12897 28064 12909 28067
rect 12676 28036 12909 28064
rect 12676 28024 12682 28036
rect 12897 28033 12909 28036
rect 12943 28033 12955 28067
rect 13164 28064 13176 28073
rect 13131 28036 13176 28064
rect 12897 28027 12955 28033
rect 13164 28027 13176 28036
rect 13170 28024 13176 28027
rect 13228 28024 13234 28076
rect 13538 28024 13544 28076
rect 13596 28064 13602 28076
rect 14292 28064 14320 28104
rect 14737 28101 14749 28104
rect 14783 28101 14795 28135
rect 18874 28132 18880 28144
rect 14737 28095 14795 28101
rect 18156 28104 18880 28132
rect 13596 28036 14320 28064
rect 13596 28024 13602 28036
rect 14458 28024 14464 28076
rect 14516 28064 14522 28076
rect 14826 28064 14832 28076
rect 14516 28036 14832 28064
rect 14516 28024 14522 28036
rect 14826 28024 14832 28036
rect 14884 28064 14890 28076
rect 14921 28067 14979 28073
rect 14921 28064 14933 28067
rect 14884 28036 14933 28064
rect 14884 28024 14890 28036
rect 14921 28033 14933 28036
rect 14967 28033 14979 28067
rect 14921 28027 14979 28033
rect 15473 28067 15531 28073
rect 15473 28033 15485 28067
rect 15519 28033 15531 28067
rect 16666 28064 16672 28076
rect 16627 28036 16672 28064
rect 15473 28027 15531 28033
rect 11790 27956 11796 28008
rect 11848 27996 11854 28008
rect 12526 27996 12532 28008
rect 11848 27968 12532 27996
rect 11848 27956 11854 27968
rect 12526 27956 12532 27968
rect 12584 27956 12590 28008
rect 14366 27956 14372 28008
rect 14424 27996 14430 28008
rect 15488 27996 15516 28027
rect 16666 28024 16672 28036
rect 16724 28024 16730 28076
rect 16850 28064 16856 28076
rect 16811 28036 16856 28064
rect 16850 28024 16856 28036
rect 16908 28024 16914 28076
rect 17862 28064 17868 28076
rect 17823 28036 17868 28064
rect 17862 28024 17868 28036
rect 17920 28024 17926 28076
rect 18046 28064 18052 28076
rect 18007 28036 18052 28064
rect 18046 28024 18052 28036
rect 18104 28024 18110 28076
rect 18156 28073 18184 28104
rect 18874 28092 18880 28104
rect 18932 28132 18938 28144
rect 18932 28104 20300 28132
rect 18932 28092 18938 28104
rect 18141 28067 18199 28073
rect 18141 28033 18153 28067
rect 18187 28033 18199 28067
rect 18414 28064 18420 28076
rect 18375 28036 18420 28064
rect 18141 28027 18199 28033
rect 18414 28024 18420 28036
rect 18472 28024 18478 28076
rect 18506 28024 18512 28076
rect 18564 28064 18570 28076
rect 20272 28073 20300 28104
rect 19429 28067 19487 28073
rect 19429 28064 19441 28067
rect 18564 28036 19441 28064
rect 18564 28024 18570 28036
rect 19429 28033 19441 28036
rect 19475 28033 19487 28067
rect 19429 28027 19487 28033
rect 20257 28067 20315 28073
rect 20257 28033 20269 28067
rect 20303 28033 20315 28067
rect 20438 28064 20444 28076
rect 20399 28036 20444 28064
rect 20257 28027 20315 28033
rect 20438 28024 20444 28036
rect 20496 28024 20502 28076
rect 20622 28024 20628 28076
rect 20680 28064 20686 28076
rect 20717 28067 20775 28073
rect 20717 28064 20729 28067
rect 20680 28036 20729 28064
rect 20680 28024 20686 28036
rect 20717 28033 20729 28036
rect 20763 28064 20775 28067
rect 21450 28064 21456 28076
rect 20763 28036 21456 28064
rect 20763 28033 20775 28036
rect 20717 28027 20775 28033
rect 21450 28024 21456 28036
rect 21508 28024 21514 28076
rect 21818 28064 21824 28076
rect 21779 28036 21824 28064
rect 21818 28024 21824 28036
rect 21876 28024 21882 28076
rect 29638 28024 29644 28076
rect 29696 28064 29702 28076
rect 29917 28067 29975 28073
rect 29917 28064 29929 28067
rect 29696 28036 29929 28064
rect 29696 28024 29702 28036
rect 29917 28033 29929 28036
rect 29963 28033 29975 28067
rect 30098 28064 30104 28076
rect 30059 28036 30104 28064
rect 29917 28027 29975 28033
rect 30098 28024 30104 28036
rect 30156 28024 30162 28076
rect 14424 27968 15516 27996
rect 14424 27956 14430 27968
rect 17954 27956 17960 28008
rect 18012 27996 18018 28008
rect 18233 27999 18291 28005
rect 18233 27996 18245 27999
rect 18012 27968 18245 27996
rect 18012 27956 18018 27968
rect 18233 27965 18245 27968
rect 18279 27965 18291 27999
rect 19518 27996 19524 28008
rect 19479 27968 19524 27996
rect 18233 27959 18291 27965
rect 19518 27956 19524 27968
rect 19576 27956 19582 28008
rect 19613 27999 19671 28005
rect 19613 27965 19625 27999
rect 19659 27965 19671 27999
rect 19613 27959 19671 27965
rect 7208 27900 7696 27928
rect 7208 27872 7236 27900
rect 12066 27888 12072 27940
rect 12124 27928 12130 27940
rect 12161 27931 12219 27937
rect 12161 27928 12173 27931
rect 12124 27900 12173 27928
rect 12124 27888 12130 27900
rect 12161 27897 12173 27900
rect 12207 27897 12219 27931
rect 12161 27891 12219 27897
rect 18598 27888 18604 27940
rect 18656 27928 18662 27940
rect 19628 27928 19656 27959
rect 20530 27928 20536 27940
rect 18656 27900 19656 27928
rect 20491 27900 20536 27928
rect 18656 27888 18662 27900
rect 20530 27888 20536 27900
rect 20588 27888 20594 27940
rect 20625 27931 20683 27937
rect 20625 27897 20637 27931
rect 20671 27928 20683 27931
rect 21174 27928 21180 27940
rect 20671 27900 21180 27928
rect 20671 27897 20683 27900
rect 20625 27891 20683 27897
rect 21174 27888 21180 27900
rect 21232 27888 21238 27940
rect 1486 27860 1492 27872
rect 1447 27832 1492 27860
rect 1486 27820 1492 27832
rect 1544 27820 1550 27872
rect 2774 27820 2780 27872
rect 2832 27860 2838 27872
rect 3053 27863 3111 27869
rect 3053 27860 3065 27863
rect 2832 27832 3065 27860
rect 2832 27820 2838 27832
rect 3053 27829 3065 27832
rect 3099 27860 3111 27863
rect 3602 27860 3608 27872
rect 3099 27832 3608 27860
rect 3099 27829 3111 27832
rect 3053 27823 3111 27829
rect 3602 27820 3608 27832
rect 3660 27820 3666 27872
rect 7190 27820 7196 27872
rect 7248 27820 7254 27872
rect 7561 27863 7619 27869
rect 7561 27829 7573 27863
rect 7607 27860 7619 27863
rect 7926 27860 7932 27872
rect 7607 27832 7932 27860
rect 7607 27829 7619 27832
rect 7561 27823 7619 27829
rect 7926 27820 7932 27832
rect 7984 27860 7990 27872
rect 8941 27863 8999 27869
rect 8941 27860 8953 27863
rect 7984 27832 8953 27860
rect 7984 27820 7990 27832
rect 8941 27829 8953 27832
rect 8987 27829 8999 27863
rect 8941 27823 8999 27829
rect 9490 27820 9496 27872
rect 9548 27860 9554 27872
rect 10965 27863 11023 27869
rect 10965 27860 10977 27863
rect 9548 27832 10977 27860
rect 9548 27820 9554 27832
rect 10965 27829 10977 27832
rect 11011 27829 11023 27863
rect 15562 27860 15568 27872
rect 15523 27832 15568 27860
rect 10965 27823 11023 27829
rect 15562 27820 15568 27832
rect 15620 27820 15626 27872
rect 16666 27820 16672 27872
rect 16724 27860 16730 27872
rect 19426 27860 19432 27872
rect 16724 27832 19432 27860
rect 16724 27820 16730 27832
rect 19426 27820 19432 27832
rect 19484 27820 19490 27872
rect 1104 27770 30820 27792
rect 1104 27718 5915 27770
rect 5967 27718 5979 27770
rect 6031 27718 6043 27770
rect 6095 27718 6107 27770
rect 6159 27718 6171 27770
rect 6223 27718 15846 27770
rect 15898 27718 15910 27770
rect 15962 27718 15974 27770
rect 16026 27718 16038 27770
rect 16090 27718 16102 27770
rect 16154 27718 25776 27770
rect 25828 27718 25840 27770
rect 25892 27718 25904 27770
rect 25956 27718 25968 27770
rect 26020 27718 26032 27770
rect 26084 27718 30820 27770
rect 1104 27696 30820 27718
rect 3326 27616 3332 27668
rect 3384 27656 3390 27668
rect 3384 27628 4292 27656
rect 3384 27616 3390 27628
rect 4264 27597 4292 27628
rect 9122 27616 9128 27668
rect 9180 27656 9186 27668
rect 9180 27628 9441 27656
rect 9180 27616 9186 27628
rect 4249 27591 4307 27597
rect 4249 27557 4261 27591
rect 4295 27557 4307 27591
rect 5810 27588 5816 27600
rect 5771 27560 5816 27588
rect 4249 27551 4307 27557
rect 5810 27548 5816 27560
rect 5868 27548 5874 27600
rect 6641 27591 6699 27597
rect 6641 27557 6653 27591
rect 6687 27588 6699 27591
rect 7466 27588 7472 27600
rect 6687 27560 7472 27588
rect 6687 27557 6699 27560
rect 6641 27551 6699 27557
rect 7466 27548 7472 27560
rect 7524 27548 7530 27600
rect 8754 27588 8760 27600
rect 7576 27560 8760 27588
rect 5736 27492 6592 27520
rect 5736 27464 5764 27492
rect 3053 27455 3111 27461
rect 3053 27421 3065 27455
rect 3099 27452 3111 27455
rect 3142 27452 3148 27464
rect 3099 27424 3148 27452
rect 3099 27421 3111 27424
rect 3053 27415 3111 27421
rect 3142 27412 3148 27424
rect 3200 27412 3206 27464
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27421 3295 27455
rect 3237 27415 3295 27421
rect 5629 27455 5687 27461
rect 5629 27421 5641 27455
rect 5675 27421 5687 27455
rect 5629 27415 5687 27421
rect 1670 27276 1676 27328
rect 1728 27316 1734 27328
rect 3145 27319 3203 27325
rect 3145 27316 3157 27319
rect 1728 27288 3157 27316
rect 1728 27276 1734 27288
rect 3145 27285 3157 27288
rect 3191 27285 3203 27319
rect 3252 27316 3280 27415
rect 4433 27387 4491 27393
rect 4433 27353 4445 27387
rect 4479 27384 4491 27387
rect 4614 27384 4620 27396
rect 4479 27356 4620 27384
rect 4479 27353 4491 27356
rect 4433 27347 4491 27353
rect 4614 27344 4620 27356
rect 4672 27344 4678 27396
rect 5644 27384 5672 27415
rect 5718 27412 5724 27464
rect 5776 27452 5782 27464
rect 5905 27455 5963 27461
rect 5776 27424 5821 27452
rect 5776 27412 5782 27424
rect 5905 27421 5917 27455
rect 5951 27452 5963 27455
rect 6362 27452 6368 27464
rect 5951 27424 6368 27452
rect 5951 27421 5963 27424
rect 5905 27415 5963 27421
rect 6362 27412 6368 27424
rect 6420 27412 6426 27464
rect 6564 27461 6592 27492
rect 6549 27455 6607 27461
rect 6549 27421 6561 27455
rect 6595 27421 6607 27455
rect 7374 27452 7380 27464
rect 7335 27424 7380 27452
rect 6549 27415 6607 27421
rect 7374 27412 7380 27424
rect 7432 27412 7438 27464
rect 7469 27455 7527 27461
rect 7469 27421 7481 27455
rect 7515 27452 7527 27455
rect 7576 27452 7604 27560
rect 8754 27548 8760 27560
rect 8812 27588 8818 27600
rect 9030 27588 9036 27600
rect 8812 27560 9036 27588
rect 8812 27548 8818 27560
rect 9030 27548 9036 27560
rect 9088 27548 9094 27600
rect 9306 27588 9312 27600
rect 9232 27560 9312 27588
rect 7653 27523 7711 27529
rect 7653 27489 7665 27523
rect 7699 27520 7711 27523
rect 8202 27520 8208 27532
rect 7699 27492 8208 27520
rect 7699 27489 7711 27492
rect 7653 27483 7711 27489
rect 8202 27480 8208 27492
rect 8260 27480 8266 27532
rect 9232 27529 9260 27560
rect 9306 27548 9312 27560
rect 9364 27548 9370 27600
rect 9217 27523 9275 27529
rect 9217 27489 9229 27523
rect 9263 27489 9275 27523
rect 9413 27520 9441 27628
rect 9490 27616 9496 27668
rect 9548 27656 9554 27668
rect 10778 27656 10784 27668
rect 9548 27628 10784 27656
rect 9548 27616 9554 27628
rect 10778 27616 10784 27628
rect 10836 27616 10842 27668
rect 11974 27656 11980 27668
rect 11348 27628 11980 27656
rect 9674 27588 9680 27600
rect 9635 27560 9680 27588
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 10689 27591 10747 27597
rect 10689 27557 10701 27591
rect 10735 27588 10747 27591
rect 11348 27588 11376 27628
rect 11974 27616 11980 27628
rect 12032 27616 12038 27668
rect 16850 27616 16856 27668
rect 16908 27656 16914 27668
rect 16945 27659 17003 27665
rect 16945 27656 16957 27659
rect 16908 27628 16957 27656
rect 16908 27616 16914 27628
rect 16945 27625 16957 27628
rect 16991 27625 17003 27659
rect 16945 27619 17003 27625
rect 17957 27659 18015 27665
rect 17957 27625 17969 27659
rect 18003 27656 18015 27659
rect 18046 27656 18052 27668
rect 18003 27628 18052 27656
rect 18003 27625 18015 27628
rect 17957 27619 18015 27625
rect 18046 27616 18052 27628
rect 18104 27616 18110 27668
rect 19429 27659 19487 27665
rect 19429 27625 19441 27659
rect 19475 27656 19487 27659
rect 19610 27656 19616 27668
rect 19475 27628 19616 27656
rect 19475 27625 19487 27628
rect 19429 27619 19487 27625
rect 19610 27616 19616 27628
rect 19668 27616 19674 27668
rect 19794 27616 19800 27668
rect 19852 27656 19858 27668
rect 19978 27656 19984 27668
rect 19852 27628 19984 27656
rect 19852 27616 19858 27628
rect 19978 27616 19984 27628
rect 20036 27616 20042 27668
rect 20441 27659 20499 27665
rect 20441 27625 20453 27659
rect 20487 27656 20499 27659
rect 20530 27656 20536 27668
rect 20487 27628 20536 27656
rect 20487 27625 20499 27628
rect 20441 27619 20499 27625
rect 20530 27616 20536 27628
rect 20588 27616 20594 27668
rect 10735 27560 11376 27588
rect 15473 27591 15531 27597
rect 10735 27557 10747 27560
rect 10689 27551 10747 27557
rect 15473 27557 15485 27591
rect 15519 27588 15531 27591
rect 19518 27588 19524 27600
rect 15519 27560 19524 27588
rect 15519 27557 15531 27560
rect 15473 27551 15531 27557
rect 19518 27548 19524 27560
rect 19576 27548 19582 27600
rect 20070 27588 20076 27600
rect 20031 27560 20076 27588
rect 20070 27548 20076 27560
rect 20128 27548 20134 27600
rect 10318 27520 10324 27532
rect 9413 27492 10324 27520
rect 9217 27483 9275 27489
rect 10318 27480 10324 27492
rect 10376 27480 10382 27532
rect 10597 27523 10655 27529
rect 10597 27489 10609 27523
rect 10643 27489 10655 27523
rect 11330 27520 11336 27532
rect 11291 27492 11336 27520
rect 10597 27483 10655 27489
rect 7515 27424 7604 27452
rect 7745 27455 7803 27461
rect 7515 27421 7527 27424
rect 7469 27415 7527 27421
rect 7745 27421 7757 27455
rect 7791 27452 7803 27455
rect 8297 27455 8355 27461
rect 8297 27452 8309 27455
rect 7791 27424 8309 27452
rect 7791 27421 7803 27424
rect 7745 27415 7803 27421
rect 8297 27421 8309 27424
rect 8343 27421 8355 27455
rect 8297 27415 8355 27421
rect 8386 27412 8392 27464
rect 8444 27452 8450 27464
rect 8444 27424 8489 27452
rect 8444 27412 8450 27424
rect 8846 27412 8852 27464
rect 8904 27452 8910 27464
rect 8941 27455 8999 27461
rect 8941 27452 8953 27455
rect 8904 27424 8953 27452
rect 8904 27412 8910 27424
rect 8941 27421 8953 27424
rect 8987 27421 8999 27455
rect 9122 27452 9128 27464
rect 9180 27461 9186 27464
rect 9087 27424 9128 27452
rect 8941 27415 8999 27421
rect 9122 27412 9128 27424
rect 9180 27415 9187 27461
rect 9309 27455 9367 27461
rect 9309 27442 9321 27455
rect 9355 27442 9367 27455
rect 9493 27455 9551 27461
rect 9180 27412 9186 27415
rect 5994 27384 6000 27396
rect 5644 27356 6000 27384
rect 5994 27344 6000 27356
rect 6052 27344 6058 27396
rect 6089 27387 6147 27393
rect 9306 27390 9312 27442
rect 9364 27390 9370 27442
rect 9493 27421 9505 27455
rect 9539 27452 9551 27455
rect 10226 27452 10232 27464
rect 9539 27424 10232 27452
rect 9539 27421 9551 27424
rect 9493 27415 9551 27421
rect 10226 27412 10232 27424
rect 10284 27412 10290 27464
rect 6089 27353 6101 27387
rect 6135 27384 6147 27387
rect 10502 27384 10508 27396
rect 6135 27356 9261 27384
rect 6135 27353 6147 27356
rect 6089 27347 6147 27353
rect 6822 27316 6828 27328
rect 3252 27288 6828 27316
rect 3145 27279 3203 27285
rect 6822 27276 6828 27288
rect 6880 27276 6886 27328
rect 7098 27276 7104 27328
rect 7156 27316 7162 27328
rect 7193 27319 7251 27325
rect 7193 27316 7205 27319
rect 7156 27288 7205 27316
rect 7156 27276 7162 27288
rect 7193 27285 7205 27288
rect 7239 27285 7251 27319
rect 9233 27316 9261 27356
rect 9508 27356 10508 27384
rect 9508 27316 9536 27356
rect 10502 27344 10508 27356
rect 10560 27344 10566 27396
rect 9233 27288 9536 27316
rect 7193 27279 7251 27285
rect 9582 27276 9588 27328
rect 9640 27316 9646 27328
rect 10612 27316 10640 27483
rect 11330 27480 11336 27492
rect 11388 27480 11394 27532
rect 14090 27480 14096 27532
rect 14148 27520 14154 27532
rect 14829 27523 14887 27529
rect 14148 27492 14688 27520
rect 14148 27480 14154 27492
rect 10778 27452 10784 27464
rect 10739 27424 10784 27452
rect 10778 27412 10784 27424
rect 10836 27412 10842 27464
rect 10870 27412 10876 27464
rect 10928 27452 10934 27464
rect 14366 27452 14372 27464
rect 10928 27424 10973 27452
rect 14327 27424 14372 27452
rect 10928 27412 10934 27424
rect 14366 27412 14372 27424
rect 14424 27412 14430 27464
rect 14660 27461 14688 27492
rect 14829 27489 14841 27523
rect 14875 27520 14887 27523
rect 15381 27523 15439 27529
rect 15381 27520 15393 27523
rect 14875 27492 15393 27520
rect 14875 27489 14887 27492
rect 14829 27483 14887 27489
rect 15381 27489 15393 27492
rect 15427 27489 15439 27523
rect 15381 27483 15439 27489
rect 15565 27523 15623 27529
rect 15565 27489 15577 27523
rect 15611 27489 15623 27523
rect 15565 27483 15623 27489
rect 16393 27523 16451 27529
rect 16393 27489 16405 27523
rect 16439 27520 16451 27523
rect 17494 27520 17500 27532
rect 16439 27492 17500 27520
rect 16439 27489 16451 27492
rect 16393 27483 16451 27489
rect 14461 27455 14519 27461
rect 14461 27421 14473 27455
rect 14507 27421 14519 27455
rect 14461 27415 14519 27421
rect 14645 27455 14703 27461
rect 14645 27421 14657 27455
rect 14691 27421 14703 27455
rect 15286 27452 15292 27464
rect 15247 27424 15292 27452
rect 14645 27415 14703 27421
rect 11422 27344 11428 27396
rect 11480 27384 11486 27396
rect 11578 27387 11636 27393
rect 11578 27384 11590 27387
rect 11480 27356 11590 27384
rect 11480 27344 11486 27356
rect 11578 27353 11590 27356
rect 11624 27353 11636 27387
rect 14476 27384 14504 27415
rect 15286 27412 15292 27424
rect 15344 27412 15350 27464
rect 14734 27384 14740 27396
rect 11578 27347 11636 27353
rect 12728 27356 14740 27384
rect 9640 27288 10640 27316
rect 9640 27276 9646 27288
rect 10778 27276 10784 27328
rect 10836 27316 10842 27328
rect 12728 27325 12756 27356
rect 14734 27344 14740 27356
rect 14792 27344 14798 27396
rect 15580 27384 15608 27483
rect 17494 27480 17500 27492
rect 17552 27520 17558 27532
rect 18509 27523 18567 27529
rect 18509 27520 18521 27523
rect 17552 27492 18521 27520
rect 17552 27480 17558 27492
rect 18509 27489 18521 27492
rect 18555 27520 18567 27523
rect 18598 27520 18604 27532
rect 18555 27492 18604 27520
rect 18555 27489 18567 27492
rect 18509 27483 18567 27489
rect 18598 27480 18604 27492
rect 18656 27480 18662 27532
rect 19794 27520 19800 27532
rect 18708 27492 19800 27520
rect 16577 27455 16635 27461
rect 16577 27421 16589 27455
rect 16623 27452 16635 27455
rect 17218 27452 17224 27464
rect 16623 27424 17224 27452
rect 16623 27421 16635 27424
rect 16577 27415 16635 27421
rect 17218 27412 17224 27424
rect 17276 27412 17282 27464
rect 18325 27455 18383 27461
rect 18325 27421 18337 27455
rect 18371 27452 18383 27455
rect 18414 27452 18420 27464
rect 18371 27424 18420 27452
rect 18371 27421 18383 27424
rect 18325 27415 18383 27421
rect 18414 27412 18420 27424
rect 18472 27412 18478 27464
rect 17586 27384 17592 27396
rect 15580 27356 17592 27384
rect 17586 27344 17592 27356
rect 17644 27384 17650 27396
rect 18708 27384 18736 27492
rect 19794 27480 19800 27492
rect 19852 27520 19858 27532
rect 19981 27523 20039 27529
rect 19981 27520 19993 27523
rect 19852 27492 19993 27520
rect 19852 27480 19858 27492
rect 19981 27489 19993 27492
rect 20027 27489 20039 27523
rect 19981 27483 20039 27489
rect 19337 27455 19395 27461
rect 19337 27421 19349 27455
rect 19383 27452 19395 27455
rect 19426 27452 19432 27464
rect 19383 27424 19432 27452
rect 19383 27421 19395 27424
rect 19337 27415 19395 27421
rect 19426 27412 19432 27424
rect 19484 27412 19490 27464
rect 20254 27452 20260 27464
rect 20215 27424 20260 27452
rect 20254 27412 20260 27424
rect 20312 27412 20318 27464
rect 21358 27452 21364 27464
rect 21319 27424 21364 27452
rect 21358 27412 21364 27424
rect 21416 27412 21422 27464
rect 21634 27452 21640 27464
rect 21595 27424 21640 27452
rect 21634 27412 21640 27424
rect 21692 27412 21698 27464
rect 29825 27455 29883 27461
rect 29825 27421 29837 27455
rect 29871 27452 29883 27455
rect 29914 27452 29920 27464
rect 29871 27424 29920 27452
rect 29871 27421 29883 27424
rect 29825 27415 29883 27421
rect 29914 27412 29920 27424
rect 29972 27412 29978 27464
rect 17644 27356 18736 27384
rect 17644 27344 17650 27356
rect 12713 27319 12771 27325
rect 12713 27316 12725 27319
rect 10836 27288 12725 27316
rect 10836 27276 10842 27288
rect 12713 27285 12725 27288
rect 12759 27285 12771 27319
rect 16482 27316 16488 27328
rect 16443 27288 16488 27316
rect 12713 27279 12771 27285
rect 16482 27276 16488 27288
rect 16540 27276 16546 27328
rect 18417 27319 18475 27325
rect 18417 27285 18429 27319
rect 18463 27316 18475 27319
rect 18598 27316 18604 27328
rect 18463 27288 18604 27316
rect 18463 27285 18475 27288
rect 18417 27279 18475 27285
rect 18598 27276 18604 27288
rect 18656 27276 18662 27328
rect 30006 27316 30012 27328
rect 29967 27288 30012 27316
rect 30006 27276 30012 27288
rect 30064 27276 30070 27328
rect 1104 27226 30820 27248
rect 1104 27174 10880 27226
rect 10932 27174 10944 27226
rect 10996 27174 11008 27226
rect 11060 27174 11072 27226
rect 11124 27174 11136 27226
rect 11188 27174 20811 27226
rect 20863 27174 20875 27226
rect 20927 27174 20939 27226
rect 20991 27174 21003 27226
rect 21055 27174 21067 27226
rect 21119 27174 30820 27226
rect 1104 27152 30820 27174
rect 6457 27115 6515 27121
rect 6457 27081 6469 27115
rect 6503 27112 6515 27115
rect 6546 27112 6552 27124
rect 6503 27084 6552 27112
rect 6503 27081 6515 27084
rect 6457 27075 6515 27081
rect 6546 27072 6552 27084
rect 6604 27072 6610 27124
rect 8570 27072 8576 27124
rect 8628 27112 8634 27124
rect 10318 27112 10324 27124
rect 8628 27084 10324 27112
rect 8628 27072 8634 27084
rect 10318 27072 10324 27084
rect 10376 27072 10382 27124
rect 10965 27115 11023 27121
rect 10965 27081 10977 27115
rect 11011 27112 11023 27115
rect 11422 27112 11428 27124
rect 11011 27084 11428 27112
rect 11011 27081 11023 27084
rect 10965 27075 11023 27081
rect 11422 27072 11428 27084
rect 11480 27072 11486 27124
rect 11790 27072 11796 27124
rect 11848 27112 11854 27124
rect 13722 27112 13728 27124
rect 11848 27084 13728 27112
rect 11848 27072 11854 27084
rect 13722 27072 13728 27084
rect 13780 27072 13786 27124
rect 16853 27115 16911 27121
rect 16853 27081 16865 27115
rect 16899 27112 16911 27115
rect 17034 27112 17040 27124
rect 16899 27084 17040 27112
rect 16899 27081 16911 27084
rect 16853 27075 16911 27081
rect 17034 27072 17040 27084
rect 17092 27072 17098 27124
rect 17218 27112 17224 27124
rect 17179 27084 17224 27112
rect 17218 27072 17224 27084
rect 17276 27072 17282 27124
rect 18138 27112 18144 27124
rect 18099 27084 18144 27112
rect 18138 27072 18144 27084
rect 18196 27072 18202 27124
rect 19521 27115 19579 27121
rect 19521 27081 19533 27115
rect 19567 27112 19579 27115
rect 21358 27112 21364 27124
rect 19567 27084 21364 27112
rect 19567 27081 19579 27084
rect 19521 27075 19579 27081
rect 21358 27072 21364 27084
rect 21416 27072 21422 27124
rect 21818 27072 21824 27124
rect 21876 27072 21882 27124
rect 29914 27112 29920 27124
rect 29875 27084 29920 27112
rect 29914 27072 29920 27084
rect 29972 27072 29978 27124
rect 7466 27004 7472 27056
rect 7524 27004 7530 27056
rect 8018 27004 8024 27056
rect 8076 27044 8082 27056
rect 8389 27047 8447 27053
rect 8389 27044 8401 27047
rect 8076 27016 8401 27044
rect 8076 27004 8082 27016
rect 8389 27013 8401 27016
rect 8435 27044 8447 27047
rect 11977 27047 12035 27053
rect 11977 27044 11989 27047
rect 8435 27016 11989 27044
rect 8435 27013 8447 27016
rect 8389 27007 8447 27013
rect 11977 27013 11989 27016
rect 12023 27013 12035 27047
rect 11977 27007 12035 27013
rect 12161 27047 12219 27053
rect 12161 27013 12173 27047
rect 12207 27044 12219 27047
rect 13354 27044 13360 27056
rect 12207 27016 13360 27044
rect 12207 27013 12219 27016
rect 12161 27007 12219 27013
rect 13354 27004 13360 27016
rect 13412 27004 13418 27056
rect 15562 27044 15568 27056
rect 15028 27016 15568 27044
rect 1670 26976 1676 26988
rect 1631 26948 1676 26976
rect 1670 26936 1676 26948
rect 1728 26936 1734 26988
rect 5534 26976 5540 26988
rect 5592 26985 5598 26988
rect 5504 26948 5540 26976
rect 5534 26936 5540 26948
rect 5592 26939 5604 26985
rect 6549 26979 6607 26985
rect 6549 26945 6561 26979
rect 6595 26976 6607 26979
rect 7006 26976 7012 26988
rect 6595 26948 7012 26976
rect 6595 26945 6607 26948
rect 6549 26939 6607 26945
rect 5592 26936 5598 26939
rect 7006 26936 7012 26948
rect 7064 26936 7070 26988
rect 7098 26936 7104 26988
rect 7156 26976 7162 26988
rect 7285 26979 7343 26985
rect 7156 26948 7201 26976
rect 7156 26936 7162 26948
rect 7285 26945 7297 26979
rect 7331 26976 7343 26979
rect 7484 26976 7512 27004
rect 7331 26948 7512 26976
rect 7653 26979 7711 26985
rect 7331 26945 7343 26948
rect 7285 26939 7343 26945
rect 7653 26945 7665 26979
rect 7699 26976 7711 26979
rect 8294 26976 8300 26988
rect 7699 26948 8300 26976
rect 7699 26945 7711 26948
rect 7653 26939 7711 26945
rect 8294 26936 8300 26948
rect 8352 26936 8358 26988
rect 8573 26979 8631 26985
rect 8573 26945 8585 26979
rect 8619 26945 8631 26979
rect 8573 26939 8631 26945
rect 5813 26911 5871 26917
rect 5813 26877 5825 26911
rect 5859 26908 5871 26911
rect 6822 26908 6828 26920
rect 5859 26880 6828 26908
rect 5859 26877 5871 26880
rect 5813 26871 5871 26877
rect 6822 26868 6828 26880
rect 6880 26868 6886 26920
rect 7377 26911 7435 26917
rect 7377 26877 7389 26911
rect 7423 26877 7435 26911
rect 7377 26871 7435 26877
rect 7469 26911 7527 26917
rect 7469 26877 7481 26911
rect 7515 26908 7527 26911
rect 7926 26908 7932 26920
rect 7515 26880 7932 26908
rect 7515 26877 7527 26880
rect 7469 26871 7527 26877
rect 1486 26840 1492 26852
rect 1447 26812 1492 26840
rect 1486 26800 1492 26812
rect 1544 26800 1550 26852
rect 7392 26840 7420 26871
rect 7926 26868 7932 26880
rect 7984 26868 7990 26920
rect 8386 26840 8392 26852
rect 7392 26812 8392 26840
rect 8386 26800 8392 26812
rect 8444 26800 8450 26852
rect 8588 26840 8616 26939
rect 8938 26936 8944 26988
rect 8996 26976 9002 26988
rect 9125 26979 9183 26985
rect 9125 26976 9137 26979
rect 8996 26948 9137 26976
rect 8996 26936 9002 26948
rect 9125 26945 9137 26948
rect 9171 26945 9183 26979
rect 9125 26939 9183 26945
rect 9214 26936 9220 26988
rect 9272 26976 9278 26988
rect 9398 26976 9404 26988
rect 9272 26948 9317 26976
rect 9359 26948 9404 26976
rect 9272 26936 9278 26948
rect 9398 26936 9404 26948
rect 9456 26936 9462 26988
rect 9493 26979 9551 26985
rect 9493 26945 9505 26979
rect 9539 26945 9551 26979
rect 9493 26939 9551 26945
rect 8662 26868 8668 26920
rect 8720 26908 8726 26920
rect 9508 26908 9536 26939
rect 9582 26936 9588 26988
rect 9640 26985 9646 26988
rect 9640 26976 9648 26985
rect 10226 26976 10232 26988
rect 9640 26948 9685 26976
rect 10187 26948 10232 26976
rect 9640 26939 9648 26948
rect 9640 26936 9646 26939
rect 10226 26936 10232 26948
rect 10284 26936 10290 26988
rect 10318 26936 10324 26988
rect 10376 26976 10382 26988
rect 10413 26979 10471 26985
rect 10413 26976 10425 26979
rect 10376 26948 10425 26976
rect 10376 26936 10382 26948
rect 10413 26945 10425 26948
rect 10459 26945 10471 26979
rect 10413 26939 10471 26945
rect 10502 26936 10508 26988
rect 10560 26976 10566 26988
rect 10778 26976 10784 26988
rect 10560 26948 10605 26976
rect 10739 26948 10784 26976
rect 10560 26936 10566 26948
rect 10778 26936 10784 26948
rect 10836 26936 10842 26988
rect 12618 26976 12624 26988
rect 12579 26948 12624 26976
rect 12618 26936 12624 26948
rect 12676 26936 12682 26988
rect 12710 26936 12716 26988
rect 12768 26976 12774 26988
rect 12877 26979 12935 26985
rect 12877 26976 12889 26979
rect 12768 26948 12889 26976
rect 12768 26936 12774 26948
rect 12877 26945 12889 26948
rect 12923 26945 12935 26979
rect 12877 26939 12935 26945
rect 13998 26936 14004 26988
rect 14056 26976 14062 26988
rect 14366 26976 14372 26988
rect 14056 26948 14372 26976
rect 14056 26936 14062 26948
rect 14366 26936 14372 26948
rect 14424 26976 14430 26988
rect 14645 26979 14703 26985
rect 14645 26976 14657 26979
rect 14424 26948 14657 26976
rect 14424 26936 14430 26948
rect 14645 26945 14657 26948
rect 14691 26945 14703 26979
rect 14918 26976 14924 26988
rect 14879 26948 14924 26976
rect 14645 26939 14703 26945
rect 14918 26936 14924 26948
rect 14976 26936 14982 26988
rect 15028 26985 15056 27016
rect 15562 27004 15568 27016
rect 15620 27004 15626 27056
rect 21082 27004 21088 27056
rect 21140 27044 21146 27056
rect 21836 27044 21864 27072
rect 21140 27016 21864 27044
rect 21140 27004 21146 27016
rect 15013 26979 15071 26985
rect 15013 26945 15025 26979
rect 15059 26945 15071 26979
rect 15013 26939 15071 26945
rect 15197 26979 15255 26985
rect 15197 26945 15209 26979
rect 15243 26976 15255 26979
rect 15657 26979 15715 26985
rect 15657 26976 15669 26979
rect 15243 26948 15669 26976
rect 15243 26945 15255 26948
rect 15197 26939 15255 26945
rect 15657 26945 15669 26948
rect 15703 26945 15715 26979
rect 15657 26939 15715 26945
rect 15841 26979 15899 26985
rect 15841 26945 15853 26979
rect 15887 26945 15899 26979
rect 15841 26939 15899 26945
rect 8720 26880 9536 26908
rect 10597 26911 10655 26917
rect 8720 26868 8726 26880
rect 10597 26877 10609 26911
rect 10643 26908 10655 26911
rect 12342 26908 12348 26920
rect 10643 26880 12348 26908
rect 10643 26877 10655 26880
rect 10597 26871 10655 26877
rect 12342 26868 12348 26880
rect 12400 26868 12406 26920
rect 14734 26908 14740 26920
rect 14695 26880 14740 26908
rect 14734 26868 14740 26880
rect 14792 26868 14798 26920
rect 15102 26868 15108 26920
rect 15160 26908 15166 26920
rect 15856 26908 15884 26939
rect 18322 26936 18328 26988
rect 18380 26976 18386 26988
rect 18509 26979 18567 26985
rect 18509 26976 18521 26979
rect 18380 26948 18521 26976
rect 18380 26936 18386 26948
rect 18509 26945 18521 26948
rect 18555 26945 18567 26979
rect 18509 26939 18567 26945
rect 19705 26979 19763 26985
rect 19705 26945 19717 26979
rect 19751 26945 19763 26979
rect 19705 26939 19763 26945
rect 19889 26979 19947 26985
rect 19889 26945 19901 26979
rect 19935 26976 19947 26979
rect 20254 26976 20260 26988
rect 19935 26948 20260 26976
rect 19935 26945 19947 26948
rect 19889 26939 19947 26945
rect 17310 26908 17316 26920
rect 15160 26880 15884 26908
rect 17271 26880 17316 26908
rect 15160 26868 15166 26880
rect 17310 26868 17316 26880
rect 17368 26868 17374 26920
rect 17494 26908 17500 26920
rect 17455 26880 17500 26908
rect 17494 26868 17500 26880
rect 17552 26868 17558 26920
rect 18598 26908 18604 26920
rect 18559 26880 18604 26908
rect 18598 26868 18604 26880
rect 18656 26868 18662 26920
rect 18690 26868 18696 26920
rect 18748 26908 18754 26920
rect 19720 26908 19748 26939
rect 20254 26936 20260 26948
rect 20312 26976 20318 26988
rect 20809 26979 20867 26985
rect 20809 26976 20821 26979
rect 20312 26948 20821 26976
rect 20312 26936 20318 26948
rect 20809 26945 20821 26948
rect 20855 26976 20867 26979
rect 21910 26976 21916 26988
rect 20855 26948 21916 26976
rect 20855 26945 20867 26948
rect 20809 26939 20867 26945
rect 21910 26936 21916 26948
rect 21968 26936 21974 26988
rect 22094 26985 22100 26988
rect 22088 26939 22100 26985
rect 22152 26976 22158 26988
rect 30098 26976 30104 26988
rect 22152 26948 22188 26976
rect 30059 26948 30104 26976
rect 22094 26936 22100 26939
rect 22152 26936 22158 26948
rect 30098 26936 30104 26948
rect 30156 26936 30162 26988
rect 20622 26908 20628 26920
rect 18748 26880 18793 26908
rect 19720 26880 20628 26908
rect 18748 26868 18754 26880
rect 20622 26868 20628 26880
rect 20680 26868 20686 26920
rect 20717 26911 20775 26917
rect 20717 26877 20729 26911
rect 20763 26877 20775 26911
rect 20717 26871 20775 26877
rect 12434 26840 12440 26852
rect 8588 26812 12440 26840
rect 12434 26800 12440 26812
rect 12492 26800 12498 26852
rect 20254 26800 20260 26852
rect 20312 26840 20318 26852
rect 20530 26840 20536 26852
rect 20312 26812 20536 26840
rect 20312 26800 20318 26812
rect 20530 26800 20536 26812
rect 20588 26840 20594 26852
rect 20732 26840 20760 26871
rect 21726 26868 21732 26920
rect 21784 26908 21790 26920
rect 21821 26911 21879 26917
rect 21821 26908 21833 26911
rect 21784 26880 21833 26908
rect 21784 26868 21790 26880
rect 21821 26877 21833 26880
rect 21867 26877 21879 26911
rect 21821 26871 21879 26877
rect 20588 26812 20760 26840
rect 20588 26800 20594 26812
rect 4433 26775 4491 26781
rect 4433 26741 4445 26775
rect 4479 26772 4491 26775
rect 4890 26772 4896 26784
rect 4479 26744 4896 26772
rect 4479 26741 4491 26744
rect 4433 26735 4491 26741
rect 4890 26732 4896 26744
rect 4948 26732 4954 26784
rect 7466 26732 7472 26784
rect 7524 26772 7530 26784
rect 7837 26775 7895 26781
rect 7837 26772 7849 26775
rect 7524 26744 7849 26772
rect 7524 26732 7530 26744
rect 7837 26741 7849 26744
rect 7883 26741 7895 26775
rect 8404 26772 8432 26800
rect 9306 26772 9312 26784
rect 8404 26744 9312 26772
rect 7837 26735 7895 26741
rect 9306 26732 9312 26744
rect 9364 26732 9370 26784
rect 9769 26775 9827 26781
rect 9769 26741 9781 26775
rect 9815 26772 9827 26775
rect 9858 26772 9864 26784
rect 9815 26744 9864 26772
rect 9815 26741 9827 26744
rect 9769 26735 9827 26741
rect 9858 26732 9864 26744
rect 9916 26732 9922 26784
rect 13998 26772 14004 26784
rect 13959 26744 14004 26772
rect 13998 26732 14004 26744
rect 14056 26732 14062 26784
rect 16025 26775 16083 26781
rect 16025 26741 16037 26775
rect 16071 26772 16083 26775
rect 16298 26772 16304 26784
rect 16071 26744 16304 26772
rect 16071 26741 16083 26744
rect 16025 26735 16083 26741
rect 16298 26732 16304 26744
rect 16356 26732 16362 26784
rect 19426 26732 19432 26784
rect 19484 26772 19490 26784
rect 20441 26775 20499 26781
rect 20441 26772 20453 26775
rect 19484 26744 20453 26772
rect 19484 26732 19490 26744
rect 20441 26741 20453 26744
rect 20487 26741 20499 26775
rect 20441 26735 20499 26741
rect 20809 26775 20867 26781
rect 20809 26741 20821 26775
rect 20855 26772 20867 26775
rect 21174 26772 21180 26784
rect 20855 26744 21180 26772
rect 20855 26741 20867 26744
rect 20809 26735 20867 26741
rect 21174 26732 21180 26744
rect 21232 26772 21238 26784
rect 21542 26772 21548 26784
rect 21232 26744 21548 26772
rect 21232 26732 21238 26744
rect 21542 26732 21548 26744
rect 21600 26732 21606 26784
rect 22002 26732 22008 26784
rect 22060 26772 22066 26784
rect 23201 26775 23259 26781
rect 23201 26772 23213 26775
rect 22060 26744 23213 26772
rect 22060 26732 22066 26744
rect 23201 26741 23213 26744
rect 23247 26741 23259 26775
rect 23201 26735 23259 26741
rect 1104 26682 30820 26704
rect 1104 26630 5915 26682
rect 5967 26630 5979 26682
rect 6031 26630 6043 26682
rect 6095 26630 6107 26682
rect 6159 26630 6171 26682
rect 6223 26630 15846 26682
rect 15898 26630 15910 26682
rect 15962 26630 15974 26682
rect 16026 26630 16038 26682
rect 16090 26630 16102 26682
rect 16154 26630 25776 26682
rect 25828 26630 25840 26682
rect 25892 26630 25904 26682
rect 25956 26630 25968 26682
rect 26020 26630 26032 26682
rect 26084 26630 30820 26682
rect 1104 26608 30820 26630
rect 7009 26571 7067 26577
rect 7009 26568 7021 26571
rect 3252 26540 7021 26568
rect 1673 26367 1731 26373
rect 1673 26333 1685 26367
rect 1719 26364 1731 26367
rect 2866 26364 2872 26376
rect 1719 26336 2872 26364
rect 1719 26333 1731 26336
rect 1673 26327 1731 26333
rect 2866 26324 2872 26336
rect 2924 26324 2930 26376
rect 3053 26367 3111 26373
rect 3053 26333 3065 26367
rect 3099 26364 3111 26367
rect 3142 26364 3148 26376
rect 3099 26336 3148 26364
rect 3099 26333 3111 26336
rect 3053 26327 3111 26333
rect 3142 26324 3148 26336
rect 3200 26324 3206 26376
rect 3252 26373 3280 26540
rect 7009 26537 7021 26540
rect 7055 26537 7067 26571
rect 8294 26568 8300 26580
rect 8255 26540 8300 26568
rect 7009 26531 7067 26537
rect 8294 26528 8300 26540
rect 8352 26528 8358 26580
rect 9677 26571 9735 26577
rect 9677 26537 9689 26571
rect 9723 26568 9735 26571
rect 9766 26568 9772 26580
rect 9723 26540 9772 26568
rect 9723 26537 9735 26540
rect 9677 26531 9735 26537
rect 9766 26528 9772 26540
rect 9824 26528 9830 26580
rect 10318 26528 10324 26580
rect 10376 26568 10382 26580
rect 12066 26568 12072 26580
rect 10376 26540 12072 26568
rect 10376 26528 10382 26540
rect 12066 26528 12072 26540
rect 12124 26528 12130 26580
rect 12621 26571 12679 26577
rect 12621 26537 12633 26571
rect 12667 26568 12679 26571
rect 12710 26568 12716 26580
rect 12667 26540 12716 26568
rect 12667 26537 12679 26540
rect 12621 26531 12679 26537
rect 12710 26528 12716 26540
rect 12768 26528 12774 26580
rect 14369 26571 14427 26577
rect 14369 26537 14381 26571
rect 14415 26568 14427 26571
rect 14734 26568 14740 26580
rect 14415 26540 14740 26568
rect 14415 26537 14427 26540
rect 14369 26531 14427 26537
rect 14734 26528 14740 26540
rect 14792 26528 14798 26580
rect 14918 26528 14924 26580
rect 14976 26568 14982 26580
rect 15105 26571 15163 26577
rect 15105 26568 15117 26571
rect 14976 26540 15117 26568
rect 14976 26528 14982 26540
rect 15105 26537 15117 26540
rect 15151 26537 15163 26571
rect 16482 26568 16488 26580
rect 16443 26540 16488 26568
rect 15105 26531 15163 26537
rect 3786 26500 3792 26512
rect 3747 26472 3792 26500
rect 3786 26460 3792 26472
rect 3844 26460 3850 26512
rect 5629 26503 5687 26509
rect 5629 26500 5641 26503
rect 5460 26472 5641 26500
rect 5460 26432 5488 26472
rect 5629 26469 5641 26472
rect 5675 26469 5687 26503
rect 11698 26500 11704 26512
rect 5629 26463 5687 26469
rect 6288 26472 8984 26500
rect 5092 26404 5488 26432
rect 3237 26367 3295 26373
rect 3237 26333 3249 26367
rect 3283 26333 3295 26367
rect 3237 26327 3295 26333
rect 4913 26367 4971 26373
rect 4913 26333 4925 26367
rect 4959 26364 4971 26367
rect 5092 26364 5120 26404
rect 5902 26392 5908 26444
rect 5960 26432 5966 26444
rect 5960 26404 6040 26432
rect 5960 26392 5966 26404
rect 4959 26336 5120 26364
rect 5169 26367 5227 26373
rect 4959 26333 4971 26336
rect 4913 26327 4971 26333
rect 5169 26333 5181 26367
rect 5215 26364 5227 26367
rect 5258 26364 5264 26376
rect 5215 26336 5264 26364
rect 5215 26333 5227 26336
rect 5169 26327 5227 26333
rect 5258 26324 5264 26336
rect 5316 26324 5322 26376
rect 5350 26324 5356 26376
rect 5408 26364 5414 26376
rect 6012 26373 6040 26404
rect 6288 26376 6316 26472
rect 7466 26432 7472 26444
rect 7427 26404 7472 26432
rect 7466 26392 7472 26404
rect 7524 26392 7530 26444
rect 7650 26432 7656 26444
rect 7611 26404 7656 26432
rect 7650 26392 7656 26404
rect 7708 26392 7714 26444
rect 8956 26376 8984 26472
rect 9324 26472 11704 26500
rect 5767 26367 5825 26373
rect 5767 26364 5779 26367
rect 5408 26336 5779 26364
rect 5408 26324 5414 26336
rect 5767 26333 5779 26336
rect 5813 26333 5825 26367
rect 5767 26327 5825 26333
rect 5997 26367 6055 26373
rect 5997 26333 6009 26367
rect 6043 26333 6055 26367
rect 5997 26327 6055 26333
rect 6086 26324 6092 26376
rect 6144 26373 6150 26376
rect 6144 26367 6183 26373
rect 6171 26333 6183 26367
rect 6144 26327 6183 26333
rect 6144 26324 6150 26327
rect 6270 26324 6276 26376
rect 6328 26364 6334 26376
rect 7377 26367 7435 26373
rect 6328 26336 6421 26364
rect 6328 26324 6334 26336
rect 7377 26333 7389 26367
rect 7423 26364 7435 26367
rect 7834 26364 7840 26376
rect 7423 26336 7840 26364
rect 7423 26333 7435 26336
rect 7377 26327 7435 26333
rect 7834 26324 7840 26336
rect 7892 26324 7898 26376
rect 8294 26324 8300 26376
rect 8352 26364 8358 26376
rect 8389 26367 8447 26373
rect 8389 26364 8401 26367
rect 8352 26336 8401 26364
rect 8352 26324 8358 26336
rect 8389 26333 8401 26336
rect 8435 26364 8447 26367
rect 8570 26364 8576 26376
rect 8435 26336 8576 26364
rect 8435 26333 8447 26336
rect 8389 26327 8447 26333
rect 8570 26324 8576 26336
rect 8628 26324 8634 26376
rect 8938 26324 8944 26376
rect 8996 26364 9002 26376
rect 9214 26373 9220 26376
rect 9033 26367 9091 26373
rect 9033 26364 9045 26367
rect 8996 26336 9045 26364
rect 8996 26324 9002 26336
rect 9033 26333 9045 26336
rect 9079 26333 9091 26367
rect 9033 26327 9091 26333
rect 9181 26367 9220 26373
rect 9181 26333 9193 26367
rect 9181 26327 9220 26333
rect 9214 26324 9220 26327
rect 9272 26324 9278 26376
rect 9324 26373 9352 26472
rect 11698 26460 11704 26472
rect 11756 26460 11762 26512
rect 12161 26435 12219 26441
rect 12161 26432 12173 26435
rect 9692 26404 12173 26432
rect 9692 26376 9720 26404
rect 12161 26401 12173 26404
rect 12207 26401 12219 26435
rect 13998 26432 14004 26444
rect 12161 26395 12219 26401
rect 12452 26404 14004 26432
rect 9309 26367 9367 26373
rect 9309 26333 9321 26367
rect 9355 26333 9367 26367
rect 9309 26327 9367 26333
rect 9490 26324 9496 26376
rect 9548 26373 9554 26376
rect 9548 26364 9556 26373
rect 9548 26336 9593 26364
rect 9548 26327 9556 26336
rect 9548 26324 9554 26327
rect 9674 26324 9680 26376
rect 9732 26324 9738 26376
rect 10321 26367 10379 26373
rect 10321 26333 10333 26367
rect 10367 26364 10379 26367
rect 10594 26364 10600 26376
rect 10367 26336 10600 26364
rect 10367 26333 10379 26336
rect 10321 26327 10379 26333
rect 10594 26324 10600 26336
rect 10652 26364 10658 26376
rect 10778 26364 10784 26376
rect 10652 26336 10784 26364
rect 10652 26324 10658 26336
rect 10778 26324 10784 26336
rect 10836 26324 10842 26376
rect 11698 26324 11704 26376
rect 11756 26364 11762 26376
rect 11885 26367 11943 26373
rect 11885 26364 11897 26367
rect 11756 26336 11897 26364
rect 11756 26324 11762 26336
rect 11885 26333 11897 26336
rect 11931 26333 11943 26367
rect 12066 26364 12072 26376
rect 12027 26336 12072 26364
rect 11885 26327 11943 26333
rect 12066 26324 12072 26336
rect 12124 26324 12130 26376
rect 12452 26373 12480 26404
rect 13998 26392 14004 26404
rect 14056 26432 14062 26444
rect 14277 26435 14335 26441
rect 14277 26432 14289 26435
rect 14056 26404 14289 26432
rect 14056 26392 14062 26404
rect 14277 26401 14289 26404
rect 14323 26401 14335 26435
rect 14277 26395 14335 26401
rect 12253 26367 12311 26373
rect 12253 26333 12265 26367
rect 12299 26333 12311 26367
rect 12253 26327 12311 26333
rect 12437 26367 12495 26373
rect 12437 26333 12449 26367
rect 12483 26333 12495 26367
rect 12437 26327 12495 26333
rect 5905 26299 5963 26305
rect 5905 26265 5917 26299
rect 5951 26296 5963 26299
rect 8110 26296 8116 26308
rect 5951 26268 8116 26296
rect 5951 26265 5963 26268
rect 5905 26259 5963 26265
rect 8110 26256 8116 26268
rect 8168 26256 8174 26308
rect 9398 26296 9404 26308
rect 9359 26268 9404 26296
rect 9398 26256 9404 26268
rect 9456 26256 9462 26308
rect 9582 26256 9588 26308
rect 9640 26296 9646 26308
rect 9640 26268 10088 26296
rect 9640 26256 9646 26268
rect 1486 26228 1492 26240
rect 1447 26200 1492 26228
rect 1486 26188 1492 26200
rect 1544 26188 1550 26240
rect 2958 26188 2964 26240
rect 3016 26228 3022 26240
rect 3145 26231 3203 26237
rect 3145 26228 3157 26231
rect 3016 26200 3157 26228
rect 3016 26188 3022 26200
rect 3145 26197 3157 26200
rect 3191 26197 3203 26231
rect 3145 26191 3203 26197
rect 4706 26188 4712 26240
rect 4764 26228 4770 26240
rect 5350 26228 5356 26240
rect 4764 26200 5356 26228
rect 4764 26188 4770 26200
rect 5350 26188 5356 26200
rect 5408 26188 5414 26240
rect 5810 26188 5816 26240
rect 5868 26228 5874 26240
rect 9766 26228 9772 26240
rect 5868 26200 9772 26228
rect 5868 26188 5874 26200
rect 9766 26188 9772 26200
rect 9824 26188 9830 26240
rect 10060 26228 10088 26268
rect 10134 26256 10140 26308
rect 10192 26296 10198 26308
rect 10229 26299 10287 26305
rect 10229 26296 10241 26299
rect 10192 26268 10241 26296
rect 10192 26256 10198 26268
rect 10229 26265 10241 26268
rect 10275 26265 10287 26299
rect 10229 26259 10287 26265
rect 11790 26228 11796 26240
rect 10060 26200 11796 26228
rect 11790 26188 11796 26200
rect 11848 26188 11854 26240
rect 12268 26228 12296 26327
rect 14090 26324 14096 26376
rect 14148 26364 14154 26376
rect 14185 26367 14243 26373
rect 14185 26364 14197 26367
rect 14148 26336 14197 26364
rect 14148 26324 14154 26336
rect 14185 26333 14197 26336
rect 14231 26333 14243 26367
rect 14752 26364 14780 26528
rect 15013 26367 15071 26373
rect 15013 26364 15025 26367
rect 14752 26336 15025 26364
rect 14185 26327 14243 26333
rect 15013 26333 15025 26336
rect 15059 26333 15071 26367
rect 15120 26364 15148 26531
rect 16482 26528 16488 26540
rect 16540 26528 16546 26580
rect 17773 26571 17831 26577
rect 17773 26537 17785 26571
rect 17819 26568 17831 26571
rect 17862 26568 17868 26580
rect 17819 26540 17868 26568
rect 17819 26537 17831 26540
rect 17773 26531 17831 26537
rect 17862 26528 17868 26540
rect 17920 26528 17926 26580
rect 19518 26528 19524 26580
rect 19576 26568 19582 26580
rect 19613 26571 19671 26577
rect 19613 26568 19625 26571
rect 19576 26540 19625 26568
rect 19576 26528 19582 26540
rect 19613 26537 19625 26540
rect 19659 26568 19671 26571
rect 20438 26568 20444 26580
rect 19659 26540 20444 26568
rect 19659 26537 19671 26540
rect 19613 26531 19671 26537
rect 20438 26528 20444 26540
rect 20496 26528 20502 26580
rect 19886 26460 19892 26512
rect 19944 26460 19950 26512
rect 20714 26460 20720 26512
rect 20772 26460 20778 26512
rect 19904 26432 19932 26460
rect 20732 26432 20760 26460
rect 20809 26435 20867 26441
rect 20809 26432 20821 26435
rect 19904 26404 20576 26432
rect 20732 26404 20821 26432
rect 20548 26376 20576 26404
rect 20809 26401 20821 26404
rect 20855 26401 20867 26435
rect 20809 26395 20867 26401
rect 20901 26435 20959 26441
rect 20901 26401 20913 26435
rect 20947 26432 20959 26435
rect 21174 26432 21180 26444
rect 20947 26404 21180 26432
rect 20947 26401 20959 26404
rect 20901 26395 20959 26401
rect 21174 26392 21180 26404
rect 21232 26392 21238 26444
rect 21726 26432 21732 26444
rect 21687 26404 21732 26432
rect 21726 26392 21732 26404
rect 21784 26392 21790 26444
rect 15657 26367 15715 26373
rect 15657 26364 15669 26367
rect 15120 26336 15669 26364
rect 15013 26327 15071 26333
rect 15657 26333 15669 26336
rect 15703 26333 15715 26367
rect 15657 26327 15715 26333
rect 15841 26367 15899 26373
rect 15841 26333 15853 26367
rect 15887 26333 15899 26367
rect 16298 26364 16304 26376
rect 16259 26336 16304 26364
rect 15841 26327 15899 26333
rect 14918 26256 14924 26308
rect 14976 26296 14982 26308
rect 15102 26296 15108 26308
rect 14976 26268 15108 26296
rect 14976 26256 14982 26268
rect 15102 26256 15108 26268
rect 15160 26296 15166 26308
rect 15856 26296 15884 26327
rect 16298 26324 16304 26336
rect 16356 26324 16362 26376
rect 16758 26324 16764 26376
rect 16816 26364 16822 26376
rect 17405 26367 17463 26373
rect 17405 26364 17417 26367
rect 16816 26336 17417 26364
rect 16816 26324 16822 26336
rect 17405 26333 17417 26336
rect 17451 26333 17463 26367
rect 18230 26364 18236 26376
rect 18191 26336 18236 26364
rect 17405 26327 17463 26333
rect 18230 26324 18236 26336
rect 18288 26324 18294 26376
rect 19426 26324 19432 26376
rect 19484 26364 19490 26376
rect 19521 26367 19579 26373
rect 19521 26364 19533 26367
rect 19484 26336 19533 26364
rect 19484 26324 19490 26336
rect 19521 26333 19533 26336
rect 19567 26333 19579 26367
rect 19521 26327 19579 26333
rect 19702 26324 19708 26376
rect 19760 26364 19766 26376
rect 19797 26367 19855 26373
rect 19797 26364 19809 26367
rect 19760 26336 19809 26364
rect 19760 26324 19766 26336
rect 19797 26333 19809 26336
rect 19843 26333 19855 26367
rect 19797 26327 19855 26333
rect 19886 26324 19892 26376
rect 19944 26364 19950 26376
rect 20530 26364 20536 26376
rect 19944 26336 19989 26364
rect 20443 26336 20536 26364
rect 19944 26324 19950 26336
rect 20530 26324 20536 26336
rect 20588 26324 20594 26376
rect 20622 26324 20628 26376
rect 20680 26364 20686 26376
rect 20717 26367 20775 26373
rect 20717 26364 20729 26367
rect 20680 26336 20729 26364
rect 20680 26324 20686 26336
rect 20717 26333 20729 26336
rect 20763 26333 20775 26367
rect 21082 26364 21088 26376
rect 20995 26336 21088 26364
rect 20717 26327 20775 26333
rect 17586 26296 17592 26308
rect 15160 26268 15884 26296
rect 17547 26268 17592 26296
rect 15160 26256 15166 26268
rect 17586 26256 17592 26268
rect 17644 26256 17650 26308
rect 17954 26256 17960 26308
rect 18012 26296 18018 26308
rect 18325 26299 18383 26305
rect 18325 26296 18337 26299
rect 18012 26268 18337 26296
rect 18012 26256 18018 26268
rect 18325 26265 18337 26268
rect 18371 26265 18383 26299
rect 20732 26296 20760 26327
rect 21082 26324 21088 26336
rect 21140 26364 21146 26376
rect 21358 26364 21364 26376
rect 21140 26336 21364 26364
rect 21140 26324 21146 26336
rect 21358 26324 21364 26336
rect 21416 26324 21422 26376
rect 21269 26299 21327 26305
rect 20732 26268 20852 26296
rect 18325 26259 18383 26265
rect 12342 26228 12348 26240
rect 12268 26200 12348 26228
rect 12342 26188 12348 26200
rect 12400 26188 12406 26240
rect 14550 26228 14556 26240
rect 14511 26200 14556 26228
rect 14550 26188 14556 26200
rect 14608 26188 14614 26240
rect 15746 26228 15752 26240
rect 15707 26200 15752 26228
rect 15746 26188 15752 26200
rect 15804 26188 15810 26240
rect 18046 26188 18052 26240
rect 18104 26228 18110 26240
rect 18230 26228 18236 26240
rect 18104 26200 18236 26228
rect 18104 26188 18110 26200
rect 18230 26188 18236 26200
rect 18288 26188 18294 26240
rect 19981 26231 20039 26237
rect 19981 26197 19993 26231
rect 20027 26228 20039 26231
rect 20714 26228 20720 26240
rect 20027 26200 20720 26228
rect 20027 26197 20039 26200
rect 19981 26191 20039 26197
rect 20714 26188 20720 26200
rect 20772 26188 20778 26240
rect 20824 26228 20852 26268
rect 21269 26265 21281 26299
rect 21315 26296 21327 26299
rect 21974 26299 22032 26305
rect 21974 26296 21986 26299
rect 21315 26268 21986 26296
rect 21315 26265 21327 26268
rect 21269 26259 21327 26265
rect 21974 26265 21986 26268
rect 22020 26265 22032 26299
rect 21974 26259 22032 26265
rect 22186 26228 22192 26240
rect 20824 26200 22192 26228
rect 22186 26188 22192 26200
rect 22244 26228 22250 26240
rect 23109 26231 23167 26237
rect 23109 26228 23121 26231
rect 22244 26200 23121 26228
rect 22244 26188 22250 26200
rect 23109 26197 23121 26200
rect 23155 26197 23167 26231
rect 23109 26191 23167 26197
rect 1104 26138 30820 26160
rect 1104 26086 10880 26138
rect 10932 26086 10944 26138
rect 10996 26086 11008 26138
rect 11060 26086 11072 26138
rect 11124 26086 11136 26138
rect 11188 26086 20811 26138
rect 20863 26086 20875 26138
rect 20927 26086 20939 26138
rect 20991 26086 21003 26138
rect 21055 26086 21067 26138
rect 21119 26086 30820 26138
rect 1104 26064 30820 26086
rect 2866 25984 2872 26036
rect 2924 26024 2930 26036
rect 3237 26027 3295 26033
rect 3237 26024 3249 26027
rect 2924 25996 3249 26024
rect 2924 25984 2930 25996
rect 3237 25993 3249 25996
rect 3283 25993 3295 26027
rect 3237 25987 3295 25993
rect 4525 26027 4583 26033
rect 4525 25993 4537 26027
rect 4571 26024 4583 26027
rect 5534 26024 5540 26036
rect 4571 25996 5540 26024
rect 4571 25993 4583 25996
rect 4525 25987 4583 25993
rect 5534 25984 5540 25996
rect 5592 25984 5598 26036
rect 6270 26024 6276 26036
rect 5644 25996 6276 26024
rect 4890 25956 4896 25968
rect 4851 25928 4896 25956
rect 4890 25916 4896 25928
rect 4948 25916 4954 25968
rect 1673 25891 1731 25897
rect 1673 25857 1685 25891
rect 1719 25888 1731 25891
rect 2958 25888 2964 25900
rect 1719 25860 2964 25888
rect 1719 25857 1731 25860
rect 1673 25851 1731 25857
rect 2958 25848 2964 25860
rect 3016 25848 3022 25900
rect 3142 25888 3148 25900
rect 3103 25860 3148 25888
rect 3142 25848 3148 25860
rect 3200 25848 3206 25900
rect 4706 25897 4712 25900
rect 3329 25891 3387 25897
rect 3329 25857 3341 25891
rect 3375 25857 3387 25891
rect 4704 25888 4712 25897
rect 4667 25860 4712 25888
rect 3329 25851 3387 25857
rect 4704 25851 4712 25860
rect 3344 25820 3372 25851
rect 4706 25848 4712 25851
rect 4764 25848 4770 25900
rect 4798 25848 4804 25900
rect 4856 25888 4862 25900
rect 5074 25888 5080 25900
rect 4856 25860 4901 25888
rect 5035 25860 5080 25888
rect 4856 25848 4862 25860
rect 5074 25848 5080 25860
rect 5132 25848 5138 25900
rect 5169 25891 5227 25897
rect 5169 25857 5181 25891
rect 5215 25888 5227 25891
rect 5644 25888 5672 25996
rect 6270 25984 6276 25996
rect 6328 25984 6334 26036
rect 6822 25984 6828 26036
rect 6880 26024 6886 26036
rect 6880 25996 8156 26024
rect 6880 25984 6886 25996
rect 5721 25959 5779 25965
rect 5721 25925 5733 25959
rect 5767 25956 5779 25959
rect 5767 25928 6868 25956
rect 5767 25925 5779 25928
rect 5721 25919 5779 25925
rect 5810 25888 5816 25900
rect 5215 25860 5672 25888
rect 5771 25860 5816 25888
rect 5215 25857 5227 25860
rect 5169 25851 5227 25857
rect 5810 25848 5816 25860
rect 5868 25848 5874 25900
rect 5902 25848 5908 25900
rect 5960 25888 5966 25900
rect 6457 25891 6515 25897
rect 6457 25888 6469 25891
rect 5960 25860 6469 25888
rect 5960 25848 5966 25860
rect 6457 25857 6469 25860
rect 6503 25857 6515 25891
rect 6730 25888 6736 25900
rect 6691 25860 6736 25888
rect 6457 25851 6515 25857
rect 6730 25848 6736 25860
rect 6788 25848 6794 25900
rect 6840 25888 6868 25928
rect 7006 25916 7012 25968
rect 7064 25956 7070 25968
rect 7561 25959 7619 25965
rect 7561 25956 7573 25959
rect 7064 25928 7573 25956
rect 7064 25916 7070 25928
rect 7561 25925 7573 25928
rect 7607 25925 7619 25959
rect 7561 25919 7619 25925
rect 7745 25959 7803 25965
rect 7745 25925 7757 25959
rect 7791 25956 7803 25959
rect 8018 25956 8024 25968
rect 7791 25928 8024 25956
rect 7791 25925 7803 25928
rect 7745 25919 7803 25925
rect 8018 25916 8024 25928
rect 8076 25916 8082 25968
rect 8128 25956 8156 25996
rect 8404 25996 9536 26024
rect 8404 25956 8432 25996
rect 8128 25928 8432 25956
rect 8665 25959 8723 25965
rect 8665 25925 8677 25959
rect 8711 25956 8723 25959
rect 9122 25956 9128 25968
rect 8711 25928 9128 25956
rect 8711 25925 8723 25928
rect 8665 25919 8723 25925
rect 9122 25916 9128 25928
rect 9180 25916 9186 25968
rect 7374 25888 7380 25900
rect 6840 25860 7380 25888
rect 7374 25848 7380 25860
rect 7432 25848 7438 25900
rect 8570 25848 8576 25900
rect 8628 25888 8634 25900
rect 9508 25897 9536 25996
rect 9766 25984 9772 26036
rect 9824 26024 9830 26036
rect 10318 26024 10324 26036
rect 9824 25996 10324 26024
rect 9824 25984 9830 25996
rect 10318 25984 10324 25996
rect 10376 26024 10382 26036
rect 10873 26027 10931 26033
rect 10873 26024 10885 26027
rect 10376 25996 10885 26024
rect 10376 25984 10382 25996
rect 10873 25993 10885 25996
rect 10919 25993 10931 26027
rect 10873 25987 10931 25993
rect 15657 26027 15715 26033
rect 15657 25993 15669 26027
rect 15703 26024 15715 26027
rect 15746 26024 15752 26036
rect 15703 25996 15752 26024
rect 15703 25993 15715 25996
rect 15657 25987 15715 25993
rect 15746 25984 15752 25996
rect 15804 25984 15810 26036
rect 17586 26024 17592 26036
rect 17547 25996 17592 26024
rect 17586 25984 17592 25996
rect 17644 25984 17650 26036
rect 19886 25984 19892 26036
rect 19944 26024 19950 26036
rect 20073 26027 20131 26033
rect 20073 26024 20085 26027
rect 19944 25996 20085 26024
rect 19944 25984 19950 25996
rect 20073 25993 20085 25996
rect 20119 25993 20131 26027
rect 21910 26024 21916 26036
rect 20073 25987 20131 25993
rect 20732 25996 21496 26024
rect 21871 25996 21916 26024
rect 13354 25956 13360 25968
rect 13315 25928 13360 25956
rect 13354 25916 13360 25928
rect 13412 25916 13418 25968
rect 14829 25959 14887 25965
rect 14829 25925 14841 25959
rect 14875 25956 14887 25959
rect 18598 25956 18604 25968
rect 14875 25928 18604 25956
rect 14875 25925 14887 25928
rect 14829 25919 14887 25925
rect 18598 25916 18604 25928
rect 18656 25916 18662 25968
rect 19429 25959 19487 25965
rect 19429 25925 19441 25959
rect 19475 25956 19487 25959
rect 19518 25956 19524 25968
rect 19475 25928 19524 25956
rect 19475 25925 19487 25928
rect 19429 25919 19487 25925
rect 19518 25916 19524 25928
rect 19576 25916 19582 25968
rect 19794 25916 19800 25968
rect 19852 25916 19858 25968
rect 9493 25891 9551 25897
rect 8628 25860 8892 25888
rect 8628 25848 8634 25860
rect 8754 25820 8760 25832
rect 3344 25792 8340 25820
rect 8715 25792 8760 25820
rect 5718 25712 5724 25764
rect 5776 25752 5782 25764
rect 8312 25761 8340 25792
rect 8754 25780 8760 25792
rect 8812 25780 8818 25832
rect 8864 25829 8892 25860
rect 9493 25857 9505 25891
rect 9539 25857 9551 25891
rect 9493 25851 9551 25857
rect 9582 25848 9588 25900
rect 9640 25848 9646 25900
rect 9766 25897 9772 25900
rect 9760 25851 9772 25897
rect 9824 25888 9830 25900
rect 9824 25860 9860 25888
rect 9766 25848 9772 25851
rect 9824 25848 9830 25860
rect 11698 25848 11704 25900
rect 11756 25888 11762 25900
rect 11977 25891 12035 25897
rect 11977 25888 11989 25891
rect 11756 25860 11989 25888
rect 11756 25848 11762 25860
rect 11977 25857 11989 25860
rect 12023 25857 12035 25891
rect 11977 25851 12035 25857
rect 12161 25891 12219 25897
rect 12161 25857 12173 25891
rect 12207 25857 12219 25891
rect 12161 25851 12219 25857
rect 8849 25823 8907 25829
rect 8849 25789 8861 25823
rect 8895 25789 8907 25823
rect 9600 25820 9628 25848
rect 8849 25783 8907 25789
rect 9508 25792 9628 25820
rect 6549 25755 6607 25761
rect 6549 25752 6561 25755
rect 5776 25724 6561 25752
rect 5776 25712 5782 25724
rect 6549 25721 6561 25724
rect 6595 25721 6607 25755
rect 6549 25715 6607 25721
rect 6641 25755 6699 25761
rect 6641 25721 6653 25755
rect 6687 25721 6699 25755
rect 6641 25715 6699 25721
rect 8297 25755 8355 25761
rect 8297 25721 8309 25755
rect 8343 25721 8355 25755
rect 8297 25715 8355 25721
rect 1486 25684 1492 25696
rect 1447 25656 1492 25684
rect 1486 25644 1492 25656
rect 1544 25644 1550 25696
rect 6270 25644 6276 25696
rect 6328 25684 6334 25696
rect 6656 25684 6684 25715
rect 6328 25656 6684 25684
rect 6917 25687 6975 25693
rect 6328 25644 6334 25656
rect 6917 25653 6929 25687
rect 6963 25684 6975 25687
rect 9508 25684 9536 25792
rect 11422 25780 11428 25832
rect 11480 25820 11486 25832
rect 12176 25820 12204 25851
rect 12250 25848 12256 25900
rect 12308 25888 12314 25900
rect 12529 25891 12587 25897
rect 12308 25860 12353 25888
rect 12308 25848 12314 25860
rect 12529 25857 12541 25891
rect 12575 25888 12587 25891
rect 12894 25888 12900 25900
rect 12575 25860 12900 25888
rect 12575 25857 12587 25860
rect 12529 25851 12587 25857
rect 12894 25848 12900 25860
rect 12952 25888 12958 25900
rect 14737 25891 14795 25897
rect 14737 25888 14749 25891
rect 12952 25860 14749 25888
rect 12952 25848 12958 25860
rect 14737 25857 14749 25860
rect 14783 25857 14795 25891
rect 14737 25851 14795 25857
rect 15749 25891 15807 25897
rect 15749 25857 15761 25891
rect 15795 25888 15807 25891
rect 16482 25888 16488 25900
rect 15795 25860 16488 25888
rect 15795 25857 15807 25860
rect 15749 25851 15807 25857
rect 16482 25848 16488 25860
rect 16540 25848 16546 25900
rect 16945 25891 17003 25897
rect 16945 25857 16957 25891
rect 16991 25888 17003 25891
rect 17034 25888 17040 25900
rect 16991 25860 17040 25888
rect 16991 25857 17003 25860
rect 16945 25851 17003 25857
rect 17034 25848 17040 25860
rect 17092 25848 17098 25900
rect 17957 25891 18015 25897
rect 17957 25857 17969 25891
rect 18003 25888 18015 25891
rect 18414 25888 18420 25900
rect 18003 25860 18420 25888
rect 18003 25857 18015 25860
rect 17957 25851 18015 25857
rect 18414 25848 18420 25860
rect 18472 25888 18478 25900
rect 18966 25888 18972 25900
rect 18472 25860 18972 25888
rect 18472 25848 18478 25860
rect 18966 25848 18972 25860
rect 19024 25848 19030 25900
rect 19812 25888 19840 25916
rect 19628 25860 19840 25888
rect 19889 25891 19947 25897
rect 12342 25820 12348 25832
rect 11480 25792 12204 25820
rect 12303 25792 12348 25820
rect 11480 25780 11486 25792
rect 12342 25780 12348 25792
rect 12400 25780 12406 25832
rect 15565 25823 15623 25829
rect 15565 25789 15577 25823
rect 15611 25820 15623 25823
rect 16850 25820 16856 25832
rect 15611 25792 16856 25820
rect 15611 25789 15623 25792
rect 15565 25783 15623 25789
rect 16850 25780 16856 25792
rect 16908 25780 16914 25832
rect 18046 25820 18052 25832
rect 18007 25792 18052 25820
rect 18046 25780 18052 25792
rect 18104 25780 18110 25832
rect 18141 25823 18199 25829
rect 18141 25789 18153 25823
rect 18187 25789 18199 25823
rect 18141 25783 18199 25789
rect 11882 25712 11888 25764
rect 11940 25752 11946 25764
rect 13173 25755 13231 25761
rect 13173 25752 13185 25755
rect 11940 25724 13185 25752
rect 11940 25712 11946 25724
rect 13173 25721 13185 25724
rect 13219 25721 13231 25755
rect 16868 25752 16896 25780
rect 17494 25752 17500 25764
rect 16868 25724 17500 25752
rect 13173 25715 13231 25721
rect 17494 25712 17500 25724
rect 17552 25752 17558 25764
rect 18156 25752 18184 25783
rect 19518 25780 19524 25832
rect 19576 25820 19582 25832
rect 19628 25820 19656 25860
rect 19889 25857 19901 25891
rect 19935 25857 19947 25891
rect 20530 25888 20536 25900
rect 20491 25860 20536 25888
rect 19889 25851 19947 25857
rect 19794 25820 19800 25832
rect 19576 25792 19656 25820
rect 19755 25792 19800 25820
rect 19576 25780 19582 25792
rect 19794 25780 19800 25792
rect 19852 25780 19858 25832
rect 19904 25820 19932 25851
rect 20530 25848 20536 25860
rect 20588 25848 20594 25900
rect 20732 25897 20760 25996
rect 21358 25956 21364 25968
rect 21100 25928 21364 25956
rect 21100 25900 21128 25928
rect 21358 25916 21364 25928
rect 21416 25916 21422 25968
rect 20717 25891 20775 25897
rect 20717 25857 20729 25891
rect 20763 25857 20775 25891
rect 20717 25851 20775 25857
rect 20806 25848 20812 25900
rect 20864 25888 20870 25900
rect 21082 25888 21088 25900
rect 20864 25860 20909 25888
rect 21043 25860 21088 25888
rect 20864 25848 20870 25860
rect 21082 25848 21088 25860
rect 21140 25848 21146 25900
rect 21468 25888 21496 25996
rect 21910 25984 21916 25996
rect 21968 25984 21974 26036
rect 22002 25888 22008 25900
rect 21468 25860 22008 25888
rect 22002 25848 22008 25860
rect 22060 25848 22066 25900
rect 29178 25848 29184 25900
rect 29236 25888 29242 25900
rect 29825 25891 29883 25897
rect 29825 25888 29837 25891
rect 29236 25860 29837 25888
rect 29236 25848 29242 25860
rect 29825 25857 29837 25860
rect 29871 25857 29883 25891
rect 29825 25851 29883 25857
rect 20901 25823 20959 25829
rect 19904 25792 20668 25820
rect 17552 25724 18184 25752
rect 17552 25712 17558 25724
rect 20640 25696 20668 25792
rect 20901 25789 20913 25823
rect 20947 25789 20959 25823
rect 20901 25783 20959 25789
rect 21269 25823 21327 25829
rect 21269 25789 21281 25823
rect 21315 25820 21327 25823
rect 22094 25820 22100 25832
rect 21315 25792 22100 25820
rect 21315 25789 21327 25792
rect 21269 25783 21327 25789
rect 20806 25712 20812 25764
rect 20864 25752 20870 25764
rect 20916 25752 20944 25783
rect 22094 25780 22100 25792
rect 22152 25780 22158 25832
rect 20864 25724 20944 25752
rect 20864 25712 20870 25724
rect 6963 25656 9536 25684
rect 12713 25687 12771 25693
rect 6963 25653 6975 25656
rect 6917 25647 6975 25653
rect 12713 25653 12725 25687
rect 12759 25684 12771 25687
rect 13998 25684 14004 25696
rect 12759 25656 14004 25684
rect 12759 25653 12771 25656
rect 12713 25647 12771 25653
rect 13998 25644 14004 25656
rect 14056 25644 14062 25696
rect 16117 25687 16175 25693
rect 16117 25653 16129 25687
rect 16163 25684 16175 25687
rect 16206 25684 16212 25696
rect 16163 25656 16212 25684
rect 16163 25653 16175 25656
rect 16117 25647 16175 25653
rect 16206 25644 16212 25656
rect 16264 25644 16270 25696
rect 17037 25687 17095 25693
rect 17037 25653 17049 25687
rect 17083 25684 17095 25687
rect 17678 25684 17684 25696
rect 17083 25656 17684 25684
rect 17083 25653 17095 25656
rect 17037 25647 17095 25653
rect 17678 25644 17684 25656
rect 17736 25644 17742 25696
rect 19610 25684 19616 25696
rect 19571 25656 19616 25684
rect 19610 25644 19616 25656
rect 19668 25684 19674 25696
rect 19978 25684 19984 25696
rect 19668 25656 19984 25684
rect 19668 25644 19674 25656
rect 19978 25644 19984 25656
rect 20036 25644 20042 25696
rect 20622 25644 20628 25696
rect 20680 25644 20686 25696
rect 30006 25684 30012 25696
rect 29967 25656 30012 25684
rect 30006 25644 30012 25656
rect 30064 25644 30070 25696
rect 1104 25594 30820 25616
rect 1104 25542 5915 25594
rect 5967 25542 5979 25594
rect 6031 25542 6043 25594
rect 6095 25542 6107 25594
rect 6159 25542 6171 25594
rect 6223 25542 15846 25594
rect 15898 25542 15910 25594
rect 15962 25542 15974 25594
rect 16026 25542 16038 25594
rect 16090 25542 16102 25594
rect 16154 25542 25776 25594
rect 25828 25542 25840 25594
rect 25892 25542 25904 25594
rect 25956 25542 25968 25594
rect 26020 25542 26032 25594
rect 26084 25542 30820 25594
rect 1104 25520 30820 25542
rect 6365 25483 6423 25489
rect 6365 25449 6377 25483
rect 6411 25480 6423 25483
rect 6411 25452 8708 25480
rect 6411 25449 6423 25452
rect 6365 25443 6423 25449
rect 4154 25372 4160 25424
rect 4212 25412 4218 25424
rect 6917 25415 6975 25421
rect 6917 25412 6929 25415
rect 4212 25384 6929 25412
rect 4212 25372 4218 25384
rect 6917 25381 6929 25384
rect 6963 25381 6975 25415
rect 8680 25412 8708 25452
rect 8956 25452 9536 25480
rect 8956 25412 8984 25452
rect 8680 25384 8984 25412
rect 6917 25375 6975 25381
rect 7466 25344 7472 25356
rect 7427 25316 7472 25344
rect 7466 25304 7472 25316
rect 7524 25344 7530 25356
rect 7650 25344 7656 25356
rect 7524 25316 7656 25344
rect 7524 25304 7530 25316
rect 7650 25304 7656 25316
rect 7708 25304 7714 25356
rect 7742 25304 7748 25356
rect 7800 25344 7806 25356
rect 8386 25344 8392 25356
rect 7800 25316 8392 25344
rect 7800 25304 7806 25316
rect 8386 25304 8392 25316
rect 8444 25344 8450 25356
rect 9401 25347 9459 25353
rect 9401 25344 9413 25347
rect 8444 25316 9413 25344
rect 8444 25304 8450 25316
rect 9401 25313 9413 25316
rect 9447 25313 9459 25347
rect 9401 25307 9459 25313
rect 6270 25276 6276 25288
rect 6231 25248 6276 25276
rect 6270 25236 6276 25248
rect 6328 25236 6334 25288
rect 7834 25236 7840 25288
rect 7892 25276 7898 25288
rect 8113 25279 8171 25285
rect 8113 25276 8125 25279
rect 7892 25248 8125 25276
rect 7892 25236 7898 25248
rect 8113 25245 8125 25248
rect 8159 25245 8171 25279
rect 8113 25239 8171 25245
rect 8754 25236 8760 25288
rect 8812 25276 8818 25288
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8812 25248 8953 25276
rect 8812 25236 8818 25248
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 9125 25279 9183 25285
rect 9125 25274 9137 25279
rect 8941 25239 8999 25245
rect 9048 25246 9137 25274
rect 5721 25211 5779 25217
rect 5721 25177 5733 25211
rect 5767 25208 5779 25211
rect 6546 25208 6552 25220
rect 5767 25180 6552 25208
rect 5767 25177 5779 25180
rect 5721 25171 5779 25177
rect 6546 25168 6552 25180
rect 6604 25168 6610 25220
rect 7282 25208 7288 25220
rect 7243 25180 7288 25208
rect 7282 25168 7288 25180
rect 7340 25168 7346 25220
rect 5626 25140 5632 25152
rect 5587 25112 5632 25140
rect 5626 25100 5632 25112
rect 5684 25100 5690 25152
rect 7374 25100 7380 25152
rect 7432 25140 7438 25152
rect 8205 25143 8263 25149
rect 7432 25112 7477 25140
rect 7432 25100 7438 25112
rect 8205 25109 8217 25143
rect 8251 25140 8263 25143
rect 8938 25140 8944 25152
rect 8251 25112 8944 25140
rect 8251 25109 8263 25112
rect 8205 25103 8263 25109
rect 8938 25100 8944 25112
rect 8996 25100 9002 25152
rect 9048 25140 9076 25246
rect 9125 25245 9137 25246
rect 9171 25245 9183 25279
rect 9125 25239 9183 25245
rect 9306 25236 9312 25288
rect 9364 25276 9370 25288
rect 9508 25285 9536 25452
rect 9858 25440 9864 25492
rect 9916 25480 9922 25492
rect 10321 25483 10379 25489
rect 10321 25480 10333 25483
rect 9916 25452 10333 25480
rect 9916 25440 9922 25452
rect 10321 25449 10333 25452
rect 10367 25480 10379 25483
rect 10410 25480 10416 25492
rect 10367 25452 10416 25480
rect 10367 25449 10379 25452
rect 10321 25443 10379 25449
rect 10410 25440 10416 25452
rect 10468 25440 10474 25492
rect 14185 25483 14243 25489
rect 14185 25449 14197 25483
rect 14231 25480 14243 25483
rect 18046 25480 18052 25492
rect 14231 25452 18052 25480
rect 14231 25449 14243 25452
rect 14185 25443 14243 25449
rect 18046 25440 18052 25452
rect 18104 25440 18110 25492
rect 19702 25480 19708 25492
rect 19663 25452 19708 25480
rect 19702 25440 19708 25452
rect 19760 25440 19766 25492
rect 20622 25480 20628 25492
rect 20583 25452 20628 25480
rect 20622 25440 20628 25452
rect 20680 25440 20686 25492
rect 20901 25483 20959 25489
rect 20901 25449 20913 25483
rect 20947 25480 20959 25483
rect 21174 25480 21180 25492
rect 20947 25452 21180 25480
rect 20947 25449 20959 25452
rect 20901 25443 20959 25449
rect 21174 25440 21180 25452
rect 21232 25440 21238 25492
rect 12618 25412 12624 25424
rect 12531 25384 12624 25412
rect 12618 25372 12624 25384
rect 12676 25412 12682 25424
rect 12676 25384 14136 25412
rect 12676 25372 12682 25384
rect 9493 25279 9551 25285
rect 9364 25248 9409 25276
rect 9364 25236 9370 25248
rect 9493 25245 9505 25279
rect 9539 25245 9551 25279
rect 9674 25276 9680 25288
rect 9635 25248 9680 25276
rect 9493 25239 9551 25245
rect 9674 25236 9680 25248
rect 9732 25236 9738 25288
rect 10413 25279 10471 25285
rect 10413 25245 10425 25279
rect 10459 25276 10471 25279
rect 10502 25276 10508 25288
rect 10459 25248 10508 25276
rect 10459 25245 10471 25248
rect 10413 25239 10471 25245
rect 10502 25236 10508 25248
rect 10560 25236 10566 25288
rect 11241 25279 11299 25285
rect 11241 25245 11253 25279
rect 11287 25276 11299 25279
rect 12710 25276 12716 25288
rect 11287 25248 12716 25276
rect 11287 25245 11299 25248
rect 11241 25239 11299 25245
rect 12710 25236 12716 25248
rect 12768 25236 12774 25288
rect 14108 25285 14136 25384
rect 14274 25372 14280 25424
rect 14332 25412 14338 25424
rect 15013 25415 15071 25421
rect 15013 25412 15025 25415
rect 14332 25384 15025 25412
rect 14332 25372 14338 25384
rect 15013 25381 15025 25384
rect 15059 25412 15071 25415
rect 21726 25412 21732 25424
rect 15059 25384 21732 25412
rect 15059 25381 15071 25384
rect 15013 25375 15071 25381
rect 21726 25372 21732 25384
rect 21784 25372 21790 25424
rect 16666 25344 16672 25356
rect 16408 25316 16672 25344
rect 14093 25279 14151 25285
rect 14093 25245 14105 25279
rect 14139 25245 14151 25279
rect 14093 25239 14151 25245
rect 15933 25279 15991 25285
rect 15933 25245 15945 25279
rect 15979 25276 15991 25279
rect 16206 25276 16212 25288
rect 15979 25248 16212 25276
rect 15979 25245 15991 25248
rect 15933 25239 15991 25245
rect 16206 25236 16212 25248
rect 16264 25236 16270 25288
rect 11508 25211 11566 25217
rect 11508 25177 11520 25211
rect 11554 25208 11566 25211
rect 11790 25208 11796 25220
rect 11554 25180 11796 25208
rect 11554 25177 11566 25180
rect 11508 25171 11566 25177
rect 11790 25168 11796 25180
rect 11848 25168 11854 25220
rect 11882 25168 11888 25220
rect 11940 25208 11946 25220
rect 14829 25211 14887 25217
rect 14829 25208 14841 25211
rect 11940 25180 14841 25208
rect 11940 25168 11946 25180
rect 14829 25177 14841 25180
rect 14875 25177 14887 25211
rect 14829 25171 14887 25177
rect 16117 25211 16175 25217
rect 16117 25177 16129 25211
rect 16163 25208 16175 25211
rect 16408 25208 16436 25316
rect 16666 25304 16672 25316
rect 16724 25304 16730 25356
rect 16850 25344 16856 25356
rect 16811 25316 16856 25344
rect 16850 25304 16856 25316
rect 16908 25304 16914 25356
rect 19797 25347 19855 25353
rect 19797 25313 19809 25347
rect 19843 25344 19855 25347
rect 19978 25344 19984 25356
rect 19843 25316 19984 25344
rect 19843 25313 19855 25316
rect 19797 25307 19855 25313
rect 19978 25304 19984 25316
rect 20036 25304 20042 25356
rect 20530 25344 20536 25356
rect 20491 25316 20536 25344
rect 20530 25304 20536 25316
rect 20588 25304 20594 25356
rect 21818 25344 21824 25356
rect 20818 25316 21824 25344
rect 16574 25236 16580 25288
rect 16632 25276 16638 25288
rect 16945 25279 17003 25285
rect 16945 25276 16957 25279
rect 16632 25248 16957 25276
rect 16632 25236 16638 25248
rect 16945 25245 16957 25248
rect 16991 25245 17003 25279
rect 19518 25276 19524 25288
rect 19479 25248 19524 25276
rect 16945 25239 17003 25245
rect 19518 25236 19524 25248
rect 19576 25236 19582 25288
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 16163 25180 16436 25208
rect 16163 25177 16175 25180
rect 16117 25171 16175 25177
rect 16482 25168 16488 25220
rect 16540 25208 16546 25220
rect 17037 25211 17095 25217
rect 17037 25208 17049 25211
rect 16540 25180 17049 25208
rect 16540 25168 16546 25180
rect 17037 25177 17049 25180
rect 17083 25177 17095 25211
rect 17037 25171 17095 25177
rect 18414 25168 18420 25220
rect 18472 25208 18478 25220
rect 18601 25211 18659 25217
rect 18601 25208 18613 25211
rect 18472 25180 18613 25208
rect 18472 25168 18478 25180
rect 18601 25177 18613 25180
rect 18647 25208 18659 25211
rect 19426 25208 19432 25220
rect 18647 25180 19432 25208
rect 18647 25177 18659 25180
rect 18601 25171 18659 25177
rect 19426 25168 19432 25180
rect 19484 25168 19490 25220
rect 19628 25208 19656 25239
rect 19702 25236 19708 25288
rect 19760 25276 19766 25288
rect 20257 25279 20315 25285
rect 20257 25276 20269 25279
rect 19760 25248 20269 25276
rect 19760 25236 19766 25248
rect 20257 25245 20269 25248
rect 20303 25245 20315 25279
rect 20257 25239 20315 25245
rect 20714 25236 20720 25288
rect 20772 25276 20778 25288
rect 20818 25276 20846 25316
rect 21818 25304 21824 25316
rect 21876 25304 21882 25356
rect 21637 25279 21695 25285
rect 20772 25248 20865 25276
rect 20772 25236 20778 25248
rect 21637 25245 21649 25279
rect 21683 25276 21695 25279
rect 22186 25276 22192 25288
rect 21683 25248 22192 25276
rect 21683 25245 21695 25248
rect 21637 25239 21695 25245
rect 22186 25236 22192 25248
rect 22244 25236 22250 25288
rect 20070 25208 20076 25220
rect 19628 25180 20076 25208
rect 20070 25168 20076 25180
rect 20128 25168 20134 25220
rect 21542 25168 21548 25220
rect 21600 25208 21606 25220
rect 21729 25211 21787 25217
rect 21729 25208 21741 25211
rect 21600 25180 21741 25208
rect 21600 25168 21606 25180
rect 21729 25177 21741 25180
rect 21775 25208 21787 25211
rect 22094 25208 22100 25220
rect 21775 25180 22100 25208
rect 21775 25177 21787 25180
rect 21729 25171 21787 25177
rect 22094 25168 22100 25180
rect 22152 25168 22158 25220
rect 11238 25140 11244 25152
rect 9048 25112 11244 25140
rect 11238 25100 11244 25112
rect 11296 25100 11302 25152
rect 15746 25140 15752 25152
rect 15707 25112 15752 25140
rect 15746 25100 15752 25112
rect 15804 25100 15810 25152
rect 17218 25100 17224 25152
rect 17276 25140 17282 25152
rect 17405 25143 17463 25149
rect 17405 25140 17417 25143
rect 17276 25112 17417 25140
rect 17276 25100 17282 25112
rect 17405 25109 17417 25112
rect 17451 25109 17463 25143
rect 17405 25103 17463 25109
rect 18046 25100 18052 25152
rect 18104 25140 18110 25152
rect 18509 25143 18567 25149
rect 18509 25140 18521 25143
rect 18104 25112 18521 25140
rect 18104 25100 18110 25112
rect 18509 25109 18521 25112
rect 18555 25109 18567 25143
rect 18509 25103 18567 25109
rect 1104 25050 30820 25072
rect 1104 24998 10880 25050
rect 10932 24998 10944 25050
rect 10996 24998 11008 25050
rect 11060 24998 11072 25050
rect 11124 24998 11136 25050
rect 11188 24998 20811 25050
rect 20863 24998 20875 25050
rect 20927 24998 20939 25050
rect 20991 24998 21003 25050
rect 21055 24998 21067 25050
rect 21119 24998 30820 25050
rect 1104 24976 30820 24998
rect 6917 24939 6975 24945
rect 6917 24905 6929 24939
rect 6963 24936 6975 24939
rect 7374 24936 7380 24948
rect 6963 24908 7380 24936
rect 6963 24905 6975 24908
rect 6917 24899 6975 24905
rect 7374 24896 7380 24908
rect 7432 24896 7438 24948
rect 7650 24936 7656 24948
rect 7484 24908 7656 24936
rect 7484 24868 7512 24908
rect 7650 24896 7656 24908
rect 7708 24896 7714 24948
rect 8110 24896 8116 24948
rect 8168 24936 8174 24948
rect 9677 24939 9735 24945
rect 8168 24908 8340 24936
rect 8168 24896 8174 24908
rect 8312 24868 8340 24908
rect 9677 24905 9689 24939
rect 9723 24936 9735 24939
rect 9766 24936 9772 24948
rect 9723 24908 9772 24936
rect 9723 24905 9735 24908
rect 9677 24899 9735 24905
rect 9766 24896 9772 24908
rect 9824 24896 9830 24948
rect 11790 24896 11796 24948
rect 11848 24936 11854 24948
rect 12253 24939 12311 24945
rect 12253 24936 12265 24939
rect 11848 24908 12265 24936
rect 11848 24896 11854 24908
rect 12253 24905 12265 24908
rect 12299 24905 12311 24939
rect 12894 24936 12900 24948
rect 12855 24908 12900 24936
rect 12253 24899 12311 24905
rect 12894 24896 12900 24908
rect 12952 24896 12958 24948
rect 17678 24936 17684 24948
rect 17639 24908 17684 24936
rect 17678 24896 17684 24908
rect 17736 24896 17742 24948
rect 19429 24939 19487 24945
rect 19429 24905 19441 24939
rect 19475 24936 19487 24939
rect 19610 24936 19616 24948
rect 19475 24908 19616 24936
rect 19475 24905 19487 24908
rect 19429 24899 19487 24905
rect 19610 24896 19616 24908
rect 19668 24896 19674 24948
rect 22186 24936 22192 24948
rect 22147 24908 22192 24936
rect 22186 24896 22192 24908
rect 22244 24936 22250 24948
rect 22244 24908 23244 24936
rect 22244 24896 22250 24908
rect 9401 24871 9459 24877
rect 9401 24868 9413 24871
rect 7392 24840 7512 24868
rect 7944 24840 8248 24868
rect 8312 24840 9413 24868
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24769 1731 24803
rect 3142 24800 3148 24812
rect 3103 24772 3148 24800
rect 1673 24763 1731 24769
rect 1688 24732 1716 24763
rect 3142 24760 3148 24772
rect 3200 24760 3206 24812
rect 3329 24803 3387 24809
rect 3329 24769 3341 24803
rect 3375 24800 3387 24803
rect 4154 24800 4160 24812
rect 3375 24772 4160 24800
rect 3375 24769 3387 24772
rect 3329 24763 3387 24769
rect 4154 24760 4160 24772
rect 4212 24760 4218 24812
rect 5534 24800 5540 24812
rect 5592 24809 5598 24812
rect 5504 24772 5540 24800
rect 5534 24760 5540 24772
rect 5592 24763 5604 24809
rect 5592 24760 5598 24763
rect 5718 24760 5724 24812
rect 5776 24800 5782 24812
rect 5813 24803 5871 24809
rect 5813 24800 5825 24803
rect 5776 24772 5825 24800
rect 5776 24760 5782 24772
rect 5813 24769 5825 24772
rect 5859 24769 5871 24803
rect 7098 24800 7104 24812
rect 7059 24772 7104 24800
rect 5813 24763 5871 24769
rect 7098 24760 7104 24772
rect 7156 24760 7162 24812
rect 7392 24809 7420 24840
rect 7377 24803 7435 24809
rect 7377 24769 7389 24803
rect 7423 24769 7435 24803
rect 7377 24763 7435 24769
rect 7469 24803 7527 24809
rect 7469 24769 7481 24803
rect 7515 24800 7527 24803
rect 7653 24801 7711 24807
rect 7515 24772 7604 24800
rect 7515 24769 7527 24772
rect 7469 24763 7527 24769
rect 3237 24735 3295 24741
rect 3237 24732 3249 24735
rect 1688 24704 3249 24732
rect 3237 24701 3249 24704
rect 3283 24701 3295 24735
rect 3237 24695 3295 24701
rect 7190 24692 7196 24744
rect 7248 24732 7254 24744
rect 7285 24735 7343 24741
rect 7285 24732 7297 24735
rect 7248 24704 7297 24732
rect 7248 24692 7254 24704
rect 7285 24701 7297 24704
rect 7331 24701 7343 24735
rect 7576 24732 7604 24772
rect 7653 24767 7665 24801
rect 7699 24798 7711 24801
rect 7944 24800 7972 24840
rect 8110 24800 8116 24812
rect 7852 24798 7972 24800
rect 7699 24772 7972 24798
rect 8071 24772 8116 24800
rect 7699 24770 7880 24772
rect 7699 24767 7711 24770
rect 7653 24761 7711 24767
rect 8110 24760 8116 24772
rect 8168 24760 8174 24812
rect 8220 24800 8248 24840
rect 9401 24837 9413 24840
rect 9447 24868 9459 24871
rect 9582 24868 9588 24880
rect 9447 24840 9588 24868
rect 9447 24837 9459 24840
rect 9401 24831 9459 24837
rect 9582 24828 9588 24840
rect 9640 24828 9646 24880
rect 15102 24828 15108 24880
rect 15160 24868 15166 24880
rect 15160 24840 15516 24868
rect 15160 24828 15166 24840
rect 8570 24800 8576 24812
rect 8220 24772 8576 24800
rect 8570 24760 8576 24772
rect 8628 24760 8634 24812
rect 8754 24760 8760 24812
rect 8812 24800 8818 24812
rect 9030 24800 9036 24812
rect 8812 24772 9036 24800
rect 8812 24760 8818 24772
rect 9030 24760 9036 24772
rect 9088 24760 9094 24812
rect 9214 24809 9220 24812
rect 9181 24803 9220 24809
rect 9181 24769 9193 24803
rect 9181 24763 9220 24769
rect 9214 24760 9220 24763
rect 9272 24760 9278 24812
rect 9309 24803 9367 24809
rect 9309 24769 9321 24803
rect 9355 24769 9367 24803
rect 9309 24763 9367 24769
rect 8205 24735 8263 24741
rect 8205 24732 8217 24735
rect 7576 24704 8217 24732
rect 7285 24695 7343 24701
rect 8205 24701 8217 24704
rect 8251 24701 8263 24735
rect 9324 24732 9352 24763
rect 9490 24760 9496 24812
rect 9548 24809 9554 24812
rect 9548 24800 9556 24809
rect 10410 24800 10416 24812
rect 9548 24772 9593 24800
rect 10371 24772 10416 24800
rect 9548 24763 9556 24772
rect 9548 24760 9554 24763
rect 10410 24760 10416 24772
rect 10468 24760 10474 24812
rect 10502 24760 10508 24812
rect 10560 24800 10566 24812
rect 10689 24803 10747 24809
rect 10560 24772 10605 24800
rect 10560 24760 10566 24772
rect 10689 24769 10701 24803
rect 10735 24800 10747 24803
rect 10778 24800 10784 24812
rect 10735 24772 10784 24800
rect 10735 24769 10747 24772
rect 10689 24763 10747 24769
rect 10778 24760 10784 24772
rect 10836 24760 10842 24812
rect 11517 24803 11575 24809
rect 11517 24769 11529 24803
rect 11563 24800 11575 24803
rect 11606 24800 11612 24812
rect 11563 24772 11612 24800
rect 11563 24769 11575 24772
rect 11517 24763 11575 24769
rect 11606 24760 11612 24772
rect 11664 24760 11670 24812
rect 11701 24803 11759 24809
rect 11701 24769 11713 24803
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 12069 24803 12127 24809
rect 12069 24769 12081 24803
rect 12115 24800 12127 24803
rect 12618 24800 12624 24812
rect 12115 24772 12624 24800
rect 12115 24769 12127 24772
rect 12069 24763 12127 24769
rect 10318 24732 10324 24744
rect 9324 24704 10324 24732
rect 8205 24695 8263 24701
rect 10318 24692 10324 24704
rect 10376 24732 10382 24744
rect 10597 24735 10655 24741
rect 10597 24732 10609 24735
rect 10376 24704 10609 24732
rect 10376 24692 10382 24704
rect 10597 24701 10609 24704
rect 10643 24701 10655 24735
rect 10597 24695 10655 24701
rect 1486 24664 1492 24676
rect 1447 24636 1492 24664
rect 1486 24624 1492 24636
rect 1544 24624 1550 24676
rect 10686 24624 10692 24676
rect 10744 24664 10750 24676
rect 10873 24667 10931 24673
rect 10873 24664 10885 24667
rect 10744 24636 10885 24664
rect 10744 24624 10750 24636
rect 10873 24633 10885 24636
rect 10919 24633 10931 24667
rect 10873 24627 10931 24633
rect 4433 24599 4491 24605
rect 4433 24565 4445 24599
rect 4479 24596 4491 24599
rect 5810 24596 5816 24608
rect 4479 24568 5816 24596
rect 4479 24565 4491 24568
rect 4433 24559 4491 24565
rect 5810 24556 5816 24568
rect 5868 24556 5874 24608
rect 7466 24556 7472 24608
rect 7524 24596 7530 24608
rect 11716 24596 11744 24763
rect 12618 24760 12624 24772
rect 12676 24760 12682 24812
rect 13998 24760 14004 24812
rect 14056 24809 14062 24812
rect 14056 24800 14068 24809
rect 14274 24800 14280 24812
rect 14056 24772 14101 24800
rect 14235 24772 14280 24800
rect 14056 24763 14068 24772
rect 14056 24760 14062 24763
rect 14274 24760 14280 24772
rect 14332 24760 14338 24812
rect 14366 24760 14372 24812
rect 14424 24800 14430 24812
rect 14737 24803 14795 24809
rect 14737 24800 14749 24803
rect 14424 24772 14749 24800
rect 14424 24760 14430 24772
rect 14737 24769 14749 24772
rect 14783 24769 14795 24803
rect 14737 24763 14795 24769
rect 14826 24760 14832 24812
rect 14884 24800 14890 24812
rect 15381 24803 15439 24809
rect 15381 24800 15393 24803
rect 14884 24772 15393 24800
rect 14884 24760 14890 24772
rect 15381 24769 15393 24772
rect 15427 24769 15439 24803
rect 15488 24800 15516 24840
rect 22002 24828 22008 24880
rect 22060 24868 22066 24880
rect 23216 24877 23244 24908
rect 23017 24871 23075 24877
rect 23017 24868 23029 24871
rect 22060 24840 23029 24868
rect 22060 24828 22066 24840
rect 16669 24803 16727 24809
rect 16669 24800 16681 24803
rect 15488 24772 16681 24800
rect 15381 24763 15439 24769
rect 16669 24769 16681 24772
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 16758 24760 16764 24812
rect 16816 24800 16822 24812
rect 18874 24800 18880 24812
rect 16816 24772 18736 24800
rect 18835 24772 18880 24800
rect 16816 24760 16822 24772
rect 11793 24735 11851 24741
rect 11793 24701 11805 24735
rect 11839 24701 11851 24735
rect 11793 24695 11851 24701
rect 11885 24735 11943 24741
rect 11885 24701 11897 24735
rect 11931 24732 11943 24735
rect 11974 24732 11980 24744
rect 11931 24704 11980 24732
rect 11931 24701 11943 24704
rect 11885 24695 11943 24701
rect 11808 24664 11836 24695
rect 11974 24692 11980 24704
rect 12032 24692 12038 24744
rect 13078 24732 13084 24744
rect 12406 24704 13084 24732
rect 12066 24664 12072 24676
rect 11808 24636 12072 24664
rect 12066 24624 12072 24636
rect 12124 24624 12130 24676
rect 12406 24596 12434 24704
rect 13078 24692 13084 24704
rect 13136 24692 13142 24744
rect 14292 24732 14320 24760
rect 15470 24732 15476 24744
rect 14292 24704 15476 24732
rect 15470 24692 15476 24704
rect 15528 24692 15534 24744
rect 16206 24692 16212 24744
rect 16264 24732 16270 24744
rect 17405 24735 17463 24741
rect 17405 24732 17417 24735
rect 16264 24704 17417 24732
rect 16264 24692 16270 24704
rect 17405 24701 17417 24704
rect 17451 24701 17463 24735
rect 17405 24695 17463 24701
rect 17589 24735 17647 24741
rect 17589 24701 17601 24735
rect 17635 24732 17647 24735
rect 18708 24732 18736 24772
rect 18874 24760 18880 24772
rect 18932 24760 18938 24812
rect 19521 24803 19579 24809
rect 19521 24769 19533 24803
rect 19567 24769 19579 24803
rect 19521 24763 19579 24769
rect 19150 24732 19156 24744
rect 17635 24704 17724 24732
rect 18708 24704 19156 24732
rect 17635 24701 17647 24704
rect 17589 24695 17647 24701
rect 17696 24676 17724 24704
rect 19150 24692 19156 24704
rect 19208 24692 19214 24744
rect 19536 24732 19564 24763
rect 19886 24760 19892 24812
rect 19944 24800 19950 24812
rect 19981 24803 20039 24809
rect 19981 24800 19993 24803
rect 19944 24772 19993 24800
rect 19944 24760 19950 24772
rect 19981 24769 19993 24772
rect 20027 24769 20039 24803
rect 19981 24763 20039 24769
rect 20622 24760 20628 24812
rect 20680 24800 20686 24812
rect 20901 24803 20959 24809
rect 20901 24800 20913 24803
rect 20680 24772 20913 24800
rect 20680 24760 20686 24772
rect 20901 24769 20913 24772
rect 20947 24769 20959 24803
rect 20901 24763 20959 24769
rect 20993 24803 21051 24809
rect 20993 24769 21005 24803
rect 21039 24769 21051 24803
rect 20993 24763 21051 24769
rect 20714 24732 20720 24744
rect 19536 24704 20720 24732
rect 20714 24692 20720 24704
rect 20772 24692 20778 24744
rect 14829 24667 14887 24673
rect 14829 24633 14841 24667
rect 14875 24664 14887 24667
rect 16390 24664 16396 24676
rect 14875 24636 16396 24664
rect 14875 24633 14887 24636
rect 14829 24627 14887 24633
rect 16390 24624 16396 24636
rect 16448 24624 16454 24676
rect 17678 24624 17684 24676
rect 17736 24624 17742 24676
rect 21008 24664 21036 24763
rect 21450 24692 21456 24744
rect 21508 24732 21514 24744
rect 21910 24732 21916 24744
rect 21508 24704 21916 24732
rect 21508 24692 21514 24704
rect 21910 24692 21916 24704
rect 21968 24732 21974 24744
rect 22388 24741 22416 24840
rect 23017 24837 23029 24840
rect 23063 24837 23075 24871
rect 23017 24831 23075 24837
rect 23201 24871 23259 24877
rect 23201 24837 23213 24871
rect 23247 24837 23259 24871
rect 23201 24831 23259 24837
rect 22281 24735 22339 24741
rect 22281 24732 22293 24735
rect 21968 24704 22293 24732
rect 21968 24692 21974 24704
rect 22281 24701 22293 24704
rect 22327 24701 22339 24735
rect 22281 24695 22339 24701
rect 22373 24735 22431 24741
rect 22373 24701 22385 24735
rect 22419 24701 22431 24735
rect 22373 24695 22431 24701
rect 22738 24664 22744 24676
rect 21008 24636 22744 24664
rect 22738 24624 22744 24636
rect 22796 24624 22802 24676
rect 7524 24568 12434 24596
rect 7524 24556 7530 24568
rect 15286 24556 15292 24608
rect 15344 24596 15350 24608
rect 15473 24599 15531 24605
rect 15473 24596 15485 24599
rect 15344 24568 15485 24596
rect 15344 24556 15350 24568
rect 15473 24565 15485 24568
rect 15519 24565 15531 24599
rect 15473 24559 15531 24565
rect 16574 24556 16580 24608
rect 16632 24596 16638 24608
rect 16761 24599 16819 24605
rect 16761 24596 16773 24599
rect 16632 24568 16773 24596
rect 16632 24556 16638 24568
rect 16761 24565 16773 24568
rect 16807 24565 16819 24599
rect 16761 24559 16819 24565
rect 17770 24556 17776 24608
rect 17828 24596 17834 24608
rect 18049 24599 18107 24605
rect 18049 24596 18061 24599
rect 17828 24568 18061 24596
rect 17828 24556 17834 24568
rect 18049 24565 18061 24568
rect 18095 24565 18107 24599
rect 18049 24559 18107 24565
rect 18598 24556 18604 24608
rect 18656 24596 18662 24608
rect 18693 24599 18751 24605
rect 18693 24596 18705 24599
rect 18656 24568 18705 24596
rect 18656 24556 18662 24568
rect 18693 24565 18705 24568
rect 18739 24565 18751 24599
rect 18693 24559 18751 24565
rect 19978 24556 19984 24608
rect 20036 24596 20042 24608
rect 20073 24599 20131 24605
rect 20073 24596 20085 24599
rect 20036 24568 20085 24596
rect 20036 24556 20042 24568
rect 20073 24565 20085 24568
rect 20119 24565 20131 24599
rect 20073 24559 20131 24565
rect 21082 24556 21088 24608
rect 21140 24596 21146 24608
rect 21821 24599 21879 24605
rect 21821 24596 21833 24599
rect 21140 24568 21833 24596
rect 21140 24556 21146 24568
rect 21821 24565 21833 24568
rect 21867 24565 21879 24599
rect 21821 24559 21879 24565
rect 23385 24599 23443 24605
rect 23385 24565 23397 24599
rect 23431 24596 23443 24599
rect 23750 24596 23756 24608
rect 23431 24568 23756 24596
rect 23431 24565 23443 24568
rect 23385 24559 23443 24565
rect 23750 24556 23756 24568
rect 23808 24556 23814 24608
rect 1104 24506 30820 24528
rect 1104 24454 5915 24506
rect 5967 24454 5979 24506
rect 6031 24454 6043 24506
rect 6095 24454 6107 24506
rect 6159 24454 6171 24506
rect 6223 24454 15846 24506
rect 15898 24454 15910 24506
rect 15962 24454 15974 24506
rect 16026 24454 16038 24506
rect 16090 24454 16102 24506
rect 16154 24454 25776 24506
rect 25828 24454 25840 24506
rect 25892 24454 25904 24506
rect 25956 24454 25968 24506
rect 26020 24454 26032 24506
rect 26084 24454 30820 24506
rect 1104 24432 30820 24454
rect 4430 24352 4436 24404
rect 4488 24392 4494 24404
rect 4706 24392 4712 24404
rect 4488 24364 4712 24392
rect 4488 24352 4494 24364
rect 4706 24352 4712 24364
rect 4764 24352 4770 24404
rect 5534 24352 5540 24404
rect 5592 24392 5598 24404
rect 5721 24395 5779 24401
rect 5721 24392 5733 24395
rect 5592 24364 5733 24392
rect 5592 24352 5598 24364
rect 5721 24361 5733 24364
rect 5767 24361 5779 24395
rect 5721 24355 5779 24361
rect 7098 24352 7104 24404
rect 7156 24392 7162 24404
rect 8205 24395 8263 24401
rect 8205 24392 8217 24395
rect 7156 24364 8217 24392
rect 7156 24352 7162 24364
rect 8205 24361 8217 24364
rect 8251 24361 8263 24395
rect 8205 24355 8263 24361
rect 8570 24352 8576 24404
rect 8628 24392 8634 24404
rect 9493 24395 9551 24401
rect 9493 24392 9505 24395
rect 8628 24364 9505 24392
rect 8628 24352 8634 24364
rect 9493 24361 9505 24364
rect 9539 24361 9551 24395
rect 9493 24355 9551 24361
rect 9674 24352 9680 24404
rect 9732 24392 9738 24404
rect 9953 24395 10011 24401
rect 9953 24392 9965 24395
rect 9732 24364 9965 24392
rect 9732 24352 9738 24364
rect 9953 24361 9965 24364
rect 9999 24361 10011 24395
rect 13173 24395 13231 24401
rect 13173 24392 13185 24395
rect 9953 24355 10011 24361
rect 10520 24364 13185 24392
rect 4724 24324 4752 24352
rect 6086 24324 6092 24336
rect 4724 24296 6092 24324
rect 6086 24284 6092 24296
rect 6144 24284 6150 24336
rect 3142 24256 3148 24268
rect 3055 24228 3148 24256
rect 3068 24197 3096 24228
rect 3142 24216 3148 24228
rect 3200 24256 3206 24268
rect 3200 24228 3924 24256
rect 3200 24216 3206 24228
rect 1673 24191 1731 24197
rect 1673 24157 1685 24191
rect 1719 24157 1731 24191
rect 1673 24151 1731 24157
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24157 3111 24191
rect 3053 24151 3111 24157
rect 3237 24191 3295 24197
rect 3237 24157 3249 24191
rect 3283 24157 3295 24191
rect 3786 24188 3792 24200
rect 3747 24160 3792 24188
rect 3237 24151 3295 24157
rect 1688 24120 1716 24151
rect 3145 24123 3203 24129
rect 3145 24120 3157 24123
rect 1688 24092 3157 24120
rect 3145 24089 3157 24092
rect 3191 24089 3203 24123
rect 3145 24083 3203 24089
rect 1486 24052 1492 24064
rect 1447 24024 1492 24052
rect 1486 24012 1492 24024
rect 1544 24012 1550 24064
rect 3252 24052 3280 24151
rect 3786 24148 3792 24160
rect 3844 24148 3850 24200
rect 3896 24188 3924 24228
rect 6178 24216 6184 24268
rect 6236 24256 6242 24268
rect 6730 24256 6736 24268
rect 6236 24228 6281 24256
rect 6380 24228 6736 24256
rect 6236 24216 6242 24228
rect 5166 24188 5172 24200
rect 3896 24160 5172 24188
rect 5166 24148 5172 24160
rect 5224 24148 5230 24200
rect 5810 24148 5816 24200
rect 5868 24188 5874 24200
rect 5905 24191 5963 24197
rect 5905 24188 5917 24191
rect 5868 24160 5917 24188
rect 5868 24148 5874 24160
rect 5905 24157 5917 24160
rect 5951 24157 5963 24191
rect 6086 24188 6092 24200
rect 6047 24160 6092 24188
rect 5905 24151 5963 24157
rect 6086 24148 6092 24160
rect 6144 24148 6150 24200
rect 6273 24191 6331 24197
rect 6273 24157 6285 24191
rect 6319 24188 6331 24191
rect 6380 24188 6408 24228
rect 6730 24216 6736 24228
rect 6788 24216 6794 24268
rect 7374 24216 7380 24268
rect 7432 24256 7438 24268
rect 7469 24259 7527 24265
rect 7469 24256 7481 24259
rect 7432 24228 7481 24256
rect 7432 24216 7438 24228
rect 7469 24225 7481 24228
rect 7515 24256 7527 24259
rect 7515 24228 7696 24256
rect 7515 24225 7527 24228
rect 7469 24219 7527 24225
rect 7668 24200 7696 24228
rect 8202 24216 8208 24268
rect 8260 24256 8266 24268
rect 9033 24259 9091 24265
rect 9033 24256 9045 24259
rect 8260 24228 9045 24256
rect 8260 24216 8266 24228
rect 9033 24225 9045 24228
rect 9079 24256 9091 24259
rect 10413 24259 10471 24265
rect 10413 24256 10425 24259
rect 9079 24228 10425 24256
rect 9079 24225 9091 24228
rect 9033 24219 9091 24225
rect 10413 24225 10425 24228
rect 10459 24225 10471 24259
rect 10413 24219 10471 24225
rect 6319 24160 6408 24188
rect 6457 24191 6515 24197
rect 6319 24157 6331 24160
rect 6273 24151 6331 24157
rect 6457 24157 6469 24191
rect 6503 24188 6515 24191
rect 6546 24188 6552 24200
rect 6503 24160 6552 24188
rect 6503 24157 6515 24160
rect 6457 24151 6515 24157
rect 6546 24148 6552 24160
rect 6604 24148 6610 24200
rect 7285 24191 7343 24197
rect 7285 24157 7297 24191
rect 7331 24188 7343 24191
rect 7558 24188 7564 24200
rect 7331 24160 7564 24188
rect 7331 24157 7343 24160
rect 7285 24151 7343 24157
rect 7558 24148 7564 24160
rect 7616 24148 7622 24200
rect 7650 24148 7656 24200
rect 7708 24148 7714 24200
rect 8297 24191 8355 24197
rect 8297 24157 8309 24191
rect 8343 24157 8355 24191
rect 8938 24188 8944 24200
rect 8899 24160 8944 24188
rect 8297 24151 8355 24157
rect 4062 24129 4068 24132
rect 4056 24083 4068 24129
rect 4120 24120 4126 24132
rect 4120 24092 4156 24120
rect 4264 24092 6960 24120
rect 4062 24080 4068 24083
rect 4120 24080 4126 24092
rect 4264 24052 4292 24092
rect 3252 24024 4292 24052
rect 4338 24012 4344 24064
rect 4396 24052 4402 24064
rect 5169 24055 5227 24061
rect 5169 24052 5181 24055
rect 4396 24024 5181 24052
rect 4396 24012 4402 24024
rect 5169 24021 5181 24024
rect 5215 24052 5227 24055
rect 6270 24052 6276 24064
rect 5215 24024 6276 24052
rect 5215 24021 5227 24024
rect 5169 24015 5227 24021
rect 6270 24012 6276 24024
rect 6328 24012 6334 24064
rect 6932 24061 6960 24092
rect 7190 24080 7196 24132
rect 7248 24120 7254 24132
rect 7926 24120 7932 24132
rect 7248 24092 7932 24120
rect 7248 24080 7254 24092
rect 7926 24080 7932 24092
rect 7984 24080 7990 24132
rect 8312 24120 8340 24151
rect 8938 24148 8944 24160
rect 8996 24148 9002 24200
rect 9122 24148 9128 24200
rect 9180 24188 9186 24200
rect 9217 24191 9275 24197
rect 9217 24188 9229 24191
rect 9180 24160 9229 24188
rect 9180 24148 9186 24160
rect 9217 24157 9229 24160
rect 9263 24157 9275 24191
rect 9217 24151 9275 24157
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24188 9367 24191
rect 9858 24188 9864 24200
rect 9355 24160 9864 24188
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 9858 24148 9864 24160
rect 9916 24148 9922 24200
rect 10134 24188 10140 24200
rect 10095 24160 10140 24188
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 10520 24197 10548 24364
rect 13173 24361 13185 24364
rect 13219 24361 13231 24395
rect 13173 24355 13231 24361
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 19702 24392 19708 24404
rect 15519 24364 19708 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 19702 24352 19708 24364
rect 19760 24352 19766 24404
rect 19794 24352 19800 24404
rect 19852 24392 19858 24404
rect 19889 24395 19947 24401
rect 19889 24392 19901 24395
rect 19852 24364 19901 24392
rect 19852 24352 19858 24364
rect 19889 24361 19901 24364
rect 19935 24361 19947 24395
rect 19889 24355 19947 24361
rect 20073 24395 20131 24401
rect 20073 24361 20085 24395
rect 20119 24361 20131 24395
rect 20073 24355 20131 24361
rect 11057 24327 11115 24333
rect 11057 24293 11069 24327
rect 11103 24324 11115 24327
rect 11238 24324 11244 24336
rect 11103 24296 11244 24324
rect 11103 24293 11115 24296
rect 11057 24287 11115 24293
rect 11238 24284 11244 24296
rect 11296 24284 11302 24336
rect 12250 24284 12256 24336
rect 12308 24284 12314 24336
rect 14366 24284 14372 24336
rect 14424 24284 14430 24336
rect 16574 24324 16580 24336
rect 15212 24296 16580 24324
rect 12161 24259 12219 24265
rect 12161 24225 12173 24259
rect 12207 24256 12219 24259
rect 12268 24256 12296 24284
rect 14384 24256 14412 24284
rect 15010 24256 15016 24268
rect 12207 24228 12296 24256
rect 12452 24228 14412 24256
rect 14844 24228 15016 24256
rect 12207 24225 12219 24228
rect 12161 24219 12219 24225
rect 10229 24191 10287 24197
rect 10229 24157 10241 24191
rect 10275 24188 10287 24191
rect 10505 24191 10563 24197
rect 10275 24160 10364 24188
rect 10275 24157 10287 24160
rect 10229 24151 10287 24157
rect 8570 24120 8576 24132
rect 8312 24092 8576 24120
rect 8570 24080 8576 24092
rect 8628 24120 8634 24132
rect 9766 24120 9772 24132
rect 8628 24092 9772 24120
rect 8628 24080 8634 24092
rect 9766 24080 9772 24092
rect 9824 24080 9830 24132
rect 6917 24055 6975 24061
rect 6917 24021 6929 24055
rect 6963 24021 6975 24055
rect 6917 24015 6975 24021
rect 7374 24012 7380 24064
rect 7432 24052 7438 24064
rect 7432 24024 7477 24052
rect 7432 24012 7438 24024
rect 9122 24012 9128 24064
rect 9180 24052 9186 24064
rect 9306 24052 9312 24064
rect 9180 24024 9312 24052
rect 9180 24012 9186 24024
rect 9306 24012 9312 24024
rect 9364 24052 9370 24064
rect 10336 24052 10364 24160
rect 10505 24157 10517 24191
rect 10551 24157 10563 24191
rect 10505 24151 10563 24157
rect 11149 24191 11207 24197
rect 11149 24157 11161 24191
rect 11195 24188 11207 24191
rect 11238 24188 11244 24200
rect 11195 24160 11244 24188
rect 11195 24157 11207 24160
rect 11149 24151 11207 24157
rect 11238 24148 11244 24160
rect 11296 24188 11302 24200
rect 11422 24188 11428 24200
rect 11296 24160 11428 24188
rect 11296 24148 11302 24160
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 11514 24148 11520 24200
rect 11572 24188 11578 24200
rect 11698 24188 11704 24200
rect 11572 24160 11704 24188
rect 11572 24148 11578 24160
rect 11698 24148 11704 24160
rect 11756 24188 11762 24200
rect 11885 24191 11943 24197
rect 11885 24188 11897 24191
rect 11756 24160 11897 24188
rect 11756 24148 11762 24160
rect 11885 24157 11897 24160
rect 11931 24157 11943 24191
rect 11885 24151 11943 24157
rect 12069 24191 12127 24197
rect 12069 24157 12081 24191
rect 12115 24157 12127 24191
rect 12069 24151 12127 24157
rect 12253 24191 12311 24197
rect 12253 24157 12265 24191
rect 12299 24188 12311 24191
rect 12342 24188 12348 24200
rect 12299 24160 12348 24188
rect 12299 24157 12311 24160
rect 12253 24151 12311 24157
rect 10686 24080 10692 24132
rect 10744 24120 10750 24132
rect 12084 24120 12112 24151
rect 12342 24148 12348 24160
rect 12400 24148 12406 24200
rect 12452 24197 12480 24228
rect 12437 24191 12495 24197
rect 12437 24157 12449 24191
rect 12483 24157 12495 24191
rect 13078 24188 13084 24200
rect 13039 24160 13084 24188
rect 12437 24151 12495 24157
rect 13078 24148 13084 24160
rect 13136 24148 13142 24200
rect 13538 24148 13544 24200
rect 13596 24188 13602 24200
rect 14185 24191 14243 24197
rect 14185 24188 14197 24191
rect 13596 24160 14197 24188
rect 13596 24148 13602 24160
rect 14185 24157 14197 24160
rect 14231 24157 14243 24191
rect 14185 24151 14243 24157
rect 14369 24191 14427 24197
rect 14369 24157 14381 24191
rect 14415 24188 14427 24191
rect 14550 24188 14556 24200
rect 14415 24160 14556 24188
rect 14415 24157 14427 24160
rect 14369 24151 14427 24157
rect 14550 24148 14556 24160
rect 14608 24148 14614 24200
rect 14844 24197 14872 24228
rect 15010 24216 15016 24228
rect 15068 24216 15074 24268
rect 14829 24191 14887 24197
rect 14829 24157 14841 24191
rect 14875 24157 14887 24191
rect 14829 24151 14887 24157
rect 14922 24191 14980 24197
rect 14922 24157 14934 24191
rect 14968 24157 14980 24191
rect 15102 24188 15108 24200
rect 15063 24160 15108 24188
rect 14922 24151 14980 24157
rect 10744 24092 12112 24120
rect 14936 24120 14964 24151
rect 15102 24148 15108 24160
rect 15160 24148 15166 24200
rect 15212 24197 15240 24296
rect 16574 24284 16580 24296
rect 16632 24284 16638 24336
rect 17604 24296 17908 24324
rect 16301 24259 16359 24265
rect 16301 24225 16313 24259
rect 16347 24256 16359 24259
rect 16758 24256 16764 24268
rect 16347 24228 16764 24256
rect 16347 24225 16359 24228
rect 16301 24219 16359 24225
rect 16758 24216 16764 24228
rect 16816 24216 16822 24268
rect 17604 24265 17632 24296
rect 17589 24259 17647 24265
rect 17589 24225 17601 24259
rect 17635 24225 17647 24259
rect 17770 24256 17776 24268
rect 17731 24228 17776 24256
rect 17589 24219 17647 24225
rect 17770 24216 17776 24228
rect 17828 24216 17834 24268
rect 17880 24256 17908 24296
rect 19334 24284 19340 24336
rect 19392 24324 19398 24336
rect 20088 24324 20116 24355
rect 19392 24296 20116 24324
rect 19392 24284 19398 24296
rect 21910 24284 21916 24336
rect 21968 24324 21974 24336
rect 22833 24327 22891 24333
rect 22833 24324 22845 24327
rect 21968 24296 22845 24324
rect 21968 24284 21974 24296
rect 22833 24293 22845 24296
rect 22879 24293 22891 24327
rect 22833 24287 22891 24293
rect 19978 24256 19984 24268
rect 17880 24228 19984 24256
rect 19978 24216 19984 24228
rect 20036 24216 20042 24268
rect 20165 24259 20223 24265
rect 20165 24225 20177 24259
rect 20211 24256 20223 24259
rect 20530 24256 20536 24268
rect 20211 24228 20536 24256
rect 20211 24225 20223 24228
rect 20165 24219 20223 24225
rect 15197 24191 15255 24197
rect 15197 24157 15209 24191
rect 15243 24157 15255 24191
rect 15197 24151 15255 24157
rect 15286 24148 15292 24200
rect 15344 24197 15350 24200
rect 15344 24188 15352 24197
rect 15344 24160 15389 24188
rect 15344 24151 15352 24160
rect 15344 24148 15350 24151
rect 15746 24148 15752 24200
rect 15804 24188 15810 24200
rect 16025 24191 16083 24197
rect 16025 24188 16037 24191
rect 15804 24160 16037 24188
rect 15804 24148 15810 24160
rect 16025 24157 16037 24160
rect 16071 24157 16083 24191
rect 16025 24151 16083 24157
rect 16114 24148 16120 24200
rect 16172 24188 16178 24200
rect 16209 24191 16267 24197
rect 16209 24188 16221 24191
rect 16172 24160 16221 24188
rect 16172 24148 16178 24160
rect 16209 24157 16221 24160
rect 16255 24157 16267 24191
rect 16209 24151 16267 24157
rect 16393 24191 16451 24197
rect 16393 24157 16405 24191
rect 16439 24157 16451 24191
rect 16574 24188 16580 24200
rect 16535 24160 16580 24188
rect 16393 24151 16451 24157
rect 15378 24120 15384 24132
rect 14936 24092 15384 24120
rect 10744 24080 10750 24092
rect 15378 24080 15384 24092
rect 15436 24080 15442 24132
rect 16408 24120 16436 24151
rect 16574 24148 16580 24160
rect 16632 24148 16638 24200
rect 17126 24188 17132 24200
rect 16684 24160 17132 24188
rect 16684 24120 16712 24160
rect 17126 24148 17132 24160
rect 17184 24188 17190 24200
rect 18782 24188 18788 24200
rect 17184 24160 18788 24188
rect 17184 24148 17190 24160
rect 18782 24148 18788 24160
rect 18840 24148 18846 24200
rect 19150 24148 19156 24200
rect 19208 24188 19214 24200
rect 19245 24191 19303 24197
rect 19245 24188 19257 24191
rect 19208 24160 19257 24188
rect 19208 24148 19214 24160
rect 19245 24157 19257 24160
rect 19291 24157 19303 24191
rect 19245 24151 19303 24157
rect 19610 24148 19616 24200
rect 19668 24188 19674 24200
rect 20180 24188 20208 24219
rect 20530 24216 20536 24228
rect 20588 24216 20594 24268
rect 21082 24256 21088 24268
rect 21043 24228 21088 24256
rect 21082 24216 21088 24228
rect 21140 24216 21146 24268
rect 19668 24160 20208 24188
rect 20257 24191 20315 24197
rect 19668 24148 19674 24160
rect 20257 24157 20269 24191
rect 20303 24188 20315 24191
rect 20622 24188 20628 24200
rect 20303 24160 20628 24188
rect 20303 24157 20315 24160
rect 20257 24151 20315 24157
rect 20622 24148 20628 24160
rect 20680 24148 20686 24200
rect 20993 24191 21051 24197
rect 20993 24157 21005 24191
rect 21039 24188 21051 24191
rect 21266 24188 21272 24200
rect 21039 24160 21272 24188
rect 21039 24157 21051 24160
rect 20993 24151 21051 24157
rect 21266 24148 21272 24160
rect 21324 24148 21330 24200
rect 21545 24191 21603 24197
rect 21545 24157 21557 24191
rect 21591 24188 21603 24191
rect 21591 24160 22324 24188
rect 21591 24157 21603 24160
rect 21545 24151 21603 24157
rect 16408 24092 16712 24120
rect 17865 24123 17923 24129
rect 17865 24089 17877 24123
rect 17911 24120 17923 24123
rect 19426 24120 19432 24132
rect 17911 24092 19432 24120
rect 17911 24089 17923 24092
rect 17865 24083 17923 24089
rect 19426 24080 19432 24092
rect 19484 24080 19490 24132
rect 20530 24080 20536 24132
rect 20588 24120 20594 24132
rect 22002 24120 22008 24132
rect 20588 24092 21496 24120
rect 21963 24092 22008 24120
rect 20588 24080 20594 24092
rect 12618 24052 12624 24064
rect 9364 24024 10364 24052
rect 12579 24024 12624 24052
rect 9364 24012 9370 24024
rect 12618 24012 12624 24024
rect 12676 24012 12682 24064
rect 14277 24055 14335 24061
rect 14277 24021 14289 24055
rect 14323 24052 14335 24055
rect 14734 24052 14740 24064
rect 14323 24024 14740 24052
rect 14323 24021 14335 24024
rect 14277 24015 14335 24021
rect 14734 24012 14740 24024
rect 14792 24012 14798 24064
rect 16666 24012 16672 24064
rect 16724 24052 16730 24064
rect 16761 24055 16819 24061
rect 16761 24052 16773 24055
rect 16724 24024 16773 24052
rect 16724 24012 16730 24024
rect 16761 24021 16773 24024
rect 16807 24021 16819 24055
rect 16761 24015 16819 24021
rect 18233 24055 18291 24061
rect 18233 24021 18245 24055
rect 18279 24052 18291 24055
rect 18782 24052 18788 24064
rect 18279 24024 18788 24052
rect 18279 24021 18291 24024
rect 18233 24015 18291 24021
rect 18782 24012 18788 24024
rect 18840 24012 18846 24064
rect 19334 24052 19340 24064
rect 19295 24024 19340 24052
rect 19334 24012 19340 24024
rect 19392 24012 19398 24064
rect 19702 24012 19708 24064
rect 19760 24052 19766 24064
rect 20622 24052 20628 24064
rect 19760 24024 20628 24052
rect 19760 24012 19766 24024
rect 20622 24012 20628 24024
rect 20680 24012 20686 24064
rect 21358 24052 21364 24064
rect 21319 24024 21364 24052
rect 21358 24012 21364 24024
rect 21416 24012 21422 24064
rect 21468 24052 21496 24092
rect 22002 24080 22008 24092
rect 22060 24080 22066 24132
rect 22094 24080 22100 24132
rect 22152 24120 22158 24132
rect 22189 24123 22247 24129
rect 22189 24120 22201 24123
rect 22152 24092 22201 24120
rect 22152 24080 22158 24092
rect 22189 24089 22201 24092
rect 22235 24089 22247 24123
rect 22296 24120 22324 24160
rect 22922 24148 22928 24200
rect 22980 24188 22986 24200
rect 23017 24191 23075 24197
rect 23017 24188 23029 24191
rect 22980 24160 23029 24188
rect 22980 24148 22986 24160
rect 23017 24157 23029 24160
rect 23063 24157 23075 24191
rect 23750 24188 23756 24200
rect 23711 24160 23756 24188
rect 23017 24151 23075 24157
rect 23750 24148 23756 24160
rect 23808 24148 23814 24200
rect 29825 24191 29883 24197
rect 29825 24157 29837 24191
rect 29871 24188 29883 24191
rect 29914 24188 29920 24200
rect 29871 24160 29920 24188
rect 29871 24157 29883 24160
rect 29825 24151 29883 24157
rect 29914 24148 29920 24160
rect 29972 24148 29978 24200
rect 22296 24092 23152 24120
rect 22189 24083 22247 24089
rect 22112 24052 22140 24080
rect 23124 24064 23152 24092
rect 22370 24052 22376 24064
rect 21468 24024 22140 24052
rect 22331 24024 22376 24052
rect 22370 24012 22376 24024
rect 22428 24012 22434 24064
rect 23106 24012 23112 24064
rect 23164 24052 23170 24064
rect 23661 24055 23719 24061
rect 23661 24052 23673 24055
rect 23164 24024 23673 24052
rect 23164 24012 23170 24024
rect 23661 24021 23673 24024
rect 23707 24021 23719 24055
rect 30006 24052 30012 24064
rect 29967 24024 30012 24052
rect 23661 24015 23719 24021
rect 30006 24012 30012 24024
rect 30064 24012 30070 24064
rect 1104 23962 30820 23984
rect 1104 23910 10880 23962
rect 10932 23910 10944 23962
rect 10996 23910 11008 23962
rect 11060 23910 11072 23962
rect 11124 23910 11136 23962
rect 11188 23910 20811 23962
rect 20863 23910 20875 23962
rect 20927 23910 20939 23962
rect 20991 23910 21003 23962
rect 21055 23910 21067 23962
rect 21119 23910 30820 23962
rect 1104 23888 30820 23910
rect 3973 23851 4031 23857
rect 3973 23817 3985 23851
rect 4019 23848 4031 23851
rect 4062 23848 4068 23860
rect 4019 23820 4068 23848
rect 4019 23817 4031 23820
rect 3973 23811 4031 23817
rect 4062 23808 4068 23820
rect 4120 23808 4126 23860
rect 6546 23848 6552 23860
rect 5644 23820 6552 23848
rect 3786 23740 3792 23792
rect 3844 23780 3850 23792
rect 5537 23783 5595 23789
rect 5537 23780 5549 23783
rect 3844 23752 5549 23780
rect 3844 23740 3850 23752
rect 5537 23749 5549 23752
rect 5583 23749 5595 23783
rect 5537 23743 5595 23749
rect 4157 23715 4215 23721
rect 4157 23681 4169 23715
rect 4203 23712 4215 23715
rect 4246 23712 4252 23724
rect 4203 23684 4252 23712
rect 4203 23681 4215 23684
rect 4157 23675 4215 23681
rect 4246 23672 4252 23684
rect 4304 23672 4310 23724
rect 4525 23715 4583 23721
rect 4525 23681 4537 23715
rect 4571 23681 4583 23715
rect 4525 23675 4583 23681
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23712 4767 23715
rect 4890 23712 4896 23724
rect 4755 23684 4896 23712
rect 4755 23681 4767 23684
rect 4709 23675 4767 23681
rect 1394 23644 1400 23656
rect 1355 23616 1400 23644
rect 1394 23604 1400 23616
rect 1452 23604 1458 23656
rect 1673 23647 1731 23653
rect 1673 23613 1685 23647
rect 1719 23644 1731 23647
rect 2130 23644 2136 23656
rect 1719 23616 2136 23644
rect 1719 23613 1731 23616
rect 1673 23607 1731 23613
rect 2130 23604 2136 23616
rect 2188 23604 2194 23656
rect 4338 23644 4344 23656
rect 4299 23616 4344 23644
rect 4338 23604 4344 23616
rect 4396 23604 4402 23656
rect 4433 23647 4491 23653
rect 4433 23613 4445 23647
rect 4479 23613 4491 23647
rect 4540 23644 4568 23675
rect 4890 23672 4896 23684
rect 4948 23712 4954 23724
rect 5644 23712 5672 23820
rect 6546 23808 6552 23820
rect 6604 23808 6610 23860
rect 6730 23808 6736 23860
rect 6788 23848 6794 23860
rect 7837 23851 7895 23857
rect 7837 23848 7849 23851
rect 6788 23820 7849 23848
rect 6788 23808 6794 23820
rect 7837 23817 7849 23820
rect 7883 23817 7895 23851
rect 10594 23848 10600 23860
rect 7837 23811 7895 23817
rect 7944 23820 10600 23848
rect 6270 23740 6276 23792
rect 6328 23780 6334 23792
rect 6564 23780 6592 23808
rect 6914 23780 6920 23792
rect 6328 23752 6491 23780
rect 6564 23752 6920 23780
rect 6328 23740 6334 23752
rect 4948 23684 5672 23712
rect 5721 23715 5779 23721
rect 4948 23672 4954 23684
rect 5721 23681 5733 23715
rect 5767 23681 5779 23715
rect 6362 23712 6368 23724
rect 6323 23684 6368 23712
rect 5721 23675 5779 23681
rect 5736 23644 5764 23675
rect 6362 23672 6368 23684
rect 6420 23672 6426 23724
rect 6463 23712 6491 23752
rect 6914 23740 6920 23752
rect 6972 23740 6978 23792
rect 7006 23740 7012 23792
rect 7064 23780 7070 23792
rect 7285 23783 7343 23789
rect 7285 23780 7297 23783
rect 7064 23752 7297 23780
rect 7064 23740 7070 23752
rect 7285 23749 7297 23752
rect 7331 23749 7343 23783
rect 7944 23780 7972 23820
rect 10594 23808 10600 23820
rect 10652 23808 10658 23860
rect 14093 23851 14151 23857
rect 14093 23817 14105 23851
rect 14139 23848 14151 23851
rect 14366 23848 14372 23860
rect 14139 23820 14372 23848
rect 14139 23817 14151 23820
rect 14093 23811 14151 23817
rect 14366 23808 14372 23820
rect 14424 23808 14430 23860
rect 14826 23808 14832 23860
rect 14884 23848 14890 23860
rect 14921 23851 14979 23857
rect 14921 23848 14933 23851
rect 14884 23820 14933 23848
rect 14884 23808 14890 23820
rect 14921 23817 14933 23820
rect 14967 23848 14979 23851
rect 15286 23848 15292 23860
rect 14967 23820 15292 23848
rect 14967 23817 14979 23820
rect 14921 23811 14979 23817
rect 15286 23808 15292 23820
rect 15344 23808 15350 23860
rect 16114 23848 16120 23860
rect 16075 23820 16120 23848
rect 16114 23808 16120 23820
rect 16172 23808 16178 23860
rect 18598 23848 18604 23860
rect 18559 23820 18604 23848
rect 18598 23808 18604 23820
rect 18656 23808 18662 23860
rect 19702 23808 19708 23860
rect 19760 23808 19766 23860
rect 29914 23848 29920 23860
rect 29875 23820 29920 23848
rect 29914 23808 29920 23820
rect 29972 23808 29978 23860
rect 8205 23783 8263 23789
rect 8205 23780 8217 23783
rect 7285 23743 7343 23749
rect 7392 23752 7972 23780
rect 8036 23752 8217 23780
rect 7392 23712 7420 23752
rect 6463 23684 7420 23712
rect 7837 23715 7895 23721
rect 7837 23681 7849 23715
rect 7883 23712 7895 23715
rect 8036 23712 8064 23752
rect 8205 23749 8217 23752
rect 8251 23749 8263 23783
rect 8205 23743 8263 23749
rect 8297 23783 8355 23789
rect 8297 23749 8309 23783
rect 8343 23780 8355 23783
rect 9122 23780 9128 23792
rect 8343 23752 9128 23780
rect 8343 23749 8355 23752
rect 8297 23743 8355 23749
rect 9122 23740 9128 23752
rect 9180 23780 9186 23792
rect 10502 23780 10508 23792
rect 9180 23752 10508 23780
rect 9180 23740 9186 23752
rect 10502 23740 10508 23752
rect 10560 23740 10566 23792
rect 10781 23783 10839 23789
rect 10781 23749 10793 23783
rect 10827 23780 10839 23783
rect 11882 23780 11888 23792
rect 10827 23752 11888 23780
rect 10827 23749 10839 23752
rect 10781 23743 10839 23749
rect 11882 23740 11888 23752
rect 11940 23740 11946 23792
rect 12250 23780 12256 23792
rect 11992 23752 12256 23780
rect 7883 23684 8064 23712
rect 8108 23715 8166 23721
rect 7883 23681 7895 23684
rect 7837 23675 7895 23681
rect 8108 23681 8120 23715
rect 8154 23681 8166 23715
rect 8108 23675 8166 23681
rect 8480 23715 8538 23721
rect 8480 23681 8492 23715
rect 8526 23681 8538 23715
rect 8480 23675 8538 23681
rect 8573 23715 8631 23721
rect 8573 23681 8585 23715
rect 8619 23712 8631 23715
rect 8754 23712 8760 23724
rect 8619 23684 8760 23712
rect 8619 23681 8631 23684
rect 8573 23675 8631 23681
rect 4540 23616 4660 23644
rect 5736 23616 7236 23644
rect 4433 23607 4491 23613
rect 4448 23508 4476 23607
rect 4632 23576 4660 23616
rect 7098 23576 7104 23588
rect 4632 23548 7104 23576
rect 7098 23536 7104 23548
rect 7156 23536 7162 23588
rect 7208 23520 7236 23616
rect 4798 23508 4804 23520
rect 4448 23480 4804 23508
rect 4798 23468 4804 23480
rect 4856 23508 4862 23520
rect 5074 23508 5080 23520
rect 4856 23480 5080 23508
rect 4856 23468 4862 23480
rect 5074 23468 5080 23480
rect 5132 23468 5138 23520
rect 6457 23511 6515 23517
rect 6457 23477 6469 23511
rect 6503 23508 6515 23511
rect 7006 23508 7012 23520
rect 6503 23480 7012 23508
rect 6503 23477 6515 23480
rect 6457 23471 6515 23477
rect 7006 23468 7012 23480
rect 7064 23468 7070 23520
rect 7190 23508 7196 23520
rect 7151 23480 7196 23508
rect 7190 23468 7196 23480
rect 7248 23468 7254 23520
rect 7929 23511 7987 23517
rect 7929 23477 7941 23511
rect 7975 23508 7987 23511
rect 8018 23508 8024 23520
rect 7975 23480 8024 23508
rect 7975 23477 7987 23480
rect 7929 23471 7987 23477
rect 8018 23468 8024 23480
rect 8076 23468 8082 23520
rect 8128 23508 8156 23675
rect 8496 23588 8524 23675
rect 8754 23672 8760 23684
rect 8812 23672 8818 23724
rect 9030 23712 9036 23724
rect 8991 23684 9036 23712
rect 9030 23672 9036 23684
rect 9088 23672 9094 23724
rect 9217 23715 9275 23721
rect 9217 23712 9229 23715
rect 9140 23684 9229 23712
rect 8938 23604 8944 23656
rect 8996 23644 9002 23656
rect 9140 23644 9168 23684
rect 9217 23681 9229 23684
rect 9263 23681 9275 23715
rect 9217 23675 9275 23681
rect 9585 23715 9643 23721
rect 9585 23681 9597 23715
rect 9631 23712 9643 23715
rect 10870 23712 10876 23724
rect 9631 23684 10876 23712
rect 9631 23681 9643 23684
rect 9585 23675 9643 23681
rect 10870 23672 10876 23684
rect 10928 23672 10934 23724
rect 11422 23672 11428 23724
rect 11480 23712 11486 23724
rect 11517 23715 11575 23721
rect 11517 23712 11529 23715
rect 11480 23684 11529 23712
rect 11480 23672 11486 23684
rect 11517 23681 11529 23684
rect 11563 23681 11575 23715
rect 11517 23675 11575 23681
rect 11701 23715 11759 23721
rect 11701 23681 11713 23715
rect 11747 23681 11759 23715
rect 11701 23675 11759 23681
rect 9309 23647 9367 23653
rect 9309 23644 9321 23647
rect 8996 23616 9168 23644
rect 9232 23616 9321 23644
rect 8996 23604 9002 23616
rect 9232 23588 9260 23616
rect 9309 23613 9321 23616
rect 9355 23613 9367 23647
rect 9309 23607 9367 23613
rect 9401 23647 9459 23653
rect 9401 23613 9413 23647
rect 9447 23644 9459 23647
rect 9490 23644 9496 23656
rect 9447 23616 9496 23644
rect 9447 23613 9459 23616
rect 9401 23607 9459 23613
rect 9490 23604 9496 23616
rect 9548 23604 9554 23656
rect 10594 23604 10600 23656
rect 10652 23644 10658 23656
rect 11716 23644 11744 23675
rect 11790 23672 11796 23724
rect 11848 23712 11854 23724
rect 11992 23712 12020 23752
rect 12250 23740 12256 23752
rect 12308 23740 12314 23792
rect 12618 23740 12624 23792
rect 12676 23780 12682 23792
rect 12958 23783 13016 23789
rect 12958 23780 12970 23783
rect 12676 23752 12970 23780
rect 12676 23740 12682 23752
rect 12958 23749 12970 23752
rect 13004 23749 13016 23783
rect 14550 23780 14556 23792
rect 14511 23752 14556 23780
rect 12958 23743 13016 23749
rect 14550 23740 14556 23752
rect 14608 23740 14614 23792
rect 15749 23783 15807 23789
rect 15749 23749 15761 23783
rect 15795 23780 15807 23783
rect 16482 23780 16488 23792
rect 15795 23752 16488 23780
rect 15795 23749 15807 23752
rect 15749 23743 15807 23749
rect 16482 23740 16488 23752
rect 16540 23740 16546 23792
rect 17402 23740 17408 23792
rect 17460 23740 17466 23792
rect 19613 23783 19671 23789
rect 19613 23749 19625 23783
rect 19659 23780 19671 23783
rect 19720 23780 19748 23808
rect 19659 23752 20852 23780
rect 19659 23749 19671 23752
rect 19613 23743 19671 23749
rect 11848 23684 12020 23712
rect 12069 23715 12127 23721
rect 11848 23672 11854 23684
rect 12069 23681 12081 23715
rect 12115 23712 12127 23715
rect 12710 23712 12716 23724
rect 12115 23684 12434 23712
rect 12671 23684 12716 23712
rect 12115 23681 12127 23684
rect 12069 23675 12127 23681
rect 10652 23616 11744 23644
rect 11885 23647 11943 23653
rect 10652 23604 10658 23616
rect 11885 23613 11897 23647
rect 11931 23644 11943 23647
rect 12250 23644 12256 23656
rect 11931 23616 12256 23644
rect 11931 23613 11943 23616
rect 11885 23607 11943 23613
rect 12250 23604 12256 23616
rect 12308 23604 12314 23656
rect 12406 23644 12434 23684
rect 12710 23672 12716 23684
rect 12768 23672 12774 23724
rect 13538 23712 13544 23724
rect 12820 23684 13544 23712
rect 12820 23644 12848 23684
rect 13538 23672 13544 23684
rect 13596 23712 13602 23724
rect 14737 23715 14795 23721
rect 14737 23712 14749 23715
rect 13596 23684 14749 23712
rect 13596 23672 13602 23684
rect 14737 23681 14749 23684
rect 14783 23681 14795 23715
rect 16666 23712 16672 23724
rect 16627 23684 16672 23712
rect 14737 23675 14795 23681
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 17034 23672 17040 23724
rect 17092 23712 17098 23724
rect 17129 23715 17187 23721
rect 17129 23712 17141 23715
rect 17092 23684 17141 23712
rect 17092 23672 17098 23684
rect 17129 23681 17141 23684
rect 17175 23681 17187 23715
rect 17420 23712 17448 23740
rect 17497 23715 17555 23721
rect 17497 23712 17509 23715
rect 17420 23684 17509 23712
rect 17129 23675 17187 23681
rect 17497 23681 17509 23684
rect 17543 23681 17555 23715
rect 18506 23712 18512 23724
rect 18467 23684 18512 23712
rect 17497 23675 17555 23681
rect 18506 23672 18512 23684
rect 18564 23672 18570 23724
rect 19705 23715 19763 23721
rect 19705 23681 19717 23715
rect 19751 23712 19763 23715
rect 19794 23712 19800 23724
rect 19751 23684 19800 23712
rect 19751 23681 19763 23684
rect 19705 23675 19763 23681
rect 19794 23672 19800 23684
rect 19852 23672 19858 23724
rect 19886 23672 19892 23724
rect 19944 23712 19950 23724
rect 20254 23712 20260 23724
rect 19944 23684 20260 23712
rect 19944 23672 19950 23684
rect 20254 23672 20260 23684
rect 20312 23712 20318 23724
rect 20395 23715 20453 23721
rect 20395 23712 20407 23715
rect 20312 23684 20407 23712
rect 20312 23672 20318 23684
rect 20395 23681 20407 23684
rect 20441 23681 20453 23715
rect 20527 23712 20533 23724
rect 20488 23684 20533 23712
rect 20395 23675 20453 23681
rect 20527 23672 20533 23684
rect 20585 23672 20591 23724
rect 20824 23721 20852 23752
rect 20625 23715 20683 23721
rect 20625 23681 20637 23715
rect 20671 23681 20683 23715
rect 20625 23675 20683 23681
rect 20809 23715 20867 23721
rect 20809 23681 20821 23715
rect 20855 23681 20867 23715
rect 20809 23675 20867 23681
rect 22189 23715 22247 23721
rect 22189 23681 22201 23715
rect 22235 23712 22247 23715
rect 22370 23712 22376 23724
rect 22235 23684 22376 23712
rect 22235 23681 22247 23684
rect 22189 23675 22247 23681
rect 12406 23616 12848 23644
rect 15102 23604 15108 23656
rect 15160 23644 15166 23656
rect 15473 23647 15531 23653
rect 15473 23644 15485 23647
rect 15160 23616 15485 23644
rect 15160 23604 15166 23616
rect 15473 23613 15485 23616
rect 15519 23613 15531 23647
rect 15654 23644 15660 23656
rect 15615 23616 15660 23644
rect 15473 23607 15531 23613
rect 15654 23604 15660 23616
rect 15712 23604 15718 23656
rect 17218 23644 17224 23656
rect 17179 23616 17224 23644
rect 17218 23604 17224 23616
rect 17276 23604 17282 23656
rect 17402 23644 17408 23656
rect 17363 23616 17408 23644
rect 17402 23604 17408 23616
rect 17460 23604 17466 23656
rect 18598 23604 18604 23656
rect 18656 23644 18662 23656
rect 18693 23647 18751 23653
rect 18693 23644 18705 23647
rect 18656 23616 18705 23644
rect 18656 23604 18662 23616
rect 18693 23613 18705 23616
rect 18739 23644 18751 23647
rect 19518 23644 19524 23656
rect 18739 23616 19524 23644
rect 18739 23613 18751 23616
rect 18693 23607 18751 23613
rect 19518 23604 19524 23616
rect 19576 23604 19582 23656
rect 19610 23604 19616 23656
rect 19668 23604 19674 23656
rect 8478 23536 8484 23588
rect 8536 23536 8542 23588
rect 9214 23536 9220 23588
rect 9272 23536 9278 23588
rect 16850 23536 16856 23588
rect 16908 23576 16914 23588
rect 19628 23576 19656 23604
rect 16908 23548 19656 23576
rect 16908 23536 16914 23548
rect 20254 23536 20260 23588
rect 20312 23576 20318 23588
rect 20640 23576 20668 23675
rect 22370 23672 22376 23684
rect 22428 23672 22434 23724
rect 23477 23715 23535 23721
rect 23477 23681 23489 23715
rect 23523 23681 23535 23715
rect 30098 23712 30104 23724
rect 30059 23684 30104 23712
rect 23477 23675 23535 23681
rect 22462 23644 22468 23656
rect 22423 23616 22468 23644
rect 22462 23604 22468 23616
rect 22520 23604 22526 23656
rect 20312 23548 20668 23576
rect 20312 23536 20318 23548
rect 22370 23536 22376 23588
rect 22428 23576 22434 23588
rect 23492 23576 23520 23675
rect 30098 23672 30104 23684
rect 30156 23672 30162 23724
rect 22428 23548 23520 23576
rect 22428 23536 22434 23548
rect 8386 23508 8392 23520
rect 8128 23480 8392 23508
rect 8386 23468 8392 23480
rect 8444 23468 8450 23520
rect 9030 23468 9036 23520
rect 9088 23508 9094 23520
rect 9582 23508 9588 23520
rect 9088 23480 9588 23508
rect 9088 23468 9094 23480
rect 9582 23468 9588 23480
rect 9640 23468 9646 23520
rect 9769 23511 9827 23517
rect 9769 23477 9781 23511
rect 9815 23508 9827 23511
rect 9858 23508 9864 23520
rect 9815 23480 9864 23508
rect 9815 23477 9827 23480
rect 9769 23471 9827 23477
rect 9858 23468 9864 23480
rect 9916 23468 9922 23520
rect 10778 23468 10784 23520
rect 10836 23508 10842 23520
rect 10873 23511 10931 23517
rect 10873 23508 10885 23511
rect 10836 23480 10885 23508
rect 10836 23468 10842 23480
rect 10873 23477 10885 23480
rect 10919 23477 10931 23511
rect 10873 23471 10931 23477
rect 12253 23511 12311 23517
rect 12253 23477 12265 23511
rect 12299 23508 12311 23511
rect 12526 23508 12532 23520
rect 12299 23480 12532 23508
rect 12299 23477 12311 23480
rect 12253 23471 12311 23477
rect 12526 23468 12532 23480
rect 12584 23468 12590 23520
rect 16298 23468 16304 23520
rect 16356 23508 16362 23520
rect 16761 23511 16819 23517
rect 16761 23508 16773 23511
rect 16356 23480 16773 23508
rect 16356 23468 16362 23480
rect 16761 23477 16773 23480
rect 16807 23477 16819 23511
rect 16761 23471 16819 23477
rect 16942 23468 16948 23520
rect 17000 23508 17006 23520
rect 17218 23508 17224 23520
rect 17000 23480 17224 23508
rect 17000 23468 17006 23480
rect 17218 23468 17224 23480
rect 17276 23468 17282 23520
rect 18138 23508 18144 23520
rect 18099 23480 18144 23508
rect 18138 23468 18144 23480
rect 18196 23468 18202 23520
rect 20162 23508 20168 23520
rect 20123 23480 20168 23508
rect 20162 23468 20168 23480
rect 20220 23468 20226 23520
rect 20714 23468 20720 23520
rect 20772 23508 20778 23520
rect 21542 23508 21548 23520
rect 20772 23480 21548 23508
rect 20772 23468 20778 23480
rect 21542 23468 21548 23480
rect 21600 23468 21606 23520
rect 22922 23468 22928 23520
rect 22980 23508 22986 23520
rect 23569 23511 23627 23517
rect 23569 23508 23581 23511
rect 22980 23480 23581 23508
rect 22980 23468 22986 23480
rect 23569 23477 23581 23480
rect 23615 23477 23627 23511
rect 23569 23471 23627 23477
rect 1104 23418 30820 23440
rect 1104 23366 5915 23418
rect 5967 23366 5979 23418
rect 6031 23366 6043 23418
rect 6095 23366 6107 23418
rect 6159 23366 6171 23418
rect 6223 23366 15846 23418
rect 15898 23366 15910 23418
rect 15962 23366 15974 23418
rect 16026 23366 16038 23418
rect 16090 23366 16102 23418
rect 16154 23366 25776 23418
rect 25828 23366 25840 23418
rect 25892 23366 25904 23418
rect 25956 23366 25968 23418
rect 26020 23366 26032 23418
rect 26084 23366 30820 23418
rect 1104 23344 30820 23366
rect 7193 23307 7251 23313
rect 7193 23273 7205 23307
rect 7239 23304 7251 23307
rect 7374 23304 7380 23316
rect 7239 23276 7380 23304
rect 7239 23273 7251 23276
rect 7193 23267 7251 23273
rect 7374 23264 7380 23276
rect 7432 23264 7438 23316
rect 8386 23264 8392 23316
rect 8444 23304 8450 23316
rect 8938 23304 8944 23316
rect 8444 23276 8944 23304
rect 8444 23264 8450 23276
rect 8938 23264 8944 23276
rect 8996 23304 9002 23316
rect 9033 23307 9091 23313
rect 9033 23304 9045 23307
rect 8996 23276 9045 23304
rect 8996 23264 9002 23276
rect 9033 23273 9045 23276
rect 9079 23273 9091 23307
rect 9033 23267 9091 23273
rect 10870 23264 10876 23316
rect 10928 23304 10934 23316
rect 11149 23307 11207 23313
rect 11149 23304 11161 23307
rect 10928 23276 11161 23304
rect 10928 23264 10934 23276
rect 11149 23273 11161 23276
rect 11195 23273 11207 23307
rect 13538 23304 13544 23316
rect 13499 23276 13544 23304
rect 11149 23267 11207 23273
rect 13538 23264 13544 23276
rect 13596 23264 13602 23316
rect 15378 23264 15384 23316
rect 15436 23304 15442 23316
rect 15749 23307 15807 23313
rect 15749 23304 15761 23307
rect 15436 23276 15761 23304
rect 15436 23264 15442 23276
rect 15749 23273 15761 23276
rect 15795 23273 15807 23307
rect 15749 23267 15807 23273
rect 17129 23307 17187 23313
rect 17129 23273 17141 23307
rect 17175 23304 17187 23307
rect 17402 23304 17408 23316
rect 17175 23276 17408 23304
rect 17175 23273 17187 23276
rect 17129 23267 17187 23273
rect 17402 23264 17408 23276
rect 17460 23264 17466 23316
rect 17865 23307 17923 23313
rect 17865 23273 17877 23307
rect 17911 23304 17923 23307
rect 18506 23304 18512 23316
rect 17911 23276 18512 23304
rect 17911 23273 17923 23276
rect 17865 23267 17923 23273
rect 18506 23264 18512 23276
rect 18564 23264 18570 23316
rect 19337 23307 19395 23313
rect 19337 23273 19349 23307
rect 19383 23304 19395 23307
rect 20162 23304 20168 23316
rect 19383 23276 20168 23304
rect 19383 23273 19395 23276
rect 19337 23267 19395 23273
rect 20162 23264 20168 23276
rect 20220 23264 20226 23316
rect 20625 23307 20683 23313
rect 20625 23273 20637 23307
rect 20671 23304 20683 23307
rect 21174 23304 21180 23316
rect 20671 23276 21180 23304
rect 20671 23273 20683 23276
rect 20625 23267 20683 23273
rect 21174 23264 21180 23276
rect 21232 23264 21238 23316
rect 22554 23304 22560 23316
rect 22066 23276 22560 23304
rect 6546 23196 6552 23248
rect 6604 23236 6610 23248
rect 6733 23239 6791 23245
rect 6733 23236 6745 23239
rect 6604 23208 6745 23236
rect 6604 23196 6610 23208
rect 6733 23205 6745 23208
rect 6779 23236 6791 23239
rect 7466 23236 7472 23248
rect 6779 23208 7472 23236
rect 6779 23205 6791 23208
rect 6733 23199 6791 23205
rect 7466 23196 7472 23208
rect 7524 23196 7530 23248
rect 7742 23236 7748 23248
rect 7576 23208 7748 23236
rect 4430 23128 4436 23180
rect 4488 23168 4494 23180
rect 4525 23171 4583 23177
rect 4525 23168 4537 23171
rect 4488 23140 4537 23168
rect 4488 23128 4494 23140
rect 4525 23137 4537 23140
rect 4571 23137 4583 23171
rect 4525 23131 4583 23137
rect 4617 23171 4675 23177
rect 4617 23137 4629 23171
rect 4663 23168 4675 23171
rect 4798 23168 4804 23180
rect 4663 23140 4804 23168
rect 4663 23137 4675 23140
rect 4617 23131 4675 23137
rect 4798 23128 4804 23140
rect 4856 23128 4862 23180
rect 1394 23100 1400 23112
rect 1355 23072 1400 23100
rect 1394 23060 1400 23072
rect 1452 23060 1458 23112
rect 4341 23103 4399 23109
rect 4341 23069 4353 23103
rect 4387 23069 4399 23103
rect 4341 23063 4399 23069
rect 4709 23103 4767 23109
rect 4709 23069 4721 23103
rect 4755 23069 4767 23103
rect 4890 23100 4896 23112
rect 4851 23072 4896 23100
rect 4709 23063 4767 23069
rect 4356 23032 4384 23063
rect 4356 23004 4568 23032
rect 4540 22976 4568 23004
rect 1578 22964 1584 22976
rect 1539 22936 1584 22964
rect 1578 22924 1584 22936
rect 1636 22924 1642 22976
rect 4154 22964 4160 22976
rect 4115 22936 4160 22964
rect 4154 22924 4160 22936
rect 4212 22924 4218 22976
rect 4522 22924 4528 22976
rect 4580 22924 4586 22976
rect 4724 22964 4752 23063
rect 4890 23060 4896 23072
rect 4948 23060 4954 23112
rect 5353 23103 5411 23109
rect 5353 23069 5365 23103
rect 5399 23100 5411 23103
rect 7374 23100 7380 23112
rect 5399 23072 5764 23100
rect 7335 23072 7380 23100
rect 5399 23069 5411 23072
rect 5353 23063 5411 23069
rect 5736 23044 5764 23072
rect 7374 23060 7380 23072
rect 7432 23060 7438 23112
rect 7576 23109 7604 23208
rect 7742 23196 7748 23208
rect 7800 23236 7806 23248
rect 8202 23236 8208 23248
rect 7800 23208 8208 23236
rect 7800 23196 7806 23208
rect 8202 23196 8208 23208
rect 8260 23196 8266 23248
rect 15010 23196 15016 23248
rect 15068 23236 15074 23248
rect 17589 23239 17647 23245
rect 17589 23236 17601 23239
rect 15068 23208 17601 23236
rect 15068 23196 15074 23208
rect 17589 23205 17601 23208
rect 17635 23236 17647 23239
rect 18046 23236 18052 23248
rect 17635 23208 18052 23236
rect 17635 23205 17647 23208
rect 17589 23199 17647 23205
rect 18046 23196 18052 23208
rect 18104 23196 18110 23248
rect 19150 23196 19156 23248
rect 19208 23236 19214 23248
rect 21913 23239 21971 23245
rect 21913 23236 21925 23239
rect 19208 23208 21925 23236
rect 19208 23196 19214 23208
rect 21913 23205 21925 23208
rect 21959 23236 21971 23239
rect 22066 23236 22094 23276
rect 22554 23264 22560 23276
rect 22612 23264 22618 23316
rect 21959 23208 22094 23236
rect 21959 23205 21971 23208
rect 21913 23199 21971 23205
rect 7650 23128 7656 23180
rect 7708 23168 7714 23180
rect 16577 23171 16635 23177
rect 7708 23140 7753 23168
rect 14844 23140 15700 23168
rect 7708 23128 7714 23140
rect 14844 23112 14872 23140
rect 7561 23103 7619 23109
rect 7561 23069 7573 23103
rect 7607 23069 7619 23103
rect 7561 23063 7619 23069
rect 7745 23103 7803 23109
rect 7745 23069 7757 23103
rect 7791 23069 7803 23103
rect 7745 23063 7803 23069
rect 7929 23103 7987 23109
rect 7929 23069 7941 23103
rect 7975 23100 7987 23103
rect 8386 23100 8392 23112
rect 7975 23072 8392 23100
rect 7975 23069 7987 23072
rect 7929 23063 7987 23069
rect 5626 23041 5632 23044
rect 5620 23032 5632 23041
rect 5587 23004 5632 23032
rect 5620 22995 5632 23004
rect 5626 22992 5632 22995
rect 5684 22992 5690 23044
rect 5718 22992 5724 23044
rect 5776 22992 5782 23044
rect 5534 22964 5540 22976
rect 4724 22936 5540 22964
rect 5534 22924 5540 22936
rect 5592 22924 5598 22976
rect 7006 22924 7012 22976
rect 7064 22964 7070 22976
rect 7760 22964 7788 23063
rect 8386 23060 8392 23072
rect 8444 23060 8450 23112
rect 8478 23060 8484 23112
rect 8536 23100 8542 23112
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8536 23072 8953 23100
rect 8536 23060 8542 23072
rect 8941 23069 8953 23072
rect 8987 23069 8999 23103
rect 8941 23063 8999 23069
rect 9030 23060 9036 23112
rect 9088 23100 9094 23112
rect 9769 23103 9827 23109
rect 9769 23100 9781 23103
rect 9088 23072 9781 23100
rect 9088 23060 9094 23072
rect 9769 23069 9781 23072
rect 9815 23069 9827 23103
rect 9769 23063 9827 23069
rect 9858 23060 9864 23112
rect 9916 23100 9922 23112
rect 10025 23103 10083 23109
rect 10025 23100 10037 23103
rect 9916 23072 10037 23100
rect 9916 23060 9922 23072
rect 10025 23069 10037 23072
rect 10071 23069 10083 23103
rect 10025 23063 10083 23069
rect 11514 23060 11520 23112
rect 11572 23100 11578 23112
rect 12161 23103 12219 23109
rect 12161 23100 12173 23103
rect 11572 23072 12173 23100
rect 11572 23060 11578 23072
rect 12161 23069 12173 23072
rect 12207 23069 12219 23103
rect 14734 23100 14740 23112
rect 14695 23072 14740 23100
rect 12161 23063 12219 23069
rect 14734 23060 14740 23072
rect 14792 23060 14798 23112
rect 14826 23060 14832 23112
rect 14884 23100 14890 23112
rect 14884 23072 14929 23100
rect 14884 23060 14890 23072
rect 15010 23060 15016 23112
rect 15068 23100 15074 23112
rect 15672 23109 15700 23140
rect 16577 23137 16589 23171
rect 16623 23168 16635 23171
rect 16758 23168 16764 23180
rect 16623 23140 16764 23168
rect 16623 23137 16635 23140
rect 16577 23131 16635 23137
rect 16758 23128 16764 23140
rect 16816 23168 16822 23180
rect 18690 23168 18696 23180
rect 16816 23140 18696 23168
rect 16816 23128 16822 23140
rect 18690 23128 18696 23140
rect 18748 23128 18754 23180
rect 15657 23103 15715 23109
rect 15068 23072 15113 23100
rect 15068 23060 15074 23072
rect 15657 23069 15669 23103
rect 15703 23069 15715 23103
rect 15657 23063 15715 23069
rect 16390 23060 16396 23112
rect 16448 23100 16454 23112
rect 16669 23103 16727 23109
rect 16669 23100 16681 23103
rect 16448 23072 16681 23100
rect 16448 23060 16454 23072
rect 16669 23069 16681 23072
rect 16715 23069 16727 23103
rect 16669 23063 16727 23069
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23100 17647 23103
rect 17681 23103 17739 23109
rect 17681 23100 17693 23103
rect 17635 23072 17693 23100
rect 17635 23069 17647 23072
rect 17589 23063 17647 23069
rect 17681 23069 17693 23072
rect 17727 23069 17739 23103
rect 17681 23063 17739 23069
rect 17865 23103 17923 23109
rect 17865 23069 17877 23103
rect 17911 23100 17923 23103
rect 18046 23100 18052 23112
rect 17911 23072 18052 23100
rect 17911 23069 17923 23072
rect 17865 23063 17923 23069
rect 18046 23060 18052 23072
rect 18104 23060 18110 23112
rect 18325 23103 18383 23109
rect 18325 23069 18337 23103
rect 18371 23069 18383 23103
rect 18325 23063 18383 23069
rect 12428 23035 12486 23041
rect 12428 23001 12440 23035
rect 12474 23032 12486 23035
rect 12526 23032 12532 23044
rect 12474 23004 12532 23032
rect 12474 23001 12486 23004
rect 12428 22995 12486 23001
rect 12526 22992 12532 23004
rect 12584 22992 12590 23044
rect 15197 23035 15255 23041
rect 15197 23001 15209 23035
rect 15243 23032 15255 23035
rect 17402 23032 17408 23044
rect 15243 23004 17408 23032
rect 15243 23001 15255 23004
rect 15197 22995 15255 23001
rect 17402 22992 17408 23004
rect 17460 22992 17466 23044
rect 18332 23032 18360 23063
rect 19150 23060 19156 23112
rect 19208 23100 19214 23112
rect 19245 23103 19303 23109
rect 19245 23100 19257 23103
rect 19208 23072 19257 23100
rect 19208 23060 19214 23072
rect 19245 23069 19257 23072
rect 19291 23069 19303 23103
rect 19518 23100 19524 23112
rect 19479 23072 19524 23100
rect 19245 23063 19303 23069
rect 19518 23060 19524 23072
rect 19576 23060 19582 23112
rect 20349 23103 20407 23109
rect 20349 23069 20361 23103
rect 20395 23069 20407 23103
rect 20349 23063 20407 23069
rect 20533 23103 20591 23109
rect 20533 23069 20545 23103
rect 20579 23100 20591 23103
rect 20622 23100 20628 23112
rect 20579 23072 20628 23100
rect 20579 23069 20591 23072
rect 20533 23063 20591 23069
rect 18414 23032 18420 23044
rect 18332 23004 18420 23032
rect 18414 22992 18420 23004
rect 18472 23032 18478 23044
rect 18598 23032 18604 23044
rect 18472 23004 18604 23032
rect 18472 22992 18478 23004
rect 18598 22992 18604 23004
rect 18656 22992 18662 23044
rect 19705 23035 19763 23041
rect 19705 23001 19717 23035
rect 19751 23032 19763 23035
rect 20364 23032 20392 23063
rect 20622 23060 20628 23072
rect 20680 23060 20686 23112
rect 20717 23103 20775 23109
rect 20717 23069 20729 23103
rect 20763 23100 20775 23103
rect 21358 23100 21364 23112
rect 20763 23072 21364 23100
rect 20763 23069 20775 23072
rect 20717 23063 20775 23069
rect 21358 23060 21364 23072
rect 21416 23060 21422 23112
rect 22281 23103 22339 23109
rect 22281 23069 22293 23103
rect 22327 23100 22339 23103
rect 22462 23100 22468 23112
rect 22327 23072 22468 23100
rect 22327 23069 22339 23072
rect 22281 23063 22339 23069
rect 22462 23060 22468 23072
rect 22520 23060 22526 23112
rect 22922 23100 22928 23112
rect 22664 23072 22928 23100
rect 19751 23004 20392 23032
rect 22097 23035 22155 23041
rect 19751 23001 19763 23004
rect 19705 22995 19763 23001
rect 22097 23001 22109 23035
rect 22143 23032 22155 23035
rect 22664 23032 22692 23072
rect 22922 23060 22928 23072
rect 22980 23060 22986 23112
rect 23106 23100 23112 23112
rect 23067 23072 23112 23100
rect 23106 23060 23112 23072
rect 23164 23060 23170 23112
rect 22143 23004 22692 23032
rect 22143 23001 22155 23004
rect 22097 22995 22155 23001
rect 22738 22992 22744 23044
rect 22796 23032 22802 23044
rect 22796 23004 22841 23032
rect 22796 22992 22802 23004
rect 7064 22936 7788 22964
rect 16761 22967 16819 22973
rect 7064 22924 7070 22936
rect 16761 22933 16773 22967
rect 16807 22964 16819 22967
rect 16942 22964 16948 22976
rect 16807 22936 16948 22964
rect 16807 22933 16819 22936
rect 16761 22927 16819 22933
rect 16942 22924 16948 22936
rect 17000 22924 17006 22976
rect 18509 22967 18567 22973
rect 18509 22933 18521 22967
rect 18555 22964 18567 22967
rect 18874 22964 18880 22976
rect 18555 22936 18880 22964
rect 18555 22933 18567 22936
rect 18509 22927 18567 22933
rect 18874 22924 18880 22936
rect 18932 22924 18938 22976
rect 1104 22874 30820 22896
rect 1104 22822 10880 22874
rect 10932 22822 10944 22874
rect 10996 22822 11008 22874
rect 11060 22822 11072 22874
rect 11124 22822 11136 22874
rect 11188 22822 20811 22874
rect 20863 22822 20875 22874
rect 20927 22822 20939 22874
rect 20991 22822 21003 22874
rect 21055 22822 21067 22874
rect 21119 22822 30820 22874
rect 1104 22800 30820 22822
rect 4522 22720 4528 22772
rect 4580 22760 4586 22772
rect 5445 22763 5503 22769
rect 5445 22760 5457 22763
rect 4580 22732 5457 22760
rect 4580 22720 4586 22732
rect 5445 22729 5457 22732
rect 5491 22729 5503 22763
rect 5445 22723 5503 22729
rect 4154 22652 4160 22704
rect 4212 22692 4218 22704
rect 4310 22695 4368 22701
rect 4310 22692 4322 22695
rect 4212 22664 4322 22692
rect 4212 22652 4218 22664
rect 4310 22661 4322 22664
rect 4356 22661 4368 22695
rect 5460 22692 5488 22723
rect 5626 22720 5632 22772
rect 5684 22760 5690 22772
rect 6365 22763 6423 22769
rect 6365 22760 6377 22763
rect 5684 22732 6377 22760
rect 5684 22720 5690 22732
rect 6365 22729 6377 22732
rect 6411 22729 6423 22763
rect 7098 22760 7104 22772
rect 6365 22723 6423 22729
rect 6932 22732 7104 22760
rect 6270 22692 6276 22704
rect 5460 22664 6276 22692
rect 4310 22655 4368 22661
rect 6270 22652 6276 22664
rect 6328 22652 6334 22704
rect 1397 22627 1455 22633
rect 1397 22593 1409 22627
rect 1443 22624 1455 22627
rect 2038 22624 2044 22636
rect 1443 22596 1900 22624
rect 1999 22596 2044 22624
rect 1443 22593 1455 22596
rect 1397 22587 1455 22593
rect 1872 22556 1900 22596
rect 2038 22584 2044 22596
rect 2096 22584 2102 22636
rect 2685 22627 2743 22633
rect 2685 22593 2697 22627
rect 2731 22624 2743 22627
rect 2774 22624 2780 22636
rect 2731 22596 2780 22624
rect 2731 22593 2743 22596
rect 2685 22587 2743 22593
rect 2774 22584 2780 22596
rect 2832 22584 2838 22636
rect 3786 22584 3792 22636
rect 3844 22624 3850 22636
rect 4065 22627 4123 22633
rect 4065 22624 4077 22627
rect 3844 22596 4077 22624
rect 3844 22584 3850 22596
rect 4065 22593 4077 22596
rect 4111 22593 4123 22627
rect 6546 22624 6552 22636
rect 6507 22596 6552 22624
rect 4065 22587 4123 22593
rect 6546 22584 6552 22596
rect 6604 22584 6610 22636
rect 6932 22633 6960 22732
rect 7098 22720 7104 22732
rect 7156 22760 7162 22772
rect 8110 22760 8116 22772
rect 7156 22732 8116 22760
rect 7156 22720 7162 22732
rect 8110 22720 8116 22732
rect 8168 22720 8174 22772
rect 9122 22760 9128 22772
rect 9083 22732 9128 22760
rect 9122 22720 9128 22732
rect 9180 22720 9186 22772
rect 9585 22763 9643 22769
rect 9585 22729 9597 22763
rect 9631 22760 9643 22763
rect 10410 22760 10416 22772
rect 9631 22732 10416 22760
rect 9631 22729 9643 22732
rect 9585 22723 9643 22729
rect 10410 22720 10416 22732
rect 10468 22720 10474 22772
rect 11422 22760 11428 22772
rect 11164 22732 11428 22760
rect 11164 22704 11192 22732
rect 11422 22720 11428 22732
rect 11480 22720 11486 22772
rect 12066 22720 12072 22772
rect 12124 22720 12130 22772
rect 12802 22760 12808 22772
rect 12406 22732 12808 22760
rect 8294 22692 8300 22704
rect 7760 22664 8300 22692
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22593 6975 22627
rect 6917 22587 6975 22593
rect 7006 22584 7012 22636
rect 7064 22624 7070 22636
rect 7760 22633 7788 22664
rect 8294 22652 8300 22664
rect 8352 22692 8358 22704
rect 9030 22692 9036 22704
rect 8352 22664 9036 22692
rect 8352 22652 8358 22664
rect 9030 22652 9036 22664
rect 9088 22652 9094 22704
rect 11146 22652 11152 22704
rect 11204 22652 11210 22704
rect 11330 22652 11336 22704
rect 11388 22692 11394 22704
rect 11882 22692 11888 22704
rect 11388 22664 11560 22692
rect 11795 22664 11888 22692
rect 11388 22652 11394 22664
rect 8018 22633 8024 22636
rect 7101 22627 7159 22633
rect 7101 22624 7113 22627
rect 7064 22596 7113 22624
rect 7064 22584 7070 22596
rect 7101 22593 7113 22596
rect 7147 22593 7159 22627
rect 7101 22587 7159 22593
rect 7745 22627 7803 22633
rect 7745 22593 7757 22627
rect 7791 22593 7803 22627
rect 8012 22624 8024 22633
rect 7979 22596 8024 22624
rect 7745 22587 7803 22593
rect 8012 22587 8024 22596
rect 8018 22584 8024 22587
rect 8076 22584 8082 22636
rect 9122 22584 9128 22636
rect 9180 22624 9186 22636
rect 9398 22624 9404 22636
rect 9180 22596 9404 22624
rect 9180 22584 9186 22596
rect 9398 22584 9404 22596
rect 9456 22584 9462 22636
rect 9950 22584 9956 22636
rect 10008 22624 10014 22636
rect 10410 22624 10416 22636
rect 10008 22596 10416 22624
rect 10008 22584 10014 22596
rect 10410 22584 10416 22596
rect 10468 22584 10474 22636
rect 10686 22624 10692 22636
rect 10744 22633 10750 22636
rect 10656 22596 10692 22624
rect 10686 22584 10692 22596
rect 10744 22587 10756 22633
rect 10744 22584 10750 22587
rect 10870 22584 10876 22636
rect 10928 22624 10934 22636
rect 10965 22627 11023 22633
rect 10965 22624 10977 22627
rect 10928 22596 10977 22624
rect 10928 22584 10934 22596
rect 10965 22593 10977 22596
rect 11011 22624 11023 22627
rect 11422 22624 11428 22636
rect 11011 22596 11428 22624
rect 11011 22593 11023 22596
rect 10965 22587 11023 22593
rect 11422 22584 11428 22596
rect 11480 22584 11486 22636
rect 11532 22633 11560 22664
rect 11808 22633 11836 22664
rect 11882 22652 11888 22664
rect 11940 22692 11946 22704
rect 12084 22692 12112 22720
rect 11940 22664 12112 22692
rect 11940 22652 11946 22664
rect 11517 22627 11575 22633
rect 11517 22593 11529 22627
rect 11563 22593 11575 22627
rect 11517 22587 11575 22593
rect 11701 22627 11759 22633
rect 11701 22593 11713 22627
rect 11747 22593 11759 22627
rect 11701 22587 11759 22593
rect 11793 22627 11851 22633
rect 11793 22593 11805 22627
rect 11839 22593 11851 22627
rect 11793 22587 11851 22593
rect 12069 22627 12127 22633
rect 12069 22593 12081 22627
rect 12115 22624 12127 22627
rect 12406 22624 12434 22732
rect 12802 22720 12808 22732
rect 12860 22720 12866 22772
rect 14829 22763 14887 22769
rect 14829 22729 14841 22763
rect 14875 22760 14887 22763
rect 15654 22760 15660 22772
rect 14875 22732 15660 22760
rect 14875 22729 14887 22732
rect 14829 22723 14887 22729
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 16574 22720 16580 22772
rect 16632 22760 16638 22772
rect 16669 22763 16727 22769
rect 16669 22760 16681 22763
rect 16632 22732 16681 22760
rect 16632 22720 16638 22732
rect 16669 22729 16681 22732
rect 16715 22729 16727 22763
rect 16669 22723 16727 22729
rect 17402 22720 17408 22772
rect 17460 22760 17466 22772
rect 18693 22763 18751 22769
rect 18693 22760 18705 22763
rect 17460 22732 18705 22760
rect 17460 22720 17466 22732
rect 18693 22729 18705 22732
rect 18739 22729 18751 22763
rect 18693 22723 18751 22729
rect 20073 22763 20131 22769
rect 20073 22729 20085 22763
rect 20119 22760 20131 22763
rect 20346 22760 20352 22772
rect 20119 22732 20352 22760
rect 20119 22729 20131 22732
rect 20073 22723 20131 22729
rect 20346 22720 20352 22732
rect 20404 22720 20410 22772
rect 22462 22720 22468 22772
rect 22520 22760 22526 22772
rect 23109 22763 23167 22769
rect 23109 22760 23121 22763
rect 22520 22732 23121 22760
rect 22520 22720 22526 22732
rect 23109 22729 23121 22732
rect 23155 22729 23167 22763
rect 23109 22723 23167 22729
rect 12526 22652 12532 22704
rect 12584 22692 12590 22704
rect 12958 22695 13016 22701
rect 12958 22692 12970 22695
rect 12584 22664 12970 22692
rect 12584 22652 12590 22664
rect 12958 22661 12970 22664
rect 13004 22661 13016 22695
rect 12958 22655 13016 22661
rect 16390 22652 16396 22704
rect 16448 22692 16454 22704
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 16448 22664 17141 22692
rect 16448 22652 16454 22664
rect 17129 22661 17141 22664
rect 17175 22661 17187 22695
rect 17129 22655 17187 22661
rect 19886 22652 19892 22704
rect 19944 22692 19950 22704
rect 20990 22692 20996 22704
rect 19944 22664 20996 22692
rect 19944 22652 19950 22664
rect 20990 22652 20996 22664
rect 21048 22652 21054 22704
rect 12710 22624 12716 22636
rect 12115 22596 12434 22624
rect 12671 22596 12716 22624
rect 12115 22593 12127 22596
rect 12069 22587 12127 22593
rect 2866 22556 2872 22568
rect 1872 22528 2872 22556
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 6362 22516 6368 22568
rect 6420 22556 6426 22568
rect 6733 22559 6791 22565
rect 6733 22556 6745 22559
rect 6420 22528 6745 22556
rect 6420 22516 6426 22528
rect 6733 22525 6745 22528
rect 6779 22525 6791 22559
rect 6733 22519 6791 22525
rect 6825 22559 6883 22565
rect 6825 22525 6837 22559
rect 6871 22525 6883 22559
rect 11716 22556 11744 22587
rect 12710 22584 12716 22596
rect 12768 22584 12774 22636
rect 14737 22627 14795 22633
rect 14737 22624 14749 22627
rect 14108 22596 14749 22624
rect 6825 22519 6883 22525
rect 10980 22528 11744 22556
rect 11885 22559 11943 22565
rect 2225 22491 2283 22497
rect 2225 22457 2237 22491
rect 2271 22488 2283 22491
rect 3970 22488 3976 22500
rect 2271 22460 3976 22488
rect 2271 22457 2283 22460
rect 2225 22451 2283 22457
rect 3970 22448 3976 22460
rect 4028 22448 4034 22500
rect 6546 22448 6552 22500
rect 6604 22488 6610 22500
rect 6840 22488 6868 22519
rect 6604 22460 6868 22488
rect 6604 22448 6610 22460
rect 1581 22423 1639 22429
rect 1581 22389 1593 22423
rect 1627 22420 1639 22423
rect 1946 22420 1952 22432
rect 1627 22392 1952 22420
rect 1627 22389 1639 22392
rect 1581 22383 1639 22389
rect 1946 22380 1952 22392
rect 2004 22380 2010 22432
rect 2869 22423 2927 22429
rect 2869 22389 2881 22423
rect 2915 22420 2927 22423
rect 4246 22420 4252 22432
rect 2915 22392 4252 22420
rect 2915 22389 2927 22392
rect 2869 22383 2927 22389
rect 4246 22380 4252 22392
rect 4304 22380 4310 22432
rect 5810 22380 5816 22432
rect 5868 22420 5874 22432
rect 10980 22420 11008 22528
rect 11885 22525 11897 22559
rect 11931 22556 11943 22559
rect 12158 22556 12164 22568
rect 11931 22528 12164 22556
rect 11931 22525 11943 22528
rect 11885 22519 11943 22525
rect 12158 22516 12164 22528
rect 12216 22516 12222 22568
rect 11514 22448 11520 22500
rect 11572 22488 11578 22500
rect 12728 22488 12756 22584
rect 11572 22460 12756 22488
rect 11572 22448 11578 22460
rect 12250 22420 12256 22432
rect 5868 22392 11008 22420
rect 12211 22392 12256 22420
rect 5868 22380 5874 22392
rect 12250 22380 12256 22392
rect 12308 22380 12314 22432
rect 13722 22380 13728 22432
rect 13780 22420 13786 22432
rect 14108 22429 14136 22596
rect 14737 22593 14749 22596
rect 14783 22593 14795 22627
rect 14737 22587 14795 22593
rect 16482 22584 16488 22636
rect 16540 22624 16546 22636
rect 16758 22624 16764 22636
rect 16540 22596 16764 22624
rect 16540 22584 16546 22596
rect 16758 22584 16764 22596
rect 16816 22624 16822 22636
rect 17037 22627 17095 22633
rect 17037 22624 17049 22627
rect 16816 22596 17049 22624
rect 16816 22584 16822 22596
rect 17037 22593 17049 22596
rect 17083 22593 17095 22627
rect 17037 22587 17095 22593
rect 18785 22627 18843 22633
rect 18785 22593 18797 22627
rect 18831 22624 18843 22627
rect 19702 22624 19708 22636
rect 18831 22596 19708 22624
rect 18831 22593 18843 22596
rect 18785 22587 18843 22593
rect 19702 22584 19708 22596
rect 19760 22624 19766 22636
rect 19981 22627 20039 22633
rect 19981 22624 19993 22627
rect 19760 22596 19993 22624
rect 19760 22584 19766 22596
rect 19981 22593 19993 22596
rect 20027 22593 20039 22627
rect 21174 22624 21180 22636
rect 21135 22596 21180 22624
rect 19981 22587 20039 22593
rect 21174 22584 21180 22596
rect 21232 22584 21238 22636
rect 23014 22584 23020 22636
rect 23072 22584 23078 22636
rect 29825 22627 29883 22633
rect 29825 22593 29837 22627
rect 29871 22624 29883 22627
rect 30190 22624 30196 22636
rect 29871 22596 30196 22624
rect 29871 22593 29883 22596
rect 29825 22587 29883 22593
rect 30190 22584 30196 22596
rect 30248 22584 30254 22636
rect 22376 22568 22428 22574
rect 15562 22516 15568 22568
rect 15620 22556 15626 22568
rect 16390 22556 16396 22568
rect 15620 22528 16396 22556
rect 15620 22516 15626 22528
rect 16390 22516 16396 22528
rect 16448 22516 16454 22568
rect 17221 22559 17279 22565
rect 17221 22556 17233 22559
rect 17144 22528 17233 22556
rect 15010 22448 15016 22500
rect 15068 22488 15074 22500
rect 16206 22488 16212 22500
rect 15068 22460 16212 22488
rect 15068 22448 15074 22460
rect 16206 22448 16212 22460
rect 16264 22448 16270 22500
rect 16482 22448 16488 22500
rect 16540 22488 16546 22500
rect 16850 22488 16856 22500
rect 16540 22460 16856 22488
rect 16540 22448 16546 22460
rect 16850 22448 16856 22460
rect 16908 22448 16914 22500
rect 14093 22423 14151 22429
rect 14093 22420 14105 22423
rect 13780 22392 14105 22420
rect 13780 22380 13786 22392
rect 14093 22389 14105 22392
rect 14139 22389 14151 22423
rect 14093 22383 14151 22389
rect 15102 22380 15108 22432
rect 15160 22420 15166 22432
rect 16666 22420 16672 22432
rect 15160 22392 16672 22420
rect 15160 22380 15166 22392
rect 16666 22380 16672 22392
rect 16724 22420 16730 22432
rect 17144 22420 17172 22528
rect 17221 22525 17233 22528
rect 17267 22556 17279 22559
rect 18046 22556 18052 22568
rect 17267 22528 18052 22556
rect 17267 22525 17279 22528
rect 17221 22519 17279 22525
rect 18046 22516 18052 22528
rect 18104 22556 18110 22568
rect 18509 22559 18567 22565
rect 18509 22556 18521 22559
rect 18104 22528 18521 22556
rect 18104 22516 18110 22528
rect 18509 22525 18521 22528
rect 18555 22556 18567 22559
rect 18874 22556 18880 22568
rect 18555 22528 18880 22556
rect 18555 22525 18567 22528
rect 18509 22519 18567 22525
rect 18874 22516 18880 22528
rect 18932 22556 18938 22568
rect 20165 22559 20223 22565
rect 20165 22556 20177 22559
rect 18932 22528 20177 22556
rect 18932 22516 18938 22528
rect 20165 22525 20177 22528
rect 20211 22525 20223 22559
rect 20165 22519 20223 22525
rect 24121 22559 24179 22565
rect 24121 22525 24133 22559
rect 24167 22556 24179 22559
rect 30098 22556 30104 22568
rect 24167 22528 30104 22556
rect 24167 22525 24179 22528
rect 24121 22519 24179 22525
rect 30098 22516 30104 22528
rect 30156 22516 30162 22568
rect 22376 22510 22428 22516
rect 19518 22448 19524 22500
rect 19576 22488 19582 22500
rect 20809 22491 20867 22497
rect 20809 22488 20821 22491
rect 19576 22460 20821 22488
rect 19576 22448 19582 22460
rect 20809 22457 20821 22460
rect 20855 22457 20867 22491
rect 20809 22451 20867 22457
rect 16724 22392 17172 22420
rect 19153 22423 19211 22429
rect 16724 22380 16730 22392
rect 19153 22389 19165 22423
rect 19199 22420 19211 22423
rect 19426 22420 19432 22432
rect 19199 22392 19432 22420
rect 19199 22389 19211 22392
rect 19153 22383 19211 22389
rect 19426 22380 19432 22392
rect 19484 22380 19490 22432
rect 19610 22420 19616 22432
rect 19571 22392 19616 22420
rect 19610 22380 19616 22392
rect 19668 22380 19674 22432
rect 30006 22420 30012 22432
rect 29967 22392 30012 22420
rect 30006 22380 30012 22392
rect 30064 22380 30070 22432
rect 1104 22330 30820 22352
rect 1104 22278 5915 22330
rect 5967 22278 5979 22330
rect 6031 22278 6043 22330
rect 6095 22278 6107 22330
rect 6159 22278 6171 22330
rect 6223 22278 15846 22330
rect 15898 22278 15910 22330
rect 15962 22278 15974 22330
rect 16026 22278 16038 22330
rect 16090 22278 16102 22330
rect 16154 22278 25776 22330
rect 25828 22278 25840 22330
rect 25892 22278 25904 22330
rect 25956 22278 25968 22330
rect 26020 22278 26032 22330
rect 26084 22278 30820 22330
rect 1104 22256 30820 22278
rect 10686 22176 10692 22228
rect 10744 22216 10750 22228
rect 10965 22219 11023 22225
rect 10965 22216 10977 22219
rect 10744 22188 10977 22216
rect 10744 22176 10750 22188
rect 10965 22185 10977 22188
rect 11011 22185 11023 22219
rect 10965 22179 11023 22185
rect 15309 22188 16804 22216
rect 8202 22108 8208 22160
rect 8260 22148 8266 22160
rect 9398 22148 9404 22160
rect 8260 22120 9404 22148
rect 8260 22108 8266 22120
rect 9398 22108 9404 22120
rect 9456 22108 9462 22160
rect 4798 22040 4804 22092
rect 4856 22080 4862 22092
rect 5261 22083 5319 22089
rect 5261 22080 5273 22083
rect 4856 22052 5273 22080
rect 4856 22040 4862 22052
rect 5261 22049 5273 22052
rect 5307 22049 5319 22083
rect 5261 22043 5319 22049
rect 5718 22040 5724 22092
rect 5776 22080 5782 22092
rect 6181 22083 6239 22089
rect 6181 22080 6193 22083
rect 5776 22052 6193 22080
rect 5776 22040 5782 22052
rect 6181 22049 6193 22052
rect 6227 22049 6239 22083
rect 8938 22080 8944 22092
rect 8899 22052 8944 22080
rect 6181 22043 6239 22049
rect 8938 22040 8944 22052
rect 8996 22040 9002 22092
rect 9217 22083 9275 22089
rect 9217 22049 9229 22083
rect 9263 22080 9275 22083
rect 9490 22080 9496 22092
rect 9263 22052 9496 22080
rect 9263 22049 9275 22052
rect 9217 22043 9275 22049
rect 9490 22040 9496 22052
rect 9548 22080 9554 22092
rect 10597 22083 10655 22089
rect 10597 22080 10609 22083
rect 9548 22052 10609 22080
rect 9548 22040 9554 22052
rect 10597 22049 10609 22052
rect 10643 22049 10655 22083
rect 11882 22080 11888 22092
rect 11843 22052 11888 22080
rect 10597 22043 10655 22049
rect 11882 22040 11888 22052
rect 11940 22040 11946 22092
rect 12345 22083 12403 22089
rect 12345 22049 12357 22083
rect 12391 22080 12403 22083
rect 12526 22080 12532 22092
rect 12391 22052 12532 22080
rect 12391 22049 12403 22052
rect 12345 22043 12403 22049
rect 12526 22040 12532 22052
rect 12584 22040 12590 22092
rect 1670 21972 1676 22024
rect 1728 22012 1734 22024
rect 1857 22015 1915 22021
rect 1857 22012 1869 22015
rect 1728 21984 1869 22012
rect 1728 21972 1734 21984
rect 1857 21981 1869 21984
rect 1903 22012 1915 22015
rect 3694 22012 3700 22024
rect 1903 21984 3700 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 3694 21972 3700 21984
rect 3752 21972 3758 22024
rect 5534 22012 5540 22024
rect 5495 21984 5540 22012
rect 5534 21972 5540 21984
rect 5592 21972 5598 22024
rect 7190 21972 7196 22024
rect 7248 22012 7254 22024
rect 8113 22015 8171 22021
rect 8113 22012 8125 22015
rect 7248 21984 8125 22012
rect 7248 21972 7254 21984
rect 8113 21981 8125 21984
rect 8159 21981 8171 22015
rect 8113 21975 8171 21981
rect 9582 21972 9588 22024
rect 9640 22012 9646 22024
rect 10229 22015 10287 22021
rect 10229 22012 10241 22015
rect 9640 21984 10241 22012
rect 9640 21972 9646 21984
rect 10229 21981 10241 21984
rect 10275 21981 10287 22015
rect 10229 21975 10287 21981
rect 10318 21972 10324 22024
rect 10376 22012 10382 22024
rect 10413 22015 10471 22021
rect 10413 22012 10425 22015
rect 10376 21984 10425 22012
rect 10376 21972 10382 21984
rect 10413 21981 10425 21984
rect 10459 21981 10471 22015
rect 10413 21975 10471 21981
rect 10505 22015 10563 22021
rect 10505 21981 10517 22015
rect 10551 21981 10563 22015
rect 10778 22012 10784 22024
rect 10739 21984 10784 22012
rect 10505 21975 10563 21981
rect 2124 21947 2182 21953
rect 2124 21913 2136 21947
rect 2170 21944 2182 21947
rect 2406 21944 2412 21956
rect 2170 21916 2412 21944
rect 2170 21913 2182 21916
rect 2124 21907 2182 21913
rect 2406 21904 2412 21916
rect 2464 21904 2470 21956
rect 6448 21947 6506 21953
rect 6448 21913 6460 21947
rect 6494 21944 6506 21947
rect 6730 21944 6736 21956
rect 6494 21916 6736 21944
rect 6494 21913 6506 21916
rect 6448 21907 6506 21913
rect 6730 21904 6736 21916
rect 6788 21904 6794 21956
rect 8294 21944 8300 21956
rect 8255 21916 8300 21944
rect 8294 21904 8300 21916
rect 8352 21904 8358 21956
rect 9214 21904 9220 21956
rect 9272 21944 9278 21956
rect 10520 21944 10548 21975
rect 10778 21972 10784 21984
rect 10836 21972 10842 22024
rect 11238 21972 11244 22024
rect 11296 22012 11302 22024
rect 11606 22012 11612 22024
rect 11296 21984 11612 22012
rect 11296 21972 11302 21984
rect 11606 21972 11612 21984
rect 11664 21972 11670 22024
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 21981 11851 22015
rect 11974 22012 11980 22024
rect 11935 21984 11980 22012
rect 11793 21975 11851 21981
rect 9272 21916 10548 21944
rect 9272 21904 9278 21916
rect 2958 21836 2964 21888
rect 3016 21876 3022 21888
rect 3237 21879 3295 21885
rect 3237 21876 3249 21879
rect 3016 21848 3249 21876
rect 3016 21836 3022 21848
rect 3237 21845 3249 21848
rect 3283 21845 3295 21879
rect 3237 21839 3295 21845
rect 7006 21836 7012 21888
rect 7064 21876 7070 21888
rect 7561 21879 7619 21885
rect 7561 21876 7573 21879
rect 7064 21848 7573 21876
rect 7064 21836 7070 21848
rect 7561 21845 7573 21848
rect 7607 21876 7619 21879
rect 7834 21876 7840 21888
rect 7607 21848 7840 21876
rect 7607 21845 7619 21848
rect 7561 21839 7619 21845
rect 7834 21836 7840 21848
rect 7892 21876 7898 21888
rect 11808 21876 11836 21975
rect 11974 21972 11980 21984
rect 12032 21972 12038 22024
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 22012 12219 22015
rect 13722 22012 13728 22024
rect 12207 21984 13728 22012
rect 12207 21981 12219 21984
rect 12161 21975 12219 21981
rect 13722 21972 13728 21984
rect 13780 21972 13786 22024
rect 15194 21972 15200 22024
rect 15252 22012 15258 22024
rect 15309 22012 15337 22188
rect 15378 22108 15384 22160
rect 15436 22148 15442 22160
rect 16669 22151 16727 22157
rect 16669 22148 16681 22151
rect 15436 22120 16681 22148
rect 15436 22108 15442 22120
rect 16669 22117 16681 22120
rect 16715 22117 16727 22151
rect 16776 22148 16804 22188
rect 17034 22176 17040 22228
rect 17092 22216 17098 22228
rect 17129 22219 17187 22225
rect 17129 22216 17141 22219
rect 17092 22188 17141 22216
rect 17092 22176 17098 22188
rect 17129 22185 17141 22188
rect 17175 22216 17187 22219
rect 18690 22216 18696 22228
rect 17175 22188 18696 22216
rect 17175 22185 17187 22188
rect 17129 22179 17187 22185
rect 18690 22176 18696 22188
rect 18748 22176 18754 22228
rect 19058 22176 19064 22228
rect 19116 22216 19122 22228
rect 21450 22216 21456 22228
rect 19116 22188 21456 22216
rect 19116 22176 19122 22188
rect 21450 22176 21456 22188
rect 21508 22176 21514 22228
rect 16776 22120 19334 22148
rect 16669 22111 16727 22117
rect 19306 22092 19334 22120
rect 19426 22108 19432 22160
rect 19484 22108 19490 22160
rect 15654 22080 15660 22092
rect 15615 22052 15660 22080
rect 15654 22040 15660 22052
rect 15712 22040 15718 22092
rect 18138 22080 18144 22092
rect 18099 22052 18144 22080
rect 18138 22040 18144 22052
rect 18196 22040 18202 22092
rect 18233 22083 18291 22089
rect 18233 22049 18245 22083
rect 18279 22049 18291 22083
rect 19306 22052 19340 22092
rect 18233 22043 18291 22049
rect 15381 22015 15439 22021
rect 15381 22012 15393 22015
rect 15252 21984 15393 22012
rect 15252 21972 15258 21984
rect 15381 21981 15393 21984
rect 15427 21981 15439 22015
rect 15381 21975 15439 21981
rect 15746 21972 15752 22024
rect 15804 22021 15810 22024
rect 15804 22012 15812 22021
rect 16482 22012 16488 22024
rect 15804 21984 16488 22012
rect 15804 21975 15812 21984
rect 15804 21972 15810 21975
rect 16482 21972 16488 21984
rect 16540 21972 16546 22024
rect 16666 22012 16672 22024
rect 16627 21984 16672 22012
rect 16666 21972 16672 21984
rect 16724 21972 16730 22024
rect 16850 22012 16856 22024
rect 16811 21984 16856 22012
rect 16850 21972 16856 21984
rect 16908 21972 16914 22024
rect 16945 22015 17003 22021
rect 16945 21981 16957 22015
rect 16991 22012 17003 22015
rect 17034 22012 17040 22024
rect 16991 21984 17040 22012
rect 16991 21981 17003 21984
rect 16945 21975 17003 21981
rect 17034 21972 17040 21984
rect 17092 21972 17098 22024
rect 17221 22015 17279 22021
rect 17221 21981 17233 22015
rect 17267 21981 17279 22015
rect 17221 21975 17279 21981
rect 15562 21944 15568 21956
rect 15523 21916 15568 21944
rect 15562 21904 15568 21916
rect 15620 21904 15626 21956
rect 15657 21947 15715 21953
rect 15657 21913 15669 21947
rect 15703 21944 15715 21947
rect 15838 21944 15844 21956
rect 15703 21916 15844 21944
rect 15703 21913 15715 21916
rect 15657 21907 15715 21913
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 7892 21848 11836 21876
rect 17236 21876 17264 21975
rect 17310 21972 17316 22024
rect 17368 22012 17374 22024
rect 17678 22012 17684 22024
rect 17368 21984 17684 22012
rect 17368 21972 17374 21984
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 18046 21972 18052 22024
rect 18104 22012 18110 22024
rect 18248 22012 18276 22043
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 19444 22021 19472 22108
rect 20990 22040 20996 22092
rect 21048 22080 21054 22092
rect 21177 22083 21235 22089
rect 21177 22080 21189 22083
rect 21048 22052 21189 22080
rect 21048 22040 21054 22052
rect 21177 22049 21189 22052
rect 21223 22080 21235 22083
rect 22002 22080 22008 22092
rect 21223 22052 22008 22080
rect 21223 22049 21235 22052
rect 21177 22043 21235 22049
rect 22002 22040 22008 22052
rect 22060 22080 22066 22092
rect 22370 22080 22376 22092
rect 22060 22052 22376 22080
rect 22060 22040 22066 22052
rect 22370 22040 22376 22052
rect 22428 22040 22434 22092
rect 18104 21984 18276 22012
rect 19429 22015 19487 22021
rect 18104 21972 18110 21984
rect 19429 21981 19441 22015
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 22012 19671 22015
rect 20438 22012 20444 22024
rect 19659 21984 20444 22012
rect 19659 21981 19671 21984
rect 19613 21975 19671 21981
rect 20438 21972 20444 21984
rect 20496 21972 20502 22024
rect 21085 22015 21143 22021
rect 21085 21981 21097 22015
rect 21131 22012 21143 22015
rect 21634 22012 21640 22024
rect 21131 21984 21640 22012
rect 21131 21981 21143 21984
rect 21085 21975 21143 21981
rect 21634 21972 21640 21984
rect 21692 21972 21698 22024
rect 22281 22015 22339 22021
rect 22281 21981 22293 22015
rect 22327 22012 22339 22015
rect 22462 22012 22468 22024
rect 22327 21984 22468 22012
rect 22327 21981 22339 21984
rect 22281 21975 22339 21981
rect 22462 21972 22468 21984
rect 22520 21972 22526 22024
rect 20993 21947 21051 21953
rect 18332 21916 19380 21944
rect 17681 21879 17739 21885
rect 17681 21876 17693 21879
rect 17236 21848 17693 21876
rect 7892 21836 7898 21848
rect 17681 21845 17693 21848
rect 17727 21845 17739 21879
rect 18046 21876 18052 21888
rect 18007 21848 18052 21876
rect 17681 21839 17739 21845
rect 18046 21836 18052 21848
rect 18104 21836 18110 21888
rect 18138 21836 18144 21888
rect 18196 21876 18202 21888
rect 18332 21876 18360 21916
rect 18196 21848 18360 21876
rect 18196 21836 18202 21848
rect 19058 21836 19064 21888
rect 19116 21876 19122 21888
rect 19245 21879 19303 21885
rect 19245 21876 19257 21879
rect 19116 21848 19257 21876
rect 19116 21836 19122 21848
rect 19245 21845 19257 21848
rect 19291 21845 19303 21879
rect 19352 21876 19380 21916
rect 20993 21913 21005 21947
rect 21039 21944 21051 21947
rect 21174 21944 21180 21956
rect 21039 21916 21180 21944
rect 21039 21913 21051 21916
rect 20993 21907 21051 21913
rect 21174 21904 21180 21916
rect 21232 21944 21238 21956
rect 22189 21947 22247 21953
rect 22189 21944 22201 21947
rect 21232 21916 22201 21944
rect 21232 21904 21238 21916
rect 22189 21913 22201 21916
rect 22235 21944 22247 21947
rect 23014 21944 23020 21956
rect 22235 21916 23020 21944
rect 22235 21913 22247 21916
rect 22189 21907 22247 21913
rect 23014 21904 23020 21916
rect 23072 21904 23078 21956
rect 20625 21879 20683 21885
rect 20625 21876 20637 21879
rect 19352 21848 20637 21876
rect 19245 21839 19303 21845
rect 20625 21845 20637 21848
rect 20671 21845 20683 21879
rect 21818 21876 21824 21888
rect 21779 21848 21824 21876
rect 20625 21839 20683 21845
rect 21818 21836 21824 21848
rect 21876 21836 21882 21888
rect 1104 21786 30820 21808
rect 1104 21734 10880 21786
rect 10932 21734 10944 21786
rect 10996 21734 11008 21786
rect 11060 21734 11072 21786
rect 11124 21734 11136 21786
rect 11188 21734 20811 21786
rect 20863 21734 20875 21786
rect 20927 21734 20939 21786
rect 20991 21734 21003 21786
rect 21055 21734 21067 21786
rect 21119 21734 30820 21786
rect 1104 21712 30820 21734
rect 4430 21632 4436 21684
rect 4488 21672 4494 21684
rect 4893 21675 4951 21681
rect 4893 21672 4905 21675
rect 4488 21644 4905 21672
rect 4488 21632 4494 21644
rect 4893 21641 4905 21644
rect 4939 21641 4951 21675
rect 4893 21635 4951 21641
rect 5721 21675 5779 21681
rect 5721 21641 5733 21675
rect 5767 21672 5779 21675
rect 7374 21672 7380 21684
rect 5767 21644 7380 21672
rect 5767 21641 5779 21644
rect 5721 21635 5779 21641
rect 7374 21632 7380 21644
rect 7432 21632 7438 21684
rect 12802 21632 12808 21684
rect 12860 21672 12866 21684
rect 12989 21675 13047 21681
rect 12989 21672 13001 21675
rect 12860 21644 13001 21672
rect 12860 21632 12866 21644
rect 12989 21641 13001 21644
rect 13035 21672 13047 21675
rect 15473 21675 15531 21681
rect 15473 21672 15485 21675
rect 13035 21644 15485 21672
rect 13035 21641 13047 21644
rect 12989 21635 13047 21641
rect 15473 21641 15485 21644
rect 15519 21641 15531 21675
rect 15473 21635 15531 21641
rect 15562 21632 15568 21684
rect 15620 21672 15626 21684
rect 15933 21675 15991 21681
rect 15933 21672 15945 21675
rect 15620 21644 15945 21672
rect 15620 21632 15626 21644
rect 15933 21641 15945 21644
rect 15979 21641 15991 21675
rect 15933 21635 15991 21641
rect 16666 21632 16672 21684
rect 16724 21672 16730 21684
rect 17405 21675 17463 21681
rect 17405 21672 17417 21675
rect 16724 21644 17417 21672
rect 16724 21632 16730 21644
rect 17405 21641 17417 21644
rect 17451 21641 17463 21675
rect 17405 21635 17463 21641
rect 19061 21675 19119 21681
rect 19061 21641 19073 21675
rect 19107 21672 19119 21675
rect 19426 21672 19432 21684
rect 19107 21644 19432 21672
rect 19107 21641 19119 21644
rect 19061 21635 19119 21641
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 7926 21604 7932 21616
rect 7887 21576 7932 21604
rect 7926 21564 7932 21576
rect 7984 21564 7990 21616
rect 9582 21604 9588 21616
rect 8036 21576 9588 21604
rect 1670 21536 1676 21548
rect 1631 21508 1676 21536
rect 1670 21496 1676 21508
rect 1728 21496 1734 21548
rect 1940 21539 1998 21545
rect 1940 21505 1952 21539
rect 1986 21536 1998 21539
rect 2222 21536 2228 21548
rect 1986 21508 2228 21536
rect 1986 21505 1998 21508
rect 1940 21499 1998 21505
rect 2222 21496 2228 21508
rect 2280 21496 2286 21548
rect 3234 21496 3240 21548
rect 3292 21536 3298 21548
rect 3697 21539 3755 21545
rect 3697 21536 3709 21539
rect 3292 21508 3709 21536
rect 3292 21496 3298 21508
rect 3697 21505 3709 21508
rect 3743 21505 3755 21539
rect 3697 21499 3755 21505
rect 4985 21539 5043 21545
rect 4985 21505 4997 21539
rect 5031 21536 5043 21539
rect 5534 21536 5540 21548
rect 5031 21508 5540 21536
rect 5031 21505 5043 21508
rect 4985 21499 5043 21505
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 5810 21536 5816 21548
rect 5771 21508 5816 21536
rect 5810 21496 5816 21508
rect 5868 21496 5874 21548
rect 6270 21496 6276 21548
rect 6328 21536 6334 21548
rect 6914 21536 6920 21548
rect 6328 21508 6920 21536
rect 6328 21496 6334 21508
rect 6914 21496 6920 21508
rect 6972 21496 6978 21548
rect 7190 21536 7196 21548
rect 7103 21508 7196 21536
rect 7190 21496 7196 21508
rect 7248 21536 7254 21548
rect 8036 21536 8064 21576
rect 9582 21564 9588 21576
rect 9640 21564 9646 21616
rect 10410 21564 10416 21616
rect 10468 21604 10474 21616
rect 10781 21607 10839 21613
rect 10781 21604 10793 21607
rect 10468 21576 10793 21604
rect 10468 21564 10474 21576
rect 10781 21573 10793 21576
rect 10827 21573 10839 21607
rect 10781 21567 10839 21573
rect 11876 21607 11934 21613
rect 11876 21573 11888 21607
rect 11922 21604 11934 21607
rect 12250 21604 12256 21616
rect 11922 21576 12256 21604
rect 11922 21573 11934 21576
rect 11876 21567 11934 21573
rect 12250 21564 12256 21576
rect 12308 21564 12314 21616
rect 15286 21564 15292 21616
rect 15344 21604 15350 21616
rect 15838 21604 15844 21616
rect 15344 21576 15844 21604
rect 15344 21564 15350 21576
rect 7248 21508 8064 21536
rect 8113 21539 8171 21545
rect 7248 21496 7254 21508
rect 8113 21505 8125 21539
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 8128 21468 8156 21499
rect 8478 21496 8484 21548
rect 8536 21536 8542 21548
rect 8665 21539 8723 21545
rect 8665 21536 8677 21539
rect 8536 21508 8677 21536
rect 8536 21496 8542 21508
rect 8665 21505 8677 21508
rect 8711 21505 8723 21539
rect 8665 21499 8723 21505
rect 8941 21539 8999 21545
rect 8941 21505 8953 21539
rect 8987 21536 8999 21539
rect 9214 21536 9220 21548
rect 8987 21508 9220 21536
rect 8987 21505 8999 21508
rect 8941 21499 8999 21505
rect 9214 21496 9220 21508
rect 9272 21496 9278 21548
rect 10137 21539 10195 21545
rect 10137 21505 10149 21539
rect 10183 21536 10195 21539
rect 10686 21536 10692 21548
rect 10183 21508 10692 21536
rect 10183 21505 10195 21508
rect 10137 21499 10195 21505
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 15580 21545 15608 21576
rect 15838 21564 15844 21576
rect 15896 21564 15902 21616
rect 17034 21564 17040 21616
rect 17092 21604 17098 21616
rect 18598 21604 18604 21616
rect 17092 21576 18604 21604
rect 17092 21564 17098 21576
rect 18598 21564 18604 21576
rect 18656 21564 18662 21616
rect 19886 21564 19892 21616
rect 19944 21604 19950 21616
rect 20073 21607 20131 21613
rect 20073 21604 20085 21607
rect 19944 21576 20085 21604
rect 19944 21564 19950 21576
rect 20073 21573 20085 21576
rect 20119 21604 20131 21607
rect 20438 21604 20444 21616
rect 20119 21576 20444 21604
rect 20119 21573 20131 21576
rect 20073 21567 20131 21573
rect 20438 21564 20444 21576
rect 20496 21564 20502 21616
rect 21542 21564 21548 21616
rect 21600 21604 21606 21616
rect 21821 21607 21879 21613
rect 21821 21604 21833 21607
rect 21600 21576 21833 21604
rect 21600 21564 21606 21576
rect 21821 21573 21833 21576
rect 21867 21573 21879 21607
rect 22002 21604 22008 21616
rect 21963 21576 22008 21604
rect 21821 21567 21879 21573
rect 22002 21564 22008 21576
rect 22060 21564 22066 21616
rect 22189 21607 22247 21613
rect 22189 21573 22201 21607
rect 22235 21604 22247 21607
rect 22462 21604 22468 21616
rect 22235 21576 22468 21604
rect 22235 21573 22247 21576
rect 22189 21567 22247 21573
rect 22462 21564 22468 21576
rect 22520 21564 22526 21616
rect 15565 21539 15623 21545
rect 15565 21505 15577 21539
rect 15611 21505 15623 21539
rect 15565 21499 15623 21505
rect 15654 21496 15660 21548
rect 15712 21536 15718 21548
rect 16669 21539 16727 21545
rect 16669 21536 16681 21539
rect 15712 21508 16681 21536
rect 15712 21496 15718 21508
rect 16669 21505 16681 21508
rect 16715 21505 16727 21539
rect 16669 21499 16727 21505
rect 16853 21539 16911 21545
rect 16853 21505 16865 21539
rect 16899 21536 16911 21539
rect 17126 21536 17132 21548
rect 16899 21508 17132 21536
rect 16899 21505 16911 21508
rect 16853 21499 16911 21505
rect 17126 21496 17132 21508
rect 17184 21496 17190 21548
rect 17221 21539 17279 21545
rect 17221 21505 17233 21539
rect 17267 21536 17279 21539
rect 17267 21508 17908 21536
rect 17267 21505 17279 21508
rect 17221 21499 17279 21505
rect 8128 21440 8984 21468
rect 8956 21412 8984 21440
rect 11514 21428 11520 21480
rect 11572 21468 11578 21480
rect 11609 21471 11667 21477
rect 11609 21468 11621 21471
rect 11572 21440 11621 21468
rect 11572 21428 11578 21440
rect 11609 21437 11621 21440
rect 11655 21437 11667 21471
rect 11609 21431 11667 21437
rect 15102 21428 15108 21480
rect 15160 21468 15166 21480
rect 15289 21471 15347 21477
rect 15289 21468 15301 21471
rect 15160 21440 15301 21468
rect 15160 21428 15166 21440
rect 15289 21437 15301 21440
rect 15335 21437 15347 21471
rect 15289 21431 15347 21437
rect 16945 21471 17003 21477
rect 16945 21437 16957 21471
rect 16991 21437 17003 21471
rect 16945 21431 17003 21437
rect 17037 21471 17095 21477
rect 17037 21437 17049 21471
rect 17083 21468 17095 21471
rect 17083 21440 17816 21468
rect 17083 21437 17095 21440
rect 17037 21431 17095 21437
rect 2774 21360 2780 21412
rect 2832 21400 2838 21412
rect 3513 21403 3571 21409
rect 3513 21400 3525 21403
rect 2832 21372 3525 21400
rect 2832 21360 2838 21372
rect 3513 21369 3525 21372
rect 3559 21369 3571 21403
rect 3513 21363 3571 21369
rect 8938 21360 8944 21412
rect 8996 21360 9002 21412
rect 10965 21403 11023 21409
rect 10965 21369 10977 21403
rect 11011 21400 11023 21403
rect 11238 21400 11244 21412
rect 11011 21372 11244 21400
rect 11011 21369 11023 21372
rect 10965 21363 11023 21369
rect 11238 21360 11244 21372
rect 11296 21360 11302 21412
rect 16960 21400 16988 21431
rect 17494 21400 17500 21412
rect 16960 21372 17500 21400
rect 17494 21360 17500 21372
rect 17552 21360 17558 21412
rect 3050 21332 3056 21344
rect 3011 21304 3056 21332
rect 3050 21292 3056 21304
rect 3108 21292 3114 21344
rect 6454 21292 6460 21344
rect 6512 21332 6518 21344
rect 7926 21332 7932 21344
rect 6512 21304 7932 21332
rect 6512 21292 6518 21304
rect 7926 21292 7932 21304
rect 7984 21292 7990 21344
rect 10042 21332 10048 21344
rect 10003 21304 10048 21332
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 17788 21332 17816 21440
rect 17880 21409 17908 21508
rect 18046 21496 18052 21548
rect 18104 21536 18110 21548
rect 18233 21539 18291 21545
rect 18233 21536 18245 21539
rect 18104 21508 18245 21536
rect 18104 21496 18110 21508
rect 18233 21505 18245 21508
rect 18279 21505 18291 21539
rect 19058 21536 19064 21548
rect 19019 21508 19064 21536
rect 18233 21499 18291 21505
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 19245 21539 19303 21545
rect 19245 21505 19257 21539
rect 19291 21505 19303 21539
rect 19245 21499 19303 21505
rect 18325 21471 18383 21477
rect 18325 21437 18337 21471
rect 18371 21468 18383 21471
rect 18414 21468 18420 21480
rect 18371 21440 18420 21468
rect 18371 21437 18383 21440
rect 18325 21431 18383 21437
rect 18414 21428 18420 21440
rect 18472 21428 18478 21480
rect 18509 21471 18567 21477
rect 18509 21437 18521 21471
rect 18555 21468 18567 21471
rect 18874 21468 18880 21480
rect 18555 21440 18880 21468
rect 18555 21437 18567 21440
rect 18509 21431 18567 21437
rect 18874 21428 18880 21440
rect 18932 21468 18938 21480
rect 19260 21468 19288 21499
rect 19334 21496 19340 21548
rect 19392 21536 19398 21548
rect 19610 21536 19616 21548
rect 19392 21508 19437 21536
rect 19571 21508 19616 21536
rect 19392 21496 19398 21508
rect 19610 21496 19616 21508
rect 19668 21496 19674 21548
rect 20257 21539 20315 21545
rect 20257 21505 20269 21539
rect 20303 21536 20315 21539
rect 20530 21536 20536 21548
rect 20303 21508 20536 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 18932 21440 19288 21468
rect 19521 21471 19579 21477
rect 18932 21428 18938 21440
rect 19521 21437 19533 21471
rect 19567 21468 19579 21471
rect 20438 21468 20444 21480
rect 19567 21440 20444 21468
rect 19567 21437 19579 21440
rect 19521 21431 19579 21437
rect 17865 21403 17923 21409
rect 17865 21369 17877 21403
rect 17911 21369 17923 21403
rect 17865 21363 17923 21369
rect 18690 21360 18696 21412
rect 18748 21400 18754 21412
rect 19536 21400 19564 21431
rect 20438 21428 20444 21440
rect 20496 21428 20502 21480
rect 18748 21372 19564 21400
rect 18748 21360 18754 21372
rect 19886 21332 19892 21344
rect 17788 21304 19892 21332
rect 19886 21292 19892 21304
rect 19944 21292 19950 21344
rect 20346 21292 20352 21344
rect 20404 21332 20410 21344
rect 20441 21335 20499 21341
rect 20441 21332 20453 21335
rect 20404 21304 20453 21332
rect 20404 21292 20410 21304
rect 20441 21301 20453 21304
rect 20487 21301 20499 21335
rect 20441 21295 20499 21301
rect 1104 21242 30820 21264
rect 1104 21190 5915 21242
rect 5967 21190 5979 21242
rect 6031 21190 6043 21242
rect 6095 21190 6107 21242
rect 6159 21190 6171 21242
rect 6223 21190 15846 21242
rect 15898 21190 15910 21242
rect 15962 21190 15974 21242
rect 16026 21190 16038 21242
rect 16090 21190 16102 21242
rect 16154 21190 25776 21242
rect 25828 21190 25840 21242
rect 25892 21190 25904 21242
rect 25956 21190 25968 21242
rect 26020 21190 26032 21242
rect 26084 21190 30820 21242
rect 1104 21168 30820 21190
rect 2222 21128 2228 21140
rect 2183 21100 2228 21128
rect 2222 21088 2228 21100
rect 2280 21088 2286 21140
rect 6546 21128 6552 21140
rect 6291 21100 6552 21128
rect 6178 21020 6184 21072
rect 6236 21020 6242 21072
rect 6196 20992 6224 21020
rect 6291 21001 6319 21100
rect 6546 21088 6552 21100
rect 6604 21088 6610 21140
rect 6730 21128 6736 21140
rect 6691 21100 6736 21128
rect 6730 21088 6736 21100
rect 6788 21088 6794 21140
rect 8478 21088 8484 21140
rect 8536 21128 8542 21140
rect 8941 21131 8999 21137
rect 8941 21128 8953 21131
rect 8536 21100 8953 21128
rect 8536 21088 8542 21100
rect 8941 21097 8953 21100
rect 8987 21097 8999 21131
rect 10410 21128 10416 21140
rect 10371 21100 10416 21128
rect 8941 21091 8999 21097
rect 10410 21088 10416 21100
rect 10468 21088 10474 21140
rect 11149 21131 11207 21137
rect 11149 21097 11161 21131
rect 11195 21128 11207 21131
rect 11330 21128 11336 21140
rect 11195 21100 11336 21128
rect 11195 21097 11207 21100
rect 11149 21091 11207 21097
rect 11330 21088 11336 21100
rect 11388 21088 11394 21140
rect 13538 21088 13544 21140
rect 13596 21128 13602 21140
rect 19245 21131 19303 21137
rect 13596 21100 18276 21128
rect 13596 21088 13602 21100
rect 7650 21020 7656 21072
rect 7708 21060 7714 21072
rect 8113 21063 8171 21069
rect 8113 21060 8125 21063
rect 7708 21032 8125 21060
rect 7708 21020 7714 21032
rect 8113 21029 8125 21032
rect 8159 21029 8171 21063
rect 8113 21023 8171 21029
rect 12618 21020 12624 21072
rect 12676 21060 12682 21072
rect 13173 21063 13231 21069
rect 13173 21060 13185 21063
rect 12676 21032 13185 21060
rect 12676 21020 12682 21032
rect 13173 21029 13185 21032
rect 13219 21029 13231 21063
rect 13173 21023 13231 21029
rect 16574 21020 16580 21072
rect 16632 21020 16638 21072
rect 17589 21063 17647 21069
rect 17589 21029 17601 21063
rect 17635 21029 17647 21063
rect 18248 21060 18276 21100
rect 19245 21097 19257 21131
rect 19291 21128 19303 21131
rect 19334 21128 19340 21140
rect 19291 21100 19340 21128
rect 19291 21097 19303 21100
rect 19245 21091 19303 21097
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 19702 21128 19708 21140
rect 19663 21100 19708 21128
rect 19702 21088 19708 21100
rect 19760 21088 19766 21140
rect 20530 21128 20536 21140
rect 20491 21100 20536 21128
rect 20530 21088 20536 21100
rect 20588 21088 20594 21140
rect 19518 21060 19524 21072
rect 18248 21032 19524 21060
rect 17589 21023 17647 21029
rect 6012 20964 6224 20992
rect 6273 20995 6331 21001
rect 1486 20924 1492 20936
rect 1447 20896 1492 20924
rect 1486 20884 1492 20896
rect 1544 20884 1550 20936
rect 1578 20884 1584 20936
rect 1636 20924 1642 20936
rect 1673 20927 1731 20933
rect 1673 20924 1685 20927
rect 1636 20896 1685 20924
rect 1636 20884 1642 20896
rect 1673 20893 1685 20896
rect 1719 20893 1731 20927
rect 1673 20887 1731 20893
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20893 1823 20927
rect 1765 20887 1823 20893
rect 1780 20856 1808 20887
rect 1854 20884 1860 20936
rect 1912 20924 1918 20936
rect 2041 20927 2099 20933
rect 1912 20896 1957 20924
rect 1912 20884 1918 20896
rect 2041 20893 2053 20927
rect 2087 20924 2099 20927
rect 3050 20924 3056 20936
rect 2087 20896 3056 20924
rect 2087 20893 2099 20896
rect 2041 20887 2099 20893
rect 3050 20884 3056 20896
rect 3108 20884 3114 20936
rect 3789 20927 3847 20933
rect 3789 20893 3801 20927
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 1596 20828 1808 20856
rect 1596 20800 1624 20828
rect 2958 20816 2964 20868
rect 3016 20856 3022 20868
rect 3804 20856 3832 20887
rect 4154 20884 4160 20936
rect 4212 20924 4218 20936
rect 6012 20933 6040 20964
rect 6273 20961 6285 20995
rect 6319 20961 6331 20995
rect 6273 20955 6331 20961
rect 6362 20952 6368 21004
rect 6420 20992 6426 21004
rect 7377 20995 7435 21001
rect 6420 20964 6465 20992
rect 6420 20952 6426 20964
rect 7377 20961 7389 20995
rect 7423 20992 7435 20995
rect 9306 20992 9312 21004
rect 7423 20964 9312 20992
rect 7423 20961 7435 20964
rect 7377 20955 7435 20961
rect 9306 20952 9312 20964
rect 9364 20952 9370 21004
rect 15010 20992 15016 21004
rect 14971 20964 15016 20992
rect 15010 20952 15016 20964
rect 15068 20952 15074 21004
rect 16485 20995 16543 21001
rect 16485 20961 16497 20995
rect 16531 20992 16543 20995
rect 16592 20992 16620 21020
rect 16531 20964 16620 20992
rect 16531 20961 16543 20964
rect 16485 20955 16543 20961
rect 16850 20952 16856 21004
rect 16908 20992 16914 21004
rect 17604 20992 17632 21023
rect 19518 21020 19524 21032
rect 19576 21020 19582 21072
rect 16908 20964 17632 20992
rect 18233 20995 18291 21001
rect 16908 20952 16914 20964
rect 18233 20961 18245 20995
rect 18279 20992 18291 20995
rect 18874 20992 18880 21004
rect 18279 20964 18880 20992
rect 18279 20961 18291 20964
rect 18233 20955 18291 20961
rect 4617 20927 4675 20933
rect 4617 20924 4629 20927
rect 4212 20896 4629 20924
rect 4212 20884 4218 20896
rect 4617 20893 4629 20896
rect 4663 20893 4675 20927
rect 4617 20887 4675 20893
rect 5997 20927 6055 20933
rect 5997 20893 6009 20927
rect 6043 20893 6055 20927
rect 6181 20927 6239 20933
rect 6181 20926 6193 20927
rect 5997 20887 6055 20893
rect 6104 20898 6193 20926
rect 3016 20828 3832 20856
rect 3881 20859 3939 20865
rect 3016 20816 3022 20828
rect 3881 20825 3893 20859
rect 3927 20856 3939 20859
rect 6104 20856 6132 20898
rect 6181 20893 6193 20898
rect 6227 20893 6239 20927
rect 6181 20887 6239 20893
rect 6549 20927 6607 20933
rect 6549 20893 6561 20927
rect 6595 20924 6607 20927
rect 7006 20924 7012 20936
rect 6595 20896 7012 20924
rect 6595 20893 6607 20896
rect 6549 20887 6607 20893
rect 7006 20884 7012 20896
rect 7064 20884 7070 20936
rect 7561 20927 7619 20933
rect 7561 20893 7573 20927
rect 7607 20924 7619 20927
rect 7607 20896 9352 20924
rect 7607 20893 7619 20896
rect 7561 20887 7619 20893
rect 9324 20868 9352 20896
rect 12894 20884 12900 20936
rect 12952 20924 12958 20936
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 12952 20896 14105 20924
rect 12952 20884 12958 20896
rect 14093 20893 14105 20896
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 15197 20927 15255 20933
rect 15197 20893 15209 20927
rect 15243 20924 15255 20927
rect 16574 20924 16580 20936
rect 15243 20896 16580 20924
rect 15243 20893 15255 20896
rect 15197 20887 15255 20893
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 18049 20927 18107 20933
rect 18049 20924 18061 20927
rect 17236 20896 18061 20924
rect 6822 20856 6828 20868
rect 3927 20828 6040 20856
rect 6104 20828 6828 20856
rect 3927 20825 3939 20828
rect 3881 20819 3939 20825
rect 1578 20748 1584 20800
rect 1636 20748 1642 20800
rect 3142 20788 3148 20800
rect 3103 20760 3148 20788
rect 3142 20748 3148 20760
rect 3200 20748 3206 20800
rect 4430 20788 4436 20800
rect 4391 20760 4436 20788
rect 4430 20748 4436 20760
rect 4488 20748 4494 20800
rect 6012 20788 6040 20828
rect 6822 20816 6828 20828
rect 6880 20856 6886 20868
rect 7282 20856 7288 20868
rect 6880 20828 7288 20856
rect 6880 20816 6886 20828
rect 7282 20816 7288 20828
rect 7340 20816 7346 20868
rect 8297 20859 8355 20865
rect 8297 20825 8309 20859
rect 8343 20856 8355 20859
rect 8478 20856 8484 20868
rect 8343 20828 8484 20856
rect 8343 20825 8355 20828
rect 8297 20819 8355 20825
rect 8478 20816 8484 20828
rect 8536 20816 8542 20868
rect 9030 20816 9036 20868
rect 9088 20856 9094 20868
rect 9125 20859 9183 20865
rect 9125 20856 9137 20859
rect 9088 20828 9137 20856
rect 9088 20816 9094 20828
rect 9125 20825 9137 20828
rect 9171 20825 9183 20859
rect 9306 20856 9312 20868
rect 9267 20828 9312 20856
rect 9125 20819 9183 20825
rect 9306 20816 9312 20828
rect 9364 20816 9370 20868
rect 10505 20859 10563 20865
rect 10505 20825 10517 20859
rect 10551 20856 10563 20859
rect 10594 20856 10600 20868
rect 10551 20828 10600 20856
rect 10551 20825 10563 20828
rect 10505 20819 10563 20825
rect 10594 20816 10600 20828
rect 10652 20816 10658 20868
rect 11241 20859 11299 20865
rect 11241 20825 11253 20859
rect 11287 20856 11299 20859
rect 11330 20856 11336 20868
rect 11287 20828 11336 20856
rect 11287 20825 11299 20828
rect 11241 20819 11299 20825
rect 11330 20816 11336 20828
rect 11388 20816 11394 20868
rect 13357 20859 13415 20865
rect 13357 20825 13369 20859
rect 13403 20856 13415 20859
rect 13446 20856 13452 20868
rect 13403 20828 13452 20856
rect 13403 20825 13415 20828
rect 13357 20819 13415 20825
rect 13446 20816 13452 20828
rect 13504 20816 13510 20868
rect 13538 20816 13544 20868
rect 13596 20856 13602 20868
rect 14185 20859 14243 20865
rect 13596 20828 13641 20856
rect 13596 20816 13602 20828
rect 14185 20825 14197 20859
rect 14231 20856 14243 20859
rect 16669 20859 16727 20865
rect 16669 20856 16681 20859
rect 14231 20828 16681 20856
rect 14231 20825 14243 20828
rect 14185 20819 14243 20825
rect 16669 20825 16681 20828
rect 16715 20856 16727 20859
rect 17236 20856 17264 20896
rect 18049 20893 18061 20896
rect 18095 20893 18107 20927
rect 18049 20887 18107 20893
rect 16715 20828 17264 20856
rect 16715 20825 16727 20828
rect 16669 20819 16727 20825
rect 17494 20816 17500 20868
rect 17552 20856 17558 20868
rect 17957 20859 18015 20865
rect 17957 20856 17969 20859
rect 17552 20828 17969 20856
rect 17552 20816 17558 20828
rect 17957 20825 17969 20828
rect 18003 20856 18015 20859
rect 18616 20856 18644 20964
rect 18874 20952 18880 20964
rect 18932 20952 18938 21004
rect 20254 20992 20260 21004
rect 19536 20964 20260 20992
rect 18690 20884 18696 20936
rect 18748 20924 18754 20936
rect 19536 20933 19564 20964
rect 20254 20952 20260 20964
rect 20312 20952 20318 21004
rect 20714 20952 20720 21004
rect 20772 20992 20778 21004
rect 20993 20995 21051 21001
rect 20993 20992 21005 20995
rect 20772 20964 21005 20992
rect 20772 20952 20778 20964
rect 20993 20961 21005 20964
rect 21039 20961 21051 20995
rect 20993 20955 21051 20961
rect 21085 20995 21143 21001
rect 21085 20961 21097 20995
rect 21131 20961 21143 20995
rect 21085 20955 21143 20961
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 18748 20896 19441 20924
rect 18748 20884 18754 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19794 20924 19800 20936
rect 19755 20896 19800 20924
rect 19521 20887 19579 20893
rect 19794 20884 19800 20896
rect 19852 20884 19858 20936
rect 21100 20924 21128 20955
rect 22370 20924 22376 20936
rect 20548 20896 22376 20924
rect 20548 20868 20576 20896
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 29822 20924 29828 20936
rect 29783 20896 29828 20924
rect 29822 20884 29828 20896
rect 29880 20884 29886 20936
rect 19610 20856 19616 20868
rect 18003 20828 18092 20856
rect 18616 20828 19616 20856
rect 18003 20825 18015 20828
rect 17957 20819 18015 20825
rect 18064 20800 18092 20828
rect 19610 20816 19616 20828
rect 19668 20856 19674 20868
rect 20530 20856 20536 20868
rect 19668 20828 20536 20856
rect 19668 20816 19674 20828
rect 20530 20816 20536 20828
rect 20588 20816 20594 20868
rect 20901 20859 20959 20865
rect 20901 20825 20913 20859
rect 20947 20856 20959 20859
rect 20947 20828 22094 20856
rect 20947 20825 20959 20828
rect 20901 20819 20959 20825
rect 7374 20788 7380 20800
rect 6012 20760 7380 20788
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 12986 20788 12992 20800
rect 9732 20760 12992 20788
rect 9732 20748 9738 20760
rect 12986 20748 12992 20760
rect 13044 20788 13050 20800
rect 15105 20791 15163 20797
rect 15105 20788 15117 20791
rect 13044 20760 15117 20788
rect 13044 20748 13050 20760
rect 15105 20757 15117 20760
rect 15151 20757 15163 20791
rect 15562 20788 15568 20800
rect 15523 20760 15568 20788
rect 15105 20751 15163 20757
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 16758 20748 16764 20800
rect 16816 20788 16822 20800
rect 17126 20788 17132 20800
rect 16816 20760 16861 20788
rect 17087 20760 17132 20788
rect 16816 20748 16822 20760
rect 17126 20748 17132 20760
rect 17184 20748 17190 20800
rect 18046 20748 18052 20800
rect 18104 20748 18110 20800
rect 18874 20748 18880 20800
rect 18932 20788 18938 20800
rect 21818 20788 21824 20800
rect 18932 20760 21824 20788
rect 18932 20748 18938 20760
rect 21818 20748 21824 20760
rect 21876 20748 21882 20800
rect 22066 20788 22094 20828
rect 22186 20788 22192 20800
rect 22066 20760 22192 20788
rect 22186 20748 22192 20760
rect 22244 20748 22250 20800
rect 30006 20788 30012 20800
rect 29967 20760 30012 20788
rect 30006 20748 30012 20760
rect 30064 20748 30070 20800
rect 1104 20698 30820 20720
rect 1104 20646 10880 20698
rect 10932 20646 10944 20698
rect 10996 20646 11008 20698
rect 11060 20646 11072 20698
rect 11124 20646 11136 20698
rect 11188 20646 20811 20698
rect 20863 20646 20875 20698
rect 20927 20646 20939 20698
rect 20991 20646 21003 20698
rect 21055 20646 21067 20698
rect 21119 20646 30820 20698
rect 1104 20624 30820 20646
rect 2406 20584 2412 20596
rect 2367 20556 2412 20584
rect 2406 20544 2412 20556
rect 2464 20544 2470 20596
rect 5534 20544 5540 20596
rect 5592 20584 5598 20596
rect 8113 20587 8171 20593
rect 8113 20584 8125 20587
rect 5592 20556 8125 20584
rect 5592 20544 5598 20556
rect 8113 20553 8125 20556
rect 8159 20553 8171 20587
rect 8113 20547 8171 20553
rect 8478 20544 8484 20596
rect 8536 20544 8542 20596
rect 8846 20544 8852 20596
rect 8904 20584 8910 20596
rect 8941 20587 8999 20593
rect 8941 20584 8953 20587
rect 8904 20556 8953 20584
rect 8904 20544 8910 20556
rect 8941 20553 8953 20556
rect 8987 20553 8999 20587
rect 8941 20547 8999 20553
rect 10134 20544 10140 20596
rect 10192 20584 10198 20596
rect 14642 20584 14648 20596
rect 10192 20556 14648 20584
rect 10192 20544 10198 20556
rect 14642 20544 14648 20556
rect 14700 20544 14706 20596
rect 15378 20584 15384 20596
rect 15339 20556 15384 20584
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 15473 20587 15531 20593
rect 15473 20553 15485 20587
rect 15519 20584 15531 20587
rect 15562 20584 15568 20596
rect 15519 20556 15568 20584
rect 15519 20553 15531 20556
rect 15473 20547 15531 20553
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 16758 20544 16764 20596
rect 16816 20584 16822 20596
rect 16853 20587 16911 20593
rect 16853 20584 16865 20587
rect 16816 20556 16865 20584
rect 16816 20544 16822 20556
rect 16853 20553 16865 20556
rect 16899 20553 16911 20587
rect 16853 20547 16911 20553
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19521 20587 19579 20593
rect 19521 20584 19533 20587
rect 19484 20556 19533 20584
rect 19484 20544 19490 20556
rect 19521 20553 19533 20556
rect 19567 20553 19579 20587
rect 19521 20547 19579 20553
rect 20622 20544 20628 20596
rect 20680 20544 20686 20596
rect 22278 20584 22284 20596
rect 22239 20556 22284 20584
rect 22278 20544 22284 20556
rect 22336 20544 22342 20596
rect 29822 20544 29828 20596
rect 29880 20584 29886 20596
rect 29917 20587 29975 20593
rect 29917 20584 29929 20587
rect 29880 20556 29929 20584
rect 29880 20544 29886 20556
rect 29917 20553 29929 20556
rect 29963 20553 29975 20587
rect 29917 20547 29975 20553
rect 4430 20516 4436 20528
rect 1872 20488 4436 20516
rect 1486 20408 1492 20460
rect 1544 20448 1550 20460
rect 1872 20457 1900 20488
rect 4430 20476 4436 20488
rect 4488 20476 4494 20528
rect 6362 20476 6368 20528
rect 6420 20516 6426 20528
rect 8297 20519 8355 20525
rect 6420 20488 7006 20516
rect 6420 20476 6426 20488
rect 1673 20451 1731 20457
rect 1673 20448 1685 20451
rect 1544 20420 1685 20448
rect 1544 20408 1550 20420
rect 1673 20417 1685 20420
rect 1719 20417 1731 20451
rect 1673 20411 1731 20417
rect 1857 20451 1915 20457
rect 1857 20417 1869 20451
rect 1903 20417 1915 20451
rect 1857 20411 1915 20417
rect 2225 20451 2283 20457
rect 2225 20417 2237 20451
rect 2271 20448 2283 20451
rect 2958 20448 2964 20460
rect 2271 20420 2964 20448
rect 2271 20417 2283 20420
rect 2225 20411 2283 20417
rect 2958 20408 2964 20420
rect 3016 20408 3022 20460
rect 3050 20408 3056 20460
rect 3108 20448 3114 20460
rect 3964 20451 4022 20457
rect 3108 20420 3153 20448
rect 3108 20408 3114 20420
rect 3964 20417 3976 20451
rect 4010 20448 4022 20451
rect 4522 20448 4528 20460
rect 4010 20420 4528 20448
rect 4010 20417 4022 20420
rect 3964 20411 4022 20417
rect 4522 20408 4528 20420
rect 4580 20408 4586 20460
rect 5537 20451 5595 20457
rect 5537 20448 5549 20451
rect 5092 20420 5549 20448
rect 1578 20340 1584 20392
rect 1636 20380 1642 20392
rect 1949 20383 2007 20389
rect 1949 20380 1961 20383
rect 1636 20352 1961 20380
rect 1636 20340 1642 20352
rect 1949 20349 1961 20352
rect 1995 20349 2007 20383
rect 1949 20343 2007 20349
rect 2041 20383 2099 20389
rect 2041 20349 2053 20383
rect 2087 20349 2099 20383
rect 3694 20380 3700 20392
rect 3655 20352 3700 20380
rect 2041 20343 2099 20349
rect 1762 20272 1768 20324
rect 1820 20312 1826 20324
rect 2056 20312 2084 20343
rect 3694 20340 3700 20352
rect 3752 20340 3758 20392
rect 1820 20284 3740 20312
rect 1820 20272 1826 20284
rect 2866 20244 2872 20256
rect 2827 20216 2872 20244
rect 2866 20204 2872 20216
rect 2924 20204 2930 20256
rect 3712 20244 3740 20284
rect 5092 20256 5120 20420
rect 5537 20417 5549 20420
rect 5583 20417 5595 20451
rect 5537 20411 5595 20417
rect 6457 20451 6515 20457
rect 6457 20417 6469 20451
rect 6503 20417 6515 20451
rect 6457 20411 6515 20417
rect 6472 20380 6500 20411
rect 6546 20408 6552 20460
rect 6604 20448 6610 20460
rect 6730 20448 6736 20460
rect 6604 20420 6649 20448
rect 6691 20420 6736 20448
rect 6604 20408 6610 20420
rect 6730 20408 6736 20420
rect 6788 20408 6794 20460
rect 6822 20408 6828 20460
rect 6880 20448 6886 20460
rect 6978 20457 7006 20488
rect 8297 20485 8309 20519
rect 8343 20516 8355 20519
rect 8496 20516 8524 20544
rect 9582 20516 9588 20528
rect 8343 20488 9588 20516
rect 8343 20485 8355 20488
rect 8297 20479 8355 20485
rect 9582 20476 9588 20488
rect 9640 20476 9646 20528
rect 18138 20516 18144 20528
rect 14568 20488 18144 20516
rect 14568 20460 14596 20488
rect 18138 20476 18144 20488
rect 18196 20476 18202 20528
rect 20640 20516 20668 20544
rect 22186 20516 22192 20528
rect 18524 20488 20668 20516
rect 22147 20488 22192 20516
rect 6963 20451 7021 20457
rect 6880 20420 6925 20448
rect 6880 20408 6886 20420
rect 6963 20417 6975 20451
rect 7009 20417 7021 20451
rect 8478 20448 8484 20460
rect 8439 20420 8484 20448
rect 6963 20411 7021 20417
rect 8478 20408 8484 20420
rect 8536 20448 8542 20460
rect 9030 20448 9036 20460
rect 8536 20420 9036 20448
rect 8536 20408 8542 20420
rect 9030 20408 9036 20420
rect 9088 20408 9094 20460
rect 9401 20451 9459 20457
rect 9401 20417 9413 20451
rect 9447 20448 9459 20451
rect 9674 20448 9680 20460
rect 9447 20420 9680 20448
rect 9447 20417 9459 20420
rect 9401 20411 9459 20417
rect 9674 20408 9680 20420
rect 9732 20408 9738 20460
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 9953 20451 10011 20457
rect 9953 20417 9965 20451
rect 9999 20448 10011 20451
rect 10594 20448 10600 20460
rect 9999 20420 10600 20448
rect 9999 20417 10011 20420
rect 9953 20411 10011 20417
rect 6638 20380 6644 20392
rect 6472 20352 6644 20380
rect 6638 20340 6644 20352
rect 6696 20380 6702 20392
rect 8754 20380 8760 20392
rect 6696 20352 8760 20380
rect 6696 20340 6702 20352
rect 8754 20340 8760 20352
rect 8812 20340 8818 20392
rect 9876 20380 9904 20411
rect 10594 20408 10600 20420
rect 10652 20408 10658 20460
rect 11238 20408 11244 20460
rect 11296 20448 11302 20460
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 11296 20420 11529 20448
rect 11296 20408 11302 20420
rect 11517 20417 11529 20420
rect 11563 20417 11575 20451
rect 11517 20411 11575 20417
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 10134 20380 10140 20392
rect 9876 20352 10140 20380
rect 10134 20340 10140 20352
rect 10192 20340 10198 20392
rect 11054 20340 11060 20392
rect 11112 20380 11118 20392
rect 11716 20380 11744 20411
rect 11790 20408 11796 20460
rect 11848 20448 11854 20460
rect 12069 20451 12127 20457
rect 11848 20420 11893 20448
rect 11848 20408 11854 20420
rect 12069 20417 12081 20451
rect 12115 20448 12127 20451
rect 12894 20448 12900 20460
rect 12115 20420 12900 20448
rect 12115 20417 12127 20420
rect 12069 20411 12127 20417
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 13446 20448 13452 20460
rect 13407 20420 13452 20448
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 13538 20408 13544 20460
rect 13596 20448 13602 20460
rect 14093 20451 14151 20457
rect 14093 20448 14105 20451
rect 13596 20420 14105 20448
rect 13596 20408 13602 20420
rect 14093 20417 14105 20420
rect 14139 20417 14151 20451
rect 14550 20448 14556 20460
rect 14463 20420 14556 20448
rect 14093 20411 14151 20417
rect 14550 20408 14556 20420
rect 14608 20408 14614 20460
rect 15010 20408 15016 20460
rect 15068 20448 15074 20460
rect 16482 20448 16488 20460
rect 15068 20420 16488 20448
rect 15068 20408 15074 20420
rect 16482 20408 16488 20420
rect 16540 20408 16546 20460
rect 16666 20448 16672 20460
rect 16627 20420 16672 20448
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 18524 20457 18552 20488
rect 22186 20476 22192 20488
rect 22244 20476 22250 20528
rect 18509 20451 18567 20457
rect 18509 20417 18521 20451
rect 18555 20417 18567 20451
rect 18690 20448 18696 20460
rect 18651 20420 18696 20448
rect 18509 20411 18567 20417
rect 11112 20352 11744 20380
rect 11885 20383 11943 20389
rect 11112 20340 11118 20352
rect 11885 20349 11897 20383
rect 11931 20380 11943 20383
rect 11974 20380 11980 20392
rect 11931 20352 11980 20380
rect 11931 20349 11943 20352
rect 11885 20343 11943 20349
rect 11974 20340 11980 20352
rect 12032 20340 12038 20392
rect 15028 20380 15056 20408
rect 15562 20380 15568 20392
rect 13556 20352 15056 20380
rect 15523 20352 15568 20380
rect 6822 20272 6828 20324
rect 6880 20312 6886 20324
rect 8938 20312 8944 20324
rect 6880 20284 8944 20312
rect 6880 20272 6886 20284
rect 8938 20272 8944 20284
rect 8996 20312 9002 20324
rect 9490 20312 9496 20324
rect 8996 20284 9496 20312
rect 8996 20272 9002 20284
rect 9490 20272 9496 20284
rect 9548 20272 9554 20324
rect 13556 20321 13584 20352
rect 15562 20340 15568 20352
rect 15620 20340 15626 20392
rect 18524 20380 18552 20411
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 19794 20448 19800 20460
rect 18800 20420 19800 20448
rect 18598 20380 18604 20392
rect 18524 20352 18604 20380
rect 18598 20340 18604 20352
rect 18656 20340 18662 20392
rect 13541 20315 13599 20321
rect 13541 20281 13553 20315
rect 13587 20281 13599 20315
rect 13541 20275 13599 20281
rect 13722 20272 13728 20324
rect 13780 20312 13786 20324
rect 14415 20315 14473 20321
rect 14415 20312 14427 20315
rect 13780 20284 14427 20312
rect 13780 20272 13786 20284
rect 14415 20281 14427 20284
rect 14461 20281 14473 20315
rect 14415 20275 14473 20281
rect 14642 20272 14648 20324
rect 14700 20312 14706 20324
rect 18800 20312 18828 20420
rect 19794 20408 19800 20420
rect 19852 20408 19858 20460
rect 20346 20448 20352 20460
rect 20307 20420 20352 20448
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 20530 20448 20536 20460
rect 20491 20420 20536 20448
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 20625 20451 20683 20457
rect 20625 20417 20637 20451
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 20901 20451 20959 20457
rect 20901 20417 20913 20451
rect 20947 20448 20959 20451
rect 30098 20448 30104 20460
rect 20947 20420 21864 20448
rect 30059 20420 30104 20448
rect 20947 20417 20959 20420
rect 20901 20411 20959 20417
rect 19613 20383 19671 20389
rect 19613 20380 19625 20383
rect 14700 20284 18828 20312
rect 19076 20352 19625 20380
rect 14700 20272 14706 20284
rect 4338 20244 4344 20256
rect 3712 20216 4344 20244
rect 4338 20204 4344 20216
rect 4396 20204 4402 20256
rect 5074 20244 5080 20256
rect 5035 20216 5080 20244
rect 5074 20204 5080 20216
rect 5132 20204 5138 20256
rect 5629 20247 5687 20253
rect 5629 20213 5641 20247
rect 5675 20244 5687 20247
rect 6362 20244 6368 20256
rect 5675 20216 6368 20244
rect 5675 20213 5687 20216
rect 5629 20207 5687 20213
rect 6362 20204 6368 20216
rect 6420 20204 6426 20256
rect 7098 20244 7104 20256
rect 7059 20216 7104 20244
rect 7098 20204 7104 20216
rect 7156 20204 7162 20256
rect 8846 20204 8852 20256
rect 8904 20244 8910 20256
rect 9125 20247 9183 20253
rect 9125 20244 9137 20247
rect 8904 20216 9137 20244
rect 8904 20204 8910 20216
rect 9125 20213 9137 20216
rect 9171 20213 9183 20247
rect 9125 20207 9183 20213
rect 10226 20204 10232 20256
rect 10284 20244 10290 20256
rect 10689 20247 10747 20253
rect 10689 20244 10701 20247
rect 10284 20216 10701 20244
rect 10284 20204 10290 20216
rect 10689 20213 10701 20216
rect 10735 20213 10747 20247
rect 12250 20244 12256 20256
rect 12211 20216 12256 20244
rect 10689 20207 10747 20213
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 14090 20204 14096 20256
rect 14148 20244 14154 20256
rect 14185 20247 14243 20253
rect 14185 20244 14197 20247
rect 14148 20216 14197 20244
rect 14148 20204 14154 20216
rect 14185 20213 14197 20216
rect 14231 20213 14243 20247
rect 14185 20207 14243 20213
rect 14277 20247 14335 20253
rect 14277 20213 14289 20247
rect 14323 20244 14335 20247
rect 14826 20244 14832 20256
rect 14323 20216 14832 20244
rect 14323 20213 14335 20216
rect 14277 20207 14335 20213
rect 14826 20204 14832 20216
rect 14884 20204 14890 20256
rect 15013 20247 15071 20253
rect 15013 20213 15025 20247
rect 15059 20244 15071 20247
rect 15102 20244 15108 20256
rect 15059 20216 15108 20244
rect 15059 20213 15071 20216
rect 15013 20207 15071 20213
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 18509 20247 18567 20253
rect 18509 20213 18521 20247
rect 18555 20244 18567 20247
rect 19076 20244 19104 20352
rect 19613 20349 19625 20352
rect 19659 20349 19671 20383
rect 19613 20343 19671 20349
rect 19705 20383 19763 20389
rect 19705 20349 19717 20383
rect 19751 20380 19763 20383
rect 19978 20380 19984 20392
rect 19751 20352 19984 20380
rect 19751 20349 19763 20352
rect 19705 20343 19763 20349
rect 19334 20272 19340 20324
rect 19392 20312 19398 20324
rect 19720 20312 19748 20343
rect 19978 20340 19984 20352
rect 20036 20340 20042 20392
rect 20162 20340 20168 20392
rect 20220 20380 20226 20392
rect 20640 20380 20668 20411
rect 20220 20352 20668 20380
rect 20220 20340 20226 20352
rect 19392 20284 19748 20312
rect 19392 20272 19398 20284
rect 20438 20272 20444 20324
rect 20496 20312 20502 20324
rect 21836 20321 21864 20420
rect 30098 20408 30104 20420
rect 30156 20408 30162 20460
rect 22370 20380 22376 20392
rect 22331 20352 22376 20380
rect 22370 20340 22376 20352
rect 22428 20340 22434 20392
rect 21821 20315 21879 20321
rect 20496 20284 20852 20312
rect 20496 20272 20502 20284
rect 18555 20216 19104 20244
rect 19153 20247 19211 20253
rect 18555 20213 18567 20216
rect 18509 20207 18567 20213
rect 19153 20213 19165 20247
rect 19199 20244 19211 20247
rect 19426 20244 19432 20256
rect 19199 20216 19432 20244
rect 19199 20213 19211 20216
rect 19153 20207 19211 20213
rect 19426 20204 19432 20216
rect 19484 20204 19490 20256
rect 20349 20247 20407 20253
rect 20349 20213 20361 20247
rect 20395 20244 20407 20247
rect 20622 20244 20628 20256
rect 20395 20216 20628 20244
rect 20395 20213 20407 20216
rect 20349 20207 20407 20213
rect 20622 20204 20628 20216
rect 20680 20204 20686 20256
rect 20824 20253 20852 20284
rect 21821 20281 21833 20315
rect 21867 20281 21879 20315
rect 21821 20275 21879 20281
rect 20809 20247 20867 20253
rect 20809 20213 20821 20247
rect 20855 20244 20867 20247
rect 21726 20244 21732 20256
rect 20855 20216 21732 20244
rect 20855 20213 20867 20216
rect 20809 20207 20867 20213
rect 21726 20204 21732 20216
rect 21784 20204 21790 20256
rect 1104 20154 30820 20176
rect 1104 20102 5915 20154
rect 5967 20102 5979 20154
rect 6031 20102 6043 20154
rect 6095 20102 6107 20154
rect 6159 20102 6171 20154
rect 6223 20102 15846 20154
rect 15898 20102 15910 20154
rect 15962 20102 15974 20154
rect 16026 20102 16038 20154
rect 16090 20102 16102 20154
rect 16154 20102 25776 20154
rect 25828 20102 25840 20154
rect 25892 20102 25904 20154
rect 25956 20102 25968 20154
rect 26020 20102 26032 20154
rect 26084 20102 30820 20154
rect 1104 20080 30820 20102
rect 4522 20040 4528 20052
rect 4483 20012 4528 20040
rect 4522 20000 4528 20012
rect 4580 20000 4586 20052
rect 5629 20043 5687 20049
rect 5629 20009 5641 20043
rect 5675 20040 5687 20043
rect 6454 20040 6460 20052
rect 5675 20012 6460 20040
rect 5675 20009 5687 20012
rect 5629 20003 5687 20009
rect 6454 20000 6460 20012
rect 6512 20000 6518 20052
rect 8386 20000 8392 20052
rect 8444 20040 8450 20052
rect 9401 20043 9459 20049
rect 9401 20040 9413 20043
rect 8444 20012 9413 20040
rect 8444 20000 8450 20012
rect 9401 20009 9413 20012
rect 9447 20009 9459 20043
rect 10502 20040 10508 20052
rect 9401 20003 9459 20009
rect 9508 20012 10508 20040
rect 4338 19932 4344 19984
rect 4396 19932 4402 19984
rect 6546 19932 6552 19984
rect 6604 19972 6610 19984
rect 7561 19975 7619 19981
rect 7561 19972 7573 19975
rect 6604 19944 7573 19972
rect 6604 19932 6610 19944
rect 7561 19941 7573 19944
rect 7607 19941 7619 19975
rect 7561 19935 7619 19941
rect 4157 19907 4215 19913
rect 4157 19873 4169 19907
rect 4203 19904 4215 19907
rect 4356 19904 4384 19932
rect 6451 19907 6509 19913
rect 6451 19904 6463 19907
rect 4203 19876 4384 19904
rect 5736 19876 6463 19904
rect 4203 19873 4215 19876
rect 4157 19867 4215 19873
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19836 1823 19839
rect 1854 19836 1860 19848
rect 1811 19808 1860 19836
rect 1811 19805 1823 19808
rect 1765 19799 1823 19805
rect 1854 19796 1860 19808
rect 1912 19836 1918 19848
rect 3694 19836 3700 19848
rect 1912 19808 3700 19836
rect 1912 19796 1918 19808
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 3789 19839 3847 19845
rect 3789 19805 3801 19839
rect 3835 19805 3847 19839
rect 3970 19836 3976 19848
rect 3931 19808 3976 19836
rect 3789 19799 3847 19805
rect 2032 19771 2090 19777
rect 2032 19737 2044 19771
rect 2078 19768 2090 19771
rect 2222 19768 2228 19780
rect 2078 19740 2228 19768
rect 2078 19737 2090 19740
rect 2032 19731 2090 19737
rect 2222 19728 2228 19740
rect 2280 19728 2286 19780
rect 3510 19728 3516 19780
rect 3568 19768 3574 19780
rect 3804 19768 3832 19799
rect 3970 19796 3976 19808
rect 4028 19796 4034 19848
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19805 4123 19839
rect 4065 19799 4123 19805
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19836 4399 19839
rect 5074 19836 5080 19848
rect 4387 19808 5080 19836
rect 4387 19805 4399 19808
rect 4341 19799 4399 19805
rect 3568 19740 3832 19768
rect 4080 19768 4108 19799
rect 5074 19796 5080 19808
rect 5132 19796 5138 19848
rect 5626 19796 5632 19848
rect 5684 19796 5690 19848
rect 5736 19845 5764 19876
rect 6451 19873 6463 19876
rect 6497 19904 6509 19907
rect 6564 19904 6592 19932
rect 9508 19904 9536 20012
rect 10502 20000 10508 20012
rect 10560 20000 10566 20052
rect 12894 20040 12900 20052
rect 12855 20012 12900 20040
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 13449 20043 13507 20049
rect 13449 20009 13461 20043
rect 13495 20040 13507 20043
rect 13538 20040 13544 20052
rect 13495 20012 13544 20040
rect 13495 20009 13507 20012
rect 13449 20003 13507 20009
rect 9861 19975 9919 19981
rect 9861 19941 9873 19975
rect 9907 19972 9919 19975
rect 10413 19975 10471 19981
rect 10413 19972 10425 19975
rect 9907 19944 10425 19972
rect 9907 19941 9919 19944
rect 9861 19935 9919 19941
rect 10413 19941 10425 19944
rect 10459 19941 10471 19975
rect 10413 19935 10471 19941
rect 10042 19904 10048 19916
rect 6497 19876 6592 19904
rect 7668 19876 9536 19904
rect 9600 19876 10048 19904
rect 6497 19873 6509 19876
rect 6451 19867 6509 19873
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19805 5779 19839
rect 5721 19799 5779 19805
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19836 6239 19839
rect 6270 19836 6276 19848
rect 6227 19808 6276 19836
rect 6227 19805 6239 19808
rect 6181 19799 6239 19805
rect 6270 19796 6276 19808
rect 6328 19796 6334 19848
rect 6365 19839 6423 19845
rect 6365 19805 6377 19839
rect 6411 19805 6423 19839
rect 6546 19836 6552 19848
rect 6507 19808 6552 19836
rect 6365 19799 6423 19805
rect 4522 19768 4528 19780
rect 4080 19740 4528 19768
rect 3568 19728 3574 19740
rect 4522 19728 4528 19740
rect 4580 19728 4586 19780
rect 5644 19768 5672 19796
rect 6380 19768 6408 19799
rect 6546 19796 6552 19808
rect 6604 19796 6610 19848
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 6914 19836 6920 19848
rect 6779 19808 6920 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 6914 19796 6920 19808
rect 6972 19796 6978 19848
rect 7668 19768 7696 19876
rect 7745 19839 7803 19845
rect 7745 19805 7757 19839
rect 7791 19836 7803 19839
rect 8478 19836 8484 19848
rect 7791 19808 8484 19836
rect 7791 19805 7803 19808
rect 7745 19799 7803 19805
rect 8478 19796 8484 19808
rect 8536 19796 8542 19848
rect 9600 19845 9628 19876
rect 10042 19864 10048 19876
rect 10100 19864 10106 19916
rect 10597 19907 10655 19913
rect 10597 19873 10609 19907
rect 10643 19904 10655 19907
rect 10778 19904 10784 19916
rect 10643 19876 10784 19904
rect 10643 19873 10655 19876
rect 10597 19867 10655 19873
rect 10778 19864 10784 19876
rect 10836 19864 10842 19916
rect 11514 19904 11520 19916
rect 11475 19876 11520 19904
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 13464 19904 13492 20003
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 13906 20000 13912 20052
rect 13964 20040 13970 20052
rect 13964 20012 16528 20040
rect 13964 20000 13970 20012
rect 13814 19932 13820 19984
rect 13872 19972 13878 19984
rect 14274 19972 14280 19984
rect 13872 19944 14280 19972
rect 13872 19932 13878 19944
rect 14274 19932 14280 19944
rect 14332 19972 14338 19984
rect 14642 19972 14648 19984
rect 14332 19944 14648 19972
rect 14332 19932 14338 19944
rect 14642 19932 14648 19944
rect 14700 19932 14706 19984
rect 15562 19932 15568 19984
rect 15620 19972 15626 19984
rect 16500 19972 16528 20012
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 16669 20043 16727 20049
rect 16669 20040 16681 20043
rect 16632 20012 16681 20040
rect 16632 20000 16638 20012
rect 16669 20009 16681 20012
rect 16715 20009 16727 20043
rect 20162 20040 20168 20052
rect 20123 20012 20168 20040
rect 16669 20003 16727 20009
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 20254 20000 20260 20052
rect 20312 20040 20318 20052
rect 20625 20043 20683 20049
rect 20625 20040 20637 20043
rect 20312 20012 20637 20040
rect 20312 20000 20318 20012
rect 20625 20009 20637 20012
rect 20671 20009 20683 20043
rect 20625 20003 20683 20009
rect 18874 19972 18880 19984
rect 15620 19944 16436 19972
rect 16500 19944 18880 19972
rect 15620 19932 15626 19944
rect 13280 19876 13492 19904
rect 9585 19839 9643 19845
rect 9585 19805 9597 19839
rect 9631 19805 9643 19839
rect 9585 19799 9643 19805
rect 9677 19839 9735 19845
rect 9677 19805 9689 19839
rect 9723 19805 9735 19839
rect 9677 19799 9735 19805
rect 5644 19740 6408 19768
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 2774 19700 2780 19712
rect 1728 19672 2780 19700
rect 1728 19660 1734 19672
rect 2774 19660 2780 19672
rect 2832 19660 2838 19712
rect 3142 19700 3148 19712
rect 3055 19672 3148 19700
rect 3142 19660 3148 19672
rect 3200 19700 3206 19712
rect 5258 19700 5264 19712
rect 3200 19672 5264 19700
rect 3200 19660 3206 19672
rect 5258 19660 5264 19672
rect 5316 19660 5322 19712
rect 6380 19700 6408 19740
rect 6564 19740 7696 19768
rect 6564 19700 6592 19740
rect 7834 19728 7840 19780
rect 7892 19768 7898 19780
rect 7929 19771 7987 19777
rect 7929 19768 7941 19771
rect 7892 19740 7941 19768
rect 7892 19728 7898 19740
rect 7929 19737 7941 19740
rect 7975 19737 7987 19771
rect 7929 19731 7987 19737
rect 8846 19728 8852 19780
rect 8904 19768 8910 19780
rect 9692 19768 9720 19799
rect 9858 19796 9864 19848
rect 9916 19836 9922 19848
rect 9953 19839 10011 19845
rect 9953 19836 9965 19839
rect 9916 19808 9965 19836
rect 9916 19796 9922 19808
rect 9953 19805 9965 19808
rect 9999 19805 10011 19839
rect 9953 19799 10011 19805
rect 10318 19796 10324 19848
rect 10376 19836 10382 19848
rect 10689 19839 10747 19845
rect 10689 19836 10701 19839
rect 10376 19808 10701 19836
rect 10376 19796 10382 19808
rect 10689 19805 10701 19808
rect 10735 19836 10747 19839
rect 10965 19839 11023 19845
rect 10965 19836 10977 19839
rect 10735 19808 10977 19836
rect 10735 19805 10747 19808
rect 10689 19799 10747 19805
rect 10965 19805 10977 19808
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 11784 19839 11842 19845
rect 11784 19805 11796 19839
rect 11830 19836 11842 19839
rect 12250 19836 12256 19848
rect 11830 19808 12256 19836
rect 11830 19805 11842 19808
rect 11784 19799 11842 19805
rect 12250 19796 12256 19808
rect 12308 19796 12314 19848
rect 8904 19740 9720 19768
rect 11057 19771 11115 19777
rect 8904 19728 8910 19740
rect 11057 19737 11069 19771
rect 11103 19768 11115 19771
rect 13280 19768 13308 19876
rect 13722 19864 13728 19916
rect 13780 19904 13786 19916
rect 14461 19907 14519 19913
rect 14461 19904 14473 19907
rect 13780 19876 14473 19904
rect 13780 19864 13786 19876
rect 14461 19873 14473 19876
rect 14507 19873 14519 19907
rect 14461 19867 14519 19873
rect 15838 19864 15844 19916
rect 15896 19904 15902 19916
rect 16025 19907 16083 19913
rect 15896 19876 15941 19904
rect 15896 19864 15902 19876
rect 16025 19873 16037 19907
rect 16071 19904 16083 19907
rect 16298 19904 16304 19916
rect 16071 19876 16304 19904
rect 16071 19873 16083 19876
rect 16025 19867 16083 19873
rect 16298 19864 16304 19876
rect 16356 19864 16362 19916
rect 16408 19904 16436 19944
rect 18874 19932 18880 19944
rect 18932 19932 18938 19984
rect 17865 19907 17923 19913
rect 17865 19904 17877 19907
rect 16408 19876 17877 19904
rect 17865 19873 17877 19876
rect 17911 19904 17923 19907
rect 19334 19904 19340 19916
rect 17911 19876 19340 19904
rect 17911 19873 17923 19876
rect 17865 19867 17923 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 20272 19904 20300 20000
rect 19444 19876 20300 19904
rect 20732 19876 21404 19904
rect 13538 19836 13544 19848
rect 13499 19808 13544 19836
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 14090 19836 14096 19848
rect 14051 19808 14096 19836
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14274 19836 14280 19848
rect 14235 19808 14280 19836
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19805 14427 19839
rect 14550 19836 14556 19848
rect 14511 19808 14556 19836
rect 14369 19799 14427 19805
rect 11103 19740 13308 19768
rect 14384 19768 14412 19799
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 15746 19836 15752 19848
rect 15707 19808 15752 19836
rect 15746 19796 15752 19808
rect 15804 19796 15810 19848
rect 15930 19836 15936 19848
rect 15891 19808 15936 19836
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 16758 19836 16764 19848
rect 16719 19808 16764 19836
rect 16758 19796 16764 19808
rect 16816 19796 16822 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19836 17739 19839
rect 17954 19836 17960 19848
rect 17727 19808 17960 19836
rect 17727 19805 17739 19808
rect 17681 19799 17739 19805
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 19444 19845 19472 19876
rect 19429 19839 19487 19845
rect 19429 19805 19441 19839
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 19886 19796 19892 19848
rect 19944 19836 19950 19848
rect 20732 19845 20760 19876
rect 21376 19848 21404 19876
rect 20349 19839 20407 19845
rect 20349 19836 20361 19839
rect 19944 19808 20361 19836
rect 19944 19796 19950 19808
rect 20349 19805 20361 19808
rect 20395 19805 20407 19839
rect 20349 19799 20407 19805
rect 20441 19839 20499 19845
rect 20441 19805 20453 19839
rect 20487 19805 20499 19839
rect 20441 19799 20499 19805
rect 20717 19839 20775 19845
rect 20717 19805 20729 19839
rect 20763 19805 20775 19839
rect 20717 19799 20775 19805
rect 19337 19771 19395 19777
rect 19337 19768 19349 19771
rect 14384 19740 19349 19768
rect 11103 19737 11115 19740
rect 11057 19731 11115 19737
rect 19337 19737 19349 19740
rect 19383 19737 19395 19771
rect 20456 19768 20484 19799
rect 20806 19796 20812 19848
rect 20864 19836 20870 19848
rect 21177 19839 21235 19845
rect 21177 19836 21189 19839
rect 20864 19808 21189 19836
rect 20864 19796 20870 19808
rect 21177 19805 21189 19808
rect 21223 19805 21235 19839
rect 21358 19836 21364 19848
rect 21319 19808 21364 19836
rect 21177 19799 21235 19805
rect 21358 19796 21364 19808
rect 21416 19796 21422 19848
rect 21082 19768 21088 19780
rect 20456 19740 21088 19768
rect 19337 19731 19395 19737
rect 21082 19728 21088 19740
rect 21140 19728 21146 19780
rect 6380 19672 6592 19700
rect 6917 19703 6975 19709
rect 6917 19669 6929 19703
rect 6963 19700 6975 19703
rect 7006 19700 7012 19712
rect 6963 19672 7012 19700
rect 6963 19669 6975 19672
rect 6917 19663 6975 19669
rect 7006 19660 7012 19672
rect 7064 19660 7070 19712
rect 8386 19660 8392 19712
rect 8444 19700 8450 19712
rect 8938 19700 8944 19712
rect 8444 19672 8944 19700
rect 8444 19660 8450 19672
rect 8938 19660 8944 19672
rect 8996 19660 9002 19712
rect 14734 19700 14740 19712
rect 14695 19672 14740 19700
rect 14734 19660 14740 19672
rect 14792 19660 14798 19712
rect 15378 19660 15384 19712
rect 15436 19700 15442 19712
rect 15565 19703 15623 19709
rect 15565 19700 15577 19703
rect 15436 19672 15577 19700
rect 15436 19660 15442 19672
rect 15565 19669 15577 19672
rect 15611 19669 15623 19703
rect 17310 19700 17316 19712
rect 17271 19672 17316 19700
rect 15565 19663 15623 19669
rect 17310 19660 17316 19672
rect 17368 19660 17374 19712
rect 17770 19660 17776 19712
rect 17828 19700 17834 19712
rect 17828 19672 17873 19700
rect 17828 19660 17834 19672
rect 20714 19660 20720 19712
rect 20772 19700 20778 19712
rect 21269 19703 21327 19709
rect 21269 19700 21281 19703
rect 20772 19672 21281 19700
rect 20772 19660 20778 19672
rect 21269 19669 21281 19672
rect 21315 19669 21327 19703
rect 21269 19663 21327 19669
rect 1104 19610 30820 19632
rect 1104 19558 10880 19610
rect 10932 19558 10944 19610
rect 10996 19558 11008 19610
rect 11060 19558 11072 19610
rect 11124 19558 11136 19610
rect 11188 19558 20811 19610
rect 20863 19558 20875 19610
rect 20927 19558 20939 19610
rect 20991 19558 21003 19610
rect 21055 19558 21067 19610
rect 21119 19558 30820 19610
rect 1104 19536 30820 19558
rect 1302 19456 1308 19508
rect 1360 19496 1366 19508
rect 1360 19468 2774 19496
rect 1360 19456 1366 19468
rect 1762 19388 1768 19440
rect 1820 19428 1826 19440
rect 2222 19428 2228 19440
rect 1820 19400 1900 19428
rect 2183 19400 2228 19428
rect 1820 19388 1826 19400
rect 1486 19360 1492 19372
rect 1447 19332 1492 19360
rect 1486 19320 1492 19332
rect 1544 19320 1550 19372
rect 1670 19360 1676 19372
rect 1631 19332 1676 19360
rect 1670 19320 1676 19332
rect 1728 19320 1734 19372
rect 1872 19369 1900 19400
rect 2222 19388 2228 19400
rect 2280 19388 2286 19440
rect 2746 19428 2774 19468
rect 6730 19456 6736 19508
rect 6788 19496 6794 19508
rect 8202 19496 8208 19508
rect 6788 19468 8208 19496
rect 6788 19456 6794 19468
rect 8202 19456 8208 19468
rect 8260 19456 8266 19508
rect 9858 19456 9864 19508
rect 9916 19496 9922 19508
rect 10410 19496 10416 19508
rect 9916 19468 10416 19496
rect 9916 19456 9922 19468
rect 10410 19456 10416 19468
rect 10468 19456 10474 19508
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 13170 19496 13176 19508
rect 12492 19468 13176 19496
rect 12492 19456 12498 19468
rect 13170 19456 13176 19468
rect 13228 19456 13234 19508
rect 13538 19456 13544 19508
rect 13596 19496 13602 19508
rect 14093 19499 14151 19505
rect 14093 19496 14105 19499
rect 13596 19468 14105 19496
rect 13596 19456 13602 19468
rect 14093 19465 14105 19468
rect 14139 19465 14151 19499
rect 16666 19496 16672 19508
rect 16627 19468 16672 19496
rect 14093 19459 14151 19465
rect 16666 19456 16672 19468
rect 16724 19456 16730 19508
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 17494 19496 17500 19508
rect 16816 19468 17500 19496
rect 16816 19456 16822 19468
rect 17494 19456 17500 19468
rect 17552 19456 17558 19508
rect 17589 19499 17647 19505
rect 17589 19465 17601 19499
rect 17635 19496 17647 19499
rect 17770 19496 17776 19508
rect 17635 19468 17776 19496
rect 17635 19465 17647 19468
rect 17589 19459 17647 19465
rect 17770 19456 17776 19468
rect 17828 19456 17834 19508
rect 18322 19456 18328 19508
rect 18380 19496 18386 19508
rect 18785 19499 18843 19505
rect 18785 19496 18797 19499
rect 18380 19468 18797 19496
rect 18380 19456 18386 19468
rect 18785 19465 18797 19468
rect 18831 19465 18843 19499
rect 18785 19459 18843 19465
rect 18966 19456 18972 19508
rect 19024 19496 19030 19508
rect 19153 19499 19211 19505
rect 19153 19496 19165 19499
rect 19024 19468 19165 19496
rect 19024 19456 19030 19468
rect 19153 19465 19165 19468
rect 19199 19465 19211 19499
rect 20714 19496 20720 19508
rect 20675 19468 20720 19496
rect 19153 19459 19211 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 30006 19496 30012 19508
rect 29967 19468 30012 19496
rect 30006 19456 30012 19468
rect 30064 19456 30070 19508
rect 11885 19431 11943 19437
rect 11885 19428 11897 19431
rect 2746 19400 11897 19428
rect 11885 19397 11897 19400
rect 11931 19397 11943 19431
rect 11885 19391 11943 19397
rect 14734 19388 14740 19440
rect 14792 19428 14798 19440
rect 15206 19431 15264 19437
rect 15206 19428 15218 19431
rect 14792 19400 15218 19428
rect 14792 19388 14798 19400
rect 15206 19397 15218 19400
rect 15252 19397 15264 19431
rect 18049 19431 18107 19437
rect 18049 19428 18061 19431
rect 15206 19391 15264 19397
rect 15304 19400 18061 19428
rect 1857 19363 1915 19369
rect 1857 19329 1869 19363
rect 1903 19329 1915 19363
rect 1857 19323 1915 19329
rect 2041 19363 2099 19369
rect 2041 19329 2053 19363
rect 2087 19360 2099 19363
rect 3510 19360 3516 19372
rect 2087 19332 2820 19360
rect 2087 19329 2099 19332
rect 2041 19323 2099 19329
rect 1578 19252 1584 19304
rect 1636 19292 1642 19304
rect 1765 19295 1823 19301
rect 1765 19292 1777 19295
rect 1636 19264 1777 19292
rect 1636 19252 1642 19264
rect 1765 19261 1777 19264
rect 1811 19292 1823 19295
rect 1811 19264 2084 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 2056 19236 2084 19264
rect 2038 19184 2044 19236
rect 2096 19184 2102 19236
rect 2792 19224 2820 19332
rect 3252 19332 3516 19360
rect 3142 19224 3148 19236
rect 2792 19196 3148 19224
rect 3142 19184 3148 19196
rect 3200 19184 3206 19236
rect 1486 19116 1492 19168
rect 1544 19156 1550 19168
rect 3252 19156 3280 19332
rect 3510 19320 3516 19332
rect 3568 19320 3574 19372
rect 3694 19320 3700 19372
rect 3752 19360 3758 19372
rect 4249 19363 4307 19369
rect 4249 19360 4261 19363
rect 3752 19332 4261 19360
rect 3752 19320 3758 19332
rect 4249 19329 4261 19332
rect 4295 19329 4307 19363
rect 4249 19323 4307 19329
rect 4516 19363 4574 19369
rect 4516 19329 4528 19363
rect 4562 19360 4574 19363
rect 4798 19360 4804 19372
rect 4562 19332 4804 19360
rect 4562 19329 4574 19332
rect 4516 19323 4574 19329
rect 4798 19320 4804 19332
rect 4856 19320 4862 19372
rect 6825 19363 6883 19369
rect 6825 19329 6837 19363
rect 6871 19360 6883 19363
rect 6914 19360 6920 19372
rect 6871 19332 6920 19360
rect 6871 19329 6883 19332
rect 6825 19323 6883 19329
rect 6914 19320 6920 19332
rect 6972 19320 6978 19372
rect 7098 19369 7104 19372
rect 7092 19360 7104 19369
rect 7059 19332 7104 19360
rect 7092 19323 7104 19332
rect 7098 19320 7104 19323
rect 7156 19320 7162 19372
rect 7926 19320 7932 19372
rect 7984 19360 7990 19372
rect 9214 19360 9220 19372
rect 7984 19332 8800 19360
rect 9127 19332 9220 19360
rect 7984 19320 7990 19332
rect 3786 19292 3792 19304
rect 3747 19264 3792 19292
rect 3786 19252 3792 19264
rect 3844 19252 3850 19304
rect 8772 19301 8800 19332
rect 9214 19320 9220 19332
rect 9272 19360 9278 19372
rect 10229 19363 10287 19369
rect 9272 19332 10180 19360
rect 9272 19320 9278 19332
rect 8757 19295 8815 19301
rect 8757 19261 8769 19295
rect 8803 19261 8815 19295
rect 8757 19255 8815 19261
rect 9306 19252 9312 19304
rect 9364 19292 9370 19304
rect 10045 19295 10103 19301
rect 10045 19292 10057 19295
rect 9364 19264 10057 19292
rect 9364 19252 9370 19264
rect 10045 19261 10057 19264
rect 10091 19261 10103 19295
rect 10152 19292 10180 19332
rect 10229 19329 10241 19363
rect 10275 19360 10287 19363
rect 10318 19360 10324 19372
rect 10275 19332 10324 19360
rect 10275 19329 10287 19332
rect 10229 19323 10287 19329
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 10410 19320 10416 19372
rect 10468 19360 10474 19372
rect 15304 19360 15332 19400
rect 18049 19397 18061 19400
rect 18095 19397 18107 19431
rect 18049 19391 18107 19397
rect 19334 19388 19340 19440
rect 19392 19428 19398 19440
rect 20622 19428 20628 19440
rect 19392 19400 19472 19428
rect 20583 19400 20628 19428
rect 19392 19388 19398 19400
rect 15470 19360 15476 19372
rect 10468 19332 10513 19360
rect 10612 19332 15332 19360
rect 15431 19332 15476 19360
rect 10468 19320 10474 19332
rect 10612 19292 10640 19332
rect 15470 19320 15476 19332
rect 15528 19320 15534 19372
rect 16758 19320 16764 19372
rect 16816 19360 16822 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16816 19332 16865 19360
rect 16816 19320 16822 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16853 19323 16911 19329
rect 16960 19332 17049 19360
rect 10152 19264 10640 19292
rect 10045 19255 10103 19261
rect 16206 19252 16212 19304
rect 16264 19292 16270 19304
rect 16960 19292 16988 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17954 19360 17960 19372
rect 17915 19332 17960 19360
rect 17037 19323 17095 19329
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 19242 19320 19248 19372
rect 19300 19360 19306 19372
rect 19300 19332 19345 19360
rect 19300 19320 19306 19332
rect 16264 19264 16988 19292
rect 18233 19295 18291 19301
rect 16264 19252 16270 19264
rect 18233 19261 18245 19295
rect 18279 19292 18291 19295
rect 18598 19292 18604 19304
rect 18279 19264 18604 19292
rect 18279 19261 18291 19264
rect 18233 19255 18291 19261
rect 6546 19184 6552 19236
rect 6604 19224 6610 19236
rect 6822 19224 6828 19236
rect 6604 19196 6828 19224
rect 6604 19184 6610 19196
rect 6822 19184 6828 19196
rect 6880 19184 6886 19236
rect 15930 19184 15936 19236
rect 15988 19184 15994 19236
rect 16482 19184 16488 19236
rect 16540 19224 16546 19236
rect 18248 19224 18276 19255
rect 18598 19252 18604 19264
rect 18656 19252 18662 19304
rect 19334 19292 19340 19304
rect 19295 19264 19340 19292
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 19444 19292 19472 19400
rect 20622 19388 20628 19400
rect 20680 19388 20686 19440
rect 29825 19363 29883 19369
rect 29825 19329 29837 19363
rect 29871 19360 29883 19363
rect 29914 19360 29920 19372
rect 29871 19332 29920 19360
rect 29871 19329 29883 19332
rect 29825 19323 29883 19329
rect 29914 19320 29920 19332
rect 29972 19320 29978 19372
rect 20809 19295 20867 19301
rect 20809 19292 20821 19295
rect 19444 19264 20821 19292
rect 20809 19261 20821 19264
rect 20855 19261 20867 19295
rect 20809 19255 20867 19261
rect 16540 19196 18276 19224
rect 19352 19224 19380 19252
rect 19610 19224 19616 19236
rect 19352 19196 19616 19224
rect 16540 19184 16546 19196
rect 19610 19184 19616 19196
rect 19668 19184 19674 19236
rect 20530 19224 20536 19236
rect 19720 19196 20536 19224
rect 5626 19156 5632 19168
rect 1544 19128 3280 19156
rect 5539 19128 5632 19156
rect 1544 19116 1550 19128
rect 5626 19116 5632 19128
rect 5684 19156 5690 19168
rect 6454 19156 6460 19168
rect 5684 19128 6460 19156
rect 5684 19116 5690 19128
rect 6454 19116 6460 19128
rect 6512 19116 6518 19168
rect 8846 19116 8852 19168
rect 8904 19156 8910 19168
rect 8941 19159 8999 19165
rect 8941 19156 8953 19159
rect 8904 19128 8953 19156
rect 8904 19116 8910 19128
rect 8941 19125 8953 19128
rect 8987 19125 8999 19159
rect 8941 19119 8999 19125
rect 14826 19116 14832 19168
rect 14884 19156 14890 19168
rect 15948 19156 15976 19184
rect 19720 19156 19748 19196
rect 20530 19184 20536 19196
rect 20588 19184 20594 19236
rect 20254 19156 20260 19168
rect 14884 19128 19748 19156
rect 20215 19128 20260 19156
rect 14884 19116 14890 19128
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 1104 19066 30820 19088
rect 1104 19014 5915 19066
rect 5967 19014 5979 19066
rect 6031 19014 6043 19066
rect 6095 19014 6107 19066
rect 6159 19014 6171 19066
rect 6223 19014 15846 19066
rect 15898 19014 15910 19066
rect 15962 19014 15974 19066
rect 16026 19014 16038 19066
rect 16090 19014 16102 19066
rect 16154 19014 25776 19066
rect 25828 19014 25840 19066
rect 25892 19014 25904 19066
rect 25956 19014 25968 19066
rect 26020 19014 26032 19066
rect 26084 19014 30820 19066
rect 1104 18992 30820 19014
rect 4798 18952 4804 18964
rect 4759 18924 4804 18952
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 5810 18912 5816 18964
rect 5868 18952 5874 18964
rect 5905 18955 5963 18961
rect 5905 18952 5917 18955
rect 5868 18924 5917 18952
rect 5868 18912 5874 18924
rect 5905 18921 5917 18924
rect 5951 18921 5963 18955
rect 10042 18952 10048 18964
rect 5905 18915 5963 18921
rect 6012 18924 10048 18952
rect 4338 18844 4344 18896
rect 4396 18884 4402 18896
rect 4396 18856 4476 18884
rect 4396 18844 4402 18856
rect 1854 18816 1860 18828
rect 1815 18788 1860 18816
rect 1854 18776 1860 18788
rect 1912 18776 1918 18828
rect 4448 18825 4476 18856
rect 4522 18844 4528 18896
rect 4580 18884 4586 18896
rect 6012 18884 6040 18924
rect 10042 18912 10048 18924
rect 10100 18912 10106 18964
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 18141 18955 18199 18961
rect 18141 18952 18153 18955
rect 18012 18924 18153 18952
rect 18012 18912 18018 18924
rect 18141 18921 18153 18924
rect 18187 18921 18199 18955
rect 18141 18915 18199 18921
rect 18690 18912 18696 18964
rect 18748 18952 18754 18964
rect 19245 18955 19303 18961
rect 19245 18952 19257 18955
rect 18748 18924 19257 18952
rect 18748 18912 18754 18924
rect 19245 18921 19257 18924
rect 19291 18921 19303 18955
rect 19245 18915 19303 18921
rect 21085 18955 21143 18961
rect 21085 18921 21097 18955
rect 21131 18952 21143 18955
rect 21358 18952 21364 18964
rect 21131 18924 21364 18952
rect 21131 18921 21143 18924
rect 21085 18915 21143 18921
rect 21358 18912 21364 18924
rect 21416 18912 21422 18964
rect 4580 18856 6040 18884
rect 4580 18844 4586 18856
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18785 4491 18819
rect 4433 18779 4491 18785
rect 4065 18751 4123 18757
rect 4065 18717 4077 18751
rect 4111 18717 4123 18751
rect 4246 18748 4252 18760
rect 4207 18720 4252 18748
rect 4065 18711 4123 18717
rect 2124 18683 2182 18689
rect 2124 18649 2136 18683
rect 2170 18680 2182 18683
rect 2498 18680 2504 18692
rect 2170 18652 2504 18680
rect 2170 18649 2182 18652
rect 2124 18643 2182 18649
rect 2498 18640 2504 18652
rect 2556 18640 2562 18692
rect 4080 18680 4108 18711
rect 4246 18708 4252 18720
rect 4304 18708 4310 18760
rect 4341 18751 4399 18757
rect 4341 18717 4353 18751
rect 4387 18748 4399 18751
rect 4540 18748 4568 18844
rect 5626 18816 5632 18828
rect 4632 18788 5632 18816
rect 4632 18757 4660 18788
rect 5626 18776 5632 18788
rect 5684 18776 5690 18828
rect 9217 18819 9275 18825
rect 9217 18785 9229 18819
rect 9263 18816 9275 18819
rect 9398 18816 9404 18828
rect 9263 18788 9404 18816
rect 9263 18785 9275 18788
rect 9217 18779 9275 18785
rect 9398 18776 9404 18788
rect 9456 18776 9462 18828
rect 11422 18816 11428 18828
rect 9508 18788 11428 18816
rect 4387 18720 4568 18748
rect 4617 18751 4675 18757
rect 4387 18717 4399 18720
rect 4341 18711 4399 18717
rect 4617 18717 4629 18751
rect 4663 18717 4675 18751
rect 5258 18748 5264 18760
rect 5219 18720 5264 18748
rect 4617 18711 4675 18717
rect 5258 18708 5264 18720
rect 5316 18708 5322 18760
rect 7285 18751 7343 18757
rect 7285 18748 7297 18751
rect 6932 18720 7297 18748
rect 6932 18692 6960 18720
rect 7285 18717 7297 18720
rect 7331 18748 7343 18751
rect 8202 18748 8208 18760
rect 7331 18720 8208 18748
rect 7331 18717 7343 18720
rect 7285 18711 7343 18717
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 8938 18748 8944 18760
rect 8899 18720 8944 18748
rect 8938 18708 8944 18720
rect 8996 18708 9002 18760
rect 9125 18751 9183 18757
rect 9125 18717 9137 18751
rect 9171 18717 9183 18751
rect 9306 18748 9312 18760
rect 9267 18720 9312 18748
rect 9125 18711 9183 18717
rect 4982 18680 4988 18692
rect 4080 18652 4988 18680
rect 4982 18640 4988 18652
rect 5040 18640 5046 18692
rect 6914 18640 6920 18692
rect 6972 18640 6978 18692
rect 7006 18640 7012 18692
rect 7064 18689 7070 18692
rect 7064 18680 7076 18689
rect 7064 18652 7109 18680
rect 7064 18643 7076 18652
rect 7064 18640 7070 18643
rect 8110 18640 8116 18692
rect 8168 18680 8174 18692
rect 8754 18680 8760 18692
rect 8168 18652 8760 18680
rect 8168 18640 8174 18652
rect 8754 18640 8760 18652
rect 8812 18680 8818 18692
rect 9140 18680 9168 18711
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 9508 18757 9536 18788
rect 11422 18776 11428 18788
rect 11480 18776 11486 18828
rect 15013 18819 15071 18825
rect 15013 18785 15025 18819
rect 15059 18816 15071 18819
rect 16482 18816 16488 18828
rect 15059 18788 16488 18816
rect 15059 18785 15071 18788
rect 15013 18779 15071 18785
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 16666 18816 16672 18828
rect 16627 18788 16672 18816
rect 16666 18776 16672 18788
rect 16724 18816 16730 18828
rect 19334 18816 19340 18828
rect 16724 18788 19340 18816
rect 16724 18776 16730 18788
rect 19334 18776 19340 18788
rect 19392 18816 19398 18828
rect 19797 18819 19855 18825
rect 19797 18816 19809 18819
rect 19392 18788 19809 18816
rect 19392 18776 19398 18788
rect 19797 18785 19809 18788
rect 19843 18816 19855 18819
rect 21637 18819 21695 18825
rect 21637 18816 21649 18819
rect 19843 18788 21649 18816
rect 19843 18785 19855 18788
rect 19797 18779 19855 18785
rect 21637 18785 21649 18788
rect 21683 18785 21695 18819
rect 21637 18779 21695 18785
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18717 9551 18751
rect 9493 18711 9551 18717
rect 10594 18708 10600 18760
rect 10652 18748 10658 18760
rect 10781 18751 10839 18757
rect 10781 18748 10793 18751
rect 10652 18720 10793 18748
rect 10652 18708 10658 18720
rect 10781 18717 10793 18720
rect 10827 18748 10839 18751
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 10827 18720 11253 18748
rect 10827 18717 10839 18720
rect 10781 18711 10839 18717
rect 11241 18717 11253 18720
rect 11287 18717 11299 18751
rect 12526 18748 12532 18760
rect 12487 18720 12532 18748
rect 11241 18711 11299 18717
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 12713 18751 12771 18757
rect 12713 18717 12725 18751
rect 12759 18748 12771 18751
rect 13998 18748 14004 18760
rect 12759 18720 14004 18748
rect 12759 18717 12771 18720
rect 12713 18711 12771 18717
rect 13998 18708 14004 18720
rect 14056 18708 14062 18760
rect 14369 18751 14427 18757
rect 14369 18717 14381 18751
rect 14415 18748 14427 18751
rect 14415 18720 15608 18748
rect 14415 18717 14427 18720
rect 14369 18711 14427 18717
rect 8812 18652 9168 18680
rect 14093 18683 14151 18689
rect 8812 18640 8818 18652
rect 14093 18649 14105 18683
rect 14139 18680 14151 18683
rect 15197 18683 15255 18689
rect 15197 18680 15209 18683
rect 14139 18652 15209 18680
rect 14139 18649 14151 18652
rect 14093 18643 14151 18649
rect 15197 18649 15209 18652
rect 15243 18649 15255 18683
rect 15580 18680 15608 18720
rect 15654 18708 15660 18760
rect 15712 18748 15718 18760
rect 16206 18748 16212 18760
rect 15712 18720 16212 18748
rect 15712 18708 15718 18720
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 18322 18748 18328 18760
rect 18283 18720 18328 18748
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 19702 18748 19708 18760
rect 19659 18720 19708 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 19702 18708 19708 18720
rect 19760 18708 19766 18760
rect 20438 18748 20444 18760
rect 20399 18720 20444 18748
rect 20438 18708 20444 18720
rect 20496 18708 20502 18760
rect 22186 18748 22192 18760
rect 22066 18720 22192 18748
rect 16942 18680 16948 18692
rect 15580 18652 16948 18680
rect 15197 18643 15255 18649
rect 16942 18640 16948 18652
rect 17000 18640 17006 18692
rect 21453 18683 21511 18689
rect 21453 18680 21465 18683
rect 20640 18652 21465 18680
rect 2314 18572 2320 18624
rect 2372 18612 2378 18624
rect 3237 18615 3295 18621
rect 3237 18612 3249 18615
rect 2372 18584 3249 18612
rect 2372 18572 2378 18584
rect 3237 18581 3249 18584
rect 3283 18612 3295 18615
rect 4154 18612 4160 18624
rect 3283 18584 4160 18612
rect 3283 18581 3295 18584
rect 3237 18575 3295 18581
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 5353 18615 5411 18621
rect 5353 18581 5365 18615
rect 5399 18612 5411 18615
rect 5810 18612 5816 18624
rect 5399 18584 5816 18612
rect 5399 18581 5411 18584
rect 5353 18575 5411 18581
rect 5810 18572 5816 18584
rect 5868 18572 5874 18624
rect 9674 18612 9680 18624
rect 9635 18584 9680 18612
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 10318 18572 10324 18624
rect 10376 18612 10382 18624
rect 10502 18612 10508 18624
rect 10376 18584 10508 18612
rect 10376 18572 10382 18584
rect 10502 18572 10508 18584
rect 10560 18572 10566 18624
rect 10597 18615 10655 18621
rect 10597 18581 10609 18615
rect 10643 18612 10655 18615
rect 10686 18612 10692 18624
rect 10643 18584 10692 18612
rect 10643 18581 10655 18584
rect 10597 18575 10655 18581
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 11238 18572 11244 18624
rect 11296 18612 11302 18624
rect 11425 18615 11483 18621
rect 11425 18612 11437 18615
rect 11296 18584 11437 18612
rect 11296 18572 11302 18584
rect 11425 18581 11437 18584
rect 11471 18581 11483 18615
rect 12618 18612 12624 18624
rect 12579 18584 12624 18612
rect 11425 18575 11483 18581
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 12894 18572 12900 18624
rect 12952 18612 12958 18624
rect 15105 18615 15163 18621
rect 15105 18612 15117 18615
rect 12952 18584 15117 18612
rect 12952 18572 12958 18584
rect 15105 18581 15117 18584
rect 15151 18581 15163 18615
rect 15105 18575 15163 18581
rect 15470 18572 15476 18624
rect 15528 18612 15534 18624
rect 15565 18615 15623 18621
rect 15565 18612 15577 18615
rect 15528 18584 15577 18612
rect 15528 18572 15534 18584
rect 15565 18581 15577 18584
rect 15611 18581 15623 18615
rect 19702 18612 19708 18624
rect 19663 18584 19708 18612
rect 15565 18575 15623 18581
rect 19702 18572 19708 18584
rect 19760 18572 19766 18624
rect 20640 18621 20668 18652
rect 21453 18649 21465 18652
rect 21499 18680 21511 18683
rect 22066 18680 22094 18720
rect 22186 18708 22192 18720
rect 22244 18708 22250 18760
rect 21499 18652 22094 18680
rect 21499 18649 21511 18652
rect 21453 18643 21511 18649
rect 20625 18615 20683 18621
rect 20625 18581 20637 18615
rect 20671 18581 20683 18615
rect 20625 18575 20683 18581
rect 21545 18615 21603 18621
rect 21545 18581 21557 18615
rect 21591 18612 21603 18615
rect 21910 18612 21916 18624
rect 21591 18584 21916 18612
rect 21591 18581 21603 18584
rect 21545 18575 21603 18581
rect 21910 18572 21916 18584
rect 21968 18572 21974 18624
rect 1104 18522 30820 18544
rect 1104 18470 10880 18522
rect 10932 18470 10944 18522
rect 10996 18470 11008 18522
rect 11060 18470 11072 18522
rect 11124 18470 11136 18522
rect 11188 18470 20811 18522
rect 20863 18470 20875 18522
rect 20927 18470 20939 18522
rect 20991 18470 21003 18522
rect 21055 18470 21067 18522
rect 21119 18470 30820 18522
rect 1104 18448 30820 18470
rect 2498 18408 2504 18420
rect 2459 18380 2504 18408
rect 2498 18368 2504 18380
rect 2556 18368 2562 18420
rect 5718 18408 5724 18420
rect 4080 18380 5724 18408
rect 2148 18312 3924 18340
rect 1486 18232 1492 18284
rect 1544 18272 1550 18284
rect 1765 18275 1823 18281
rect 1765 18272 1777 18275
rect 1544 18244 1777 18272
rect 1544 18232 1550 18244
rect 1765 18241 1777 18244
rect 1811 18241 1823 18275
rect 1946 18272 1952 18284
rect 1907 18244 1952 18272
rect 1765 18235 1823 18241
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 2148 18281 2176 18312
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18241 2191 18275
rect 2314 18272 2320 18284
rect 2275 18244 2320 18272
rect 2133 18235 2191 18241
rect 2038 18204 2044 18216
rect 1999 18176 2044 18204
rect 2038 18164 2044 18176
rect 2096 18164 2102 18216
rect 1946 18096 1952 18148
rect 2004 18136 2010 18148
rect 2148 18136 2176 18235
rect 2314 18232 2320 18244
rect 2372 18232 2378 18284
rect 3510 18272 3516 18284
rect 3471 18244 3516 18272
rect 3510 18232 3516 18244
rect 3568 18232 3574 18284
rect 3694 18272 3700 18284
rect 3655 18244 3700 18272
rect 3694 18232 3700 18244
rect 3752 18232 3758 18284
rect 3896 18213 3924 18312
rect 4080 18281 4108 18380
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 9950 18368 9956 18420
rect 10008 18408 10014 18420
rect 10229 18411 10287 18417
rect 10229 18408 10241 18411
rect 10008 18380 10241 18408
rect 10008 18368 10014 18380
rect 10229 18377 10241 18380
rect 10275 18377 10287 18411
rect 12894 18408 12900 18420
rect 10229 18371 10287 18377
rect 12406 18380 12900 18408
rect 4338 18300 4344 18352
rect 4396 18340 4402 18352
rect 4709 18343 4767 18349
rect 4709 18340 4721 18343
rect 4396 18312 4721 18340
rect 4396 18300 4402 18312
rect 4709 18309 4721 18312
rect 4755 18309 4767 18343
rect 4709 18303 4767 18309
rect 5442 18300 5448 18352
rect 5500 18340 5506 18352
rect 5500 18312 6408 18340
rect 5500 18300 5506 18312
rect 4065 18275 4123 18281
rect 4065 18241 4077 18275
rect 4111 18241 4123 18275
rect 4890 18272 4896 18284
rect 4851 18244 4896 18272
rect 4065 18235 4123 18241
rect 4890 18232 4896 18244
rect 4948 18272 4954 18284
rect 6380 18281 6408 18312
rect 8662 18300 8668 18352
rect 8720 18340 8726 18352
rect 12406 18340 12434 18380
rect 12894 18368 12900 18380
rect 12952 18368 12958 18420
rect 15470 18408 15476 18420
rect 15431 18380 15476 18408
rect 15470 18368 15476 18380
rect 15528 18368 15534 18420
rect 18966 18408 18972 18420
rect 18927 18380 18972 18408
rect 18966 18368 18972 18380
rect 19024 18368 19030 18420
rect 19521 18411 19579 18417
rect 19521 18377 19533 18411
rect 19567 18408 19579 18411
rect 19610 18408 19616 18420
rect 19567 18380 19616 18408
rect 19567 18377 19579 18380
rect 19521 18371 19579 18377
rect 19610 18368 19616 18380
rect 19668 18368 19674 18420
rect 20438 18368 20444 18420
rect 20496 18408 20502 18420
rect 20901 18411 20959 18417
rect 20901 18408 20913 18411
rect 20496 18380 20913 18408
rect 20496 18368 20502 18380
rect 20901 18377 20913 18380
rect 20947 18377 20959 18411
rect 21910 18408 21916 18420
rect 21871 18380 21916 18408
rect 20901 18371 20959 18377
rect 21910 18368 21916 18380
rect 21968 18368 21974 18420
rect 13906 18340 13912 18352
rect 8720 18312 9076 18340
rect 8720 18300 8726 18312
rect 9048 18284 9076 18312
rect 10336 18312 12434 18340
rect 13867 18312 13912 18340
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 4948 18244 5641 18272
rect 4948 18232 4954 18244
rect 5629 18241 5641 18244
rect 5675 18241 5687 18275
rect 5629 18235 5687 18241
rect 6365 18275 6423 18281
rect 6365 18241 6377 18275
rect 6411 18241 6423 18275
rect 6365 18235 6423 18241
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 7009 18275 7067 18281
rect 7009 18272 7021 18275
rect 6512 18244 7021 18272
rect 6512 18232 6518 18244
rect 7009 18241 7021 18244
rect 7055 18241 7067 18275
rect 8938 18272 8944 18284
rect 8899 18244 8944 18272
rect 7009 18235 7067 18241
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 9030 18232 9036 18284
rect 9088 18272 9094 18284
rect 9125 18275 9183 18281
rect 9125 18272 9137 18275
rect 9088 18244 9137 18272
rect 9088 18232 9094 18244
rect 9125 18241 9137 18244
rect 9171 18241 9183 18275
rect 9125 18235 9183 18241
rect 9217 18275 9275 18281
rect 9217 18241 9229 18275
rect 9263 18272 9275 18275
rect 9398 18272 9404 18284
rect 9263 18244 9404 18272
rect 9263 18241 9275 18244
rect 9217 18235 9275 18241
rect 9398 18232 9404 18244
rect 9456 18232 9462 18284
rect 10336 18281 10364 18312
rect 13906 18300 13912 18312
rect 13964 18340 13970 18352
rect 14550 18340 14556 18352
rect 13964 18312 14556 18340
rect 13964 18300 13970 18312
rect 14550 18300 14556 18312
rect 14608 18300 14614 18352
rect 15378 18340 15384 18352
rect 15339 18312 15384 18340
rect 15378 18300 15384 18312
rect 15436 18300 15442 18352
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18272 9551 18275
rect 10321 18275 10379 18281
rect 10321 18272 10333 18275
rect 9539 18244 10333 18272
rect 9539 18241 9551 18244
rect 9493 18235 9551 18241
rect 10321 18241 10333 18244
rect 10367 18241 10379 18275
rect 11773 18275 11831 18281
rect 11773 18272 11785 18275
rect 10321 18235 10379 18241
rect 10704 18244 11785 18272
rect 3789 18207 3847 18213
rect 3789 18204 3801 18207
rect 2004 18108 2176 18136
rect 3712 18176 3801 18204
rect 3712 18136 3740 18176
rect 3789 18173 3801 18176
rect 3835 18173 3847 18207
rect 3789 18167 3847 18173
rect 3881 18207 3939 18213
rect 3881 18173 3893 18207
rect 3927 18204 3939 18207
rect 5445 18207 5503 18213
rect 5445 18204 5457 18207
rect 3927 18176 5457 18204
rect 3927 18173 3939 18176
rect 3881 18167 3939 18173
rect 5445 18173 5457 18176
rect 5491 18173 5503 18207
rect 9306 18204 9312 18216
rect 9219 18176 9312 18204
rect 5445 18167 5503 18173
rect 9306 18164 9312 18176
rect 9364 18204 9370 18216
rect 9677 18207 9735 18213
rect 9364 18176 9536 18204
rect 9364 18164 9370 18176
rect 9508 18148 9536 18176
rect 9677 18173 9689 18207
rect 9723 18204 9735 18207
rect 10704 18204 10732 18244
rect 11773 18241 11785 18244
rect 11819 18241 11831 18275
rect 11773 18235 11831 18241
rect 13633 18275 13691 18281
rect 13633 18241 13645 18275
rect 13679 18272 13691 18275
rect 14274 18272 14280 18284
rect 13679 18244 14280 18272
rect 13679 18241 13691 18244
rect 13633 18235 13691 18241
rect 14274 18232 14280 18244
rect 14332 18272 14338 18284
rect 14826 18272 14832 18284
rect 14332 18244 14832 18272
rect 14332 18232 14338 18244
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 17218 18272 17224 18284
rect 17179 18244 17224 18272
rect 17218 18232 17224 18244
rect 17276 18232 17282 18284
rect 18230 18232 18236 18284
rect 18288 18272 18294 18284
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 18288 18244 18337 18272
rect 18288 18232 18294 18244
rect 18325 18241 18337 18244
rect 18371 18241 18383 18275
rect 18325 18235 18383 18241
rect 19061 18275 19119 18281
rect 19061 18241 19073 18275
rect 19107 18272 19119 18275
rect 19334 18272 19340 18284
rect 19107 18244 19340 18272
rect 19107 18241 19119 18244
rect 19061 18235 19119 18241
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 19702 18272 19708 18284
rect 19664 18244 19708 18272
rect 19702 18232 19708 18244
rect 19760 18232 19766 18284
rect 19797 18275 19855 18281
rect 19797 18241 19809 18275
rect 19843 18241 19855 18275
rect 19797 18235 19855 18241
rect 20073 18275 20131 18281
rect 20073 18241 20085 18275
rect 20119 18272 20131 18275
rect 20162 18272 20168 18284
rect 20119 18244 20168 18272
rect 20119 18241 20131 18244
rect 20073 18235 20131 18241
rect 11514 18204 11520 18216
rect 9723 18176 10732 18204
rect 11475 18176 11520 18204
rect 9723 18173 9735 18176
rect 9677 18167 9735 18173
rect 11514 18164 11520 18176
rect 11572 18164 11578 18216
rect 15562 18204 15568 18216
rect 15523 18176 15568 18204
rect 15562 18164 15568 18176
rect 15620 18164 15626 18216
rect 17494 18204 17500 18216
rect 17455 18176 17500 18204
rect 17494 18164 17500 18176
rect 17552 18164 17558 18216
rect 18046 18204 18052 18216
rect 18007 18176 18052 18204
rect 18046 18164 18052 18176
rect 18104 18164 18110 18216
rect 19352 18204 19380 18232
rect 19812 18204 19840 18235
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 20530 18272 20536 18284
rect 20491 18244 20536 18272
rect 20530 18232 20536 18244
rect 20588 18232 20594 18284
rect 20714 18272 20720 18284
rect 20627 18244 20720 18272
rect 20714 18232 20720 18244
rect 20772 18272 20778 18284
rect 21174 18272 21180 18284
rect 20772 18244 21180 18272
rect 20772 18232 20778 18244
rect 21174 18232 21180 18244
rect 21232 18232 21238 18284
rect 22002 18272 22008 18284
rect 21963 18244 22008 18272
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 29822 18272 29828 18284
rect 29783 18244 29828 18272
rect 29822 18232 29828 18244
rect 29880 18232 29886 18284
rect 19352 18176 19840 18204
rect 4430 18136 4436 18148
rect 3712 18108 4436 18136
rect 2004 18096 2010 18108
rect 4430 18096 4436 18108
rect 4488 18096 4494 18148
rect 4540 18108 7236 18136
rect 4246 18068 4252 18080
rect 4207 18040 4252 18068
rect 4246 18028 4252 18040
rect 4304 18028 4310 18080
rect 4338 18028 4344 18080
rect 4396 18068 4402 18080
rect 4540 18068 4568 18108
rect 6454 18068 6460 18080
rect 4396 18040 4568 18068
rect 6415 18040 6460 18068
rect 4396 18028 4402 18040
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 6730 18028 6736 18080
rect 6788 18068 6794 18080
rect 7101 18071 7159 18077
rect 7101 18068 7113 18071
rect 6788 18040 7113 18068
rect 6788 18028 6794 18040
rect 7101 18037 7113 18040
rect 7147 18037 7159 18071
rect 7208 18068 7236 18108
rect 9490 18096 9496 18148
rect 9548 18096 9554 18148
rect 13446 18096 13452 18148
rect 13504 18136 13510 18148
rect 13722 18136 13728 18148
rect 13504 18108 13728 18136
rect 13504 18096 13510 18108
rect 13722 18096 13728 18108
rect 13780 18096 13786 18148
rect 10502 18068 10508 18080
rect 7208 18040 10508 18068
rect 7101 18031 7159 18037
rect 10502 18028 10508 18040
rect 10560 18068 10566 18080
rect 10686 18068 10692 18080
rect 10560 18040 10692 18068
rect 10560 18028 10566 18040
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 13814 18068 13820 18080
rect 13775 18040 13820 18068
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 15010 18068 15016 18080
rect 14971 18040 15016 18068
rect 15010 18028 15016 18040
rect 15068 18028 15074 18080
rect 19978 18068 19984 18080
rect 19939 18040 19984 18068
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 30006 18068 30012 18080
rect 29967 18040 30012 18068
rect 30006 18028 30012 18040
rect 30064 18028 30070 18080
rect 1104 17978 30820 18000
rect 1104 17926 5915 17978
rect 5967 17926 5979 17978
rect 6031 17926 6043 17978
rect 6095 17926 6107 17978
rect 6159 17926 6171 17978
rect 6223 17926 15846 17978
rect 15898 17926 15910 17978
rect 15962 17926 15974 17978
rect 16026 17926 16038 17978
rect 16090 17926 16102 17978
rect 16154 17926 25776 17978
rect 25828 17926 25840 17978
rect 25892 17926 25904 17978
rect 25956 17926 25968 17978
rect 26020 17926 26032 17978
rect 26084 17926 30820 17978
rect 1104 17904 30820 17926
rect 2961 17867 3019 17873
rect 2961 17833 2973 17867
rect 3007 17864 3019 17867
rect 3694 17864 3700 17876
rect 3007 17836 3700 17864
rect 3007 17833 3019 17836
rect 2961 17827 3019 17833
rect 3694 17824 3700 17836
rect 3752 17824 3758 17876
rect 11149 17867 11207 17873
rect 11149 17833 11161 17867
rect 11195 17864 11207 17867
rect 11422 17864 11428 17876
rect 11195 17836 11428 17864
rect 11195 17833 11207 17836
rect 11149 17827 11207 17833
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 12986 17864 12992 17876
rect 12947 17836 12992 17864
rect 12986 17824 12992 17836
rect 13044 17824 13050 17876
rect 13998 17824 14004 17876
rect 14056 17864 14062 17876
rect 14737 17867 14795 17873
rect 14737 17864 14749 17867
rect 14056 17836 14749 17864
rect 14056 17824 14062 17836
rect 14737 17833 14749 17836
rect 14783 17833 14795 17867
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 14737 17827 14795 17833
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15381 17867 15439 17873
rect 15381 17833 15393 17867
rect 15427 17864 15439 17867
rect 15746 17864 15752 17876
rect 15427 17836 15752 17864
rect 15427 17833 15439 17836
rect 15381 17827 15439 17833
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 16669 17867 16727 17873
rect 16669 17833 16681 17867
rect 16715 17864 16727 17867
rect 16942 17864 16948 17876
rect 16715 17836 16948 17864
rect 16715 17833 16727 17836
rect 16669 17827 16727 17833
rect 16942 17824 16948 17836
rect 17000 17824 17006 17876
rect 17129 17867 17187 17873
rect 17129 17833 17141 17867
rect 17175 17864 17187 17867
rect 17494 17864 17500 17876
rect 17175 17836 17500 17864
rect 17175 17833 17187 17836
rect 17129 17827 17187 17833
rect 17494 17824 17500 17836
rect 17552 17824 17558 17876
rect 19334 17864 19340 17876
rect 19295 17836 19340 17864
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 20257 17867 20315 17873
rect 20257 17833 20269 17867
rect 20303 17864 20315 17867
rect 20714 17864 20720 17876
rect 20303 17836 20720 17864
rect 20303 17833 20315 17836
rect 20257 17827 20315 17833
rect 20714 17824 20720 17836
rect 20772 17824 20778 17876
rect 29822 17824 29828 17876
rect 29880 17864 29886 17876
rect 29917 17867 29975 17873
rect 29917 17864 29929 17867
rect 29880 17836 29929 17864
rect 29880 17824 29886 17836
rect 29917 17833 29929 17836
rect 29963 17833 29975 17867
rect 29917 17827 29975 17833
rect 6270 17756 6276 17808
rect 6328 17756 6334 17808
rect 8938 17796 8944 17808
rect 7668 17768 8944 17796
rect 2038 17728 2044 17740
rect 1999 17700 2044 17728
rect 2038 17688 2044 17700
rect 2096 17688 2102 17740
rect 2866 17728 2872 17740
rect 2148 17700 2872 17728
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17629 1823 17663
rect 1946 17660 1952 17672
rect 1907 17632 1952 17660
rect 1765 17623 1823 17629
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17524 1639 17527
rect 1670 17524 1676 17536
rect 1627 17496 1676 17524
rect 1627 17493 1639 17496
rect 1581 17487 1639 17493
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 1780 17524 1808 17623
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 2148 17669 2176 17700
rect 2866 17688 2872 17700
rect 2924 17688 2930 17740
rect 3786 17728 3792 17740
rect 3699 17700 3792 17728
rect 3786 17688 3792 17700
rect 3844 17728 3850 17740
rect 4338 17728 4344 17740
rect 3844 17700 4344 17728
rect 3844 17688 3850 17700
rect 4338 17688 4344 17700
rect 4396 17688 4402 17740
rect 6288 17728 6316 17756
rect 6641 17731 6699 17737
rect 6641 17728 6653 17731
rect 6288 17700 6653 17728
rect 6641 17697 6653 17700
rect 6687 17697 6699 17731
rect 6641 17691 6699 17697
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17629 2191 17663
rect 2133 17623 2191 17629
rect 2317 17663 2375 17669
rect 2317 17629 2329 17663
rect 2363 17629 2375 17663
rect 2317 17623 2375 17629
rect 2332 17592 2360 17623
rect 2774 17620 2780 17672
rect 2832 17660 2838 17672
rect 4065 17663 4123 17669
rect 2832 17632 2877 17660
rect 2832 17620 2838 17632
rect 4065 17629 4077 17663
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 2866 17592 2872 17604
rect 2332 17564 2872 17592
rect 2866 17552 2872 17564
rect 2924 17592 2930 17604
rect 3510 17592 3516 17604
rect 2924 17564 3516 17592
rect 2924 17552 2930 17564
rect 3510 17552 3516 17564
rect 3568 17592 3574 17604
rect 4080 17592 4108 17623
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 5353 17663 5411 17669
rect 5353 17660 5365 17663
rect 4212 17632 5365 17660
rect 4212 17620 4218 17632
rect 5353 17629 5365 17632
rect 5399 17629 5411 17663
rect 5353 17623 5411 17629
rect 6270 17620 6276 17672
rect 6328 17660 6334 17672
rect 6365 17663 6423 17669
rect 6365 17660 6377 17663
rect 6328 17632 6377 17660
rect 6328 17620 6334 17632
rect 6365 17629 6377 17632
rect 6411 17629 6423 17663
rect 6656 17660 6684 17691
rect 7668 17669 7696 17768
rect 8938 17756 8944 17768
rect 8996 17756 9002 17808
rect 13446 17756 13452 17808
rect 13504 17796 13510 17808
rect 14461 17799 14519 17805
rect 14461 17796 14473 17799
rect 13504 17768 14473 17796
rect 13504 17756 13510 17768
rect 14461 17765 14473 17768
rect 14507 17765 14519 17799
rect 14461 17759 14519 17765
rect 15194 17756 15200 17808
rect 15252 17756 15258 17808
rect 17218 17796 17224 17808
rect 15488 17768 17224 17796
rect 7929 17731 7987 17737
rect 7929 17697 7941 17731
rect 7975 17728 7987 17731
rect 8110 17728 8116 17740
rect 7975 17700 8116 17728
rect 7975 17697 7987 17700
rect 7929 17691 7987 17697
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 9769 17731 9827 17737
rect 9769 17728 9781 17731
rect 8352 17700 9781 17728
rect 8352 17688 8358 17700
rect 9769 17697 9781 17700
rect 9815 17697 9827 17731
rect 9769 17691 9827 17697
rect 13814 17688 13820 17740
rect 13872 17728 13878 17740
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 13872 17700 14289 17728
rect 13872 17688 13878 17700
rect 14277 17697 14289 17700
rect 14323 17697 14335 17731
rect 14277 17691 14335 17697
rect 14369 17731 14427 17737
rect 14369 17697 14381 17731
rect 14415 17728 14427 17731
rect 15212 17728 15240 17756
rect 15488 17737 15516 17768
rect 17218 17756 17224 17768
rect 17276 17796 17282 17808
rect 18325 17799 18383 17805
rect 17276 17768 17356 17796
rect 17276 17756 17282 17768
rect 14415 17700 15240 17728
rect 15473 17731 15531 17737
rect 14415 17697 14427 17700
rect 14369 17691 14427 17697
rect 15473 17697 15485 17731
rect 15519 17697 15531 17731
rect 15473 17691 15531 17697
rect 16117 17731 16175 17737
rect 16117 17697 16129 17731
rect 16163 17728 16175 17731
rect 16666 17728 16672 17740
rect 16163 17700 16672 17728
rect 16163 17697 16175 17700
rect 16117 17691 16175 17697
rect 16666 17688 16672 17700
rect 16724 17688 16730 17740
rect 17328 17737 17356 17768
rect 18325 17765 18337 17799
rect 18371 17796 18383 17799
rect 19242 17796 19248 17808
rect 18371 17768 19248 17796
rect 18371 17765 18383 17768
rect 18325 17759 18383 17765
rect 19242 17756 19248 17768
rect 19300 17756 19306 17808
rect 19978 17796 19984 17808
rect 19536 17768 19984 17796
rect 17313 17731 17371 17737
rect 17313 17697 17325 17731
rect 17359 17697 17371 17731
rect 17313 17691 17371 17697
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17728 17831 17731
rect 18046 17728 18052 17740
rect 17819 17700 18052 17728
rect 17819 17697 17831 17700
rect 17773 17691 17831 17697
rect 18046 17688 18052 17700
rect 18104 17688 18110 17740
rect 19536 17672 19564 17768
rect 19978 17756 19984 17768
rect 20036 17796 20042 17808
rect 20165 17799 20223 17805
rect 20165 17796 20177 17799
rect 20036 17768 20177 17796
rect 20036 17756 20042 17768
rect 20165 17765 20177 17768
rect 20211 17765 20223 17799
rect 20165 17759 20223 17765
rect 19610 17688 19616 17740
rect 19668 17728 19674 17740
rect 20349 17731 20407 17737
rect 20349 17728 20361 17731
rect 19668 17700 20361 17728
rect 19668 17688 19674 17700
rect 20349 17697 20361 17700
rect 20395 17697 20407 17731
rect 20349 17691 20407 17697
rect 7653 17663 7711 17669
rect 7653 17660 7665 17663
rect 6656 17632 7665 17660
rect 6365 17623 6423 17629
rect 7653 17629 7665 17632
rect 7699 17629 7711 17663
rect 7653 17623 7711 17629
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17629 7895 17663
rect 7837 17623 7895 17629
rect 8021 17663 8079 17669
rect 8021 17629 8033 17663
rect 8067 17629 8079 17663
rect 8021 17623 8079 17629
rect 8205 17663 8263 17669
rect 8205 17629 8217 17663
rect 8251 17660 8263 17663
rect 9214 17660 9220 17672
rect 8251 17632 9220 17660
rect 8251 17629 8263 17632
rect 8205 17623 8263 17629
rect 3568 17564 4108 17592
rect 3568 17552 3574 17564
rect 2406 17524 2412 17536
rect 1780 17496 2412 17524
rect 2406 17484 2412 17496
rect 2464 17484 2470 17536
rect 5445 17527 5503 17533
rect 5445 17493 5457 17527
rect 5491 17524 5503 17527
rect 5626 17524 5632 17536
rect 5491 17496 5632 17524
rect 5491 17493 5503 17496
rect 5445 17487 5503 17493
rect 5626 17484 5632 17496
rect 5684 17484 5690 17536
rect 7852 17524 7880 17623
rect 8036 17592 8064 17623
rect 9214 17620 9220 17632
rect 9272 17620 9278 17672
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 10025 17663 10083 17669
rect 10025 17660 10037 17663
rect 9732 17632 10037 17660
rect 9732 17620 9738 17632
rect 10025 17629 10037 17632
rect 10071 17629 10083 17663
rect 10025 17623 10083 17629
rect 11514 17620 11520 17672
rect 11572 17660 11578 17672
rect 11609 17663 11667 17669
rect 11609 17660 11621 17663
rect 11572 17632 11621 17660
rect 11572 17620 11578 17632
rect 11609 17629 11621 17632
rect 11655 17660 11667 17663
rect 11655 17632 12020 17660
rect 11655 17629 11667 17632
rect 11609 17623 11667 17629
rect 11992 17604 12020 17632
rect 13906 17620 13912 17672
rect 13964 17660 13970 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13964 17632 14105 17660
rect 13964 17620 13970 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14550 17660 14556 17672
rect 14511 17632 14556 17660
rect 14093 17623 14151 17629
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 15197 17663 15255 17669
rect 15197 17629 15209 17663
rect 15243 17660 15255 17663
rect 16206 17660 16212 17672
rect 15243 17632 16212 17660
rect 15243 17629 15255 17632
rect 15197 17623 15255 17629
rect 16206 17620 16212 17632
rect 16264 17620 16270 17672
rect 16301 17663 16359 17669
rect 16301 17629 16313 17663
rect 16347 17660 16359 17663
rect 16850 17660 16856 17672
rect 16347 17632 16856 17660
rect 16347 17629 16359 17632
rect 16301 17623 16359 17629
rect 16850 17620 16856 17632
rect 16908 17620 16914 17672
rect 17405 17663 17463 17669
rect 17405 17629 17417 17663
rect 17451 17660 17463 17663
rect 17678 17660 17684 17672
rect 17451 17632 17684 17660
rect 17451 17629 17463 17632
rect 17405 17623 17463 17629
rect 17678 17620 17684 17632
rect 17736 17620 17742 17672
rect 18230 17660 18236 17672
rect 18191 17632 18236 17660
rect 18230 17620 18236 17632
rect 18288 17620 18294 17672
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17660 19487 17663
rect 19518 17660 19524 17672
rect 19475 17632 19524 17660
rect 19475 17629 19487 17632
rect 19429 17623 19487 17629
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17660 20131 17663
rect 20162 17660 20168 17672
rect 20119 17632 20168 17660
rect 20119 17629 20131 17632
rect 20073 17623 20131 17629
rect 20162 17620 20168 17632
rect 20220 17660 20226 17672
rect 20993 17663 21051 17669
rect 20993 17660 21005 17663
rect 20220 17632 21005 17660
rect 20220 17620 20226 17632
rect 20993 17629 21005 17632
rect 21039 17629 21051 17663
rect 30098 17660 30104 17672
rect 30059 17632 30104 17660
rect 20993 17623 21051 17629
rect 30098 17620 30104 17632
rect 30156 17620 30162 17672
rect 9490 17592 9496 17604
rect 8036 17564 9496 17592
rect 9490 17552 9496 17564
rect 9548 17552 9554 17604
rect 9858 17552 9864 17604
rect 9916 17592 9922 17604
rect 11854 17595 11912 17601
rect 11854 17592 11866 17595
rect 9916 17564 11866 17592
rect 9916 17552 9922 17564
rect 11854 17561 11866 17564
rect 11900 17561 11912 17595
rect 11854 17555 11912 17561
rect 11974 17552 11980 17604
rect 12032 17552 12038 17604
rect 19702 17552 19708 17604
rect 19760 17592 19766 17604
rect 20901 17595 20959 17601
rect 20901 17592 20913 17595
rect 19760 17564 20913 17592
rect 19760 17552 19766 17564
rect 20901 17561 20913 17564
rect 20947 17561 20959 17595
rect 20901 17555 20959 17561
rect 8202 17524 8208 17536
rect 7852 17496 8208 17524
rect 8202 17484 8208 17496
rect 8260 17484 8266 17536
rect 8386 17524 8392 17536
rect 8347 17496 8392 17524
rect 8386 17484 8392 17496
rect 8444 17484 8450 17536
rect 13630 17484 13636 17536
rect 13688 17524 13694 17536
rect 16022 17524 16028 17536
rect 13688 17496 16028 17524
rect 13688 17484 13694 17496
rect 16022 17484 16028 17496
rect 16080 17484 16086 17536
rect 1104 17434 30820 17456
rect 1104 17382 10880 17434
rect 10932 17382 10944 17434
rect 10996 17382 11008 17434
rect 11060 17382 11072 17434
rect 11124 17382 11136 17434
rect 11188 17382 20811 17434
rect 20863 17382 20875 17434
rect 20927 17382 20939 17434
rect 20991 17382 21003 17434
rect 21055 17382 21067 17434
rect 21119 17382 30820 17434
rect 1104 17360 30820 17382
rect 8665 17323 8723 17329
rect 8665 17289 8677 17323
rect 8711 17320 8723 17323
rect 9214 17320 9220 17332
rect 8711 17292 9220 17320
rect 8711 17289 8723 17292
rect 8665 17283 8723 17289
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 9858 17320 9864 17332
rect 9819 17292 9864 17320
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 15194 17280 15200 17332
rect 15252 17320 15258 17332
rect 15841 17323 15899 17329
rect 15841 17320 15853 17323
rect 15252 17292 15853 17320
rect 15252 17280 15258 17292
rect 15841 17289 15853 17292
rect 15887 17320 15899 17323
rect 16298 17320 16304 17332
rect 15887 17292 16304 17320
rect 15887 17289 15899 17292
rect 15841 17283 15899 17289
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 16761 17323 16819 17329
rect 16761 17289 16773 17323
rect 16807 17320 16819 17323
rect 16850 17320 16856 17332
rect 16807 17292 16856 17320
rect 16807 17289 16819 17292
rect 16761 17283 16819 17289
rect 16850 17280 16856 17292
rect 16908 17280 16914 17332
rect 17681 17323 17739 17329
rect 17681 17289 17693 17323
rect 17727 17320 17739 17323
rect 18046 17320 18052 17332
rect 17727 17292 18052 17320
rect 17727 17289 17739 17292
rect 17681 17283 17739 17289
rect 18046 17280 18052 17292
rect 18104 17280 18110 17332
rect 21266 17320 21272 17332
rect 19444 17292 21272 17320
rect 2314 17212 2320 17264
rect 2372 17252 2378 17264
rect 6825 17255 6883 17261
rect 2372 17224 4108 17252
rect 2372 17212 2378 17224
rect 4080 17196 4108 17224
rect 6825 17221 6837 17255
rect 6871 17252 6883 17255
rect 7190 17252 7196 17264
rect 6871 17224 7196 17252
rect 6871 17221 6883 17224
rect 6825 17215 6883 17221
rect 7190 17212 7196 17224
rect 7248 17212 7254 17264
rect 7552 17255 7610 17261
rect 7552 17221 7564 17255
rect 7598 17252 7610 17255
rect 8386 17252 8392 17264
rect 7598 17224 8392 17252
rect 7598 17221 7610 17224
rect 7552 17215 7610 17221
rect 8386 17212 8392 17224
rect 8444 17212 8450 17264
rect 12244 17255 12302 17261
rect 12244 17221 12256 17255
rect 12290 17252 12302 17255
rect 12618 17252 12624 17264
rect 12290 17224 12624 17252
rect 12290 17221 12302 17224
rect 12244 17215 12302 17221
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 14568 17224 15700 17252
rect 1670 17193 1676 17196
rect 1664 17184 1676 17193
rect 1631 17156 1676 17184
rect 1664 17147 1676 17156
rect 1670 17144 1676 17147
rect 1728 17144 1734 17196
rect 3234 17184 3240 17196
rect 3195 17156 3240 17184
rect 3234 17144 3240 17156
rect 3292 17144 3298 17196
rect 4062 17184 4068 17196
rect 3975 17156 4068 17184
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 4338 17193 4344 17196
rect 4332 17147 4344 17193
rect 4396 17184 4402 17196
rect 4396 17156 4432 17184
rect 4338 17144 4344 17147
rect 4396 17144 4402 17156
rect 6270 17144 6276 17196
rect 6328 17184 6334 17196
rect 6641 17187 6699 17193
rect 6641 17184 6653 17187
rect 6328 17156 6653 17184
rect 6328 17144 6334 17156
rect 6641 17153 6653 17156
rect 6687 17153 6699 17187
rect 7208 17184 7236 17212
rect 7926 17184 7932 17196
rect 7208 17156 7932 17184
rect 6641 17147 6699 17153
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9125 17187 9183 17193
rect 9125 17184 9137 17187
rect 8996 17156 9137 17184
rect 8996 17144 9002 17156
rect 9125 17153 9137 17156
rect 9171 17153 9183 17187
rect 9125 17147 9183 17153
rect 9214 17144 9220 17196
rect 9272 17184 9278 17196
rect 9309 17187 9367 17193
rect 9309 17184 9321 17187
rect 9272 17156 9321 17184
rect 9272 17144 9278 17156
rect 9309 17153 9321 17156
rect 9355 17153 9367 17187
rect 9309 17147 9367 17153
rect 9677 17187 9735 17193
rect 9677 17153 9689 17187
rect 9723 17184 9735 17187
rect 9766 17184 9772 17196
rect 9723 17156 9772 17184
rect 9723 17153 9735 17156
rect 9677 17147 9735 17153
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 13814 17184 13820 17196
rect 13775 17156 13820 17184
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 14568 17193 14596 17224
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17153 14611 17187
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 14553 17147 14611 17153
rect 14660 17156 14749 17184
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17085 1455 17119
rect 1397 17079 1455 17085
rect 1412 16980 1440 17079
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7285 17119 7343 17125
rect 7285 17116 7297 17119
rect 7248 17088 7297 17116
rect 7248 17076 7254 17088
rect 7285 17085 7297 17088
rect 7331 17085 7343 17119
rect 9398 17116 9404 17128
rect 9359 17088 9404 17116
rect 7285 17079 7343 17085
rect 9398 17076 9404 17088
rect 9456 17076 9462 17128
rect 9490 17076 9496 17128
rect 9548 17116 9554 17128
rect 11974 17116 11980 17128
rect 9548 17088 9593 17116
rect 11935 17088 11980 17116
rect 9548 17076 9554 17088
rect 11974 17076 11980 17088
rect 12032 17076 12038 17128
rect 2406 17008 2412 17060
rect 2464 17048 2470 17060
rect 2777 17051 2835 17057
rect 2777 17048 2789 17051
rect 2464 17020 2789 17048
rect 2464 17008 2470 17020
rect 2777 17017 2789 17020
rect 2823 17048 2835 17051
rect 2823 17020 4099 17048
rect 2823 17017 2835 17020
rect 2777 17011 2835 17017
rect 2314 16980 2320 16992
rect 1412 16952 2320 16980
rect 2314 16940 2320 16952
rect 2372 16940 2378 16992
rect 3421 16983 3479 16989
rect 3421 16949 3433 16983
rect 3467 16980 3479 16983
rect 3970 16980 3976 16992
rect 3467 16952 3976 16980
rect 3467 16949 3479 16952
rect 3421 16943 3479 16949
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 4071 16980 4099 17020
rect 4706 16980 4712 16992
rect 4071 16952 4712 16980
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 4798 16940 4804 16992
rect 4856 16980 4862 16992
rect 5442 16980 5448 16992
rect 4856 16952 5448 16980
rect 4856 16940 4862 16952
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 6638 16940 6644 16992
rect 6696 16980 6702 16992
rect 8386 16980 8392 16992
rect 6696 16952 8392 16980
rect 6696 16940 6702 16952
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 10042 16940 10048 16992
rect 10100 16980 10106 16992
rect 10318 16980 10324 16992
rect 10100 16952 10324 16980
rect 10100 16940 10106 16952
rect 10318 16940 10324 16952
rect 10376 16940 10382 16992
rect 13357 16983 13415 16989
rect 13357 16949 13369 16983
rect 13403 16980 13415 16983
rect 13814 16980 13820 16992
rect 13403 16952 13820 16980
rect 13403 16949 13415 16952
rect 13357 16943 13415 16949
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 13906 16940 13912 16992
rect 13964 16980 13970 16992
rect 14660 16980 14688 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 15102 17184 15108 17196
rect 15063 17156 15108 17184
rect 14737 17147 14795 17153
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 14829 17119 14887 17125
rect 14829 17116 14841 17119
rect 14752 17088 14841 17116
rect 14752 17060 14780 17088
rect 14829 17085 14841 17088
rect 14875 17085 14887 17119
rect 14829 17079 14887 17085
rect 14918 17076 14924 17128
rect 14976 17116 14982 17128
rect 15672 17116 15700 17224
rect 15746 17212 15752 17264
rect 15804 17252 15810 17264
rect 15804 17224 16712 17252
rect 15804 17212 15810 17224
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17184 15991 17187
rect 16022 17184 16028 17196
rect 15979 17156 16028 17184
rect 15979 17153 15991 17156
rect 15933 17147 15991 17153
rect 16022 17144 16028 17156
rect 16080 17144 16086 17196
rect 16684 17193 16712 17224
rect 17218 17212 17224 17264
rect 17276 17252 17282 17264
rect 17313 17255 17371 17261
rect 17313 17252 17325 17255
rect 17276 17224 17325 17252
rect 17276 17212 17282 17224
rect 17313 17221 17325 17224
rect 17359 17252 17371 17255
rect 17586 17252 17592 17264
rect 17359 17224 17592 17252
rect 17359 17221 17371 17224
rect 17313 17215 17371 17221
rect 17586 17212 17592 17224
rect 17644 17212 17650 17264
rect 16669 17187 16727 17193
rect 16669 17153 16681 17187
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 17497 17187 17555 17193
rect 17497 17153 17509 17187
rect 17543 17184 17555 17187
rect 17678 17184 17684 17196
rect 17543 17156 17684 17184
rect 17543 17153 17555 17156
rect 17497 17147 17555 17153
rect 17678 17144 17684 17156
rect 17736 17144 17742 17196
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17184 19119 17187
rect 19242 17184 19248 17196
rect 19107 17156 19248 17184
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 19242 17144 19248 17156
rect 19300 17184 19306 17196
rect 19444 17184 19472 17292
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 19794 17252 19800 17264
rect 19536 17224 19800 17252
rect 19536 17193 19564 17224
rect 19794 17212 19800 17224
rect 19852 17212 19858 17264
rect 19300 17156 19472 17184
rect 19521 17187 19579 17193
rect 19300 17144 19306 17156
rect 19521 17153 19533 17187
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 19610 17144 19616 17196
rect 19668 17184 19674 17196
rect 19705 17187 19763 17193
rect 19705 17184 19717 17187
rect 19668 17156 19717 17184
rect 19668 17144 19674 17156
rect 19705 17153 19717 17156
rect 19751 17153 19763 17187
rect 19705 17147 19763 17153
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17184 20131 17187
rect 20254 17184 20260 17196
rect 20119 17156 20260 17184
rect 20119 17153 20131 17156
rect 20073 17147 20131 17153
rect 20254 17144 20260 17156
rect 20312 17144 20318 17196
rect 17862 17116 17868 17128
rect 14976 17088 15021 17116
rect 15672 17088 17868 17116
rect 14976 17076 14982 17088
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 19797 17119 19855 17125
rect 19797 17116 19809 17119
rect 19720 17088 19809 17116
rect 19720 17060 19748 17088
rect 19797 17085 19809 17088
rect 19843 17085 19855 17119
rect 19797 17079 19855 17085
rect 19886 17076 19892 17128
rect 19944 17116 19950 17128
rect 19944 17088 19989 17116
rect 19944 17076 19950 17088
rect 14734 17008 14740 17060
rect 14792 17008 14798 17060
rect 16758 17048 16764 17060
rect 14936 17020 16764 17048
rect 14936 16980 14964 17020
rect 16758 17008 16764 17020
rect 16816 17008 16822 17060
rect 19702 17008 19708 17060
rect 19760 17008 19766 17060
rect 13964 16952 14009 16980
rect 14660 16952 14964 16980
rect 13964 16940 13970 16952
rect 15102 16940 15108 16992
rect 15160 16980 15166 16992
rect 15289 16983 15347 16989
rect 15289 16980 15301 16983
rect 15160 16952 15301 16980
rect 15160 16940 15166 16952
rect 15289 16949 15301 16952
rect 15335 16949 15347 16983
rect 18966 16980 18972 16992
rect 18927 16952 18972 16980
rect 15289 16943 15347 16949
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 19978 16980 19984 16992
rect 19392 16952 19984 16980
rect 19392 16940 19398 16952
rect 19978 16940 19984 16952
rect 20036 16940 20042 16992
rect 20257 16983 20315 16989
rect 20257 16949 20269 16983
rect 20303 16980 20315 16983
rect 20714 16980 20720 16992
rect 20303 16952 20720 16980
rect 20303 16949 20315 16952
rect 20257 16943 20315 16949
rect 20714 16940 20720 16952
rect 20772 16940 20778 16992
rect 1104 16890 30820 16912
rect 1104 16838 5915 16890
rect 5967 16838 5979 16890
rect 6031 16838 6043 16890
rect 6095 16838 6107 16890
rect 6159 16838 6171 16890
rect 6223 16838 15846 16890
rect 15898 16838 15910 16890
rect 15962 16838 15974 16890
rect 16026 16838 16038 16890
rect 16090 16838 16102 16890
rect 16154 16838 25776 16890
rect 25828 16838 25840 16890
rect 25892 16838 25904 16890
rect 25956 16838 25968 16890
rect 26020 16838 26032 16890
rect 26084 16838 30820 16890
rect 1104 16816 30820 16838
rect 6270 16776 6276 16788
rect 6231 16748 6276 16776
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 7190 16776 7196 16788
rect 6840 16748 7196 16776
rect 4154 16708 4160 16720
rect 2746 16680 4160 16708
rect 2133 16643 2191 16649
rect 2133 16609 2145 16643
rect 2179 16640 2191 16643
rect 2746 16640 2774 16680
rect 4154 16668 4160 16680
rect 4212 16668 4218 16720
rect 2179 16612 2774 16640
rect 2179 16609 2191 16612
rect 2133 16603 2191 16609
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 6840 16649 6868 16748
rect 7190 16736 7196 16748
rect 7248 16776 7254 16788
rect 10042 16776 10048 16788
rect 7248 16748 10048 16776
rect 7248 16736 7254 16748
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 18230 16736 18236 16788
rect 18288 16776 18294 16788
rect 18325 16779 18383 16785
rect 18325 16776 18337 16779
rect 18288 16748 18337 16776
rect 18288 16736 18294 16748
rect 18325 16745 18337 16748
rect 18371 16745 18383 16779
rect 18325 16739 18383 16745
rect 19245 16779 19303 16785
rect 19245 16745 19257 16779
rect 19291 16776 19303 16779
rect 19334 16776 19340 16788
rect 19291 16748 19340 16776
rect 19291 16745 19303 16748
rect 19245 16739 19303 16745
rect 19334 16736 19340 16748
rect 19392 16736 19398 16788
rect 13262 16708 13268 16720
rect 13223 16680 13268 16708
rect 13262 16668 13268 16680
rect 13320 16668 13326 16720
rect 19794 16708 19800 16720
rect 19628 16680 19800 16708
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 4120 16612 4353 16640
rect 4120 16600 4126 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 6825 16643 6883 16649
rect 6825 16609 6837 16643
rect 6871 16609 6883 16643
rect 6825 16603 6883 16609
rect 8110 16600 8116 16652
rect 8168 16640 8174 16652
rect 9217 16643 9275 16649
rect 9217 16640 9229 16643
rect 8168 16612 9229 16640
rect 8168 16600 8174 16612
rect 9217 16609 9229 16612
rect 9263 16640 9275 16643
rect 9398 16640 9404 16652
rect 9263 16612 9404 16640
rect 9263 16609 9275 16612
rect 9217 16603 9275 16609
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 13394 16643 13452 16649
rect 13394 16609 13406 16643
rect 13440 16640 13452 16643
rect 13814 16640 13820 16652
rect 13440 16612 13820 16640
rect 13440 16609 13452 16612
rect 13394 16603 13452 16609
rect 1394 16572 1400 16584
rect 1355 16544 1400 16572
rect 1394 16532 1400 16544
rect 1452 16532 1458 16584
rect 2038 16532 2044 16584
rect 2096 16572 2102 16584
rect 2409 16575 2467 16581
rect 2409 16572 2421 16575
rect 2096 16544 2421 16572
rect 2096 16532 2102 16544
rect 2409 16541 2421 16544
rect 2455 16541 2467 16575
rect 2409 16535 2467 16541
rect 4246 16532 4252 16584
rect 4304 16572 4310 16584
rect 4597 16575 4655 16581
rect 4597 16572 4609 16575
rect 4304 16544 4609 16572
rect 4304 16532 4310 16544
rect 4597 16541 4609 16544
rect 4643 16541 4655 16575
rect 4597 16535 4655 16541
rect 6181 16575 6239 16581
rect 6181 16541 6193 16575
rect 6227 16572 6239 16575
rect 6638 16572 6644 16584
rect 6227 16544 6644 16572
rect 6227 16541 6239 16544
rect 6181 16535 6239 16541
rect 6638 16532 6644 16544
rect 6696 16532 6702 16584
rect 8941 16575 8999 16581
rect 8941 16541 8953 16575
rect 8987 16572 8999 16575
rect 9122 16572 9128 16584
rect 8987 16544 9128 16572
rect 8987 16541 8999 16544
rect 8941 16535 8999 16541
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 10226 16532 10232 16584
rect 10284 16572 10290 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 10284 16544 11989 16572
rect 10284 16532 10290 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16572 12403 16575
rect 13078 16572 13084 16584
rect 12391 16544 13084 16572
rect 12391 16541 12403 16544
rect 12345 16535 12403 16541
rect 13078 16532 13084 16544
rect 13136 16532 13142 16584
rect 13188 16572 13216 16603
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 14458 16600 14464 16652
rect 14516 16640 14522 16652
rect 14829 16643 14887 16649
rect 14829 16640 14841 16643
rect 14516 16612 14841 16640
rect 14516 16600 14522 16612
rect 14829 16609 14841 16612
rect 14875 16640 14887 16643
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 14875 16612 16957 16640
rect 14875 16609 14887 16612
rect 14829 16603 14887 16609
rect 16945 16609 16957 16612
rect 16991 16640 17003 16643
rect 19334 16640 19340 16652
rect 16991 16612 19340 16640
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 19628 16649 19656 16680
rect 19794 16668 19800 16680
rect 19852 16668 19858 16720
rect 19613 16643 19671 16649
rect 19613 16609 19625 16643
rect 19659 16609 19671 16643
rect 20162 16640 20168 16652
rect 19613 16603 19671 16609
rect 19904 16612 20168 16640
rect 19904 16584 19932 16612
rect 20162 16600 20168 16612
rect 20220 16600 20226 16652
rect 13630 16572 13636 16584
rect 13188 16544 13636 16572
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 15102 16572 15108 16584
rect 15063 16544 15108 16572
rect 15102 16532 15108 16544
rect 15160 16532 15166 16584
rect 16485 16575 16543 16581
rect 16485 16541 16497 16575
rect 16531 16572 16543 16575
rect 16758 16572 16764 16584
rect 16531 16544 16764 16572
rect 16531 16541 16543 16544
rect 16485 16535 16543 16541
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 17218 16572 17224 16584
rect 17179 16544 17224 16572
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 19426 16572 19432 16584
rect 19387 16544 19432 16572
rect 19426 16532 19432 16544
rect 19484 16532 19490 16584
rect 19693 16572 19699 16584
rect 19751 16581 19757 16584
rect 19660 16544 19699 16572
rect 19693 16532 19699 16544
rect 19751 16535 19760 16581
rect 19793 16575 19851 16581
rect 19793 16541 19805 16575
rect 19839 16572 19851 16575
rect 19886 16572 19892 16584
rect 19839 16544 19892 16572
rect 19839 16541 19851 16544
rect 19793 16535 19851 16541
rect 19751 16532 19757 16535
rect 19886 16532 19892 16544
rect 19944 16532 19950 16584
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16572 20039 16575
rect 20254 16572 20260 16584
rect 20027 16544 20260 16572
rect 20027 16541 20039 16544
rect 19981 16535 20039 16541
rect 20254 16532 20260 16544
rect 20312 16532 20318 16584
rect 20622 16572 20628 16584
rect 20583 16544 20628 16572
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 20881 16575 20939 16581
rect 20881 16572 20893 16575
rect 20772 16544 20893 16572
rect 20772 16532 20778 16544
rect 20881 16541 20893 16544
rect 20927 16541 20939 16575
rect 20881 16535 20939 16541
rect 29825 16575 29883 16581
rect 29825 16541 29837 16575
rect 29871 16572 29883 16575
rect 29914 16572 29920 16584
rect 29871 16544 29920 16572
rect 29871 16541 29883 16544
rect 29825 16535 29883 16541
rect 29914 16532 29920 16544
rect 29972 16532 29978 16584
rect 7092 16507 7150 16513
rect 7092 16473 7104 16507
rect 7138 16504 7150 16507
rect 7190 16504 7196 16516
rect 7138 16476 7196 16504
rect 7138 16473 7150 16476
rect 7092 16467 7150 16473
rect 7190 16464 7196 16476
rect 7248 16464 7254 16516
rect 12805 16507 12863 16513
rect 12805 16504 12817 16507
rect 7852 16476 12817 16504
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16436 1639 16439
rect 2222 16436 2228 16448
rect 1627 16408 2228 16436
rect 1627 16405 1639 16408
rect 1581 16399 1639 16405
rect 2222 16396 2228 16408
rect 2280 16396 2286 16448
rect 5718 16436 5724 16448
rect 5679 16408 5724 16436
rect 5718 16396 5724 16408
rect 5776 16436 5782 16448
rect 6822 16436 6828 16448
rect 5776 16408 6828 16436
rect 5776 16396 5782 16408
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7852 16436 7880 16476
rect 12805 16473 12817 16476
rect 12851 16473 12863 16507
rect 12805 16467 12863 16473
rect 13541 16507 13599 16513
rect 13541 16473 13553 16507
rect 13587 16504 13599 16507
rect 13722 16504 13728 16516
rect 13587 16476 13728 16504
rect 13587 16473 13599 16476
rect 13541 16467 13599 16473
rect 13722 16464 13728 16476
rect 13780 16464 13786 16516
rect 6972 16408 7880 16436
rect 8205 16439 8263 16445
rect 6972 16396 6978 16408
rect 8205 16405 8217 16439
rect 8251 16436 8263 16439
rect 8570 16436 8576 16448
rect 8251 16408 8576 16436
rect 8251 16405 8263 16408
rect 8205 16399 8263 16405
rect 8570 16396 8576 16408
rect 8628 16396 8634 16448
rect 12526 16396 12532 16448
rect 12584 16436 12590 16448
rect 18046 16436 18052 16448
rect 12584 16408 18052 16436
rect 12584 16396 12590 16408
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 19610 16396 19616 16448
rect 19668 16436 19674 16448
rect 22002 16436 22008 16448
rect 19668 16408 22008 16436
rect 19668 16396 19674 16408
rect 22002 16396 22008 16408
rect 22060 16396 22066 16448
rect 30006 16436 30012 16448
rect 29967 16408 30012 16436
rect 30006 16396 30012 16408
rect 30064 16396 30070 16448
rect 1104 16346 30820 16368
rect 1104 16294 10880 16346
rect 10932 16294 10944 16346
rect 10996 16294 11008 16346
rect 11060 16294 11072 16346
rect 11124 16294 11136 16346
rect 11188 16294 20811 16346
rect 20863 16294 20875 16346
rect 20927 16294 20939 16346
rect 20991 16294 21003 16346
rect 21055 16294 21067 16346
rect 21119 16294 30820 16346
rect 1104 16272 30820 16294
rect 7190 16232 7196 16244
rect 7151 16204 7196 16232
rect 7190 16192 7196 16204
rect 7248 16192 7254 16244
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 7742 16232 7748 16244
rect 7340 16204 7748 16232
rect 7340 16192 7346 16204
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 7926 16192 7932 16244
rect 7984 16232 7990 16244
rect 13446 16232 13452 16244
rect 7984 16204 9628 16232
rect 13407 16204 13452 16232
rect 7984 16192 7990 16204
rect 2774 16124 2780 16176
rect 2832 16164 2838 16176
rect 3786 16164 3792 16176
rect 2832 16136 3792 16164
rect 2832 16124 2838 16136
rect 3786 16124 3792 16136
rect 3844 16124 3850 16176
rect 8570 16164 8576 16176
rect 7484 16136 8576 16164
rect 7484 16120 7512 16136
rect 8570 16124 8576 16136
rect 8628 16124 8634 16176
rect 1210 16056 1216 16108
rect 1268 16096 1274 16108
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 1268 16068 1409 16096
rect 1268 16056 1274 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 2584 16099 2642 16105
rect 2584 16065 2596 16099
rect 2630 16096 2642 16099
rect 2866 16096 2872 16108
rect 2630 16068 2872 16096
rect 2630 16065 2642 16068
rect 2584 16059 2642 16065
rect 2866 16056 2872 16068
rect 2924 16056 2930 16108
rect 4430 16096 4436 16108
rect 4391 16068 4436 16096
rect 4430 16056 4436 16068
rect 4488 16056 4494 16108
rect 4706 16056 4712 16108
rect 4764 16096 4770 16108
rect 5445 16099 5503 16105
rect 5445 16096 5457 16099
rect 4764 16068 5457 16096
rect 4764 16056 4770 16068
rect 5445 16065 5457 16068
rect 5491 16065 5503 16099
rect 5445 16059 5503 16065
rect 6270 16056 6276 16108
rect 6328 16096 6334 16108
rect 6549 16099 6607 16105
rect 6549 16096 6561 16099
rect 6328 16068 6561 16096
rect 6328 16056 6334 16068
rect 6549 16065 6561 16068
rect 6595 16096 6607 16099
rect 6914 16096 6920 16108
rect 6595 16068 6920 16096
rect 6595 16065 6607 16068
rect 6549 16059 6607 16065
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7392 16105 7512 16120
rect 7377 16099 7512 16105
rect 7377 16065 7389 16099
rect 7423 16092 7512 16099
rect 7423 16065 7435 16092
rect 7377 16059 7435 16065
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 7926 16096 7932 16108
rect 7800 16068 7845 16096
rect 7887 16068 7932 16096
rect 7800 16056 7806 16068
rect 7926 16056 7932 16068
rect 7984 16056 7990 16108
rect 9033 16099 9091 16105
rect 9033 16096 9045 16099
rect 8680 16068 9045 16096
rect 2314 16028 2320 16040
rect 2275 16000 2320 16028
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 4154 16028 4160 16040
rect 4067 16000 4160 16028
rect 4154 15988 4160 16000
rect 4212 16028 4218 16040
rect 4522 16028 4528 16040
rect 4212 16000 4528 16028
rect 4212 15988 4218 16000
rect 4522 15988 4528 16000
rect 4580 16028 4586 16040
rect 6638 16028 6644 16040
rect 4580 16000 6644 16028
rect 4580 15988 4586 16000
rect 6638 15988 6644 16000
rect 6696 15988 6702 16040
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 7561 16031 7619 16037
rect 7561 16028 7573 16031
rect 7156 16000 7573 16028
rect 7156 15988 7162 16000
rect 7561 15997 7573 16000
rect 7607 15997 7619 16031
rect 7561 15991 7619 15997
rect 7659 16031 7717 16037
rect 7659 15997 7671 16031
rect 7705 16028 7717 16031
rect 8110 16028 8116 16040
rect 7705 16000 8116 16028
rect 7705 15997 7717 16000
rect 7659 15991 7717 15997
rect 8110 15988 8116 16000
rect 8168 15988 8174 16040
rect 8680 16028 8708 16068
rect 9033 16065 9045 16068
rect 9079 16096 9091 16099
rect 9490 16096 9496 16108
rect 9079 16068 9496 16096
rect 9079 16065 9091 16068
rect 9033 16059 9091 16065
rect 9490 16056 9496 16068
rect 9548 16056 9554 16108
rect 9600 16096 9628 16204
rect 13446 16192 13452 16204
rect 13504 16192 13510 16244
rect 13538 16192 13544 16244
rect 13596 16232 13602 16244
rect 14461 16235 14519 16241
rect 14461 16232 14473 16235
rect 13596 16204 14473 16232
rect 13596 16192 13602 16204
rect 14461 16201 14473 16204
rect 14507 16201 14519 16235
rect 15194 16232 15200 16244
rect 14461 16195 14519 16201
rect 14568 16204 15200 16232
rect 9950 16124 9956 16176
rect 10008 16164 10014 16176
rect 10778 16164 10784 16176
rect 10008 16136 10784 16164
rect 10008 16124 10014 16136
rect 10612 16105 10640 16136
rect 10778 16124 10784 16136
rect 10836 16124 10842 16176
rect 14568 16164 14596 16204
rect 15194 16192 15200 16204
rect 15252 16192 15258 16244
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 17276 16204 17417 16232
rect 17276 16192 17282 16204
rect 17405 16201 17417 16204
rect 17451 16201 17463 16235
rect 18598 16232 18604 16244
rect 17405 16195 17463 16201
rect 18524 16204 18604 16232
rect 13924 16136 14596 16164
rect 10045 16099 10103 16105
rect 10045 16096 10057 16099
rect 9600 16068 10057 16096
rect 10045 16065 10057 16068
rect 10091 16065 10103 16099
rect 10045 16059 10103 16065
rect 10229 16099 10287 16105
rect 10229 16065 10241 16099
rect 10275 16096 10287 16099
rect 10597 16099 10655 16105
rect 10275 16068 10539 16096
rect 10275 16065 10287 16068
rect 10229 16059 10287 16065
rect 8266 16000 8708 16028
rect 8757 16031 8815 16037
rect 3694 15960 3700 15972
rect 3607 15932 3700 15960
rect 3694 15920 3700 15932
rect 3752 15960 3758 15972
rect 7466 15960 7472 15972
rect 3752 15932 7472 15960
rect 3752 15920 3758 15932
rect 7466 15920 7472 15932
rect 7524 15920 7530 15972
rect 7926 15920 7932 15972
rect 7984 15960 7990 15972
rect 8266 15960 8294 16000
rect 8757 15997 8769 16031
rect 8803 15997 8815 16031
rect 8757 15991 8815 15997
rect 7984 15932 8294 15960
rect 8772 15960 8800 15991
rect 9122 15988 9128 16040
rect 9180 16028 9186 16040
rect 10321 16031 10379 16037
rect 10321 16028 10333 16031
rect 9180 16000 10333 16028
rect 9180 15988 9186 16000
rect 10321 15997 10333 16000
rect 10367 15997 10379 16031
rect 10321 15991 10379 15997
rect 10413 16031 10471 16037
rect 10413 15997 10425 16031
rect 10459 15997 10471 16031
rect 10413 15991 10471 15997
rect 9398 15960 9404 15972
rect 8772 15932 9404 15960
rect 7984 15920 7990 15932
rect 9398 15920 9404 15932
rect 9456 15960 9462 15972
rect 10428 15960 10456 15991
rect 9456 15932 10456 15960
rect 9456 15920 9462 15932
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 2958 15892 2964 15904
rect 1627 15864 2964 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 2958 15852 2964 15864
rect 3016 15852 3022 15904
rect 5537 15895 5595 15901
rect 5537 15861 5549 15895
rect 5583 15892 5595 15895
rect 5718 15892 5724 15904
rect 5583 15864 5724 15892
rect 5583 15861 5595 15864
rect 5537 15855 5595 15861
rect 5718 15852 5724 15864
rect 5776 15852 5782 15904
rect 6638 15892 6644 15904
rect 6599 15864 6644 15892
rect 6638 15852 6644 15864
rect 6696 15852 6702 15904
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 10511 15892 10539 16068
rect 10597 16065 10609 16099
rect 10643 16065 10655 16099
rect 10597 16059 10655 16065
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16065 12403 16099
rect 12526 16096 12532 16108
rect 12487 16068 12532 16096
rect 12345 16059 12403 16065
rect 12360 15960 12388 16059
rect 12526 16056 12532 16068
rect 12584 16056 12590 16108
rect 13630 16096 13636 16108
rect 13591 16068 13636 16096
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 13814 16096 13820 16108
rect 13775 16068 13820 16096
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 13924 16105 13952 16136
rect 14918 16124 14924 16176
rect 14976 16164 14982 16176
rect 18524 16173 18552 16204
rect 18598 16192 18604 16204
rect 18656 16192 18662 16244
rect 18690 16192 18696 16244
rect 18748 16232 18754 16244
rect 20254 16232 20260 16244
rect 18748 16204 20260 16232
rect 18748 16192 18754 16204
rect 20254 16192 20260 16204
rect 20312 16192 20318 16244
rect 18509 16167 18567 16173
rect 14976 16136 17080 16164
rect 14976 16124 14982 16136
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16065 13967 16099
rect 14642 16096 14648 16108
rect 14603 16068 14648 16096
rect 13909 16059 13967 16065
rect 14642 16056 14648 16068
rect 14700 16056 14706 16108
rect 14826 16096 14832 16108
rect 14787 16068 14832 16096
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 16666 16096 16672 16108
rect 16579 16068 16672 16096
rect 16666 16056 16672 16068
rect 16724 16056 16730 16108
rect 16850 16096 16856 16108
rect 16811 16068 16856 16096
rect 16850 16056 16856 16068
rect 16908 16056 16914 16108
rect 17052 16105 17080 16136
rect 18509 16133 18521 16167
rect 18555 16133 18567 16167
rect 18509 16127 18567 16133
rect 19978 16124 19984 16176
rect 20036 16164 20042 16176
rect 20134 16167 20192 16173
rect 20134 16164 20146 16167
rect 20036 16136 20146 16164
rect 20036 16124 20042 16136
rect 20134 16133 20146 16136
rect 20180 16133 20192 16167
rect 20134 16127 20192 16133
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16096 17279 16099
rect 17310 16096 17316 16108
rect 17267 16068 17316 16096
rect 17267 16065 17279 16068
rect 17221 16059 17279 16065
rect 14550 15988 14556 16040
rect 14608 16028 14614 16040
rect 16684 16028 16712 16056
rect 16942 16028 16948 16040
rect 14608 16000 16712 16028
rect 16903 16000 16948 16028
rect 14608 15988 14614 16000
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 17052 16028 17080 16059
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 18046 16056 18052 16108
rect 18104 16096 18110 16108
rect 18233 16099 18291 16105
rect 18233 16096 18245 16099
rect 18104 16068 18245 16096
rect 18104 16056 18110 16068
rect 18233 16065 18245 16068
rect 18279 16065 18291 16099
rect 18233 16059 18291 16065
rect 18371 16099 18429 16105
rect 18371 16065 18383 16099
rect 18417 16096 18429 16099
rect 18417 16068 18493 16096
rect 18417 16065 18429 16068
rect 18371 16059 18429 16065
rect 17862 16028 17868 16040
rect 17052 16000 17868 16028
rect 17862 15988 17868 16000
rect 17920 15988 17926 16040
rect 13262 15960 13268 15972
rect 12360 15932 13268 15960
rect 13262 15920 13268 15932
rect 13320 15960 13326 15972
rect 13722 15960 13728 15972
rect 13320 15932 13728 15960
rect 13320 15920 13326 15932
rect 13722 15920 13728 15932
rect 13780 15920 13786 15972
rect 14734 15920 14740 15972
rect 14792 15960 14798 15972
rect 16960 15960 16988 15988
rect 14792 15932 16988 15960
rect 18465 15960 18493 16068
rect 18598 16056 18604 16108
rect 18656 16096 18662 16108
rect 18739 16099 18797 16105
rect 18656 16068 18701 16096
rect 18656 16056 18662 16068
rect 18739 16065 18751 16099
rect 18785 16096 18797 16099
rect 18966 16096 18972 16108
rect 18785 16068 18972 16096
rect 18785 16065 18797 16068
rect 18739 16059 18797 16065
rect 18966 16056 18972 16068
rect 19024 16056 19030 16108
rect 20622 16096 20628 16108
rect 19904 16068 20628 16096
rect 19242 16028 19248 16040
rect 18616 16000 19248 16028
rect 18616 15960 18644 16000
rect 19242 15988 19248 16000
rect 19300 15988 19306 16040
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 19904 16037 19932 16068
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 19889 16031 19947 16037
rect 19889 16028 19901 16031
rect 19392 16000 19901 16028
rect 19392 15988 19398 16000
rect 19889 15997 19901 16000
rect 19935 15997 19947 16031
rect 19889 15991 19947 15997
rect 18465 15932 18644 15960
rect 14792 15920 14798 15932
rect 19058 15920 19064 15972
rect 19116 15960 19122 15972
rect 19702 15960 19708 15972
rect 19116 15932 19708 15960
rect 19116 15920 19122 15932
rect 19702 15920 19708 15932
rect 19760 15920 19766 15972
rect 10468 15864 10539 15892
rect 10468 15852 10474 15864
rect 10686 15852 10692 15904
rect 10744 15892 10750 15904
rect 10781 15895 10839 15901
rect 10781 15892 10793 15895
rect 10744 15864 10793 15892
rect 10744 15852 10750 15864
rect 10781 15861 10793 15864
rect 10827 15861 10839 15895
rect 10781 15855 10839 15861
rect 12250 15852 12256 15904
rect 12308 15892 12314 15904
rect 12345 15895 12403 15901
rect 12345 15892 12357 15895
rect 12308 15864 12357 15892
rect 12308 15852 12314 15864
rect 12345 15861 12357 15864
rect 12391 15861 12403 15895
rect 12345 15855 12403 15861
rect 18877 15895 18935 15901
rect 18877 15861 18889 15895
rect 18923 15892 18935 15895
rect 19518 15892 19524 15904
rect 18923 15864 19524 15892
rect 18923 15861 18935 15864
rect 18877 15855 18935 15861
rect 19518 15852 19524 15864
rect 19576 15852 19582 15904
rect 19886 15852 19892 15904
rect 19944 15892 19950 15904
rect 21269 15895 21327 15901
rect 21269 15892 21281 15895
rect 19944 15864 21281 15892
rect 19944 15852 19950 15864
rect 21269 15861 21281 15864
rect 21315 15861 21327 15895
rect 21269 15855 21327 15861
rect 1104 15802 30820 15824
rect 1104 15750 5915 15802
rect 5967 15750 5979 15802
rect 6031 15750 6043 15802
rect 6095 15750 6107 15802
rect 6159 15750 6171 15802
rect 6223 15750 15846 15802
rect 15898 15750 15910 15802
rect 15962 15750 15974 15802
rect 16026 15750 16038 15802
rect 16090 15750 16102 15802
rect 16154 15750 25776 15802
rect 25828 15750 25840 15802
rect 25892 15750 25904 15802
rect 25956 15750 25968 15802
rect 26020 15750 26032 15802
rect 26084 15750 30820 15802
rect 1104 15728 30820 15750
rect 2774 15688 2780 15700
rect 2148 15660 2780 15688
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15444 1458 15496
rect 2148 15493 2176 15660
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 4338 15648 4344 15700
rect 4396 15688 4402 15700
rect 4525 15691 4583 15697
rect 4525 15688 4537 15691
rect 4396 15660 4537 15688
rect 4396 15648 4402 15660
rect 4525 15657 4537 15660
rect 4571 15657 4583 15691
rect 4525 15651 4583 15657
rect 5828 15660 6040 15688
rect 2424 15592 3096 15620
rect 2424 15561 2452 15592
rect 3068 15564 3096 15592
rect 3142 15580 3148 15632
rect 3200 15620 3206 15632
rect 3200 15592 5028 15620
rect 3200 15580 3206 15592
rect 2409 15555 2467 15561
rect 2409 15521 2421 15555
rect 2455 15521 2467 15555
rect 2866 15552 2872 15564
rect 2827 15524 2872 15552
rect 2409 15515 2467 15521
rect 2866 15512 2872 15524
rect 2924 15512 2930 15564
rect 3050 15512 3056 15564
rect 3108 15552 3114 15564
rect 4062 15552 4068 15564
rect 3108 15524 4068 15552
rect 3108 15512 3114 15524
rect 4062 15512 4068 15524
rect 4120 15552 4126 15564
rect 4430 15552 4436 15564
rect 4120 15524 4436 15552
rect 4120 15512 4126 15524
rect 4430 15512 4436 15524
rect 4488 15512 4494 15564
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15453 2191 15487
rect 2133 15447 2191 15453
rect 2222 15444 2228 15496
rect 2280 15484 2286 15496
rect 2321 15487 2379 15493
rect 2321 15484 2333 15487
rect 2280 15456 2333 15484
rect 2280 15444 2286 15456
rect 2321 15453 2333 15456
rect 2367 15453 2379 15487
rect 2321 15447 2379 15453
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15484 2559 15487
rect 2685 15487 2743 15493
rect 2547 15456 2636 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 1946 15376 1952 15428
rect 2004 15416 2010 15428
rect 2608 15416 2636 15456
rect 2685 15453 2697 15487
rect 2731 15482 2743 15487
rect 3694 15484 3700 15496
rect 2792 15482 3700 15484
rect 2731 15456 3700 15482
rect 2731 15454 2820 15456
rect 2731 15453 2743 15454
rect 2685 15447 2743 15453
rect 3694 15444 3700 15456
rect 3752 15444 3758 15496
rect 3786 15444 3792 15496
rect 3844 15484 3850 15496
rect 3970 15484 3976 15496
rect 3844 15456 3889 15484
rect 3931 15456 3976 15484
rect 3844 15444 3850 15456
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15484 4399 15487
rect 4798 15484 4804 15496
rect 4387 15456 4804 15484
rect 4387 15453 4399 15456
rect 4341 15447 4399 15453
rect 4172 15416 4200 15447
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 5000 15493 5028 15592
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15453 5043 15487
rect 4985 15447 5043 15453
rect 5350 15444 5356 15496
rect 5408 15484 5414 15496
rect 5828 15493 5856 15660
rect 5902 15580 5908 15632
rect 5960 15580 5966 15632
rect 6012 15620 6040 15660
rect 6638 15648 6644 15700
rect 6696 15688 6702 15700
rect 6696 15660 7052 15688
rect 6696 15648 6702 15660
rect 6730 15620 6736 15632
rect 6012 15592 6736 15620
rect 6730 15580 6736 15592
rect 6788 15580 6794 15632
rect 6822 15580 6828 15632
rect 6880 15580 6886 15632
rect 7024 15620 7052 15660
rect 7098 15648 7104 15700
rect 7156 15688 7162 15700
rect 7926 15688 7932 15700
rect 7156 15660 7932 15688
rect 7156 15648 7162 15660
rect 7926 15648 7932 15660
rect 7984 15648 7990 15700
rect 9306 15648 9312 15700
rect 9364 15688 9370 15700
rect 11425 15691 11483 15697
rect 11425 15688 11437 15691
rect 9364 15660 11437 15688
rect 9364 15648 9370 15660
rect 11425 15657 11437 15660
rect 11471 15657 11483 15691
rect 11425 15651 11483 15657
rect 13357 15691 13415 15697
rect 13357 15657 13369 15691
rect 13403 15688 13415 15691
rect 13630 15688 13636 15700
rect 13403 15660 13636 15688
rect 13403 15657 13415 15660
rect 13357 15651 13415 15657
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 15746 15688 15752 15700
rect 14752 15660 15752 15688
rect 9766 15620 9772 15632
rect 7024 15592 9772 15620
rect 9766 15580 9772 15592
rect 9824 15580 9830 15632
rect 5920 15493 5948 15580
rect 6840 15552 6868 15580
rect 9306 15552 9312 15564
rect 6840 15524 8156 15552
rect 5629 15487 5687 15493
rect 5629 15484 5641 15487
rect 5408 15456 5641 15484
rect 5408 15444 5414 15456
rect 5629 15453 5641 15456
rect 5675 15453 5687 15487
rect 5629 15447 5687 15453
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15453 5871 15487
rect 5813 15447 5871 15453
rect 5899 15487 5957 15493
rect 5899 15453 5911 15487
rect 5945 15453 5957 15487
rect 5899 15447 5957 15453
rect 5997 15487 6055 15493
rect 5997 15453 6009 15487
rect 6043 15484 6055 15487
rect 6086 15484 6092 15496
rect 6043 15456 6092 15484
rect 6043 15453 6055 15456
rect 5997 15447 6055 15453
rect 6086 15444 6092 15456
rect 6144 15444 6150 15496
rect 6181 15487 6239 15493
rect 6181 15453 6193 15487
rect 6227 15484 6239 15487
rect 6454 15484 6460 15496
rect 6227 15456 6460 15484
rect 6227 15453 6239 15456
rect 6181 15447 6239 15453
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15453 6883 15487
rect 7466 15484 7472 15496
rect 7427 15456 7472 15484
rect 6825 15447 6883 15453
rect 2004 15388 4200 15416
rect 2004 15376 2010 15388
rect 5258 15376 5264 15428
rect 5316 15416 5322 15428
rect 6840 15416 6868 15447
rect 7466 15444 7472 15456
rect 7524 15444 7530 15496
rect 8128 15493 8156 15524
rect 9232 15524 9312 15552
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15453 8171 15487
rect 8386 15484 8392 15496
rect 8113 15447 8171 15453
rect 8220 15456 8392 15484
rect 5316 15388 6868 15416
rect 5316 15376 5322 15388
rect 7926 15376 7932 15428
rect 7984 15416 7990 15428
rect 8220 15416 8248 15456
rect 8386 15444 8392 15456
rect 8444 15484 8450 15496
rect 9122 15493 9128 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8444 15456 8953 15484
rect 8444 15444 8450 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9089 15487 9128 15493
rect 9089 15453 9101 15487
rect 9089 15447 9128 15453
rect 9122 15444 9128 15447
rect 9180 15444 9186 15496
rect 9232 15493 9260 15524
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 14752 15552 14780 15660
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 16117 15691 16175 15697
rect 16117 15657 16129 15691
rect 16163 15688 16175 15691
rect 16206 15688 16212 15700
rect 16163 15660 16212 15688
rect 16163 15657 16175 15660
rect 16117 15651 16175 15657
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 17034 15648 17040 15700
rect 17092 15688 17098 15700
rect 17129 15691 17187 15697
rect 17129 15688 17141 15691
rect 17092 15660 17141 15688
rect 17092 15648 17098 15660
rect 17129 15657 17141 15660
rect 17175 15657 17187 15691
rect 17678 15688 17684 15700
rect 17639 15660 17684 15688
rect 17129 15651 17187 15657
rect 17144 15620 17172 15651
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 17770 15648 17776 15700
rect 17828 15688 17834 15700
rect 20714 15688 20720 15700
rect 17828 15660 20720 15688
rect 17828 15648 17834 15660
rect 20714 15648 20720 15660
rect 20772 15688 20778 15700
rect 21085 15691 21143 15697
rect 21085 15688 21097 15691
rect 20772 15660 21097 15688
rect 20772 15648 20778 15660
rect 21085 15657 21097 15660
rect 21131 15657 21143 15691
rect 29914 15688 29920 15700
rect 29875 15660 29920 15688
rect 21085 15651 21143 15657
rect 29914 15648 29920 15660
rect 29972 15648 29978 15700
rect 30098 15648 30104 15700
rect 30156 15648 30162 15700
rect 18598 15620 18604 15632
rect 17144 15592 18604 15620
rect 18598 15580 18604 15592
rect 18656 15580 18662 15632
rect 19702 15580 19708 15632
rect 19760 15620 19766 15632
rect 20257 15623 20315 15629
rect 20257 15620 20269 15623
rect 19760 15592 20269 15620
rect 19760 15580 19766 15592
rect 20257 15589 20269 15592
rect 20303 15589 20315 15623
rect 20257 15583 20315 15589
rect 14660 15524 14780 15552
rect 14829 15555 14887 15561
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15453 9275 15487
rect 9217 15447 9275 15453
rect 9398 15444 9404 15496
rect 9456 15493 9462 15496
rect 9456 15484 9464 15493
rect 10042 15484 10048 15496
rect 9456 15456 9501 15484
rect 10003 15456 10048 15484
rect 9456 15447 9464 15456
rect 9456 15444 9462 15447
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 11974 15484 11980 15496
rect 11935 15456 11980 15484
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 12250 15493 12256 15496
rect 12244 15484 12256 15493
rect 12211 15456 12256 15484
rect 12244 15447 12256 15456
rect 12250 15444 12256 15447
rect 12308 15444 12314 15496
rect 13078 15444 13084 15496
rect 13136 15484 13142 15496
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 13136 15456 14473 15484
rect 13136 15444 13142 15456
rect 14461 15453 14473 15456
rect 14507 15484 14519 15487
rect 14550 15484 14556 15496
rect 14507 15456 14556 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 14660 15493 14688 15524
rect 14829 15521 14841 15555
rect 14875 15552 14887 15555
rect 14918 15552 14924 15564
rect 14875 15524 14924 15552
rect 14875 15521 14887 15524
rect 14829 15515 14887 15521
rect 14918 15512 14924 15524
rect 14976 15512 14982 15564
rect 16850 15512 16856 15564
rect 16908 15552 16914 15564
rect 17494 15552 17500 15564
rect 16908 15524 17500 15552
rect 16908 15512 16914 15524
rect 17494 15512 17500 15524
rect 17552 15552 17558 15564
rect 17773 15555 17831 15561
rect 17773 15552 17785 15555
rect 17552 15524 17785 15552
rect 17552 15512 17558 15524
rect 17773 15521 17785 15524
rect 17819 15552 17831 15555
rect 18230 15552 18236 15564
rect 17819 15524 18236 15552
rect 17819 15521 17831 15524
rect 17773 15515 17831 15521
rect 18230 15512 18236 15524
rect 18288 15512 18294 15564
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 15010 15484 15016 15496
rect 14792 15456 14837 15484
rect 14971 15456 15016 15484
rect 14792 15444 14798 15456
rect 15010 15444 15016 15456
rect 15068 15444 15074 15496
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 16209 15487 16267 15493
rect 16209 15484 16221 15487
rect 15804 15456 16221 15484
rect 15804 15444 15810 15456
rect 16209 15453 16221 15456
rect 16255 15453 16267 15487
rect 16209 15447 16267 15453
rect 17586 15444 17592 15496
rect 17644 15484 17650 15496
rect 17681 15487 17739 15493
rect 17681 15484 17693 15487
rect 17644 15456 17693 15484
rect 17644 15444 17650 15456
rect 17681 15453 17693 15456
rect 17727 15453 17739 15487
rect 19426 15484 19432 15496
rect 17681 15447 17739 15453
rect 18248 15456 19432 15484
rect 18248 15428 18276 15456
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 19610 15484 19616 15496
rect 19571 15456 19616 15484
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15484 19855 15487
rect 19886 15484 19892 15496
rect 19843 15456 19892 15484
rect 19843 15453 19855 15456
rect 19797 15447 19855 15453
rect 19886 15444 19892 15456
rect 19944 15444 19950 15496
rect 21269 15487 21327 15493
rect 21269 15453 21281 15487
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 7984 15388 8248 15416
rect 7984 15376 7990 15388
rect 8294 15376 8300 15428
rect 8352 15416 8358 15428
rect 9309 15419 9367 15425
rect 9309 15416 9321 15419
rect 8352 15388 9321 15416
rect 8352 15376 8358 15388
rect 9309 15385 9321 15388
rect 9355 15385 9367 15419
rect 10290 15419 10348 15425
rect 10290 15416 10302 15419
rect 9309 15379 9367 15385
rect 9600 15388 10302 15416
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 4062 15348 4068 15360
rect 1627 15320 4068 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 5077 15351 5135 15357
rect 5077 15317 5089 15351
rect 5123 15348 5135 15351
rect 6270 15348 6276 15360
rect 5123 15320 6276 15348
rect 5123 15317 5135 15320
rect 5077 15311 5135 15317
rect 6270 15308 6276 15320
rect 6328 15308 6334 15360
rect 6365 15351 6423 15357
rect 6365 15317 6377 15351
rect 6411 15348 6423 15351
rect 6822 15348 6828 15360
rect 6411 15320 6828 15348
rect 6411 15317 6423 15320
rect 6365 15311 6423 15317
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 6917 15351 6975 15357
rect 6917 15317 6929 15351
rect 6963 15348 6975 15351
rect 7098 15348 7104 15360
rect 6963 15320 7104 15348
rect 6963 15317 6975 15320
rect 6917 15311 6975 15317
rect 7098 15308 7104 15320
rect 7156 15308 7162 15360
rect 7558 15348 7564 15360
rect 7519 15320 7564 15348
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 7650 15308 7656 15360
rect 7708 15348 7714 15360
rect 9600 15357 9628 15388
rect 10290 15385 10302 15388
rect 10336 15385 10348 15419
rect 10290 15379 10348 15385
rect 10778 15376 10784 15428
rect 10836 15416 10842 15428
rect 16574 15416 16580 15428
rect 10836 15388 16580 15416
rect 10836 15376 10842 15388
rect 16574 15376 16580 15388
rect 16632 15376 16638 15428
rect 17037 15419 17095 15425
rect 17037 15385 17049 15419
rect 17083 15416 17095 15419
rect 17770 15416 17776 15428
rect 17083 15388 17776 15416
rect 17083 15385 17095 15388
rect 17037 15379 17095 15385
rect 17770 15376 17776 15388
rect 17828 15376 17834 15428
rect 18230 15416 18236 15428
rect 18064 15388 18236 15416
rect 8205 15351 8263 15357
rect 8205 15348 8217 15351
rect 7708 15320 8217 15348
rect 7708 15308 7714 15320
rect 8205 15317 8217 15320
rect 8251 15317 8263 15351
rect 8205 15311 8263 15317
rect 9585 15351 9643 15357
rect 9585 15317 9597 15351
rect 9631 15317 9643 15351
rect 15194 15348 15200 15360
rect 15155 15320 15200 15348
rect 9585 15311 9643 15317
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 18064 15357 18092 15388
rect 18230 15376 18236 15388
rect 18288 15376 18294 15428
rect 19242 15376 19248 15428
rect 19300 15416 19306 15428
rect 20441 15419 20499 15425
rect 20441 15416 20453 15419
rect 19300 15388 20453 15416
rect 19300 15376 19306 15388
rect 20441 15385 20453 15388
rect 20487 15385 20499 15419
rect 21284 15416 21312 15447
rect 21542 15444 21548 15496
rect 21600 15484 21606 15496
rect 22005 15487 22063 15493
rect 22005 15484 22017 15487
rect 21600 15456 22017 15484
rect 21600 15444 21606 15456
rect 22005 15453 22017 15456
rect 22051 15453 22063 15487
rect 29914 15484 29920 15496
rect 29875 15456 29920 15484
rect 22005 15447 22063 15453
rect 29914 15444 29920 15456
rect 29972 15444 29978 15496
rect 30116 15493 30144 15648
rect 30101 15487 30159 15493
rect 30101 15453 30113 15487
rect 30147 15484 30159 15487
rect 30282 15484 30288 15496
rect 30147 15456 30288 15484
rect 30147 15453 30159 15456
rect 30101 15447 30159 15453
rect 30282 15444 30288 15456
rect 30340 15444 30346 15496
rect 22738 15416 22744 15428
rect 21284 15388 22744 15416
rect 20441 15379 20499 15385
rect 22738 15376 22744 15388
rect 22796 15376 22802 15428
rect 18049 15351 18107 15357
rect 18049 15317 18061 15351
rect 18095 15317 18107 15351
rect 18049 15311 18107 15317
rect 18138 15308 18144 15360
rect 18196 15348 18202 15360
rect 19429 15351 19487 15357
rect 19429 15348 19441 15351
rect 18196 15320 19441 15348
rect 18196 15308 18202 15320
rect 19429 15317 19441 15320
rect 19475 15317 19487 15351
rect 21818 15348 21824 15360
rect 21779 15320 21824 15348
rect 19429 15311 19487 15317
rect 21818 15308 21824 15320
rect 21876 15308 21882 15360
rect 1104 15258 30820 15280
rect 1104 15206 10880 15258
rect 10932 15206 10944 15258
rect 10996 15206 11008 15258
rect 11060 15206 11072 15258
rect 11124 15206 11136 15258
rect 11188 15206 20811 15258
rect 20863 15206 20875 15258
rect 20927 15206 20939 15258
rect 20991 15206 21003 15258
rect 21055 15206 21067 15258
rect 21119 15206 30820 15258
rect 1104 15184 30820 15206
rect 5258 15144 5264 15156
rect 3252 15116 5264 15144
rect 2774 15036 2780 15088
rect 2832 15036 2838 15088
rect 2958 15076 2964 15088
rect 2884 15048 2964 15076
rect 1397 15011 1455 15017
rect 1397 14977 1409 15011
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2685 15011 2743 15017
rect 2685 14977 2697 15011
rect 2731 15008 2743 15011
rect 2792 15008 2820 15036
rect 2884 15017 2912 15048
rect 2958 15036 2964 15048
rect 3016 15036 3022 15088
rect 3252 15017 3280 15116
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 6086 15104 6092 15156
rect 6144 15144 6150 15156
rect 6730 15144 6736 15156
rect 6144 15116 6736 15144
rect 6144 15104 6150 15116
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 8846 15144 8852 15156
rect 8759 15116 8852 15144
rect 8846 15104 8852 15116
rect 8904 15144 8910 15156
rect 9398 15144 9404 15156
rect 8904 15116 9404 15144
rect 8904 15104 8910 15116
rect 9398 15104 9404 15116
rect 9456 15104 9462 15156
rect 9490 15104 9496 15156
rect 9548 15144 9554 15156
rect 14001 15147 14059 15153
rect 9548 15116 12434 15144
rect 9548 15104 9554 15116
rect 3421 15079 3479 15085
rect 3421 15045 3433 15079
rect 3467 15076 3479 15079
rect 4126 15079 4184 15085
rect 4126 15076 4138 15079
rect 3467 15048 4138 15076
rect 3467 15045 3479 15048
rect 3421 15039 3479 15045
rect 4126 15045 4138 15048
rect 4172 15045 4184 15079
rect 4126 15039 4184 15045
rect 4246 15036 4252 15088
rect 4304 15036 4310 15088
rect 5534 15036 5540 15088
rect 5592 15076 5598 15088
rect 12069 15079 12127 15085
rect 12069 15076 12081 15079
rect 5592 15048 12081 15076
rect 5592 15036 5598 15048
rect 12069 15045 12081 15048
rect 12115 15045 12127 15079
rect 12406 15076 12434 15116
rect 14001 15113 14013 15147
rect 14047 15144 14059 15147
rect 14642 15144 14648 15156
rect 14047 15116 14648 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 14642 15104 14648 15116
rect 14700 15104 14706 15156
rect 15562 15104 15568 15156
rect 15620 15144 15626 15156
rect 16758 15144 16764 15156
rect 15620 15116 16764 15144
rect 15620 15104 15626 15116
rect 16758 15104 16764 15116
rect 16816 15104 16822 15156
rect 17862 15104 17868 15156
rect 17920 15144 17926 15156
rect 19061 15147 19119 15153
rect 19061 15144 19073 15147
rect 17920 15116 19073 15144
rect 17920 15104 17926 15116
rect 19061 15113 19073 15116
rect 19107 15144 19119 15147
rect 19794 15144 19800 15156
rect 19107 15116 19800 15144
rect 19107 15113 19119 15116
rect 19061 15107 19119 15113
rect 19794 15104 19800 15116
rect 19852 15104 19858 15156
rect 29178 15104 29184 15156
rect 29236 15144 29242 15156
rect 29273 15147 29331 15153
rect 29273 15144 29285 15147
rect 29236 15116 29285 15144
rect 29236 15104 29242 15116
rect 29273 15113 29285 15116
rect 29319 15113 29331 15147
rect 29273 15107 29331 15113
rect 14728 15079 14786 15085
rect 12406 15048 14688 15076
rect 12069 15039 12127 15045
rect 2731 14980 2820 15008
rect 2869 15011 2927 15017
rect 2731 14977 2743 14980
rect 2685 14971 2743 14977
rect 2869 14977 2881 15011
rect 2915 14977 2927 15011
rect 2869 14971 2927 14977
rect 3237 15011 3295 15017
rect 3237 14977 3249 15011
rect 3283 14977 3295 15011
rect 4264 15008 4292 15036
rect 3237 14971 3295 14977
rect 3804 14980 4292 15008
rect 1210 14900 1216 14952
rect 1268 14940 1274 14952
rect 1412 14940 1440 14971
rect 1268 14912 1440 14940
rect 2240 14940 2268 14971
rect 2774 14940 2780 14952
rect 2240 14912 2780 14940
rect 1268 14900 1274 14912
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 2958 14940 2964 14952
rect 2919 14912 2964 14940
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 3053 14943 3111 14949
rect 3053 14909 3065 14943
rect 3099 14940 3111 14943
rect 3804 14940 3832 14980
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 5316 14980 6377 15008
rect 5316 14968 5322 14980
rect 6365 14977 6377 14980
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 6454 14968 6460 15020
rect 6512 15008 6518 15020
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 6512 14980 6561 15008
rect 6512 14968 6518 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6730 15008 6736 15020
rect 6691 14980 6736 15008
rect 6549 14971 6607 14977
rect 6730 14968 6736 14980
rect 6788 14968 6794 15020
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7558 15008 7564 15020
rect 6963 14980 7564 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 15008 8815 15011
rect 9122 15008 9128 15020
rect 8803 14980 9128 15008
rect 8803 14977 8815 14980
rect 8757 14971 8815 14977
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 10686 14968 10692 15020
rect 10744 15017 10750 15020
rect 10744 15008 10756 15017
rect 10965 15011 11023 15017
rect 10744 14980 10789 15008
rect 10744 14971 10756 14980
rect 10965 14977 10977 15011
rect 11011 15008 11023 15011
rect 11974 15008 11980 15020
rect 11011 14980 11980 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 10744 14968 10750 14971
rect 11974 14968 11980 14980
rect 12032 15008 12038 15020
rect 12434 15008 12440 15020
rect 12032 14980 12440 15008
rect 12032 14968 12038 14980
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 12526 14968 12532 15020
rect 12584 15008 12590 15020
rect 12710 15008 12716 15020
rect 12584 14980 12629 15008
rect 12671 14980 12716 15008
rect 12584 14968 12590 14980
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 13541 15011 13599 15017
rect 13541 14977 13553 15011
rect 13587 15008 13599 15011
rect 13630 15008 13636 15020
rect 13587 14980 13636 15008
rect 13587 14977 13599 14980
rect 13541 14971 13599 14977
rect 13630 14968 13636 14980
rect 13688 14968 13694 15020
rect 13814 15008 13820 15020
rect 13775 14980 13820 15008
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14660 15008 14688 15048
rect 14728 15045 14740 15079
rect 14774 15076 14786 15079
rect 15194 15076 15200 15088
rect 14774 15048 15200 15076
rect 14774 15045 14786 15048
rect 14728 15039 14786 15045
rect 15194 15036 15200 15048
rect 15252 15036 15258 15088
rect 15746 15036 15752 15088
rect 15804 15076 15810 15088
rect 16853 15079 16911 15085
rect 16853 15076 16865 15079
rect 15804 15048 16865 15076
rect 15804 15036 15810 15048
rect 16853 15045 16865 15048
rect 16899 15045 16911 15079
rect 16853 15039 16911 15045
rect 16942 15036 16948 15088
rect 17000 15076 17006 15088
rect 17037 15079 17095 15085
rect 17037 15076 17049 15079
rect 17000 15048 17049 15076
rect 17000 15036 17006 15048
rect 17037 15045 17049 15048
rect 17083 15076 17095 15079
rect 17586 15076 17592 15088
rect 17083 15048 17592 15076
rect 17083 15045 17095 15048
rect 17037 15039 17095 15045
rect 17586 15036 17592 15048
rect 17644 15036 17650 15088
rect 17954 15036 17960 15088
rect 18012 15076 18018 15088
rect 18049 15079 18107 15085
rect 18049 15076 18061 15079
rect 18012 15048 18061 15076
rect 18012 15036 18018 15048
rect 18049 15045 18061 15048
rect 18095 15076 18107 15079
rect 18138 15076 18144 15088
rect 18095 15048 18144 15076
rect 18095 15045 18107 15048
rect 18049 15039 18107 15045
rect 18138 15036 18144 15048
rect 18196 15036 18202 15088
rect 18230 15036 18236 15088
rect 18288 15076 18294 15088
rect 18966 15076 18972 15088
rect 18288 15048 18333 15076
rect 18927 15048 18972 15076
rect 18288 15036 18294 15048
rect 18966 15036 18972 15048
rect 19024 15036 19030 15088
rect 21821 15079 21879 15085
rect 21821 15045 21833 15079
rect 21867 15076 21879 15079
rect 22738 15076 22744 15088
rect 21867 15048 22744 15076
rect 21867 15045 21879 15048
rect 21821 15039 21879 15045
rect 22738 15036 22744 15048
rect 22796 15036 22802 15088
rect 16574 15008 16580 15020
rect 14660 14980 16580 15008
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 16669 15011 16727 15017
rect 16669 14977 16681 15011
rect 16715 15008 16727 15011
rect 16758 15008 16764 15020
rect 16715 14980 16764 15008
rect 16715 14977 16727 14980
rect 16669 14971 16727 14977
rect 16758 14968 16764 14980
rect 16816 14968 16822 15020
rect 20438 14968 20444 15020
rect 20496 15008 20502 15020
rect 20533 15011 20591 15017
rect 20533 15008 20545 15011
rect 20496 14980 20545 15008
rect 20496 14968 20502 14980
rect 20533 14977 20545 14980
rect 20579 14977 20591 15011
rect 20533 14971 20591 14977
rect 20622 14968 20628 15020
rect 20680 15008 20686 15020
rect 20680 14980 20725 15008
rect 20680 14968 20686 14980
rect 21450 14968 21456 15020
rect 21508 15008 21514 15020
rect 21910 15008 21916 15020
rect 21508 14980 21916 15008
rect 21508 14968 21514 14980
rect 21910 14968 21916 14980
rect 21968 15008 21974 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21968 14980 22017 15008
rect 21968 14968 21974 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 29178 15008 29184 15020
rect 29139 14980 29184 15008
rect 22005 14971 22063 14977
rect 29178 14968 29184 14980
rect 29236 14968 29242 15020
rect 29365 15011 29423 15017
rect 29365 14977 29377 15011
rect 29411 14977 29423 15011
rect 29822 15008 29828 15020
rect 29783 14980 29828 15008
rect 29365 14971 29423 14977
rect 3099 14912 3832 14940
rect 3881 14943 3939 14949
rect 3099 14909 3111 14912
rect 3053 14903 3111 14909
rect 3881 14909 3893 14943
rect 3927 14909 3939 14943
rect 3881 14903 3939 14909
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14909 6699 14943
rect 9674 14940 9680 14952
rect 6641 14903 6699 14909
rect 7024 14912 9680 14940
rect 1486 14832 1492 14884
rect 1544 14872 1550 14884
rect 2314 14872 2320 14884
rect 1544 14844 2320 14872
rect 1544 14832 1550 14844
rect 2314 14832 2320 14844
rect 2372 14872 2378 14884
rect 3896 14872 3924 14903
rect 2372 14844 3924 14872
rect 2372 14832 2378 14844
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14804 1639 14807
rect 1854 14804 1860 14816
rect 1627 14776 1860 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 1946 14764 1952 14816
rect 2004 14804 2010 14816
rect 2041 14807 2099 14813
rect 2041 14804 2053 14807
rect 2004 14776 2053 14804
rect 2004 14764 2010 14776
rect 2041 14773 2053 14776
rect 2087 14773 2099 14807
rect 3896 14804 3924 14844
rect 5902 14832 5908 14884
rect 5960 14872 5966 14884
rect 6362 14872 6368 14884
rect 5960 14844 6368 14872
rect 5960 14832 5966 14844
rect 6362 14832 6368 14844
rect 6420 14872 6426 14884
rect 6656 14872 6684 14903
rect 6420 14844 6684 14872
rect 6420 14832 6426 14844
rect 6822 14832 6828 14884
rect 6880 14872 6886 14884
rect 7024 14872 7052 14912
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 12802 14940 12808 14952
rect 12763 14912 12808 14940
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 14458 14940 14464 14952
rect 14419 14912 14464 14940
rect 14458 14900 14464 14912
rect 14516 14900 14522 14952
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 17402 14940 17408 14952
rect 15528 14912 17408 14940
rect 15528 14900 15534 14912
rect 17402 14900 17408 14912
rect 17460 14900 17466 14952
rect 20254 14940 20260 14952
rect 20215 14912 20260 14940
rect 20254 14900 20260 14912
rect 20312 14900 20318 14952
rect 29380 14940 29408 14971
rect 29822 14968 29828 14980
rect 29880 14968 29886 15020
rect 30282 14940 30288 14952
rect 29380 14912 30288 14940
rect 30282 14900 30288 14912
rect 30340 14900 30346 14952
rect 6880 14844 7052 14872
rect 7101 14875 7159 14881
rect 6880 14832 6886 14844
rect 7101 14841 7113 14875
rect 7147 14872 7159 14875
rect 17865 14875 17923 14881
rect 17865 14872 17877 14875
rect 7147 14844 10088 14872
rect 7147 14841 7159 14844
rect 7101 14835 7159 14841
rect 5166 14804 5172 14816
rect 3896 14776 5172 14804
rect 2041 14767 2099 14773
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 9490 14804 9496 14816
rect 6512 14776 9496 14804
rect 6512 14764 6518 14776
rect 9490 14764 9496 14776
rect 9548 14764 9554 14816
rect 9585 14807 9643 14813
rect 9585 14773 9597 14807
rect 9631 14804 9643 14807
rect 9950 14804 9956 14816
rect 9631 14776 9956 14804
rect 9631 14773 9643 14776
rect 9585 14767 9643 14773
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10060 14804 10088 14844
rect 15396 14844 17877 14872
rect 12342 14804 12348 14816
rect 10060 14776 12348 14804
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 12526 14764 12532 14816
rect 12584 14804 12590 14816
rect 13633 14807 13691 14813
rect 13633 14804 13645 14807
rect 12584 14776 13645 14804
rect 12584 14764 12590 14776
rect 13633 14773 13645 14776
rect 13679 14804 13691 14807
rect 13722 14804 13728 14816
rect 13679 14776 13728 14804
rect 13679 14773 13691 14776
rect 13633 14767 13691 14773
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 14642 14764 14648 14816
rect 14700 14804 14706 14816
rect 14826 14804 14832 14816
rect 14700 14776 14832 14804
rect 14700 14764 14706 14776
rect 14826 14764 14832 14776
rect 14884 14804 14890 14816
rect 15396 14804 15424 14844
rect 17865 14841 17877 14844
rect 17911 14841 17923 14875
rect 17865 14835 17923 14841
rect 20809 14875 20867 14881
rect 20809 14841 20821 14875
rect 20855 14872 20867 14875
rect 29638 14872 29644 14884
rect 20855 14844 29644 14872
rect 20855 14841 20867 14844
rect 20809 14835 20867 14841
rect 29638 14832 29644 14844
rect 29696 14832 29702 14884
rect 14884 14776 15424 14804
rect 14884 14764 14890 14776
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 15804 14776 15853 14804
rect 15804 14764 15810 14776
rect 15841 14773 15853 14776
rect 15887 14773 15899 14807
rect 15841 14767 15899 14773
rect 19150 14764 19156 14816
rect 19208 14804 19214 14816
rect 20349 14807 20407 14813
rect 20349 14804 20361 14807
rect 19208 14776 20361 14804
rect 19208 14764 19214 14776
rect 20349 14773 20361 14776
rect 20395 14773 20407 14807
rect 20349 14767 20407 14773
rect 22189 14807 22247 14813
rect 22189 14773 22201 14807
rect 22235 14804 22247 14807
rect 22278 14804 22284 14816
rect 22235 14776 22284 14804
rect 22235 14773 22247 14776
rect 22189 14767 22247 14773
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 30006 14804 30012 14816
rect 29967 14776 30012 14804
rect 30006 14764 30012 14776
rect 30064 14764 30070 14816
rect 1104 14714 30820 14736
rect 1104 14662 5915 14714
rect 5967 14662 5979 14714
rect 6031 14662 6043 14714
rect 6095 14662 6107 14714
rect 6159 14662 6171 14714
rect 6223 14662 15846 14714
rect 15898 14662 15910 14714
rect 15962 14662 15974 14714
rect 16026 14662 16038 14714
rect 16090 14662 16102 14714
rect 16154 14662 25776 14714
rect 25828 14662 25840 14714
rect 25892 14662 25904 14714
rect 25956 14662 25968 14714
rect 26020 14662 26032 14714
rect 26084 14662 30820 14714
rect 1104 14640 30820 14662
rect 2869 14603 2927 14609
rect 2869 14569 2881 14603
rect 2915 14600 2927 14603
rect 3142 14600 3148 14612
rect 2915 14572 3148 14600
rect 2915 14569 2927 14572
rect 2869 14563 2927 14569
rect 3142 14560 3148 14572
rect 3200 14560 3206 14612
rect 6454 14600 6460 14612
rect 6415 14572 6460 14600
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 7653 14603 7711 14609
rect 7653 14569 7665 14603
rect 7699 14600 7711 14603
rect 11882 14600 11888 14612
rect 7699 14572 11888 14600
rect 7699 14569 7711 14572
rect 7653 14563 7711 14569
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 11977 14603 12035 14609
rect 11977 14569 11989 14603
rect 12023 14600 12035 14603
rect 12710 14600 12716 14612
rect 12023 14572 12716 14600
rect 12023 14569 12035 14572
rect 11977 14563 12035 14569
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 14553 14603 14611 14609
rect 14553 14600 14565 14603
rect 14332 14572 14565 14600
rect 14332 14560 14338 14572
rect 14553 14569 14565 14572
rect 14599 14569 14611 14603
rect 14553 14563 14611 14569
rect 16117 14603 16175 14609
rect 16117 14569 16129 14603
rect 16163 14569 16175 14603
rect 16117 14563 16175 14569
rect 6086 14492 6092 14544
rect 6144 14532 6150 14544
rect 6730 14532 6736 14544
rect 6144 14504 6736 14532
rect 6144 14492 6150 14504
rect 6730 14492 6736 14504
rect 6788 14532 6794 14544
rect 8110 14532 8116 14544
rect 6788 14504 8116 14532
rect 6788 14492 6794 14504
rect 8110 14492 8116 14504
rect 8168 14492 8174 14544
rect 9950 14492 9956 14544
rect 10008 14532 10014 14544
rect 10321 14535 10379 14541
rect 10321 14532 10333 14535
rect 10008 14504 10333 14532
rect 10008 14492 10014 14504
rect 10321 14501 10333 14504
rect 10367 14532 10379 14535
rect 10778 14532 10784 14544
rect 10367 14504 10784 14532
rect 10367 14501 10379 14504
rect 10321 14495 10379 14501
rect 10778 14492 10784 14504
rect 10836 14492 10842 14544
rect 16022 14492 16028 14544
rect 16080 14532 16086 14544
rect 16132 14532 16160 14563
rect 16298 14560 16304 14612
rect 16356 14600 16362 14612
rect 22097 14603 22155 14609
rect 22097 14600 22109 14603
rect 16356 14572 22109 14600
rect 16356 14560 16362 14572
rect 22097 14569 22109 14572
rect 22143 14569 22155 14603
rect 22097 14563 22155 14569
rect 28997 14603 29055 14609
rect 28997 14569 29009 14603
rect 29043 14600 29055 14603
rect 29822 14600 29828 14612
rect 29043 14572 29828 14600
rect 29043 14569 29055 14572
rect 28997 14563 29055 14569
rect 29822 14560 29828 14572
rect 29880 14560 29886 14612
rect 16080 14504 16160 14532
rect 16080 14492 16086 14504
rect 16574 14492 16580 14544
rect 16632 14532 16638 14544
rect 19797 14535 19855 14541
rect 19797 14532 19809 14535
rect 16632 14504 19809 14532
rect 16632 14492 16638 14504
rect 19797 14501 19809 14504
rect 19843 14501 19855 14535
rect 19797 14495 19855 14501
rect 20257 14535 20315 14541
rect 20257 14501 20269 14535
rect 20303 14532 20315 14535
rect 29914 14532 29920 14544
rect 20303 14504 29920 14532
rect 20303 14501 20315 14504
rect 20257 14495 20315 14501
rect 29914 14492 29920 14504
rect 29972 14492 29978 14544
rect 30098 14532 30104 14544
rect 30024 14504 30104 14532
rect 5166 14464 5172 14476
rect 5127 14436 5172 14464
rect 5166 14424 5172 14436
rect 5224 14424 5230 14476
rect 6454 14464 6460 14476
rect 5736 14436 6460 14464
rect 1486 14396 1492 14408
rect 1447 14368 1492 14396
rect 1486 14356 1492 14368
rect 1544 14356 1550 14408
rect 2590 14356 2596 14408
rect 2648 14396 2654 14408
rect 5534 14396 5540 14408
rect 2648 14368 5540 14396
rect 2648 14356 2654 14368
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5736 14405 5764 14436
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 7006 14424 7012 14476
rect 7064 14464 7070 14476
rect 7285 14467 7343 14473
rect 7285 14464 7297 14467
rect 7064 14436 7297 14464
rect 7064 14424 7070 14436
rect 7285 14433 7297 14436
rect 7331 14464 7343 14467
rect 8294 14464 8300 14476
rect 7331 14436 8300 14464
rect 7331 14433 7343 14436
rect 7285 14427 7343 14433
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 12526 14424 12532 14476
rect 12584 14464 12590 14476
rect 12713 14467 12771 14473
rect 12713 14464 12725 14467
rect 12584 14436 12725 14464
rect 12584 14424 12590 14436
rect 12713 14433 12725 14436
rect 12759 14433 12771 14467
rect 13630 14464 13636 14476
rect 12713 14427 12771 14433
rect 13372 14436 13636 14464
rect 5721 14399 5779 14405
rect 5721 14365 5733 14399
rect 5767 14365 5779 14399
rect 5721 14359 5779 14365
rect 5810 14356 5816 14408
rect 5868 14396 5874 14408
rect 5905 14399 5963 14405
rect 5905 14396 5917 14399
rect 5868 14368 5917 14396
rect 5868 14356 5874 14368
rect 5905 14365 5917 14368
rect 5951 14365 5963 14399
rect 5905 14359 5963 14365
rect 5997 14399 6055 14405
rect 5997 14365 6009 14399
rect 6043 14365 6055 14399
rect 5997 14359 6055 14365
rect 1394 14288 1400 14340
rect 1452 14328 1458 14340
rect 1734 14331 1792 14337
rect 1734 14328 1746 14331
rect 1452 14300 1746 14328
rect 1452 14288 1458 14300
rect 1734 14297 1746 14300
rect 1780 14297 1792 14331
rect 1734 14291 1792 14297
rect 2406 14288 2412 14340
rect 2464 14328 2470 14340
rect 2464 14300 4568 14328
rect 2464 14288 2470 14300
rect 3786 14260 3792 14272
rect 3747 14232 3792 14260
rect 3786 14220 3792 14232
rect 3844 14220 3850 14272
rect 4540 14260 4568 14300
rect 4614 14288 4620 14340
rect 4672 14328 4678 14340
rect 4902 14331 4960 14337
rect 4902 14328 4914 14331
rect 4672 14300 4914 14328
rect 4672 14288 4678 14300
rect 4902 14297 4914 14300
rect 4948 14297 4960 14331
rect 6012 14328 6040 14359
rect 6086 14356 6092 14408
rect 6144 14396 6150 14408
rect 6270 14396 6276 14408
rect 6144 14368 6189 14396
rect 6231 14368 6276 14396
rect 6144 14356 6150 14368
rect 6270 14356 6276 14368
rect 6328 14356 6334 14408
rect 6638 14356 6644 14408
rect 6696 14396 6702 14408
rect 6917 14399 6975 14405
rect 6917 14396 6929 14399
rect 6696 14368 6929 14396
rect 6696 14356 6702 14368
rect 6917 14365 6929 14368
rect 6963 14365 6975 14399
rect 7098 14396 7104 14408
rect 7059 14368 7104 14396
rect 6917 14359 6975 14365
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14365 7251 14399
rect 7193 14359 7251 14365
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14396 7527 14399
rect 8018 14396 8024 14408
rect 7515 14368 8024 14396
rect 7515 14365 7527 14368
rect 7469 14359 7527 14365
rect 6012 14300 6316 14328
rect 4902 14291 4960 14297
rect 6288 14272 6316 14300
rect 6178 14260 6184 14272
rect 4540 14232 6184 14260
rect 6178 14220 6184 14232
rect 6236 14220 6242 14272
rect 6270 14220 6276 14272
rect 6328 14220 6334 14272
rect 7098 14220 7104 14272
rect 7156 14260 7162 14272
rect 7208 14260 7236 14359
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 8941 14399 8999 14405
rect 8941 14365 8953 14399
rect 8987 14396 8999 14399
rect 10042 14396 10048 14408
rect 8987 14368 10048 14396
rect 8987 14365 8999 14368
rect 8941 14359 8999 14365
rect 10042 14356 10048 14368
rect 10100 14356 10106 14408
rect 11790 14396 11796 14408
rect 11751 14368 11796 14396
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 13372 14405 13400 14436
rect 13630 14424 13636 14436
rect 13688 14424 13694 14476
rect 16114 14464 16120 14476
rect 16075 14436 16120 14464
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 18138 14464 18144 14476
rect 18099 14436 18144 14464
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 18230 14424 18236 14476
rect 18288 14464 18294 14476
rect 18288 14436 18460 14464
rect 18288 14424 18294 14436
rect 13357 14399 13415 14405
rect 12406 14368 13308 14396
rect 8110 14288 8116 14340
rect 8168 14328 8174 14340
rect 8205 14331 8263 14337
rect 8205 14328 8217 14331
rect 8168 14300 8217 14328
rect 8168 14288 8174 14300
rect 8205 14297 8217 14300
rect 8251 14297 8263 14331
rect 8205 14291 8263 14297
rect 8662 14288 8668 14340
rect 8720 14328 8726 14340
rect 9186 14331 9244 14337
rect 9186 14328 9198 14331
rect 8720 14300 9198 14328
rect 8720 14288 8726 14300
rect 9186 14297 9198 14300
rect 9232 14297 9244 14331
rect 12406 14328 12434 14368
rect 9186 14291 9244 14297
rect 9324 14300 12434 14328
rect 12529 14331 12587 14337
rect 8297 14263 8355 14269
rect 8297 14260 8309 14263
rect 7156 14232 8309 14260
rect 7156 14220 7162 14232
rect 8297 14229 8309 14232
rect 8343 14260 8355 14263
rect 9324 14260 9352 14300
rect 12529 14297 12541 14331
rect 12575 14328 12587 14331
rect 12894 14328 12900 14340
rect 12575 14300 12900 14328
rect 12575 14297 12587 14300
rect 12529 14291 12587 14297
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 13280 14328 13308 14368
rect 13357 14365 13369 14399
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 13814 14396 13820 14408
rect 13587 14368 13820 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 14642 14396 14648 14408
rect 14603 14368 14648 14396
rect 14642 14356 14648 14368
rect 14700 14356 14706 14408
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14396 15439 14399
rect 15930 14396 15936 14408
rect 15427 14368 15936 14396
rect 15427 14365 15439 14368
rect 15381 14359 15439 14365
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 16025 14399 16083 14405
rect 16025 14365 16037 14399
rect 16071 14396 16083 14399
rect 16758 14396 16764 14408
rect 16071 14368 16764 14396
rect 16071 14365 16083 14368
rect 16025 14359 16083 14365
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 16942 14396 16948 14408
rect 16903 14368 16948 14396
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 17129 14399 17187 14405
rect 17129 14365 17141 14399
rect 17175 14365 17187 14399
rect 17310 14396 17316 14408
rect 17271 14368 17316 14396
rect 17129 14359 17187 14365
rect 15102 14328 15108 14340
rect 13280 14300 15108 14328
rect 15102 14288 15108 14300
rect 15160 14288 15166 14340
rect 16301 14331 16359 14337
rect 16301 14297 16313 14331
rect 16347 14328 16359 14331
rect 17144 14328 17172 14359
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 17494 14396 17500 14408
rect 17455 14368 17500 14396
rect 17494 14356 17500 14368
rect 17552 14356 17558 14408
rect 17862 14356 17868 14408
rect 17920 14356 17926 14408
rect 18046 14356 18052 14408
rect 18104 14396 18110 14408
rect 18322 14396 18328 14408
rect 18104 14368 18149 14396
rect 18283 14368 18328 14396
rect 18104 14356 18110 14368
rect 18322 14356 18328 14368
rect 18380 14356 18386 14408
rect 18432 14405 18460 14436
rect 18984 14436 20024 14464
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14396 18475 14399
rect 18598 14396 18604 14408
rect 18463 14368 18604 14396
rect 18463 14365 18475 14368
rect 18417 14359 18475 14365
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 17880 14328 17908 14356
rect 18984 14328 19012 14436
rect 19996 14405 20024 14436
rect 20622 14424 20628 14476
rect 20680 14464 20686 14476
rect 30024 14473 30052 14504
rect 30098 14492 30104 14504
rect 30156 14492 30162 14544
rect 30009 14467 30067 14473
rect 20680 14436 22324 14464
rect 20680 14424 20686 14436
rect 19705 14399 19763 14405
rect 19705 14365 19717 14399
rect 19751 14365 19763 14399
rect 19705 14359 19763 14365
rect 19981 14399 20039 14405
rect 19981 14365 19993 14399
rect 20027 14365 20039 14399
rect 19981 14359 20039 14365
rect 20073 14399 20131 14405
rect 20073 14365 20085 14399
rect 20119 14396 20131 14399
rect 20530 14396 20536 14408
rect 20119 14368 20536 14396
rect 20119 14365 20131 14368
rect 20073 14359 20131 14365
rect 16347 14300 17908 14328
rect 18432 14300 19012 14328
rect 19720 14328 19748 14359
rect 20530 14356 20536 14368
rect 20588 14356 20594 14408
rect 20714 14396 20720 14408
rect 20675 14368 20720 14396
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 22296 14405 22324 14436
rect 30009 14433 30021 14467
rect 30055 14433 30067 14467
rect 30009 14427 30067 14433
rect 20993 14399 21051 14405
rect 20993 14365 21005 14399
rect 21039 14396 21051 14399
rect 22005 14399 22063 14405
rect 22005 14396 22017 14399
rect 21039 14368 22017 14396
rect 21039 14365 21051 14368
rect 20993 14359 21051 14365
rect 22005 14365 22017 14368
rect 22051 14365 22063 14399
rect 22005 14359 22063 14365
rect 22281 14399 22339 14405
rect 22281 14365 22293 14399
rect 22327 14365 22339 14399
rect 22281 14359 22339 14365
rect 20254 14328 20260 14340
rect 19720 14300 20260 14328
rect 16347 14297 16359 14300
rect 16301 14291 16359 14297
rect 8343 14232 9352 14260
rect 8343 14229 8355 14232
rect 8297 14223 8355 14229
rect 12710 14220 12716 14272
rect 12768 14260 12774 14272
rect 13173 14263 13231 14269
rect 13173 14260 13185 14263
rect 12768 14232 13185 14260
rect 12768 14220 12774 14232
rect 13173 14229 13185 14232
rect 13219 14229 13231 14263
rect 13173 14223 13231 14229
rect 15289 14263 15347 14269
rect 15289 14229 15301 14263
rect 15335 14260 15347 14263
rect 15470 14260 15476 14272
rect 15335 14232 15476 14260
rect 15335 14229 15347 14232
rect 15289 14223 15347 14229
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 15838 14260 15844 14272
rect 15799 14232 15844 14260
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 16206 14220 16212 14272
rect 16264 14260 16270 14272
rect 16316 14260 16344 14291
rect 17310 14260 17316 14272
rect 16264 14232 16344 14260
rect 17271 14232 17316 14260
rect 16264 14220 16270 14232
rect 17310 14220 17316 14232
rect 17368 14220 17374 14272
rect 17862 14220 17868 14272
rect 17920 14260 17926 14272
rect 18432 14260 18460 14300
rect 20254 14288 20260 14300
rect 20312 14328 20318 14340
rect 21008 14328 21036 14359
rect 22370 14356 22376 14408
rect 22428 14396 22434 14408
rect 28813 14399 28871 14405
rect 22428 14368 22473 14396
rect 22428 14356 22434 14368
rect 28813 14365 28825 14399
rect 28859 14396 28871 14399
rect 29914 14396 29920 14408
rect 28859 14368 29500 14396
rect 29875 14368 29920 14396
rect 28859 14365 28871 14368
rect 28813 14359 28871 14365
rect 20312 14300 21036 14328
rect 22557 14331 22615 14337
rect 20312 14288 20318 14300
rect 22557 14297 22569 14331
rect 22603 14328 22615 14331
rect 29178 14328 29184 14340
rect 22603 14300 29184 14328
rect 22603 14297 22615 14300
rect 22557 14291 22615 14297
rect 29178 14288 29184 14300
rect 29236 14288 29242 14340
rect 29472 14328 29500 14368
rect 29914 14356 29920 14368
rect 29972 14356 29978 14408
rect 30101 14399 30159 14405
rect 30101 14365 30113 14399
rect 30147 14396 30159 14399
rect 30282 14396 30288 14408
rect 30147 14368 30288 14396
rect 30147 14365 30159 14368
rect 30101 14359 30159 14365
rect 30116 14328 30144 14359
rect 30282 14356 30288 14368
rect 30340 14356 30346 14408
rect 29472 14300 30144 14328
rect 18598 14260 18604 14272
rect 17920 14232 18460 14260
rect 18559 14232 18604 14260
rect 17920 14220 17926 14232
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 22462 14220 22468 14272
rect 22520 14260 22526 14272
rect 28074 14260 28080 14272
rect 22520 14232 28080 14260
rect 22520 14220 22526 14232
rect 28074 14220 28080 14232
rect 28132 14220 28138 14272
rect 1104 14170 30820 14192
rect 1104 14118 10880 14170
rect 10932 14118 10944 14170
rect 10996 14118 11008 14170
rect 11060 14118 11072 14170
rect 11124 14118 11136 14170
rect 11188 14118 20811 14170
rect 20863 14118 20875 14170
rect 20927 14118 20939 14170
rect 20991 14118 21003 14170
rect 21055 14118 21067 14170
rect 21119 14118 30820 14170
rect 1104 14096 30820 14118
rect 1394 14056 1400 14068
rect 1355 14028 1400 14056
rect 1394 14016 1400 14028
rect 1452 14016 1458 14068
rect 4614 14056 4620 14068
rect 4575 14028 4620 14056
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 7558 14056 7564 14068
rect 7519 14028 7564 14056
rect 7558 14016 7564 14028
rect 7616 14016 7622 14068
rect 8018 14016 8024 14068
rect 8076 14016 8082 14068
rect 8312 14028 9251 14056
rect 3142 13988 3148 14000
rect 1596 13960 3148 13988
rect 1596 13929 1624 13960
rect 3142 13948 3148 13960
rect 3200 13948 3206 14000
rect 3786 13948 3792 14000
rect 3844 13988 3850 14000
rect 8036 13988 8064 14016
rect 8312 13997 8340 14028
rect 8297 13991 8355 13997
rect 3844 13960 4476 13988
rect 8036 13960 8156 13988
rect 3844 13948 3850 13960
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13889 1639 13923
rect 1946 13920 1952 13932
rect 1907 13892 1952 13920
rect 1581 13883 1639 13889
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 3881 13923 3939 13929
rect 2179 13892 2774 13920
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 1670 13812 1676 13864
rect 1728 13852 1734 13864
rect 1765 13855 1823 13861
rect 1765 13852 1777 13855
rect 1728 13824 1777 13852
rect 1728 13812 1734 13824
rect 1765 13821 1777 13824
rect 1811 13821 1823 13855
rect 1765 13815 1823 13821
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13821 1915 13855
rect 1857 13815 1915 13821
rect 1872 13784 1900 13815
rect 2406 13812 2412 13864
rect 2464 13852 2470 13864
rect 2593 13855 2651 13861
rect 2593 13852 2605 13855
rect 2464 13824 2605 13852
rect 2464 13812 2470 13824
rect 2593 13821 2605 13824
rect 2639 13821 2651 13855
rect 2746 13852 2774 13892
rect 3881 13889 3893 13923
rect 3927 13889 3939 13923
rect 4062 13920 4068 13932
rect 4023 13892 4068 13920
rect 3881 13883 3939 13889
rect 2869 13855 2927 13861
rect 2869 13852 2881 13855
rect 2746 13824 2881 13852
rect 2593 13815 2651 13821
rect 2869 13821 2881 13824
rect 2915 13852 2927 13855
rect 3326 13852 3332 13864
rect 2915 13824 3332 13852
rect 2915 13821 2927 13824
rect 2869 13815 2927 13821
rect 3326 13812 3332 13824
rect 3384 13852 3390 13864
rect 3896 13852 3924 13883
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4246 13920 4252 13932
rect 4207 13892 4252 13920
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 4448 13929 4476 13960
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13889 4491 13923
rect 4433 13883 4491 13889
rect 5169 13923 5227 13929
rect 5169 13889 5181 13923
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 4154 13852 4160 13864
rect 3384 13824 3924 13852
rect 4115 13824 4160 13852
rect 3384 13812 3390 13824
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 5184 13852 5212 13883
rect 6730 13880 6736 13932
rect 6788 13920 6794 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6788 13892 6837 13920
rect 6788 13880 6794 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 7006 13920 7012 13932
rect 6967 13892 7012 13920
rect 6825 13883 6883 13889
rect 7006 13880 7012 13892
rect 7064 13880 7070 13932
rect 7098 13880 7104 13932
rect 7156 13920 7162 13932
rect 7374 13920 7380 13932
rect 7156 13892 7201 13920
rect 7335 13892 7380 13920
rect 7156 13880 7162 13892
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 8128 13929 8156 13960
rect 8297 13957 8309 13991
rect 8343 13957 8355 13991
rect 9122 13988 9128 14000
rect 9083 13960 9128 13988
rect 8297 13951 8355 13957
rect 9122 13948 9128 13960
rect 9180 13948 9186 14000
rect 9223 13988 9251 14028
rect 9582 14016 9588 14068
rect 9640 14056 9646 14068
rect 17770 14056 17776 14068
rect 9640 14028 17776 14056
rect 9640 14016 9646 14028
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 18598 14016 18604 14068
rect 18656 14056 18662 14068
rect 22462 14056 22468 14068
rect 18656 14028 22468 14056
rect 18656 14016 18662 14028
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 30009 14059 30067 14065
rect 30009 14025 30021 14059
rect 30055 14056 30067 14059
rect 30190 14056 30196 14068
rect 30055 14028 30196 14056
rect 30055 14025 30067 14028
rect 30009 14019 30067 14025
rect 30190 14016 30196 14028
rect 30248 14016 30254 14068
rect 9950 13988 9956 14000
rect 9223 13960 9956 13988
rect 9950 13948 9956 13960
rect 10008 13948 10014 14000
rect 14737 13991 14795 13997
rect 10060 13960 14688 13988
rect 8021 13923 8079 13929
rect 8021 13889 8033 13923
rect 8067 13889 8079 13923
rect 8128 13923 8199 13929
rect 8128 13894 8153 13923
rect 8137 13892 8153 13894
rect 8021 13883 8079 13889
rect 8141 13889 8153 13892
rect 8187 13889 8199 13923
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 8141 13883 8199 13889
rect 8312 13892 8401 13920
rect 4264 13824 5212 13852
rect 5261 13855 5319 13861
rect 1872 13756 2636 13784
rect 2608 13728 2636 13756
rect 2958 13744 2964 13796
rect 3016 13784 3022 13796
rect 4264 13784 4292 13824
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 6362 13852 6368 13864
rect 5307 13824 6368 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 6362 13812 6368 13824
rect 6420 13812 6426 13864
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 6972 13824 7205 13852
rect 6972 13812 6978 13824
rect 7193 13821 7205 13824
rect 7239 13821 7251 13855
rect 7193 13815 7251 13821
rect 7558 13812 7564 13864
rect 7616 13852 7622 13864
rect 7926 13852 7932 13864
rect 7616 13824 7932 13852
rect 7616 13812 7622 13824
rect 7926 13812 7932 13824
rect 7984 13852 7990 13864
rect 8045 13852 8073 13883
rect 7984 13824 8073 13852
rect 7984 13812 7990 13824
rect 3016 13756 4292 13784
rect 3016 13744 3022 13756
rect 2590 13676 2596 13728
rect 2648 13676 2654 13728
rect 8312 13716 8340 13892
rect 8389 13889 8401 13892
rect 8435 13889 8447 13923
rect 8389 13883 8447 13889
rect 8486 13923 8544 13929
rect 8486 13889 8498 13923
rect 8532 13922 8544 13923
rect 8532 13920 8616 13922
rect 8846 13920 8852 13932
rect 8532 13894 8852 13920
rect 8532 13889 8544 13894
rect 8588 13892 8852 13894
rect 8486 13883 8544 13889
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9306 13920 9312 13932
rect 9267 13892 9312 13920
rect 9306 13880 9312 13892
rect 9364 13880 9370 13932
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13920 9551 13923
rect 9582 13920 9588 13932
rect 9539 13892 9588 13920
rect 9539 13889 9551 13892
rect 9493 13883 9551 13889
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 10060 13920 10088 13960
rect 9732 13892 10088 13920
rect 10229 13923 10287 13929
rect 9732 13880 9738 13892
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10778 13920 10784 13932
rect 10275 13892 10784 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 9766 13812 9772 13864
rect 9824 13852 9830 13864
rect 10244 13852 10272 13883
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13920 12679 13923
rect 13262 13920 13268 13932
rect 12667 13892 13268 13920
rect 12667 13889 12679 13892
rect 12621 13883 12679 13889
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 13354 13880 13360 13932
rect 13412 13920 13418 13932
rect 13722 13920 13728 13932
rect 13412 13892 13457 13920
rect 13683 13892 13728 13920
rect 13412 13880 13418 13892
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 14550 13920 14556 13932
rect 14511 13892 14556 13920
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 14660 13920 14688 13960
rect 14737 13957 14749 13991
rect 14783 13988 14795 13991
rect 15378 13988 15384 14000
rect 14783 13960 15384 13988
rect 14783 13957 14795 13960
rect 14737 13951 14795 13957
rect 15378 13948 15384 13960
rect 15436 13988 15442 14000
rect 15838 13988 15844 14000
rect 15436 13960 15844 13988
rect 15436 13948 15442 13960
rect 15838 13948 15844 13960
rect 15896 13948 15902 14000
rect 19150 13988 19156 14000
rect 15948 13960 19156 13988
rect 15562 13920 15568 13932
rect 14660 13892 14780 13920
rect 15523 13892 15568 13920
rect 9824 13824 10272 13852
rect 9824 13812 9830 13824
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 14369 13855 14427 13861
rect 12492 13824 12537 13852
rect 12492 13812 12498 13824
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 14642 13852 14648 13864
rect 14415 13824 14648 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 14752 13852 14780 13892
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 15948 13852 15976 13960
rect 19150 13948 19156 13960
rect 19208 13948 19214 14000
rect 19334 13948 19340 14000
rect 19392 13988 19398 14000
rect 22370 13988 22376 14000
rect 19392 13960 19840 13988
rect 19392 13948 19398 13960
rect 16022 13880 16028 13932
rect 16080 13920 16086 13932
rect 16761 13923 16819 13929
rect 16761 13920 16773 13923
rect 16080 13892 16773 13920
rect 16080 13880 16086 13892
rect 16761 13889 16773 13892
rect 16807 13889 16819 13923
rect 16942 13920 16948 13932
rect 16903 13892 16948 13920
rect 16761 13883 16819 13889
rect 14752 13824 15976 13852
rect 16776 13852 16804 13883
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 17494 13920 17500 13932
rect 17455 13892 17500 13920
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 17954 13880 17960 13932
rect 18012 13920 18018 13932
rect 18782 13920 18788 13932
rect 18012 13892 18788 13920
rect 18012 13880 18018 13892
rect 18782 13880 18788 13892
rect 18840 13880 18846 13932
rect 19518 13880 19524 13932
rect 19576 13929 19582 13932
rect 19812 13929 19840 13960
rect 20732 13960 22376 13988
rect 19576 13920 19588 13929
rect 19797 13923 19855 13929
rect 19576 13892 19621 13920
rect 19576 13883 19588 13892
rect 19797 13889 19809 13923
rect 19843 13889 19855 13923
rect 19797 13883 19855 13889
rect 19576 13880 19582 13883
rect 20530 13880 20536 13932
rect 20588 13920 20594 13932
rect 20732 13929 20760 13960
rect 22370 13948 22376 13960
rect 22428 13948 22434 14000
rect 20717 13923 20775 13929
rect 20717 13920 20729 13923
rect 20588 13892 20729 13920
rect 20588 13880 20594 13892
rect 20717 13889 20729 13892
rect 20763 13889 20775 13923
rect 22278 13920 22284 13932
rect 22239 13892 22284 13920
rect 20717 13883 20775 13889
rect 22278 13880 22284 13892
rect 22336 13880 22342 13932
rect 28074 13880 28080 13932
rect 28132 13920 28138 13932
rect 29917 13923 29975 13929
rect 29917 13920 29929 13923
rect 28132 13892 29929 13920
rect 28132 13880 28138 13892
rect 29917 13889 29929 13892
rect 29963 13889 29975 13923
rect 29917 13883 29975 13889
rect 30101 13923 30159 13929
rect 30101 13889 30113 13923
rect 30147 13920 30159 13923
rect 30282 13920 30288 13932
rect 30147 13892 30288 13920
rect 30147 13889 30159 13892
rect 30101 13883 30159 13889
rect 30282 13880 30288 13892
rect 30340 13880 30346 13932
rect 17678 13852 17684 13864
rect 16776 13824 17684 13852
rect 17678 13812 17684 13824
rect 17736 13852 17742 13864
rect 17736 13824 18460 13852
rect 17736 13812 17742 13824
rect 8662 13784 8668 13796
rect 8623 13756 8668 13784
rect 8662 13744 8668 13756
rect 8720 13744 8726 13796
rect 8846 13744 8852 13796
rect 8904 13784 8910 13796
rect 18432 13793 18460 13824
rect 19978 13812 19984 13864
rect 20036 13852 20042 13864
rect 20441 13855 20499 13861
rect 20441 13852 20453 13855
rect 20036 13824 20453 13852
rect 20036 13812 20042 13824
rect 20441 13821 20453 13824
rect 20487 13852 20499 13855
rect 21542 13852 21548 13864
rect 20487 13824 21548 13852
rect 20487 13821 20499 13824
rect 20441 13815 20499 13821
rect 21542 13812 21548 13824
rect 21600 13812 21606 13864
rect 22557 13855 22615 13861
rect 22557 13821 22569 13855
rect 22603 13852 22615 13855
rect 29638 13852 29644 13864
rect 22603 13824 29644 13852
rect 22603 13821 22615 13824
rect 22557 13815 22615 13821
rect 29638 13812 29644 13824
rect 29696 13812 29702 13864
rect 16669 13787 16727 13793
rect 16669 13784 16681 13787
rect 8904 13756 16681 13784
rect 8904 13744 8910 13756
rect 16669 13753 16681 13756
rect 16715 13753 16727 13787
rect 16669 13747 16727 13753
rect 18417 13787 18475 13793
rect 18417 13753 18429 13787
rect 18463 13753 18475 13787
rect 18417 13747 18475 13753
rect 8570 13716 8576 13728
rect 8312 13688 8576 13716
rect 8570 13676 8576 13688
rect 8628 13676 8634 13728
rect 9122 13676 9128 13728
rect 9180 13716 9186 13728
rect 9306 13716 9312 13728
rect 9180 13688 9312 13716
rect 9180 13676 9186 13688
rect 9306 13676 9312 13688
rect 9364 13676 9370 13728
rect 9674 13676 9680 13728
rect 9732 13716 9738 13728
rect 10134 13716 10140 13728
rect 9732 13688 10140 13716
rect 9732 13676 9738 13688
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 10318 13676 10324 13728
rect 10376 13716 10382 13728
rect 10413 13719 10471 13725
rect 10413 13716 10425 13719
rect 10376 13688 10425 13716
rect 10376 13676 10382 13688
rect 10413 13685 10425 13688
rect 10459 13685 10471 13719
rect 10413 13679 10471 13685
rect 14550 13676 14556 13728
rect 14608 13716 14614 13728
rect 15286 13716 15292 13728
rect 14608 13688 15292 13716
rect 14608 13676 14614 13688
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 18322 13676 18328 13728
rect 18380 13716 18386 13728
rect 21818 13716 21824 13728
rect 18380 13688 21824 13716
rect 18380 13676 18386 13688
rect 21818 13676 21824 13688
rect 21876 13676 21882 13728
rect 1104 13626 30820 13648
rect 1104 13574 5915 13626
rect 5967 13574 5979 13626
rect 6031 13574 6043 13626
rect 6095 13574 6107 13626
rect 6159 13574 6171 13626
rect 6223 13574 15846 13626
rect 15898 13574 15910 13626
rect 15962 13574 15974 13626
rect 16026 13574 16038 13626
rect 16090 13574 16102 13626
rect 16154 13574 25776 13626
rect 25828 13574 25840 13626
rect 25892 13574 25904 13626
rect 25956 13574 25968 13626
rect 26020 13574 26032 13626
rect 26084 13574 30820 13626
rect 1104 13552 30820 13574
rect 4246 13512 4252 13524
rect 4207 13484 4252 13512
rect 4246 13472 4252 13484
rect 4304 13472 4310 13524
rect 4706 13472 4712 13524
rect 4764 13512 4770 13524
rect 4985 13515 5043 13521
rect 4985 13512 4997 13515
rect 4764 13484 4997 13512
rect 4764 13472 4770 13484
rect 4985 13481 4997 13484
rect 5031 13512 5043 13515
rect 5442 13512 5448 13524
rect 5031 13484 5448 13512
rect 5031 13481 5043 13484
rect 4985 13475 5043 13481
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 6549 13515 6607 13521
rect 6549 13481 6561 13515
rect 6595 13512 6607 13515
rect 6595 13484 11744 13512
rect 6595 13481 6607 13484
rect 6549 13475 6607 13481
rect 1857 13447 1915 13453
rect 1857 13413 1869 13447
rect 1903 13444 1915 13447
rect 7006 13444 7012 13456
rect 1903 13416 7012 13444
rect 1903 13413 1915 13416
rect 1857 13407 1915 13413
rect 7006 13404 7012 13416
rect 7064 13404 7070 13456
rect 8478 13404 8484 13456
rect 8536 13444 8542 13456
rect 9122 13444 9128 13456
rect 8536 13416 9128 13444
rect 8536 13404 8542 13416
rect 9122 13404 9128 13416
rect 9180 13404 9186 13456
rect 11609 13447 11667 13453
rect 11609 13413 11621 13447
rect 11655 13413 11667 13447
rect 11716 13444 11744 13484
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11848 13484 12081 13512
rect 11848 13472 11854 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 16209 13515 16267 13521
rect 16209 13512 16221 13515
rect 15344 13484 16221 13512
rect 15344 13472 15350 13484
rect 16209 13481 16221 13484
rect 16255 13481 16267 13515
rect 16209 13475 16267 13481
rect 17405 13515 17463 13521
rect 17405 13481 17417 13515
rect 17451 13512 17463 13515
rect 18046 13512 18052 13524
rect 17451 13484 18052 13512
rect 17451 13481 17463 13484
rect 17405 13475 17463 13481
rect 18046 13472 18052 13484
rect 18104 13512 18110 13524
rect 19337 13515 19395 13521
rect 19337 13512 19349 13515
rect 18104 13484 19349 13512
rect 18104 13472 18110 13484
rect 19337 13481 19349 13484
rect 19383 13481 19395 13515
rect 19337 13475 19395 13481
rect 20346 13472 20352 13524
rect 20404 13512 20410 13524
rect 20404 13484 20576 13512
rect 20404 13472 20410 13484
rect 20548 13456 20576 13484
rect 19886 13444 19892 13456
rect 11716 13416 19892 13444
rect 11609 13407 11667 13413
rect 3786 13376 3792 13388
rect 1964 13348 3792 13376
rect 1964 13317 1992 13348
rect 3786 13336 3792 13348
rect 3844 13336 3850 13388
rect 5626 13336 5632 13388
rect 5684 13376 5690 13388
rect 6181 13379 6239 13385
rect 5684 13348 6040 13376
rect 5684 13336 5690 13348
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13277 2007 13311
rect 1949 13271 2007 13277
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13277 2467 13311
rect 2409 13271 2467 13277
rect 2424 13172 2452 13271
rect 2590 13268 2596 13320
rect 2648 13308 2654 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2648 13280 2697 13308
rect 2648 13268 2654 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4764 13280 4905 13308
rect 4764 13268 4770 13280
rect 4893 13277 4905 13280
rect 4939 13308 4951 13311
rect 5074 13308 5080 13320
rect 4939 13280 5080 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 6012 13317 6040 13348
rect 6181 13345 6193 13379
rect 6227 13376 6239 13379
rect 8389 13379 8447 13385
rect 6227 13348 8340 13376
rect 6227 13345 6239 13348
rect 6181 13339 6239 13345
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 5997 13311 6055 13317
rect 5997 13277 6009 13311
rect 6043 13277 6055 13311
rect 5997 13271 6055 13277
rect 6092 13311 6150 13317
rect 6092 13277 6104 13311
rect 6138 13277 6150 13311
rect 6092 13271 6150 13277
rect 4341 13243 4399 13249
rect 4341 13209 4353 13243
rect 4387 13240 4399 13243
rect 4798 13240 4804 13252
rect 4387 13212 4804 13240
rect 4387 13209 4399 13212
rect 4341 13203 4399 13209
rect 4798 13200 4804 13212
rect 4856 13200 4862 13252
rect 5828 13240 5856 13271
rect 5902 13240 5908 13252
rect 5828 13212 5908 13240
rect 5902 13200 5908 13212
rect 5960 13200 5966 13252
rect 6104 13184 6132 13271
rect 4522 13172 4528 13184
rect 2424 13144 4528 13172
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 6086 13132 6092 13184
rect 6144 13132 6150 13184
rect 6196 13172 6224 13339
rect 6362 13308 6368 13320
rect 6323 13280 6368 13308
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 8110 13308 8116 13320
rect 8071 13280 8116 13308
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 8312 13308 8340 13348
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 11624 13376 11652 13407
rect 19886 13404 19892 13416
rect 19944 13404 19950 13456
rect 20530 13404 20536 13456
rect 20588 13404 20594 13456
rect 12437 13379 12495 13385
rect 12437 13376 12449 13379
rect 8435 13348 10364 13376
rect 11624 13348 12449 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 8312 13280 9720 13308
rect 7374 13200 7380 13252
rect 7432 13240 7438 13252
rect 8754 13240 8760 13252
rect 7432 13212 8760 13240
rect 7432 13200 7438 13212
rect 8754 13200 8760 13212
rect 8812 13200 8818 13252
rect 9401 13243 9459 13249
rect 9401 13209 9413 13243
rect 9447 13240 9459 13243
rect 9582 13240 9588 13252
rect 9447 13212 9588 13240
rect 9447 13209 9459 13212
rect 9401 13203 9459 13209
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 6270 13172 6276 13184
rect 6196 13144 6276 13172
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 8846 13172 8852 13184
rect 6880 13144 8852 13172
rect 6880 13132 6886 13144
rect 8846 13132 8852 13144
rect 8904 13132 8910 13184
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 9493 13175 9551 13181
rect 9493 13172 9505 13175
rect 8996 13144 9505 13172
rect 8996 13132 9002 13144
rect 9493 13141 9505 13144
rect 9539 13141 9551 13175
rect 9692 13172 9720 13280
rect 10042 13268 10048 13320
rect 10100 13308 10106 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 10100 13280 10241 13308
rect 10100 13268 10106 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 10336 13308 10364 13348
rect 12437 13345 12449 13348
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 15746 13376 15752 13388
rect 15344 13348 15752 13376
rect 15344 13336 15350 13348
rect 15746 13336 15752 13348
rect 15804 13376 15810 13388
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 15804 13348 16313 13376
rect 15804 13336 15810 13348
rect 16301 13345 16313 13348
rect 16347 13345 16359 13379
rect 16301 13339 16359 13345
rect 17218 13336 17224 13388
rect 17276 13376 17282 13388
rect 17589 13379 17647 13385
rect 17589 13376 17601 13379
rect 17276 13348 17601 13376
rect 17276 13336 17282 13348
rect 17589 13345 17601 13348
rect 17635 13345 17647 13379
rect 17589 13339 17647 13345
rect 17678 13336 17684 13388
rect 17736 13376 17742 13388
rect 18230 13376 18236 13388
rect 17736 13348 18236 13376
rect 17736 13336 17742 13348
rect 12253 13311 12311 13317
rect 10336 13280 11560 13308
rect 10229 13271 10287 13277
rect 10496 13243 10554 13249
rect 10496 13209 10508 13243
rect 10542 13240 10554 13243
rect 11422 13240 11428 13252
rect 10542 13212 11428 13240
rect 10542 13209 10554 13212
rect 10496 13203 10554 13209
rect 11422 13200 11428 13212
rect 11480 13200 11486 13252
rect 11532 13240 11560 13280
rect 12253 13277 12265 13311
rect 12299 13308 12311 13311
rect 12342 13308 12348 13320
rect 12299 13280 12348 13308
rect 12299 13277 12311 13280
rect 12253 13271 12311 13277
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 13354 13308 13360 13320
rect 12676 13280 13360 13308
rect 12676 13268 12682 13280
rect 13354 13268 13360 13280
rect 13412 13308 13418 13320
rect 13449 13311 13507 13317
rect 13449 13308 13461 13311
rect 13412 13280 13461 13308
rect 13412 13268 13418 13280
rect 13449 13277 13461 13280
rect 13495 13277 13507 13311
rect 13449 13271 13507 13277
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13308 13599 13311
rect 14274 13308 14280 13320
rect 13587 13280 14280 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 15378 13308 15384 13320
rect 15339 13280 15384 13308
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 15562 13308 15568 13320
rect 15488 13280 15568 13308
rect 14461 13243 14519 13249
rect 14461 13240 14473 13243
rect 11532 13212 14473 13240
rect 14461 13209 14473 13212
rect 14507 13240 14519 13243
rect 15010 13240 15016 13252
rect 14507 13212 15016 13240
rect 14507 13209 14519 13212
rect 14461 13203 14519 13209
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 15197 13243 15255 13249
rect 15197 13209 15209 13243
rect 15243 13240 15255 13243
rect 15488 13240 15516 13280
rect 15562 13268 15568 13280
rect 15620 13268 15626 13320
rect 16206 13308 16212 13320
rect 16167 13280 16212 13308
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 17405 13311 17463 13317
rect 17405 13277 17417 13311
rect 17451 13308 17463 13311
rect 17497 13311 17555 13317
rect 17497 13308 17509 13311
rect 17451 13280 17509 13308
rect 17451 13277 17463 13280
rect 17405 13271 17463 13277
rect 17497 13277 17509 13280
rect 17543 13277 17555 13311
rect 17770 13308 17776 13320
rect 17731 13280 17776 13308
rect 17497 13271 17555 13277
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 17880 13317 17908 13348
rect 18230 13336 18236 13348
rect 18288 13336 18294 13388
rect 19610 13336 19616 13388
rect 19668 13376 19674 13388
rect 20349 13379 20407 13385
rect 20349 13376 20361 13379
rect 19668 13348 20361 13376
rect 19668 13336 19674 13348
rect 20349 13345 20361 13348
rect 20395 13345 20407 13379
rect 20548 13376 20576 13404
rect 20548 13348 20668 13376
rect 20349 13339 20407 13345
rect 17865 13311 17923 13317
rect 17865 13277 17877 13311
rect 17911 13277 17923 13311
rect 19334 13308 19340 13320
rect 17865 13271 17923 13277
rect 17972 13280 19340 13308
rect 17972 13240 18000 13280
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 19521 13311 19579 13317
rect 19521 13277 19533 13311
rect 19567 13308 19579 13311
rect 19978 13308 19984 13320
rect 19567 13280 19984 13308
rect 19567 13277 19579 13280
rect 19521 13271 19579 13277
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 20254 13308 20260 13320
rect 20215 13280 20260 13308
rect 20254 13268 20260 13280
rect 20312 13268 20318 13320
rect 20530 13308 20536 13320
rect 20491 13280 20536 13308
rect 20530 13268 20536 13280
rect 20588 13268 20594 13320
rect 20640 13317 20668 13348
rect 20625 13311 20683 13317
rect 20625 13277 20637 13311
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 29546 13308 29552 13320
rect 20855 13280 29552 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 29546 13268 29552 13280
rect 29604 13268 29610 13320
rect 29822 13308 29828 13320
rect 29783 13280 29828 13308
rect 29822 13268 29828 13280
rect 29880 13268 29886 13320
rect 15243 13212 15516 13240
rect 15580 13212 18000 13240
rect 18049 13243 18107 13249
rect 15243 13209 15255 13212
rect 15197 13203 15255 13209
rect 14369 13175 14427 13181
rect 14369 13172 14381 13175
rect 9692 13144 14381 13172
rect 9493 13135 9551 13141
rect 14369 13141 14381 13144
rect 14415 13172 14427 13175
rect 15580 13172 15608 13212
rect 18049 13209 18061 13243
rect 18095 13240 18107 13243
rect 29914 13240 29920 13252
rect 18095 13212 29920 13240
rect 18095 13209 18107 13212
rect 18049 13203 18107 13209
rect 29914 13200 29920 13212
rect 29972 13200 29978 13252
rect 14415 13144 15608 13172
rect 16577 13175 16635 13181
rect 14415 13141 14427 13144
rect 14369 13135 14427 13141
rect 16577 13141 16589 13175
rect 16623 13172 16635 13175
rect 16942 13172 16948 13184
rect 16623 13144 16948 13172
rect 16623 13141 16635 13144
rect 16577 13135 16635 13141
rect 16942 13132 16948 13144
rect 17000 13172 17006 13184
rect 17678 13172 17684 13184
rect 17000 13144 17684 13172
rect 17000 13132 17006 13144
rect 17678 13132 17684 13144
rect 17736 13132 17742 13184
rect 30006 13172 30012 13184
rect 29967 13144 30012 13172
rect 30006 13132 30012 13144
rect 30064 13132 30070 13184
rect 1104 13082 30820 13104
rect 1104 13030 10880 13082
rect 10932 13030 10944 13082
rect 10996 13030 11008 13082
rect 11060 13030 11072 13082
rect 11124 13030 11136 13082
rect 11188 13030 20811 13082
rect 20863 13030 20875 13082
rect 20927 13030 20939 13082
rect 20991 13030 21003 13082
rect 21055 13030 21067 13082
rect 21119 13030 30820 13082
rect 1104 13008 30820 13030
rect 2869 12971 2927 12977
rect 2869 12937 2881 12971
rect 2915 12968 2927 12971
rect 2958 12968 2964 12980
rect 2915 12940 2964 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 4614 12968 4620 12980
rect 4527 12940 4620 12968
rect 4614 12928 4620 12940
rect 4672 12968 4678 12980
rect 5166 12968 5172 12980
rect 4672 12940 5172 12968
rect 4672 12928 4678 12940
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 5534 12928 5540 12980
rect 5592 12928 5598 12980
rect 5626 12928 5632 12980
rect 5684 12968 5690 12980
rect 7466 12968 7472 12980
rect 5684 12940 7472 12968
rect 5684 12928 5690 12940
rect 7466 12928 7472 12940
rect 7524 12928 7530 12980
rect 9125 12971 9183 12977
rect 9125 12937 9137 12971
rect 9171 12937 9183 12971
rect 9125 12931 9183 12937
rect 4982 12860 4988 12912
rect 5040 12900 5046 12912
rect 5445 12903 5503 12909
rect 5040 12872 5396 12900
rect 5040 12860 5046 12872
rect 1578 12792 1584 12844
rect 1636 12832 1642 12844
rect 1745 12835 1803 12841
rect 1745 12832 1757 12835
rect 1636 12804 1757 12832
rect 1636 12792 1642 12804
rect 1745 12801 1757 12804
rect 1791 12801 1803 12835
rect 3326 12832 3332 12844
rect 3287 12804 3332 12832
rect 1745 12795 1803 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 3510 12832 3516 12844
rect 3471 12804 3516 12832
rect 3510 12792 3516 12804
rect 3568 12792 3574 12844
rect 3881 12835 3939 12841
rect 3881 12801 3893 12835
rect 3927 12832 3939 12835
rect 4522 12832 4528 12844
rect 3927 12804 4528 12832
rect 3927 12801 3939 12804
rect 3881 12795 3939 12801
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12801 4767 12835
rect 5261 12835 5319 12841
rect 5261 12832 5273 12835
rect 4709 12795 4767 12801
rect 5184 12804 5273 12832
rect 1486 12764 1492 12776
rect 1447 12736 1492 12764
rect 1486 12724 1492 12736
rect 1544 12724 1550 12776
rect 2590 12724 2596 12776
rect 2648 12764 2654 12776
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 2648 12736 3617 12764
rect 2648 12724 2654 12736
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 3697 12767 3755 12773
rect 3697 12733 3709 12767
rect 3743 12764 3755 12767
rect 4246 12764 4252 12776
rect 3743 12736 4252 12764
rect 3743 12733 3755 12736
rect 3697 12727 3755 12733
rect 3712 12696 3740 12727
rect 4246 12724 4252 12736
rect 4304 12724 4310 12776
rect 2746 12668 3740 12696
rect 4724 12696 4752 12795
rect 5184 12776 5212 12804
rect 5261 12801 5273 12804
rect 5307 12801 5319 12835
rect 5368 12834 5396 12872
rect 5445 12869 5457 12903
rect 5491 12900 5503 12903
rect 5552 12900 5580 12928
rect 6822 12900 6828 12912
rect 5491 12872 5580 12900
rect 5680 12872 6828 12900
rect 5491 12869 5503 12872
rect 5445 12863 5503 12869
rect 5680 12841 5708 12872
rect 6822 12860 6828 12872
rect 6880 12860 6886 12912
rect 8757 12903 8815 12909
rect 8757 12869 8769 12903
rect 8803 12900 8815 12903
rect 8846 12900 8852 12912
rect 8803 12872 8852 12900
rect 8803 12869 8815 12872
rect 8757 12863 8815 12869
rect 8846 12860 8852 12872
rect 8904 12860 8910 12912
rect 8957 12903 9015 12909
rect 8957 12900 8969 12903
rect 8956 12869 8969 12900
rect 9003 12869 9015 12903
rect 9140 12900 9168 12931
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 11609 12971 11667 12977
rect 11609 12968 11621 12971
rect 11480 12940 11621 12968
rect 11480 12928 11486 12940
rect 11609 12937 11621 12940
rect 11655 12937 11667 12971
rect 12802 12968 12808 12980
rect 12763 12940 12808 12968
rect 11609 12931 11667 12937
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 13722 12968 13728 12980
rect 13188 12940 13728 12968
rect 13188 12900 13216 12940
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 15562 12928 15568 12980
rect 15620 12968 15626 12980
rect 16298 12968 16304 12980
rect 15620 12940 16304 12968
rect 15620 12928 15626 12940
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 17586 12968 17592 12980
rect 16684 12940 17592 12968
rect 9140 12872 11560 12900
rect 8956 12863 9015 12869
rect 5537 12835 5595 12841
rect 5368 12832 5488 12834
rect 5537 12832 5549 12835
rect 5368 12806 5549 12832
rect 5460 12804 5549 12806
rect 5261 12795 5319 12801
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 5665 12835 5723 12841
rect 5665 12801 5677 12835
rect 5711 12801 5723 12835
rect 5665 12795 5723 12801
rect 6086 12792 6092 12844
rect 6144 12832 6150 12844
rect 6362 12832 6368 12844
rect 6144 12804 6368 12832
rect 6144 12792 6150 12804
rect 6362 12792 6368 12804
rect 6420 12832 6426 12844
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 6420 12804 7297 12832
rect 6420 12792 6426 12804
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 8018 12832 8024 12844
rect 7607 12804 8024 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 8018 12792 8024 12804
rect 8076 12832 8082 12844
rect 8113 12835 8171 12841
rect 8113 12832 8125 12835
rect 8076 12804 8125 12832
rect 8076 12792 8082 12804
rect 8113 12801 8125 12804
rect 8159 12801 8171 12835
rect 8956 12832 8984 12863
rect 9766 12832 9772 12844
rect 8956 12804 9772 12832
rect 8113 12795 8171 12801
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 10060 12841 10088 12872
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12801 10103 12835
rect 10778 12832 10784 12844
rect 10739 12804 10784 12832
rect 10045 12795 10103 12801
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 11532 12841 11560 12872
rect 12406 12872 13216 12900
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 5166 12764 5172 12776
rect 5079 12736 5172 12764
rect 5166 12724 5172 12736
rect 5224 12764 5230 12776
rect 5224 12736 9812 12764
rect 5224 12724 5230 12736
rect 5810 12696 5816 12708
rect 4724 12668 5816 12696
rect 1670 12588 1676 12640
rect 1728 12628 1734 12640
rect 2746 12628 2774 12668
rect 5810 12656 5816 12668
rect 5868 12656 5874 12708
rect 5902 12656 5908 12708
rect 5960 12696 5966 12708
rect 7926 12696 7932 12708
rect 5960 12668 7932 12696
rect 5960 12656 5966 12668
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 8294 12696 8300 12708
rect 8255 12668 8300 12696
rect 8294 12656 8300 12668
rect 8352 12656 8358 12708
rect 9677 12699 9735 12705
rect 9677 12696 9689 12699
rect 8404 12668 9689 12696
rect 4062 12628 4068 12640
rect 1728 12600 2774 12628
rect 4023 12600 4068 12628
rect 1728 12588 1734 12600
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 7098 12628 7104 12640
rect 5307 12600 7104 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 7742 12588 7748 12640
rect 7800 12628 7806 12640
rect 8404 12628 8432 12668
rect 9677 12665 9689 12668
rect 9723 12665 9735 12699
rect 9677 12659 9735 12665
rect 8938 12628 8944 12640
rect 7800 12600 8432 12628
rect 8899 12600 8944 12628
rect 7800 12588 7806 12600
rect 8938 12588 8944 12600
rect 8996 12588 9002 12640
rect 9784 12628 9812 12736
rect 10318 12724 10324 12776
rect 10376 12764 10382 12776
rect 11716 12764 11744 12795
rect 10376 12736 11744 12764
rect 10376 12724 10382 12736
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 10965 12699 11023 12705
rect 10965 12696 10977 12699
rect 10836 12668 10977 12696
rect 10836 12656 10842 12668
rect 10965 12665 10977 12668
rect 11011 12665 11023 12699
rect 10965 12659 11023 12665
rect 12406 12628 12434 12872
rect 13262 12860 13268 12912
rect 13320 12900 13326 12912
rect 13449 12903 13507 12909
rect 13449 12900 13461 12903
rect 13320 12872 13461 12900
rect 13320 12860 13326 12872
rect 13449 12869 13461 12872
rect 13495 12900 13507 12903
rect 14737 12903 14795 12909
rect 14737 12900 14749 12903
rect 13495 12872 14749 12900
rect 13495 12869 13507 12872
rect 13449 12863 13507 12869
rect 14737 12869 14749 12872
rect 14783 12869 14795 12903
rect 14737 12863 14795 12869
rect 15657 12903 15715 12909
rect 15657 12869 15669 12903
rect 15703 12900 15715 12903
rect 16390 12900 16396 12912
rect 15703 12872 16396 12900
rect 15703 12869 15715 12872
rect 15657 12863 15715 12869
rect 16390 12860 16396 12872
rect 16448 12860 16454 12912
rect 12621 12835 12679 12841
rect 12621 12801 12633 12835
rect 12667 12832 12679 12835
rect 12710 12832 12716 12844
rect 12667 12804 12716 12832
rect 12667 12801 12679 12804
rect 12621 12795 12679 12801
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 13630 12832 13636 12844
rect 13591 12804 13636 12832
rect 13630 12792 13636 12804
rect 13688 12792 13694 12844
rect 15010 12792 15016 12844
rect 15068 12832 15074 12844
rect 16684 12841 16712 12940
rect 17586 12928 17592 12940
rect 17644 12928 17650 12980
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 19058 12968 19064 12980
rect 18095 12940 19064 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 19058 12928 19064 12940
rect 19116 12968 19122 12980
rect 19116 12940 19196 12968
rect 19116 12928 19122 12940
rect 19168 12909 19196 12940
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19794 12968 19800 12980
rect 19392 12940 19800 12968
rect 19392 12928 19398 12940
rect 19794 12928 19800 12940
rect 19852 12928 19858 12980
rect 29822 12928 29828 12980
rect 29880 12968 29886 12980
rect 30009 12971 30067 12977
rect 30009 12968 30021 12971
rect 29880 12940 30021 12968
rect 29880 12928 29886 12940
rect 30009 12937 30021 12940
rect 30055 12937 30067 12971
rect 30009 12931 30067 12937
rect 17221 12903 17279 12909
rect 17221 12869 17233 12903
rect 17267 12900 17279 12903
rect 19153 12903 19211 12909
rect 17267 12872 19104 12900
rect 17267 12869 17279 12872
rect 17221 12863 17279 12869
rect 15381 12835 15439 12841
rect 15381 12832 15393 12835
rect 15068 12804 15393 12832
rect 15068 12792 15074 12804
rect 15381 12801 15393 12804
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 16669 12835 16727 12841
rect 16669 12801 16681 12835
rect 16715 12801 16727 12835
rect 16942 12832 16948 12844
rect 16903 12804 16948 12832
rect 16669 12795 16727 12801
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 17034 12792 17040 12844
rect 17092 12832 17098 12844
rect 17092 12804 17137 12832
rect 17092 12792 17098 12804
rect 17494 12792 17500 12844
rect 17552 12792 17558 12844
rect 17678 12832 17684 12844
rect 17639 12804 17684 12832
rect 17678 12792 17684 12804
rect 17736 12792 17742 12844
rect 18414 12792 18420 12844
rect 18472 12832 18478 12844
rect 18509 12835 18567 12841
rect 18509 12832 18521 12835
rect 18472 12804 18521 12832
rect 18472 12792 18478 12804
rect 18509 12801 18521 12804
rect 18555 12801 18567 12835
rect 18509 12795 18567 12801
rect 18598 12792 18604 12844
rect 18656 12832 18662 12844
rect 19076 12832 19104 12872
rect 19153 12869 19165 12903
rect 19199 12869 19211 12903
rect 28994 12900 29000 12912
rect 19153 12863 19211 12869
rect 19260 12872 29000 12900
rect 19260 12832 19288 12872
rect 28994 12860 29000 12872
rect 29052 12860 29058 12912
rect 18656 12804 18701 12832
rect 19076 12804 19288 12832
rect 19337 12835 19395 12841
rect 18656 12792 18662 12804
rect 19337 12801 19349 12835
rect 19383 12801 19395 12835
rect 19337 12795 19395 12801
rect 19981 12835 20039 12841
rect 19981 12801 19993 12835
rect 20027 12832 20039 12835
rect 20162 12832 20168 12844
rect 20027 12804 20168 12832
rect 20027 12801 20039 12804
rect 19981 12795 20039 12801
rect 17512 12764 17540 12792
rect 17773 12767 17831 12773
rect 17773 12764 17785 12767
rect 17512 12736 17785 12764
rect 17773 12733 17785 12736
rect 17819 12733 17831 12767
rect 18616 12764 18644 12792
rect 19352 12764 19380 12795
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 20257 12835 20315 12841
rect 20257 12801 20269 12835
rect 20303 12801 20315 12835
rect 20257 12795 20315 12801
rect 18616 12736 19380 12764
rect 17773 12727 17831 12733
rect 19886 12724 19892 12776
rect 19944 12764 19950 12776
rect 20073 12767 20131 12773
rect 20073 12764 20085 12767
rect 19944 12736 20085 12764
rect 19944 12724 19950 12736
rect 20073 12733 20085 12736
rect 20119 12733 20131 12767
rect 20073 12727 20131 12733
rect 17494 12656 17500 12708
rect 17552 12696 17558 12708
rect 20272 12696 20300 12795
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 29917 12835 29975 12841
rect 29917 12832 29929 12835
rect 20404 12804 20449 12832
rect 26206 12804 29929 12832
rect 20404 12792 20410 12804
rect 17552 12668 20300 12696
rect 20533 12699 20591 12705
rect 17552 12656 17558 12668
rect 20533 12665 20545 12699
rect 20579 12696 20591 12699
rect 26206 12696 26234 12804
rect 29917 12801 29929 12804
rect 29963 12801 29975 12835
rect 29917 12795 29975 12801
rect 30101 12835 30159 12841
rect 30101 12801 30113 12835
rect 30147 12832 30159 12835
rect 30282 12832 30288 12844
rect 30147 12804 30288 12832
rect 30147 12801 30159 12804
rect 30101 12795 30159 12801
rect 30282 12792 30288 12804
rect 30340 12792 30346 12844
rect 20579 12668 26234 12696
rect 20579 12665 20591 12668
rect 20533 12659 20591 12665
rect 9784 12600 12434 12628
rect 14458 12588 14464 12640
rect 14516 12628 14522 12640
rect 14829 12631 14887 12637
rect 14829 12628 14841 12631
rect 14516 12600 14841 12628
rect 14516 12588 14522 12600
rect 14829 12597 14841 12600
rect 14875 12597 14887 12631
rect 16758 12628 16764 12640
rect 16719 12600 16764 12628
rect 14829 12591 14887 12597
rect 16758 12588 16764 12600
rect 16816 12588 16822 12640
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 17681 12631 17739 12637
rect 17681 12628 17693 12631
rect 17460 12600 17693 12628
rect 17460 12588 17466 12600
rect 17681 12597 17693 12600
rect 17727 12597 17739 12631
rect 19518 12628 19524 12640
rect 19479 12600 19524 12628
rect 17681 12591 17739 12597
rect 19518 12588 19524 12600
rect 19576 12588 19582 12640
rect 1104 12538 30820 12560
rect 1104 12486 5915 12538
rect 5967 12486 5979 12538
rect 6031 12486 6043 12538
rect 6095 12486 6107 12538
rect 6159 12486 6171 12538
rect 6223 12486 15846 12538
rect 15898 12486 15910 12538
rect 15962 12486 15974 12538
rect 16026 12486 16038 12538
rect 16090 12486 16102 12538
rect 16154 12486 25776 12538
rect 25828 12486 25840 12538
rect 25892 12486 25904 12538
rect 25956 12486 25968 12538
rect 26020 12486 26032 12538
rect 26084 12486 30820 12538
rect 1104 12464 30820 12486
rect 1578 12424 1584 12436
rect 1539 12396 1584 12424
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 6546 12384 6552 12436
rect 6604 12384 6610 12436
rect 6641 12427 6699 12433
rect 6641 12393 6653 12427
rect 6687 12424 6699 12427
rect 14274 12424 14280 12436
rect 6687 12396 14044 12424
rect 6687 12393 6699 12396
rect 6641 12387 6699 12393
rect 1854 12316 1860 12368
rect 1912 12356 1918 12368
rect 2958 12356 2964 12368
rect 1912 12328 2176 12356
rect 1912 12316 1918 12328
rect 1670 12248 1676 12300
rect 1728 12288 1734 12300
rect 1949 12291 2007 12297
rect 1949 12288 1961 12291
rect 1728 12260 1961 12288
rect 1728 12248 1734 12260
rect 1949 12257 1961 12260
rect 1995 12257 2007 12291
rect 1949 12251 2007 12257
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12189 1823 12223
rect 2038 12220 2044 12232
rect 1999 12192 2044 12220
rect 1765 12183 1823 12189
rect 1780 12152 1808 12183
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 2148 12229 2176 12328
rect 2240 12328 2964 12356
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 2240 12152 2268 12328
rect 2958 12316 2964 12328
rect 3016 12316 3022 12368
rect 6178 12316 6184 12368
rect 6236 12356 6242 12368
rect 6564 12356 6592 12384
rect 8018 12356 8024 12368
rect 6236 12328 6592 12356
rect 7392 12328 8024 12356
rect 6236 12316 6242 12328
rect 2866 12288 2872 12300
rect 2332 12260 2872 12288
rect 2332 12229 2360 12260
rect 2866 12248 2872 12260
rect 2924 12288 2930 12300
rect 3326 12288 3332 12300
rect 2924 12260 3332 12288
rect 2924 12248 2930 12260
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 6270 12288 6276 12300
rect 5776 12260 6132 12288
rect 6231 12260 6276 12288
rect 5776 12248 5782 12260
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12189 2375 12223
rect 2317 12183 2375 12189
rect 2774 12180 2780 12232
rect 2832 12220 2838 12232
rect 3789 12223 3847 12229
rect 2832 12192 2877 12220
rect 2832 12180 2838 12192
rect 3789 12189 3801 12223
rect 3835 12220 3847 12223
rect 4614 12220 4620 12232
rect 3835 12192 4620 12220
rect 3835 12189 3847 12192
rect 3789 12183 3847 12189
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 6104 12229 6132 12260
rect 6270 12248 6276 12260
rect 6328 12248 6334 12300
rect 7392 12297 7420 12328
rect 8018 12316 8024 12328
rect 8076 12316 8082 12368
rect 10226 12356 10232 12368
rect 8220 12328 10232 12356
rect 7377 12291 7435 12297
rect 7377 12257 7389 12291
rect 7423 12257 7435 12291
rect 7377 12251 7435 12257
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12288 7527 12291
rect 8110 12288 8116 12300
rect 7515 12260 8116 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 5905 12223 5963 12229
rect 5905 12189 5917 12223
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 6089 12223 6147 12229
rect 6089 12189 6101 12223
rect 6135 12189 6147 12223
rect 6089 12183 6147 12189
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12189 6239 12223
rect 6454 12220 6460 12232
rect 6415 12192 6460 12220
rect 6181 12183 6239 12189
rect 4062 12161 4068 12164
rect 1780 12124 2268 12152
rect 4056 12115 4068 12161
rect 4120 12152 4126 12164
rect 4120 12124 4156 12152
rect 4062 12112 4068 12115
rect 4120 12112 4126 12124
rect 5718 12112 5724 12164
rect 5776 12152 5782 12164
rect 5920 12152 5948 12183
rect 5776 12124 5948 12152
rect 6196 12152 6224 12183
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 7098 12220 7104 12232
rect 7059 12192 7104 12220
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 7282 12220 7288 12232
rect 7243 12192 7288 12220
rect 7282 12180 7288 12192
rect 7340 12180 7346 12232
rect 7650 12220 7656 12232
rect 7611 12192 7656 12220
rect 7650 12180 7656 12192
rect 7708 12180 7714 12232
rect 7742 12180 7748 12232
rect 7800 12220 7806 12232
rect 8220 12220 8248 12328
rect 10226 12316 10232 12328
rect 10284 12316 10290 12368
rect 9030 12248 9036 12300
rect 9088 12288 9094 12300
rect 9674 12288 9680 12300
rect 9088 12260 9680 12288
rect 9088 12248 9094 12260
rect 7800 12192 8248 12220
rect 7800 12180 7806 12192
rect 8294 12180 8300 12232
rect 8352 12220 8358 12232
rect 9416 12229 9444 12260
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 13078 12248 13084 12300
rect 13136 12288 13142 12300
rect 13265 12291 13323 12297
rect 13265 12288 13277 12291
rect 13136 12260 13277 12288
rect 13136 12248 13142 12260
rect 13265 12257 13277 12260
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 9401 12223 9459 12229
rect 8352 12192 9352 12220
rect 8352 12180 8358 12192
rect 6362 12152 6368 12164
rect 6196 12124 6368 12152
rect 5776 12112 5782 12124
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 7558 12112 7564 12164
rect 7616 12152 7622 12164
rect 8754 12152 8760 12164
rect 7616 12124 8760 12152
rect 7616 12112 7622 12124
rect 8754 12112 8760 12124
rect 8812 12112 8818 12164
rect 9214 12152 9220 12164
rect 9175 12124 9220 12152
rect 9214 12112 9220 12124
rect 9272 12112 9278 12164
rect 9324 12152 9352 12192
rect 9401 12189 9413 12223
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12220 9643 12223
rect 10318 12220 10324 12232
rect 9631 12192 10324 12220
rect 9631 12189 9643 12192
rect 9585 12183 9643 12189
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10965 12223 11023 12229
rect 10965 12189 10977 12223
rect 11011 12220 11023 12223
rect 12434 12220 12440 12232
rect 11011 12192 12440 12220
rect 11011 12189 11023 12192
rect 10965 12183 11023 12189
rect 12434 12180 12440 12192
rect 12492 12180 12498 12232
rect 12802 12220 12808 12232
rect 12763 12192 12808 12220
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 12986 12220 12992 12232
rect 12947 12192 12992 12220
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12189 13231 12223
rect 13354 12220 13360 12232
rect 13315 12192 13360 12220
rect 13173 12183 13231 12189
rect 9674 12152 9680 12164
rect 9324 12124 9680 12152
rect 9674 12112 9680 12124
rect 9732 12112 9738 12164
rect 11238 12161 11244 12164
rect 9968 12124 11192 12152
rect 2961 12087 3019 12093
rect 2961 12053 2973 12087
rect 3007 12084 3019 12087
rect 3510 12084 3516 12096
rect 3007 12056 3516 12084
rect 3007 12053 3019 12056
rect 2961 12047 3019 12053
rect 3510 12044 3516 12056
rect 3568 12044 3574 12096
rect 4522 12044 4528 12096
rect 4580 12084 4586 12096
rect 5169 12087 5227 12093
rect 5169 12084 5181 12087
rect 4580 12056 5181 12084
rect 4580 12044 4586 12056
rect 5169 12053 5181 12056
rect 5215 12084 5227 12087
rect 5442 12084 5448 12096
rect 5215 12056 5448 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 7837 12087 7895 12093
rect 7837 12053 7849 12087
rect 7883 12084 7895 12087
rect 9968 12084 9996 12124
rect 10134 12084 10140 12096
rect 7883 12056 9996 12084
rect 10095 12056 10140 12084
rect 7883 12053 7895 12056
rect 7837 12047 7895 12053
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 11164 12084 11192 12124
rect 11232 12115 11244 12161
rect 11296 12152 11302 12164
rect 11296 12124 11332 12152
rect 11238 12112 11244 12115
rect 11296 12112 11302 12124
rect 11514 12112 11520 12164
rect 11572 12152 11578 12164
rect 11572 12124 12664 12152
rect 11572 12112 11578 12124
rect 11606 12084 11612 12096
rect 11164 12056 11612 12084
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 12345 12087 12403 12093
rect 12345 12053 12357 12087
rect 12391 12084 12403 12087
rect 12526 12084 12532 12096
rect 12391 12056 12532 12084
rect 12391 12053 12403 12056
rect 12345 12047 12403 12053
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 12636 12084 12664 12124
rect 12710 12112 12716 12164
rect 12768 12152 12774 12164
rect 13188 12152 13216 12183
rect 13354 12180 13360 12192
rect 13412 12180 13418 12232
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 13814 12220 13820 12232
rect 13587 12192 13820 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 13814 12180 13820 12192
rect 13872 12180 13878 12232
rect 14016 12220 14044 12396
rect 14108 12396 14280 12424
rect 14108 12297 14136 12396
rect 14274 12384 14280 12396
rect 14332 12424 14338 12436
rect 14458 12424 14464 12436
rect 14332 12396 14464 12424
rect 14332 12384 14338 12396
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 17218 12384 17224 12436
rect 17276 12424 17282 12436
rect 17865 12427 17923 12433
rect 17865 12424 17877 12427
rect 17276 12396 17877 12424
rect 17276 12384 17282 12396
rect 17865 12393 17877 12396
rect 17911 12393 17923 12427
rect 17865 12387 17923 12393
rect 15194 12316 15200 12368
rect 15252 12356 15258 12368
rect 19610 12356 19616 12368
rect 15252 12328 19616 12356
rect 15252 12316 15258 12328
rect 19610 12316 19616 12328
rect 19668 12316 19674 12368
rect 14093 12291 14151 12297
rect 14093 12257 14105 12291
rect 14139 12257 14151 12291
rect 16758 12288 16764 12300
rect 14093 12251 14151 12257
rect 15120 12260 16764 12288
rect 15120 12220 15148 12260
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 18509 12291 18567 12297
rect 18509 12257 18521 12291
rect 18555 12288 18567 12291
rect 21174 12288 21180 12300
rect 18555 12260 21180 12288
rect 18555 12257 18567 12260
rect 18509 12251 18567 12257
rect 21174 12248 21180 12260
rect 21232 12248 21238 12300
rect 14016 12192 15148 12220
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12189 15991 12223
rect 16206 12220 16212 12232
rect 16167 12192 16212 12220
rect 15933 12183 15991 12189
rect 12768 12124 13216 12152
rect 14360 12155 14418 12161
rect 12768 12112 12774 12124
rect 14360 12121 14372 12155
rect 14406 12152 14418 12155
rect 14826 12152 14832 12164
rect 14406 12124 14832 12152
rect 14406 12121 14418 12124
rect 14360 12115 14418 12121
rect 14826 12112 14832 12124
rect 14884 12112 14890 12164
rect 14918 12112 14924 12164
rect 14976 12152 14982 12164
rect 15948 12152 15976 12183
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 17990 12223 18048 12229
rect 17990 12189 18002 12223
rect 18036 12189 18048 12223
rect 17990 12183 18048 12189
rect 18005 12152 18033 12183
rect 18230 12180 18236 12232
rect 18288 12220 18294 12232
rect 18417 12223 18475 12229
rect 18417 12220 18429 12223
rect 18288 12192 18429 12220
rect 18288 12180 18294 12192
rect 18417 12189 18429 12192
rect 18463 12189 18475 12223
rect 18417 12183 18475 12189
rect 19610 12180 19616 12232
rect 19668 12220 19674 12232
rect 20533 12223 20591 12229
rect 20533 12220 20545 12223
rect 19668 12192 20545 12220
rect 19668 12180 19674 12192
rect 20533 12189 20545 12192
rect 20579 12220 20591 12223
rect 21910 12220 21916 12232
rect 20579 12192 21916 12220
rect 20579 12189 20591 12192
rect 20533 12183 20591 12189
rect 21910 12180 21916 12192
rect 21968 12180 21974 12232
rect 28994 12180 29000 12232
rect 29052 12220 29058 12232
rect 29917 12223 29975 12229
rect 29917 12220 29929 12223
rect 29052 12192 29929 12220
rect 29052 12180 29058 12192
rect 29917 12189 29929 12192
rect 29963 12189 29975 12223
rect 29917 12183 29975 12189
rect 30101 12223 30159 12229
rect 30101 12189 30113 12223
rect 30147 12220 30159 12223
rect 30282 12220 30288 12232
rect 30147 12192 30288 12220
rect 30147 12189 30159 12192
rect 30101 12183 30159 12189
rect 14976 12124 15976 12152
rect 16045 12124 18033 12152
rect 14976 12112 14982 12124
rect 14550 12084 14556 12096
rect 12636 12056 14556 12084
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 15470 12084 15476 12096
rect 15383 12056 15476 12084
rect 15470 12044 15476 12056
rect 15528 12084 15534 12096
rect 16045 12084 16073 12124
rect 19058 12112 19064 12164
rect 19116 12152 19122 12164
rect 19245 12155 19303 12161
rect 19245 12152 19257 12155
rect 19116 12124 19257 12152
rect 19116 12112 19122 12124
rect 19245 12121 19257 12124
rect 19291 12121 19303 12155
rect 19245 12115 19303 12121
rect 19429 12155 19487 12161
rect 19429 12121 19441 12155
rect 19475 12152 19487 12155
rect 20070 12152 20076 12164
rect 19475 12124 20076 12152
rect 19475 12121 19487 12124
rect 19429 12115 19487 12121
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 29178 12112 29184 12164
rect 29236 12152 29242 12164
rect 30116 12152 30144 12183
rect 30282 12180 30288 12192
rect 30340 12180 30346 12232
rect 29236 12124 30144 12152
rect 29236 12112 29242 12124
rect 15528 12056 16073 12084
rect 15528 12044 15534 12056
rect 16390 12044 16396 12096
rect 16448 12084 16454 12096
rect 18049 12087 18107 12093
rect 18049 12084 18061 12087
rect 16448 12056 18061 12084
rect 16448 12044 16454 12056
rect 18049 12053 18061 12056
rect 18095 12084 18107 12087
rect 18506 12084 18512 12096
rect 18095 12056 18512 12084
rect 18095 12053 18107 12056
rect 18049 12047 18107 12053
rect 18506 12044 18512 12056
rect 18564 12044 18570 12096
rect 19613 12087 19671 12093
rect 19613 12053 19625 12087
rect 19659 12084 19671 12087
rect 19794 12084 19800 12096
rect 19659 12056 19800 12084
rect 19659 12053 19671 12056
rect 19613 12047 19671 12053
rect 19794 12044 19800 12056
rect 19852 12044 19858 12096
rect 29822 12044 29828 12096
rect 29880 12084 29886 12096
rect 30009 12087 30067 12093
rect 30009 12084 30021 12087
rect 29880 12056 30021 12084
rect 29880 12044 29886 12056
rect 30009 12053 30021 12056
rect 30055 12053 30067 12087
rect 30009 12047 30067 12053
rect 1104 11994 30820 12016
rect 1104 11942 10880 11994
rect 10932 11942 10944 11994
rect 10996 11942 11008 11994
rect 11060 11942 11072 11994
rect 11124 11942 11136 11994
rect 11188 11942 20811 11994
rect 20863 11942 20875 11994
rect 20927 11942 20939 11994
rect 20991 11942 21003 11994
rect 21055 11942 21067 11994
rect 21119 11942 30820 11994
rect 1104 11920 30820 11942
rect 4982 11880 4988 11892
rect 2976 11852 4988 11880
rect 2866 11812 2872 11824
rect 2424 11784 2872 11812
rect 1394 11744 1400 11756
rect 1355 11716 1400 11744
rect 1394 11704 1400 11716
rect 1452 11704 1458 11756
rect 2424 11753 2452 11784
rect 2866 11772 2872 11784
rect 2924 11772 2930 11824
rect 2976 11753 3004 11852
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 10965 11883 11023 11889
rect 5132 11852 6500 11880
rect 5132 11840 5138 11852
rect 4614 11812 4620 11824
rect 3620 11784 4620 11812
rect 3620 11753 3648 11784
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 5442 11772 5448 11824
rect 5500 11812 5506 11824
rect 5500 11784 6408 11812
rect 5500 11772 5506 11784
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11713 2467 11747
rect 2409 11707 2467 11713
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11713 2651 11747
rect 2593 11707 2651 11713
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11713 3019 11747
rect 2961 11707 3019 11713
rect 3605 11747 3663 11753
rect 3605 11713 3617 11747
rect 3651 11713 3663 11747
rect 3861 11747 3919 11753
rect 3861 11744 3873 11747
rect 3605 11707 3663 11713
rect 3712 11716 3873 11744
rect 2608 11676 2636 11707
rect 1596 11648 2636 11676
rect 2685 11679 2743 11685
rect 1596 11617 1624 11648
rect 2685 11645 2697 11679
rect 2731 11645 2743 11679
rect 2685 11639 2743 11645
rect 1581 11611 1639 11617
rect 1581 11577 1593 11611
rect 1627 11577 1639 11611
rect 1581 11571 1639 11577
rect 1946 11568 1952 11620
rect 2004 11608 2010 11620
rect 2590 11608 2596 11620
rect 2004 11580 2596 11608
rect 2004 11568 2010 11580
rect 2590 11568 2596 11580
rect 2648 11608 2654 11620
rect 2700 11608 2728 11639
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 3145 11679 3203 11685
rect 2832 11648 2877 11676
rect 2832 11636 2838 11648
rect 3145 11645 3157 11679
rect 3191 11676 3203 11679
rect 3712 11676 3740 11716
rect 3861 11713 3873 11716
rect 3907 11713 3919 11747
rect 3861 11707 3919 11713
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11744 5687 11747
rect 5810 11744 5816 11756
rect 5675 11716 5816 11744
rect 5675 11713 5687 11716
rect 5629 11707 5687 11713
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 6380 11753 6408 11784
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6472 11744 6500 11852
rect 7392 11852 10539 11880
rect 7006 11744 7012 11756
rect 6472 11716 7012 11744
rect 6365 11707 6423 11713
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 7392 11753 7420 11852
rect 10042 11812 10048 11824
rect 8220 11784 10048 11812
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11713 7435 11747
rect 7558 11744 7564 11756
rect 7519 11716 7564 11744
rect 7377 11707 7435 11713
rect 7208 11676 7236 11707
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 8220 11753 8248 11784
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 8205 11747 8263 11753
rect 8205 11744 8217 11747
rect 7852 11716 8217 11744
rect 3191 11648 3740 11676
rect 4908 11648 7236 11676
rect 7285 11679 7343 11685
rect 3191 11645 3203 11648
rect 3145 11639 3203 11645
rect 2648 11580 2728 11608
rect 2648 11568 2654 11580
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 4908 11540 4936 11648
rect 7285 11645 7297 11679
rect 7331 11676 7343 11679
rect 7742 11676 7748 11688
rect 7331 11648 7748 11676
rect 7331 11645 7343 11648
rect 7285 11639 7343 11645
rect 7742 11636 7748 11648
rect 7800 11636 7806 11688
rect 5813 11611 5871 11617
rect 5813 11577 5825 11611
rect 5859 11608 5871 11611
rect 7852 11608 7880 11716
rect 8205 11713 8217 11716
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 8472 11747 8530 11753
rect 8472 11713 8484 11747
rect 8518 11744 8530 11747
rect 10134 11744 10140 11756
rect 8518 11716 10140 11744
rect 8518 11713 8530 11716
rect 8472 11707 8530 11713
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10244 11676 10272 11707
rect 10318 11704 10324 11756
rect 10376 11746 10382 11756
rect 10413 11747 10471 11753
rect 10413 11746 10425 11747
rect 10376 11718 10425 11746
rect 10376 11704 10382 11718
rect 10413 11713 10425 11718
rect 10459 11713 10471 11747
rect 10511 11746 10539 11852
rect 10965 11849 10977 11883
rect 11011 11880 11023 11883
rect 11238 11880 11244 11892
rect 11011 11852 11244 11880
rect 11011 11849 11023 11852
rect 10965 11843 11023 11849
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 12986 11840 12992 11892
rect 13044 11880 13050 11892
rect 13817 11883 13875 11889
rect 13817 11880 13829 11883
rect 13044 11852 13829 11880
rect 13044 11840 13050 11852
rect 13817 11849 13829 11852
rect 13863 11880 13875 11883
rect 14182 11880 14188 11892
rect 13863 11852 14188 11880
rect 13863 11849 13875 11852
rect 13817 11843 13875 11849
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 15657 11883 15715 11889
rect 15657 11849 15669 11883
rect 15703 11880 15715 11883
rect 17586 11880 17592 11892
rect 15703 11852 17592 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 12704 11815 12762 11821
rect 12704 11781 12716 11815
rect 12750 11812 12762 11815
rect 12802 11812 12808 11824
rect 12750 11784 12808 11812
rect 12750 11781 12762 11784
rect 12704 11775 12762 11781
rect 12802 11772 12808 11784
rect 12860 11772 12866 11824
rect 13446 11772 13452 11824
rect 13504 11812 13510 11824
rect 15672 11812 15700 11843
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 17862 11880 17868 11892
rect 17823 11852 17868 11880
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 18138 11840 18144 11892
rect 18196 11880 18202 11892
rect 18325 11883 18383 11889
rect 18325 11880 18337 11883
rect 18196 11852 18337 11880
rect 18196 11840 18202 11852
rect 18325 11849 18337 11852
rect 18371 11849 18383 11883
rect 18506 11880 18512 11892
rect 18467 11852 18512 11880
rect 18325 11843 18383 11849
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 20530 11880 20536 11892
rect 20491 11852 20536 11880
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 21174 11880 21180 11892
rect 21135 11852 21180 11880
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 18230 11812 18236 11824
rect 13504 11784 15700 11812
rect 16500 11784 18236 11812
rect 13504 11772 13510 11784
rect 10597 11747 10655 11753
rect 10511 11744 10548 11746
rect 10597 11744 10609 11747
rect 10511 11718 10609 11744
rect 10520 11716 10609 11718
rect 10413 11707 10471 11713
rect 10597 11713 10609 11716
rect 10643 11744 10655 11747
rect 10781 11747 10839 11753
rect 10643 11716 10741 11744
rect 10643 11713 10655 11716
rect 10597 11707 10655 11713
rect 10502 11676 10508 11688
rect 10008 11648 10272 11676
rect 10463 11648 10508 11676
rect 10008 11636 10014 11648
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 10713 11676 10741 11716
rect 10781 11713 10793 11747
rect 10827 11744 10839 11747
rect 12526 11744 12532 11756
rect 10827 11716 12532 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 12526 11704 12532 11716
rect 12584 11744 12590 11756
rect 13906 11744 13912 11756
rect 12584 11716 13912 11744
rect 12584 11704 12590 11716
rect 13906 11704 13912 11716
rect 13964 11704 13970 11756
rect 14274 11744 14280 11756
rect 14235 11716 14280 11744
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 14366 11704 14372 11756
rect 14424 11744 14430 11756
rect 14533 11747 14591 11753
rect 14533 11744 14545 11747
rect 14424 11716 14545 11744
rect 14424 11704 14430 11716
rect 14533 11713 14545 11716
rect 14579 11713 14591 11747
rect 14533 11707 14591 11713
rect 11238 11676 11244 11688
rect 10713 11648 11244 11676
rect 11238 11636 11244 11648
rect 11296 11636 11302 11688
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 12492 11648 12537 11676
rect 12492 11636 12498 11648
rect 8202 11608 8208 11620
rect 5859 11580 8208 11608
rect 5859 11577 5871 11580
rect 5813 11571 5871 11577
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 11514 11608 11520 11620
rect 9140 11580 11520 11608
rect 6454 11540 6460 11552
rect 2188 11512 4936 11540
rect 6415 11512 6460 11540
rect 2188 11500 2194 11512
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 7742 11540 7748 11552
rect 7703 11512 7748 11540
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 9140 11540 9168 11580
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 15654 11568 15660 11620
rect 15712 11608 15718 11620
rect 16390 11608 16396 11620
rect 15712 11580 16396 11608
rect 15712 11568 15718 11580
rect 16390 11568 16396 11580
rect 16448 11568 16454 11620
rect 8076 11512 9168 11540
rect 8076 11500 8082 11512
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 9456 11512 9597 11540
rect 9456 11500 9462 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 16500 11540 16528 11784
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 17512 11753 17540 11784
rect 18230 11772 18236 11784
rect 18288 11812 18294 11824
rect 18288 11784 18920 11812
rect 18288 11772 18294 11784
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 16632 11716 17141 11744
rect 16632 11704 16638 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 17313 11747 17371 11753
rect 17313 11713 17325 11747
rect 17359 11713 17371 11747
rect 17313 11707 17371 11713
rect 17497 11747 17555 11753
rect 17497 11713 17509 11747
rect 17543 11713 17555 11747
rect 17678 11744 17684 11756
rect 17639 11716 17684 11744
rect 17497 11707 17555 11713
rect 17328 11608 17356 11707
rect 17678 11704 17684 11716
rect 17736 11704 17742 11756
rect 17770 11704 17776 11756
rect 17828 11744 17834 11756
rect 18892 11753 18920 11784
rect 19886 11772 19892 11824
rect 19944 11812 19950 11824
rect 19944 11784 20208 11812
rect 19944 11772 19950 11784
rect 18450 11747 18508 11753
rect 18450 11744 18462 11747
rect 17828 11716 18462 11744
rect 17828 11704 17834 11716
rect 18450 11713 18462 11716
rect 18496 11713 18508 11747
rect 18450 11707 18508 11713
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11713 18935 11747
rect 18877 11707 18935 11713
rect 19518 11704 19524 11756
rect 19576 11744 19582 11756
rect 19797 11747 19855 11753
rect 19797 11744 19809 11747
rect 19576 11716 19809 11744
rect 19576 11704 19582 11716
rect 19797 11713 19809 11716
rect 19843 11713 19855 11747
rect 19978 11744 19984 11756
rect 19939 11716 19984 11744
rect 19797 11707 19855 11713
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20180 11753 20208 11784
rect 20165 11747 20223 11753
rect 20165 11713 20177 11747
rect 20211 11713 20223 11747
rect 20346 11744 20352 11756
rect 20307 11716 20352 11744
rect 20165 11707 20223 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 21177 11747 21235 11753
rect 21177 11713 21189 11747
rect 21223 11744 21235 11747
rect 21358 11744 21364 11756
rect 21223 11716 21364 11744
rect 21223 11713 21235 11716
rect 21177 11707 21235 11713
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 29178 11744 29184 11756
rect 29139 11716 29184 11744
rect 29178 11704 29184 11716
rect 29236 11704 29242 11756
rect 29825 11747 29883 11753
rect 29825 11744 29837 11747
rect 29380 11716 29837 11744
rect 17402 11636 17408 11688
rect 17460 11676 17466 11688
rect 18969 11679 19027 11685
rect 17460 11648 17505 11676
rect 17460 11636 17466 11648
rect 18969 11645 18981 11679
rect 19015 11676 19027 11679
rect 19702 11676 19708 11688
rect 19015 11648 19708 11676
rect 19015 11645 19027 11648
rect 18969 11639 19027 11645
rect 19702 11636 19708 11648
rect 19760 11636 19766 11688
rect 20070 11676 20076 11688
rect 20031 11648 20076 11676
rect 20070 11636 20076 11648
rect 20128 11636 20134 11688
rect 18046 11608 18052 11620
rect 17328 11580 18052 11608
rect 18046 11568 18052 11580
rect 18104 11568 18110 11620
rect 29380 11617 29408 11716
rect 29825 11713 29837 11716
rect 29871 11713 29883 11747
rect 29825 11707 29883 11713
rect 29365 11611 29423 11617
rect 29365 11577 29377 11611
rect 29411 11577 29423 11611
rect 29365 11571 29423 11577
rect 9732 11512 16528 11540
rect 9732 11500 9738 11512
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 22094 11540 22100 11552
rect 17184 11512 22100 11540
rect 17184 11500 17190 11512
rect 22094 11500 22100 11512
rect 22152 11500 22158 11552
rect 30006 11540 30012 11552
rect 29967 11512 30012 11540
rect 30006 11500 30012 11512
rect 30064 11500 30070 11552
rect 1104 11450 30820 11472
rect 1104 11398 5915 11450
rect 5967 11398 5979 11450
rect 6031 11398 6043 11450
rect 6095 11398 6107 11450
rect 6159 11398 6171 11450
rect 6223 11398 15846 11450
rect 15898 11398 15910 11450
rect 15962 11398 15974 11450
rect 16026 11398 16038 11450
rect 16090 11398 16102 11450
rect 16154 11398 25776 11450
rect 25828 11398 25840 11450
rect 25892 11398 25904 11450
rect 25956 11398 25968 11450
rect 26020 11398 26032 11450
rect 26084 11398 30820 11450
rect 1104 11376 30820 11398
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 6270 11336 6276 11348
rect 5776 11308 6276 11336
rect 5776 11296 5782 11308
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 6914 11336 6920 11348
rect 6827 11308 6920 11336
rect 6914 11296 6920 11308
rect 6972 11336 6978 11348
rect 7558 11336 7564 11348
rect 6972 11308 7564 11336
rect 6972 11296 6978 11308
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 7650 11296 7656 11348
rect 7708 11336 7714 11348
rect 9398 11336 9404 11348
rect 7708 11308 9260 11336
rect 9359 11308 9404 11336
rect 7708 11296 7714 11308
rect 4890 11228 4896 11280
rect 4948 11268 4954 11280
rect 9232 11268 9260 11308
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 11146 11336 11152 11348
rect 10428 11308 11152 11336
rect 10428 11268 10456 11308
rect 11146 11296 11152 11308
rect 11204 11296 11210 11348
rect 13078 11336 13084 11348
rect 11532 11308 13084 11336
rect 11532 11268 11560 11308
rect 13078 11296 13084 11308
rect 13136 11296 13142 11348
rect 13541 11339 13599 11345
rect 13541 11305 13553 11339
rect 13587 11336 13599 11339
rect 14366 11336 14372 11348
rect 13587 11308 14372 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 14826 11336 14832 11348
rect 14787 11308 14832 11336
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 16393 11339 16451 11345
rect 16393 11305 16405 11339
rect 16439 11336 16451 11339
rect 16942 11336 16948 11348
rect 16439 11308 16948 11336
rect 16439 11305 16451 11308
rect 16393 11299 16451 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 17678 11296 17684 11348
rect 17736 11336 17742 11348
rect 18601 11339 18659 11345
rect 18601 11336 18613 11339
rect 17736 11308 18613 11336
rect 17736 11296 17742 11308
rect 18601 11305 18613 11308
rect 18647 11305 18659 11339
rect 18601 11299 18659 11305
rect 20438 11296 20444 11348
rect 20496 11336 20502 11348
rect 20533 11339 20591 11345
rect 20533 11336 20545 11339
rect 20496 11308 20545 11336
rect 20496 11296 20502 11308
rect 20533 11305 20545 11308
rect 20579 11305 20591 11339
rect 20533 11299 20591 11305
rect 4948 11240 7328 11268
rect 9232 11240 10456 11268
rect 11164 11240 11560 11268
rect 4948 11228 4954 11240
rect 5350 11200 5356 11212
rect 5311 11172 5356 11200
rect 5350 11160 5356 11172
rect 5408 11160 5414 11212
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 5166 11132 5172 11144
rect 5127 11104 5172 11132
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 5445 11135 5503 11141
rect 5445 11132 5457 11135
rect 5276 11104 5457 11132
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 5276 11064 5304 11104
rect 5445 11101 5457 11104
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 5534 11092 5540 11144
rect 5592 11141 5598 11144
rect 5592 11135 5631 11141
rect 5619 11132 5631 11135
rect 6822 11132 6828 11144
rect 5619 11104 6828 11132
rect 5619 11101 5631 11104
rect 5592 11095 5631 11101
rect 5592 11092 5598 11095
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 7300 11132 7328 11240
rect 8757 11203 8815 11209
rect 8757 11169 8769 11203
rect 8803 11200 8815 11203
rect 8803 11172 9536 11200
rect 8803 11169 8815 11172
rect 8757 11163 8815 11169
rect 7650 11132 7656 11144
rect 7300 11104 7656 11132
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 7742 11092 7748 11144
rect 7800 11132 7806 11144
rect 8030 11135 8088 11141
rect 8030 11132 8042 11135
rect 7800 11104 8042 11132
rect 7800 11092 7806 11104
rect 8030 11101 8042 11104
rect 8076 11101 8088 11135
rect 8030 11095 8088 11101
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 8297 11135 8355 11141
rect 8297 11132 8309 11135
rect 8260 11104 8309 11132
rect 8260 11092 8266 11104
rect 8297 11101 8309 11104
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8628 11104 8953 11132
rect 8628 11092 8634 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 9272 11104 9321 11132
rect 9272 11092 9278 11104
rect 9309 11101 9321 11104
rect 9355 11132 9367 11135
rect 9398 11132 9404 11144
rect 9355 11104 9404 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 9508 11141 9536 11172
rect 10778 11160 10784 11212
rect 10836 11200 10842 11212
rect 11164 11209 11192 11240
rect 11606 11228 11612 11280
rect 11664 11268 11670 11280
rect 12802 11268 12808 11280
rect 11664 11240 12808 11268
rect 11664 11228 11670 11240
rect 12802 11228 12808 11240
rect 12860 11228 12866 11280
rect 13814 11268 13820 11280
rect 12912 11240 13820 11268
rect 11149 11203 11207 11209
rect 11149 11200 11161 11203
rect 10836 11172 11161 11200
rect 10836 11160 10842 11172
rect 11149 11169 11161 11172
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 11514 11200 11520 11212
rect 11296 11172 11520 11200
rect 11296 11160 11302 11172
rect 11514 11160 11520 11172
rect 11572 11200 11578 11212
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 11572 11172 12357 11200
rect 11572 11160 11578 11172
rect 12345 11169 12357 11172
rect 12391 11200 12403 11203
rect 12710 11200 12716 11212
rect 12391 11172 12716 11200
rect 12391 11169 12403 11172
rect 12345 11163 12403 11169
rect 12710 11160 12716 11172
rect 12768 11160 12774 11212
rect 12912 11200 12940 11240
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 13906 11228 13912 11280
rect 13964 11268 13970 11280
rect 17034 11268 17040 11280
rect 13964 11240 17040 11268
rect 13964 11228 13970 11240
rect 17034 11228 17040 11240
rect 17092 11228 17098 11280
rect 19978 11228 19984 11280
rect 20036 11268 20042 11280
rect 21085 11271 21143 11277
rect 21085 11268 21097 11271
rect 20036 11240 21097 11268
rect 20036 11228 20042 11240
rect 21085 11237 21097 11240
rect 21131 11237 21143 11271
rect 21085 11231 21143 11237
rect 13078 11200 13084 11212
rect 12820 11172 12940 11200
rect 13039 11172 13084 11200
rect 12820 11141 12848 11172
rect 13078 11160 13084 11172
rect 13136 11200 13142 11212
rect 14366 11200 14372 11212
rect 13136 11172 14372 11200
rect 13136 11160 13142 11172
rect 14366 11160 14372 11172
rect 14424 11160 14430 11212
rect 16853 11203 16911 11209
rect 16853 11200 16865 11203
rect 15672 11172 16865 11200
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11101 9551 11135
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 9493 11095 9551 11101
rect 10060 11104 10885 11132
rect 2924 11036 5304 11064
rect 2924 11024 2930 11036
rect 5350 11024 5356 11076
rect 5408 11064 5414 11076
rect 5408 11036 5453 11064
rect 5408 11024 5414 11036
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 9950 11064 9956 11076
rect 7064 11036 9956 11064
rect 7064 11024 7070 11036
rect 9950 11024 9956 11036
rect 10008 11064 10014 11076
rect 10060 11064 10088 11104
rect 10873 11101 10885 11104
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 11057 11135 11115 11141
rect 11057 11101 11069 11135
rect 11103 11132 11115 11135
rect 11408 11135 11466 11141
rect 11103 11104 11376 11132
rect 11103 11101 11115 11104
rect 11057 11095 11115 11101
rect 10008 11036 10088 11064
rect 10008 11024 10014 11036
rect 1581 10999 1639 11005
rect 1581 10965 1593 10999
rect 1627 10996 1639 10999
rect 1670 10996 1676 11008
rect 1627 10968 1676 10996
rect 1627 10965 1639 10968
rect 1581 10959 1639 10965
rect 1670 10956 1676 10968
rect 1728 10956 1734 11008
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 8757 10999 8815 11005
rect 8757 10996 8769 10999
rect 7524 10968 8769 10996
rect 7524 10956 7530 10968
rect 8757 10965 8769 10968
rect 8803 10965 8815 10999
rect 9122 10996 9128 11008
rect 9083 10968 9128 10996
rect 8757 10959 8815 10965
rect 9122 10956 9128 10968
rect 9180 10956 9186 11008
rect 10060 10996 10088 11036
rect 10137 11067 10195 11073
rect 10137 11033 10149 11067
rect 10183 11064 10195 11067
rect 10502 11064 10508 11076
rect 10183 11036 10508 11064
rect 10183 11033 10195 11036
rect 10137 11027 10195 11033
rect 10502 11024 10508 11036
rect 10560 11024 10566 11076
rect 11348 11008 11376 11104
rect 11408 11101 11420 11135
rect 11454 11132 11466 11135
rect 12805 11135 12863 11141
rect 11454 11130 11468 11132
rect 11532 11130 12756 11132
rect 11454 11104 12756 11130
rect 11454 11102 11560 11104
rect 11454 11101 11466 11102
rect 11408 11095 11466 11101
rect 12728 11076 12756 11104
rect 12805 11101 12817 11135
rect 12851 11101 12863 11135
rect 12986 11132 12992 11144
rect 12947 11104 12992 11132
rect 12805 11095 12863 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13173 11135 13231 11141
rect 13173 11101 13185 11135
rect 13219 11101 13231 11135
rect 13173 11095 13231 11101
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 13446 11132 13452 11144
rect 13403 11104 13452 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 12158 11024 12164 11076
rect 12216 11064 12222 11076
rect 12216 11036 12261 11064
rect 12216 11024 12222 11036
rect 12710 11024 12716 11076
rect 12768 11024 12774 11076
rect 13078 11024 13084 11076
rect 13136 11064 13142 11076
rect 13188 11064 13216 11095
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13964 11104 14105 11132
rect 13964 11092 13970 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14274 11132 14280 11144
rect 14235 11104 14280 11132
rect 14093 11095 14151 11101
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14458 11132 14464 11144
rect 14419 11104 14464 11132
rect 14458 11092 14464 11104
rect 14516 11092 14522 11144
rect 14656 11135 14714 11141
rect 14656 11101 14668 11135
rect 14702 11132 14714 11135
rect 15470 11132 15476 11144
rect 14702 11104 15476 11132
rect 14702 11101 14714 11104
rect 14656 11095 14714 11101
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 15672 11141 15700 11172
rect 16853 11169 16865 11172
rect 16899 11169 16911 11203
rect 17773 11203 17831 11209
rect 17773 11200 17785 11203
rect 16853 11163 16911 11169
rect 16960 11172 17785 11200
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 15746 11092 15752 11144
rect 15804 11132 15810 11144
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 15804 11104 15853 11132
rect 15804 11092 15810 11104
rect 15841 11101 15853 11104
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11101 15991 11135
rect 15933 11095 15991 11101
rect 13136 11036 13216 11064
rect 13136 11024 13142 11036
rect 15194 11024 15200 11076
rect 15252 11064 15258 11076
rect 15948 11064 15976 11095
rect 16022 11092 16028 11144
rect 16080 11132 16086 11144
rect 16206 11132 16212 11144
rect 16080 11104 16125 11132
rect 16167 11104 16212 11132
rect 16080 11092 16086 11104
rect 16206 11092 16212 11104
rect 16264 11092 16270 11144
rect 16390 11092 16396 11144
rect 16448 11132 16454 11144
rect 16960 11132 16988 11172
rect 17773 11169 17785 11172
rect 17819 11169 17831 11203
rect 17773 11163 17831 11169
rect 19886 11160 19892 11212
rect 19944 11200 19950 11212
rect 20165 11203 20223 11209
rect 20165 11200 20177 11203
rect 19944 11172 20177 11200
rect 19944 11160 19950 11172
rect 20165 11169 20177 11172
rect 20211 11169 20223 11203
rect 20165 11163 20223 11169
rect 17310 11135 17316 11144
rect 16448 11104 16988 11132
rect 17257 11129 17316 11135
rect 16448 11092 16454 11104
rect 16868 11073 16896 11104
rect 17257 11095 17269 11129
rect 17303 11095 17316 11129
rect 17257 11092 17316 11095
rect 17368 11092 17374 11144
rect 17954 11132 17960 11144
rect 17915 11104 17960 11132
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 18509 11135 18567 11141
rect 18509 11101 18521 11135
rect 18555 11132 18567 11135
rect 18874 11132 18880 11144
rect 18555 11104 18880 11132
rect 18555 11101 18567 11104
rect 18509 11095 18567 11101
rect 18874 11092 18880 11104
rect 18932 11092 18938 11144
rect 19794 11132 19800 11144
rect 19755 11104 19800 11132
rect 19794 11092 19800 11104
rect 19852 11092 19858 11144
rect 19981 11135 20039 11141
rect 19981 11101 19993 11135
rect 20027 11101 20039 11135
rect 19981 11095 20039 11101
rect 17257 11089 17315 11092
rect 16853 11067 16911 11073
rect 15252 11036 16804 11064
rect 15252 11024 15258 11036
rect 10229 10999 10287 11005
rect 10229 10996 10241 10999
rect 10060 10968 10241 10996
rect 10229 10965 10241 10968
rect 10275 10965 10287 10999
rect 10229 10959 10287 10965
rect 11330 10956 11336 11008
rect 11388 10956 11394 11008
rect 11609 10999 11667 11005
rect 11609 10965 11621 10999
rect 11655 10996 11667 10999
rect 11882 10996 11888 11008
rect 11655 10968 11888 10996
rect 11655 10965 11667 10968
rect 11609 10959 11667 10965
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 15838 10956 15844 11008
rect 15896 10996 15902 11008
rect 16574 10996 16580 11008
rect 15896 10968 16580 10996
rect 15896 10956 15902 10968
rect 16574 10956 16580 10968
rect 16632 10956 16638 11008
rect 16776 10996 16804 11036
rect 16853 11033 16865 11067
rect 16899 11033 16911 11067
rect 17034 11064 17040 11076
rect 16995 11036 17040 11064
rect 16853 11027 16911 11033
rect 17034 11024 17040 11036
rect 17092 11024 17098 11076
rect 17126 11024 17132 11076
rect 17184 11064 17190 11076
rect 19996 11064 20024 11095
rect 20070 11092 20076 11144
rect 20128 11132 20134 11144
rect 20128 11104 20173 11132
rect 20128 11092 20134 11104
rect 20254 11092 20260 11144
rect 20312 11132 20318 11144
rect 20349 11135 20407 11141
rect 20349 11132 20361 11135
rect 20312 11104 20361 11132
rect 20312 11092 20318 11104
rect 20349 11101 20361 11104
rect 20395 11101 20407 11135
rect 20349 11095 20407 11101
rect 21177 11135 21235 11141
rect 21177 11101 21189 11135
rect 21223 11132 21235 11135
rect 21726 11132 21732 11144
rect 21223 11104 21732 11132
rect 21223 11101 21235 11104
rect 21177 11095 21235 11101
rect 21726 11092 21732 11104
rect 21784 11092 21790 11144
rect 20714 11064 20720 11076
rect 17184 11036 17229 11064
rect 19996 11036 20720 11064
rect 17184 11024 17190 11036
rect 20714 11024 20720 11036
rect 20772 11024 20778 11076
rect 17218 10996 17224 11008
rect 16776 10968 17224 10996
rect 17218 10956 17224 10968
rect 17276 10996 17282 11008
rect 17402 10996 17408 11008
rect 17276 10968 17408 10996
rect 17276 10956 17282 10968
rect 17402 10956 17408 10968
rect 17460 10956 17466 11008
rect 1104 10906 30820 10928
rect 1104 10854 10880 10906
rect 10932 10854 10944 10906
rect 10996 10854 11008 10906
rect 11060 10854 11072 10906
rect 11124 10854 11136 10906
rect 11188 10854 20811 10906
rect 20863 10854 20875 10906
rect 20927 10854 20939 10906
rect 20991 10854 21003 10906
rect 21055 10854 21067 10906
rect 21119 10854 30820 10906
rect 1104 10832 30820 10854
rect 2866 10792 2872 10804
rect 2827 10764 2872 10792
rect 2866 10752 2872 10764
rect 2924 10752 2930 10804
rect 6825 10795 6883 10801
rect 5000 10764 5396 10792
rect 5000 10736 5028 10764
rect 4982 10684 4988 10736
rect 5040 10684 5046 10736
rect 5077 10727 5135 10733
rect 5077 10693 5089 10727
rect 5123 10724 5135 10727
rect 5166 10724 5172 10736
rect 5123 10696 5172 10724
rect 5123 10693 5135 10696
rect 5077 10687 5135 10693
rect 5166 10684 5172 10696
rect 5224 10684 5230 10736
rect 5368 10733 5396 10764
rect 6825 10761 6837 10795
rect 6871 10792 6883 10795
rect 7282 10792 7288 10804
rect 6871 10764 7288 10792
rect 6871 10761 6883 10764
rect 6825 10755 6883 10761
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10134 10792 10140 10804
rect 10008 10764 10140 10792
rect 10008 10752 10014 10764
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 12158 10792 12164 10804
rect 11296 10764 12164 10792
rect 11296 10752 11302 10764
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 15105 10795 15163 10801
rect 15105 10761 15117 10795
rect 15151 10792 15163 10795
rect 16206 10792 16212 10804
rect 15151 10764 16212 10792
rect 15151 10761 15163 10764
rect 15105 10755 15163 10761
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 17310 10752 17316 10804
rect 17368 10752 17374 10804
rect 17494 10792 17500 10804
rect 17455 10764 17500 10792
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 18046 10792 18052 10804
rect 18007 10764 18052 10792
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 19886 10752 19892 10804
rect 19944 10752 19950 10804
rect 20441 10795 20499 10801
rect 20441 10761 20453 10795
rect 20487 10792 20499 10795
rect 20622 10792 20628 10804
rect 20487 10764 20628 10792
rect 20487 10761 20499 10764
rect 20441 10755 20499 10761
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 20993 10795 21051 10801
rect 20993 10792 21005 10795
rect 20772 10764 21005 10792
rect 20772 10752 20778 10764
rect 20993 10761 21005 10764
rect 21039 10761 21051 10795
rect 20993 10755 21051 10761
rect 5353 10727 5411 10733
rect 5353 10693 5365 10727
rect 5399 10693 5411 10727
rect 5353 10687 5411 10693
rect 5810 10684 5816 10736
rect 5868 10724 5874 10736
rect 7377 10727 7435 10733
rect 7377 10724 7389 10727
rect 5868 10696 7389 10724
rect 5868 10684 5874 10696
rect 7377 10693 7389 10696
rect 7423 10693 7435 10727
rect 7377 10687 7435 10693
rect 8573 10727 8631 10733
rect 8573 10693 8585 10727
rect 8619 10724 8631 10727
rect 10778 10724 10784 10736
rect 8619 10696 10784 10724
rect 8619 10693 8631 10696
rect 8573 10687 8631 10693
rect 10778 10684 10784 10696
rect 10836 10724 10842 10736
rect 11701 10727 11759 10733
rect 11701 10724 11713 10727
rect 10836 10696 11713 10724
rect 10836 10684 10842 10696
rect 11701 10693 11713 10696
rect 11747 10693 11759 10727
rect 11701 10687 11759 10693
rect 1486 10656 1492 10668
rect 1447 10628 1492 10656
rect 1486 10616 1492 10628
rect 1544 10616 1550 10668
rect 1756 10659 1814 10665
rect 1756 10625 1768 10659
rect 1802 10656 1814 10659
rect 2222 10656 2228 10668
rect 1802 10628 2228 10656
rect 1802 10625 1814 10628
rect 1756 10619 1814 10625
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 4890 10616 4896 10668
rect 4948 10656 4954 10668
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 4948 10628 5273 10656
rect 4948 10616 4954 10628
rect 5261 10625 5273 10628
rect 5307 10625 5319 10659
rect 5442 10656 5448 10668
rect 5500 10665 5506 10668
rect 5408 10628 5448 10656
rect 5261 10619 5319 10625
rect 5442 10616 5448 10628
rect 5500 10619 5508 10665
rect 6914 10656 6920 10668
rect 6875 10628 6920 10656
rect 5500 10616 5506 10619
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7834 10656 7840 10668
rect 7607 10628 7840 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 7834 10616 7840 10628
rect 7892 10656 7898 10668
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 7892 10628 8401 10656
rect 7892 10616 7898 10628
rect 8389 10625 8401 10628
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 8846 10616 8852 10668
rect 8904 10656 8910 10668
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 8904 10628 9137 10656
rect 8904 10616 8910 10628
rect 9125 10625 9137 10628
rect 9171 10656 9183 10659
rect 9217 10659 9275 10665
rect 9217 10656 9229 10659
rect 9171 10628 9229 10656
rect 9171 10625 9183 10628
rect 9125 10619 9183 10625
rect 9217 10625 9229 10628
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10656 9459 10659
rect 9447 10628 10088 10656
rect 9447 10625 9459 10628
rect 9401 10619 9459 10625
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 7800 10560 9597 10588
rect 7800 10548 7806 10560
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 10060 10588 10088 10628
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10318 10656 10324 10668
rect 10192 10628 10237 10656
rect 10279 10628 10324 10656
rect 10192 10616 10198 10628
rect 10318 10616 10324 10628
rect 10376 10616 10382 10668
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10656 10747 10659
rect 11606 10656 11612 10668
rect 10735 10628 11612 10656
rect 10735 10625 10747 10628
rect 10689 10619 10747 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12176 10656 12204 10752
rect 14277 10727 14335 10733
rect 14277 10693 14289 10727
rect 14323 10724 14335 10727
rect 15746 10724 15752 10736
rect 14323 10696 15752 10724
rect 14323 10693 14335 10696
rect 14277 10687 14335 10693
rect 15746 10684 15752 10696
rect 15804 10684 15810 10736
rect 17328 10724 17356 10752
rect 16592 10696 17356 10724
rect 19904 10724 19932 10752
rect 19904 10696 20116 10724
rect 12345 10659 12403 10665
rect 12345 10656 12357 10659
rect 12176 10628 12357 10656
rect 12345 10625 12357 10628
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 12621 10659 12679 10665
rect 12621 10625 12633 10659
rect 12667 10656 12679 10659
rect 13078 10656 13084 10668
rect 12667 10628 13084 10656
rect 12667 10625 12679 10628
rect 12621 10619 12679 10625
rect 13078 10616 13084 10628
rect 13136 10656 13142 10668
rect 13998 10656 14004 10668
rect 13136 10628 14004 10656
rect 13136 10616 13142 10628
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 14182 10656 14188 10668
rect 14143 10628 14188 10656
rect 14182 10616 14188 10628
rect 14240 10616 14246 10668
rect 15194 10656 15200 10668
rect 15155 10628 15200 10656
rect 15194 10616 15200 10628
rect 15252 10616 15258 10668
rect 15654 10656 15660 10668
rect 15615 10628 15660 10656
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 15841 10659 15899 10665
rect 15841 10625 15853 10659
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 16061 10659 16119 10665
rect 16061 10625 16073 10659
rect 16107 10656 16119 10659
rect 16592 10656 16620 10696
rect 16107 10628 16620 10656
rect 16107 10625 16119 10628
rect 16061 10619 16119 10625
rect 10060 10560 10180 10588
rect 9585 10551 9643 10557
rect 10152 10532 10180 10560
rect 10226 10548 10232 10600
rect 10284 10588 10290 10600
rect 10413 10591 10471 10597
rect 10413 10588 10425 10591
rect 10284 10560 10425 10588
rect 10284 10548 10290 10560
rect 10413 10557 10425 10560
rect 10459 10557 10471 10591
rect 10413 10551 10471 10557
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10588 10563 10591
rect 11514 10588 11520 10600
rect 10551 10560 11520 10588
rect 10551 10557 10563 10560
rect 10505 10551 10563 10557
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 15746 10588 15752 10600
rect 15707 10560 15752 10588
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 5077 10523 5135 10529
rect 5077 10489 5089 10523
rect 5123 10520 5135 10523
rect 5258 10520 5264 10532
rect 5123 10492 5264 10520
rect 5123 10489 5135 10492
rect 5077 10483 5135 10489
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 10134 10480 10140 10532
rect 10192 10480 10198 10532
rect 11885 10523 11943 10529
rect 11885 10489 11897 10523
rect 11931 10520 11943 10523
rect 13630 10520 13636 10532
rect 11931 10492 13636 10520
rect 11931 10489 11943 10492
rect 11885 10483 11943 10489
rect 13630 10480 13636 10492
rect 13688 10520 13694 10532
rect 14550 10520 14556 10532
rect 13688 10492 14556 10520
rect 13688 10480 13694 10492
rect 14550 10480 14556 10492
rect 14608 10480 14614 10532
rect 15856 10520 15884 10619
rect 15764 10492 15884 10520
rect 9125 10455 9183 10461
rect 9125 10421 9137 10455
rect 9171 10452 9183 10455
rect 9674 10452 9680 10464
rect 9171 10424 9680 10452
rect 9171 10421 9183 10424
rect 9125 10415 9183 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 10870 10452 10876 10464
rect 10831 10424 10876 10452
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 13446 10412 13452 10464
rect 13504 10452 13510 10464
rect 15764 10452 15792 10492
rect 13504 10424 15792 10452
rect 15948 10452 15976 10619
rect 16666 10616 16672 10668
rect 16724 10656 16730 10668
rect 16761 10659 16819 10665
rect 16761 10656 16773 10659
rect 16724 10628 16773 10656
rect 16724 10616 16730 10628
rect 16761 10625 16773 10628
rect 16807 10625 16819 10659
rect 16942 10656 16948 10668
rect 16903 10628 16948 10656
rect 16761 10619 16819 10625
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17218 10656 17224 10668
rect 17083 10628 17224 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 17313 10659 17371 10665
rect 17313 10625 17325 10659
rect 17359 10656 17371 10659
rect 17494 10656 17500 10668
rect 17359 10628 17500 10656
rect 17359 10625 17371 10628
rect 17313 10619 17371 10625
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 17957 10659 18015 10665
rect 17957 10656 17969 10659
rect 17644 10628 17969 10656
rect 17644 10616 17650 10628
rect 17957 10625 17969 10628
rect 18003 10625 18015 10659
rect 18782 10656 18788 10668
rect 18743 10628 18788 10656
rect 17957 10619 18015 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 19705 10659 19763 10665
rect 19705 10656 19717 10659
rect 19260 10628 19717 10656
rect 19260 10597 19288 10628
rect 19705 10625 19717 10628
rect 19751 10625 19763 10659
rect 19886 10656 19892 10668
rect 19847 10628 19892 10656
rect 19705 10619 19763 10625
rect 19886 10616 19892 10628
rect 19944 10616 19950 10668
rect 20088 10665 20116 10696
rect 20073 10659 20131 10665
rect 20073 10625 20085 10659
rect 20119 10625 20131 10659
rect 20254 10656 20260 10668
rect 20215 10628 20260 10656
rect 20073 10619 20131 10625
rect 20254 10616 20260 10628
rect 20312 10616 20318 10668
rect 21085 10659 21143 10665
rect 21085 10625 21097 10659
rect 21131 10656 21143 10659
rect 21174 10656 21180 10668
rect 21131 10628 21180 10656
rect 21131 10625 21143 10628
rect 21085 10619 21143 10625
rect 21174 10616 21180 10628
rect 21232 10616 21238 10668
rect 17129 10591 17187 10597
rect 17129 10557 17141 10591
rect 17175 10557 17187 10591
rect 17129 10551 17187 10557
rect 19245 10591 19303 10597
rect 19245 10557 19257 10591
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10557 20039 10591
rect 19981 10551 20039 10557
rect 16022 10480 16028 10532
rect 16080 10520 16086 10532
rect 17144 10520 17172 10551
rect 19996 10520 20024 10551
rect 20070 10520 20076 10532
rect 16080 10492 20076 10520
rect 16080 10480 16086 10492
rect 20070 10480 20076 10492
rect 20128 10480 20134 10532
rect 17862 10452 17868 10464
rect 15948 10424 17868 10452
rect 13504 10412 13510 10424
rect 17862 10412 17868 10424
rect 17920 10412 17926 10464
rect 19058 10452 19064 10464
rect 19019 10424 19064 10452
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 1104 10362 30820 10384
rect 1104 10310 5915 10362
rect 5967 10310 5979 10362
rect 6031 10310 6043 10362
rect 6095 10310 6107 10362
rect 6159 10310 6171 10362
rect 6223 10310 15846 10362
rect 15898 10310 15910 10362
rect 15962 10310 15974 10362
rect 16026 10310 16038 10362
rect 16090 10310 16102 10362
rect 16154 10310 25776 10362
rect 25828 10310 25840 10362
rect 25892 10310 25904 10362
rect 25956 10310 25968 10362
rect 26020 10310 26032 10362
rect 26084 10310 30820 10362
rect 1104 10288 30820 10310
rect 2222 10248 2228 10260
rect 2183 10220 2228 10248
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 9309 10251 9367 10257
rect 9309 10217 9321 10251
rect 9355 10248 9367 10251
rect 9490 10248 9496 10260
rect 9355 10220 9496 10248
rect 9355 10217 9367 10220
rect 9309 10211 9367 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 11606 10248 11612 10260
rect 11567 10220 11612 10248
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 12434 10248 12440 10260
rect 11808 10220 12440 10248
rect 1486 10140 1492 10192
rect 1544 10180 1550 10192
rect 1544 10152 3832 10180
rect 1544 10140 1550 10152
rect 1765 10115 1823 10121
rect 1765 10081 1777 10115
rect 1811 10112 1823 10115
rect 1946 10112 1952 10124
rect 1811 10084 1952 10112
rect 1811 10081 1823 10084
rect 1765 10075 1823 10081
rect 1946 10072 1952 10084
rect 2004 10072 2010 10124
rect 2866 10112 2872 10124
rect 2056 10084 2872 10112
rect 1486 10044 1492 10056
rect 1447 10016 1492 10044
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 2056 10053 2084 10084
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 3804 10121 3832 10152
rect 3789 10115 3847 10121
rect 3789 10081 3801 10115
rect 3835 10081 3847 10115
rect 3789 10075 3847 10081
rect 6273 10115 6331 10121
rect 6273 10081 6285 10115
rect 6319 10112 6331 10115
rect 6638 10112 6644 10124
rect 6319 10084 6644 10112
rect 6319 10081 6331 10084
rect 6273 10075 6331 10081
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 10042 10072 10048 10124
rect 10100 10112 10106 10124
rect 10229 10115 10287 10121
rect 10229 10112 10241 10115
rect 10100 10084 10241 10112
rect 10100 10072 10106 10084
rect 10229 10081 10241 10084
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10013 2099 10047
rect 2041 10007 2099 10013
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10044 2743 10047
rect 2774 10044 2780 10056
rect 2731 10016 2780 10044
rect 2731 10013 2743 10016
rect 2685 10007 2743 10013
rect 1872 9976 1900 10007
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 5810 10004 5816 10056
rect 5868 10044 5874 10056
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 5868 10016 6193 10044
rect 5868 10004 5874 10016
rect 6181 10013 6193 10016
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6370 10025 6428 10031
rect 6370 9991 6382 10025
rect 6416 9991 6428 10025
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 6880 10016 7113 10044
rect 6880 10004 6886 10016
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 10496 10047 10554 10053
rect 7883 10042 9449 10044
rect 9600 10042 10456 10044
rect 7883 10016 10456 10042
rect 7883 10013 7895 10016
rect 9421 10014 9628 10016
rect 7837 10007 7895 10013
rect 1872 9948 2728 9976
rect 2700 9920 2728 9948
rect 3326 9936 3332 9988
rect 3384 9976 3390 9988
rect 4034 9979 4092 9985
rect 4034 9976 4046 9979
rect 3384 9948 4046 9976
rect 3384 9936 3390 9948
rect 4034 9945 4046 9948
rect 4080 9945 4092 9979
rect 5994 9976 6000 9988
rect 5955 9948 6000 9976
rect 4034 9939 4092 9945
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 6370 9985 6428 9991
rect 6273 9979 6331 9985
rect 6273 9945 6285 9979
rect 6319 9945 6331 9979
rect 6273 9939 6331 9945
rect 2682 9868 2688 9920
rect 2740 9868 2746 9920
rect 2866 9908 2872 9920
rect 2827 9880 2872 9908
rect 2866 9868 2872 9880
rect 2924 9868 2930 9920
rect 3142 9868 3148 9920
rect 3200 9908 3206 9920
rect 4982 9908 4988 9920
rect 3200 9880 4988 9908
rect 3200 9868 3206 9880
rect 4982 9868 4988 9880
rect 5040 9908 5046 9920
rect 5169 9911 5227 9917
rect 5169 9908 5181 9911
rect 5040 9880 5181 9908
rect 5040 9868 5046 9880
rect 5169 9877 5181 9880
rect 5215 9877 5227 9911
rect 5169 9871 5227 9877
rect 5258 9868 5264 9920
rect 5316 9908 5322 9920
rect 6288 9908 6316 9939
rect 5316 9880 6316 9908
rect 6380 9908 6408 9985
rect 6917 9979 6975 9985
rect 6917 9976 6929 9979
rect 6564 9948 6929 9976
rect 6454 9908 6460 9920
rect 6380 9880 6460 9908
rect 5316 9868 5322 9880
rect 6454 9868 6460 9880
rect 6512 9908 6518 9920
rect 6564 9908 6592 9948
rect 6917 9945 6929 9948
rect 6963 9945 6975 9979
rect 7650 9976 7656 9988
rect 7611 9948 7656 9976
rect 6917 9939 6975 9945
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 9493 9979 9551 9985
rect 9493 9945 9505 9979
rect 9539 9945 9551 9979
rect 9674 9976 9680 9988
rect 9635 9948 9680 9976
rect 9493 9939 9551 9945
rect 6512 9880 6592 9908
rect 9508 9908 9536 9939
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 10428 9976 10456 10016
rect 10496 10013 10508 10047
rect 10542 10044 10554 10047
rect 10870 10044 10876 10056
rect 10542 10016 10876 10044
rect 10542 10013 10554 10016
rect 10496 10007 10554 10013
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 11808 10044 11836 10220
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 13446 10248 13452 10260
rect 12768 10220 13452 10248
rect 12768 10208 12774 10220
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 17494 10248 17500 10260
rect 13556 10220 15148 10248
rect 17455 10220 17500 10248
rect 11882 10072 11888 10124
rect 11940 10112 11946 10124
rect 11940 10084 12204 10112
rect 11940 10072 11946 10084
rect 12069 10047 12127 10053
rect 12069 10044 12081 10047
rect 11808 10016 12081 10044
rect 12069 10013 12081 10016
rect 12115 10013 12127 10047
rect 12069 10007 12127 10013
rect 12176 10038 12204 10084
rect 12325 10047 12383 10053
rect 12325 10044 12337 10047
rect 12268 10038 12337 10044
rect 12176 10016 12337 10038
rect 12176 10010 12296 10016
rect 12325 10013 12337 10016
rect 12371 10013 12383 10047
rect 12325 10007 12383 10013
rect 12618 9976 12624 9988
rect 10428 9948 12624 9976
rect 12618 9936 12624 9948
rect 12676 9936 12682 9988
rect 13556 9976 13584 10220
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14458 10112 14464 10124
rect 14056 10084 14464 10112
rect 14056 10072 14062 10084
rect 14458 10072 14464 10084
rect 14516 10072 14522 10124
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13964 10016 14105 10044
rect 13964 10004 13970 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 13464 9948 13584 9976
rect 10226 9908 10232 9920
rect 9508 9880 10232 9908
rect 6512 9868 6518 9880
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 11606 9868 11612 9920
rect 11664 9908 11670 9920
rect 13464 9908 13492 9948
rect 11664 9880 13492 9908
rect 11664 9868 11670 9880
rect 13538 9868 13544 9920
rect 13596 9908 13602 9920
rect 14292 9908 14320 10007
rect 14366 10004 14372 10056
rect 14424 10044 14430 10056
rect 14642 10044 14648 10056
rect 14424 10016 14469 10044
rect 14603 10016 14648 10044
rect 14424 10004 14430 10016
rect 14642 10004 14648 10016
rect 14700 10044 14706 10056
rect 15010 10044 15016 10056
rect 14700 10016 15016 10044
rect 14700 10004 14706 10016
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 15120 10044 15148 10220
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 19886 10208 19892 10260
rect 19944 10248 19950 10260
rect 20349 10251 20407 10257
rect 20349 10248 20361 10251
rect 19944 10220 20361 10248
rect 19944 10208 19950 10220
rect 20349 10217 20361 10220
rect 20395 10217 20407 10251
rect 28626 10248 28632 10260
rect 20349 10211 20407 10217
rect 20456 10220 28632 10248
rect 18230 10140 18236 10192
rect 18288 10180 18294 10192
rect 18509 10183 18567 10189
rect 18509 10180 18521 10183
rect 18288 10152 18521 10180
rect 18288 10140 18294 10152
rect 18509 10149 18521 10152
rect 18555 10149 18567 10183
rect 18509 10143 18567 10149
rect 16666 10112 16672 10124
rect 16627 10084 16672 10112
rect 16666 10072 16672 10084
rect 16724 10072 16730 10124
rect 17310 10112 17316 10124
rect 16796 10084 17316 10112
rect 16796 10053 16824 10084
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 18690 10112 18696 10124
rect 18340 10084 18696 10112
rect 16577 10047 16635 10053
rect 16577 10044 16589 10047
rect 15120 10016 16589 10044
rect 16577 10013 16589 10016
rect 16623 10013 16635 10047
rect 16577 10007 16635 10013
rect 16781 10047 16839 10053
rect 16781 10013 16793 10047
rect 16827 10013 16839 10047
rect 17402 10044 17408 10056
rect 17363 10016 17408 10044
rect 16781 10007 16839 10013
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 18340 10053 18368 10084
rect 18690 10072 18696 10084
rect 18748 10112 18754 10124
rect 20456 10112 20484 10220
rect 28626 10208 28632 10220
rect 28684 10208 28690 10260
rect 18748 10084 20484 10112
rect 18748 10072 18754 10084
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 18601 10047 18659 10053
rect 18601 10013 18613 10047
rect 18647 10044 18659 10047
rect 18782 10044 18788 10056
rect 18647 10016 18788 10044
rect 18647 10013 18659 10016
rect 18601 10007 18659 10013
rect 18782 10004 18788 10016
rect 18840 10044 18846 10056
rect 19242 10044 19248 10056
rect 18840 10016 19248 10044
rect 18840 10004 18846 10016
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 20441 10047 20499 10053
rect 20441 10013 20453 10047
rect 20487 10044 20499 10047
rect 20714 10044 20720 10056
rect 20487 10016 20720 10044
rect 20487 10013 20499 10016
rect 20441 10007 20499 10013
rect 20714 10004 20720 10016
rect 20772 10004 20778 10056
rect 21818 10004 21824 10056
rect 21876 10044 21882 10056
rect 22465 10047 22523 10053
rect 22465 10044 22477 10047
rect 21876 10016 22477 10044
rect 21876 10004 21882 10016
rect 22465 10013 22477 10016
rect 22511 10013 22523 10047
rect 29822 10044 29828 10056
rect 29783 10016 29828 10044
rect 22465 10007 22523 10013
rect 29822 10004 29828 10016
rect 29880 10004 29886 10056
rect 14550 9936 14556 9988
rect 14608 9976 14614 9988
rect 15381 9979 15439 9985
rect 15381 9976 15393 9979
rect 14608 9948 15393 9976
rect 14608 9936 14614 9948
rect 15381 9945 15393 9948
rect 15427 9945 15439 9979
rect 15562 9976 15568 9988
rect 15523 9948 15568 9976
rect 15381 9939 15439 9945
rect 15562 9936 15568 9948
rect 15620 9936 15626 9988
rect 16390 9976 16396 9988
rect 16351 9948 16396 9976
rect 16390 9936 16396 9948
rect 16448 9936 16454 9988
rect 16669 9979 16727 9985
rect 16669 9945 16681 9979
rect 16715 9976 16727 9979
rect 22220 9979 22278 9985
rect 16715 9948 21128 9976
rect 16715 9945 16727 9948
rect 16669 9939 16727 9945
rect 14826 9908 14832 9920
rect 13596 9880 14320 9908
rect 14787 9880 14832 9908
rect 13596 9868 13602 9880
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 18138 9908 18144 9920
rect 18099 9880 18144 9908
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 21100 9917 21128 9948
rect 22220 9945 22232 9979
rect 22266 9976 22278 9979
rect 22554 9976 22560 9988
rect 22266 9948 22560 9976
rect 22266 9945 22278 9948
rect 22220 9939 22278 9945
rect 22554 9936 22560 9948
rect 22612 9936 22618 9988
rect 21085 9911 21143 9917
rect 21085 9877 21097 9911
rect 21131 9908 21143 9911
rect 21266 9908 21272 9920
rect 21131 9880 21272 9908
rect 21131 9877 21143 9880
rect 21085 9871 21143 9877
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 30006 9908 30012 9920
rect 29967 9880 30012 9908
rect 30006 9868 30012 9880
rect 30064 9868 30070 9920
rect 1104 9818 30820 9840
rect 1104 9766 10880 9818
rect 10932 9766 10944 9818
rect 10996 9766 11008 9818
rect 11060 9766 11072 9818
rect 11124 9766 11136 9818
rect 11188 9766 20811 9818
rect 20863 9766 20875 9818
rect 20927 9766 20939 9818
rect 20991 9766 21003 9818
rect 21055 9766 21067 9818
rect 21119 9766 30820 9818
rect 1104 9744 30820 9766
rect 3326 9704 3332 9716
rect 3287 9676 3332 9704
rect 3326 9664 3332 9676
rect 3384 9664 3390 9716
rect 4430 9664 4436 9716
rect 4488 9664 4494 9716
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6052 9676 6960 9704
rect 6052 9664 6058 9676
rect 2866 9636 2872 9648
rect 2792 9608 2872 9636
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 1486 9528 1492 9580
rect 1544 9568 1550 9580
rect 2314 9568 2320 9580
rect 1544 9540 2320 9568
rect 1544 9528 1550 9540
rect 2314 9528 2320 9540
rect 2372 9568 2378 9580
rect 2792 9577 2820 9608
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 2593 9571 2651 9577
rect 2593 9568 2605 9571
rect 2372 9540 2605 9568
rect 2372 9528 2378 9540
rect 2593 9537 2605 9540
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9537 2835 9571
rect 3142 9568 3148 9580
rect 3103 9540 3148 9568
rect 2777 9531 2835 9537
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 3510 9528 3516 9580
rect 3568 9568 3574 9580
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 3568 9540 4077 9568
rect 3568 9528 3574 9540
rect 4065 9537 4077 9540
rect 4111 9537 4123 9571
rect 4246 9568 4252 9580
rect 4207 9540 4252 9568
rect 4065 9531 4123 9537
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 4448 9577 4476 9664
rect 6932 9645 6960 9676
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 12342 9704 12348 9716
rect 10560 9676 12348 9704
rect 10560 9664 10566 9676
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 14458 9664 14464 9716
rect 14516 9704 14522 9716
rect 14516 9676 15056 9704
rect 14516 9664 14522 9676
rect 6917 9639 6975 9645
rect 6917 9636 6929 9639
rect 6827 9608 6929 9636
rect 6917 9605 6929 9608
rect 6963 9636 6975 9639
rect 7650 9636 7656 9648
rect 6963 9608 7656 9636
rect 6963 9605 6975 9608
rect 6917 9599 6975 9605
rect 6544 9593 6602 9599
rect 7650 9596 7656 9608
rect 7708 9596 7714 9648
rect 10689 9639 10747 9645
rect 10689 9605 10701 9639
rect 10735 9636 10747 9639
rect 10778 9636 10784 9648
rect 10735 9608 10784 9636
rect 10735 9605 10747 9608
rect 10689 9599 10747 9605
rect 10778 9596 10784 9608
rect 10836 9596 10842 9648
rect 10873 9639 10931 9645
rect 10873 9605 10885 9639
rect 10919 9636 10931 9639
rect 13170 9636 13176 9648
rect 10919 9608 13176 9636
rect 10919 9605 10931 9608
rect 10873 9599 10931 9605
rect 13170 9596 13176 9608
rect 13228 9596 13234 9648
rect 13262 9596 13268 9648
rect 13320 9636 13326 9648
rect 13906 9636 13912 9648
rect 13320 9608 13912 9636
rect 13320 9596 13326 9608
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 14032 9639 14090 9645
rect 14032 9605 14044 9639
rect 14078 9636 14090 9639
rect 14734 9636 14740 9648
rect 14078 9608 14740 9636
rect 14078 9605 14090 9608
rect 14032 9599 14090 9605
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 4798 9568 4804 9580
rect 4663 9540 4804 9568
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 4798 9528 4804 9540
rect 4856 9568 4862 9580
rect 5350 9568 5356 9580
rect 4856 9540 5356 9568
rect 4856 9528 4862 9540
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 5442 9528 5448 9580
rect 5500 9568 5506 9580
rect 5500 9540 5545 9568
rect 6544 9559 6556 9593
rect 6590 9559 6602 9593
rect 6544 9553 6602 9559
rect 6641 9571 6699 9577
rect 5500 9528 5506 9540
rect 2869 9503 2927 9509
rect 2869 9500 2881 9503
rect 2608 9472 2881 9500
rect 2608 9444 2636 9472
rect 2869 9469 2881 9472
rect 2915 9469 2927 9503
rect 2869 9463 2927 9469
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9469 3019 9503
rect 2961 9463 3019 9469
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 2590 9392 2596 9444
rect 2648 9392 2654 9444
rect 2682 9392 2688 9444
rect 2740 9432 2746 9444
rect 2976 9432 3004 9463
rect 2740 9404 3004 9432
rect 2740 9392 2746 9404
rect 4246 9392 4252 9444
rect 4304 9432 4310 9444
rect 4356 9432 4384 9463
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 5132 9472 5273 9500
rect 5132 9460 5138 9472
rect 5261 9469 5273 9472
rect 5307 9469 5319 9503
rect 5261 9463 5319 9469
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 6559 9500 6587 9553
rect 6641 9537 6653 9571
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9568 6791 9571
rect 6822 9568 6828 9580
rect 6779 9540 6828 9568
rect 6779 9537 6791 9540
rect 6733 9531 6791 9537
rect 6512 9472 6587 9500
rect 6512 9460 6518 9472
rect 6656 9432 6684 9531
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 7466 9528 7472 9580
rect 7524 9568 7530 9580
rect 8938 9568 8944 9580
rect 7524 9540 8944 9568
rect 7524 9528 7530 9540
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9548 9540 9965 9568
rect 9548 9528 9554 9540
rect 9953 9537 9965 9540
rect 9999 9568 10011 9571
rect 10042 9568 10048 9580
rect 9999 9540 10048 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 14910 9571 14968 9577
rect 14910 9568 14922 9571
rect 14844 9540 14922 9568
rect 8294 9500 8300 9512
rect 8255 9472 8300 9500
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 9674 9500 9680 9512
rect 8619 9472 9680 9500
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 12161 9503 12219 9509
rect 12161 9469 12173 9503
rect 12207 9469 12219 9503
rect 12161 9463 12219 9469
rect 4304 9404 4384 9432
rect 4448 9404 6684 9432
rect 4304 9392 4310 9404
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 2498 9364 2504 9376
rect 1627 9336 2504 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 4448 9364 4476 9404
rect 6730 9392 6736 9444
rect 6788 9432 6794 9444
rect 6917 9435 6975 9441
rect 6917 9432 6929 9435
rect 6788 9404 6929 9432
rect 6788 9392 6794 9404
rect 6917 9401 6929 9404
rect 6963 9401 6975 9435
rect 12176 9432 12204 9463
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 12434 9500 12440 9512
rect 12400 9472 12440 9500
rect 12400 9460 12406 9472
rect 12434 9460 12440 9472
rect 12492 9500 12498 9512
rect 14277 9503 14335 9509
rect 12492 9472 12537 9500
rect 12492 9460 12498 9472
rect 14277 9469 14289 9503
rect 14323 9500 14335 9503
rect 14550 9500 14556 9512
rect 14323 9472 14556 9500
rect 14323 9469 14335 9472
rect 14277 9463 14335 9469
rect 14550 9460 14556 9472
rect 14608 9460 14614 9512
rect 14844 9500 14872 9540
rect 14910 9537 14922 9540
rect 14956 9537 14968 9571
rect 15028 9568 15056 9676
rect 15286 9674 15292 9716
rect 15212 9664 15292 9674
rect 15344 9664 15350 9716
rect 18414 9704 18420 9716
rect 15948 9676 16160 9704
rect 15212 9646 15332 9664
rect 15105 9571 15163 9577
rect 15105 9568 15117 9571
rect 15028 9540 15117 9568
rect 14910 9531 14968 9537
rect 15105 9537 15117 9540
rect 15151 9537 15163 9571
rect 15212 9570 15240 9646
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 15948 9636 15976 9676
rect 15712 9608 15976 9636
rect 16132 9636 16160 9676
rect 17788 9676 18420 9704
rect 17788 9636 17816 9676
rect 18414 9664 18420 9676
rect 18472 9664 18478 9716
rect 19242 9704 19248 9716
rect 19203 9676 19248 9704
rect 19242 9664 19248 9676
rect 19300 9664 19306 9716
rect 19797 9707 19855 9713
rect 19797 9673 19809 9707
rect 19843 9704 19855 9707
rect 20254 9704 20260 9716
rect 19843 9676 20260 9704
rect 19843 9673 19855 9676
rect 19797 9667 19855 9673
rect 20254 9664 20260 9676
rect 20312 9664 20318 9716
rect 16132 9608 17816 9636
rect 17880 9608 20944 9636
rect 15712 9596 15718 9608
rect 15289 9571 15347 9577
rect 15289 9570 15301 9571
rect 15212 9542 15301 9570
rect 15105 9531 15163 9537
rect 15289 9537 15301 9542
rect 15335 9537 15347 9571
rect 15470 9568 15476 9580
rect 15431 9540 15476 9568
rect 15289 9531 15347 9537
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 15925 9571 15983 9577
rect 15925 9568 15937 9571
rect 15764 9540 15937 9568
rect 15197 9503 15255 9509
rect 14844 9472 14964 9500
rect 13262 9432 13268 9444
rect 12176 9404 13268 9432
rect 6917 9395 6975 9401
rect 13262 9392 13268 9404
rect 13320 9392 13326 9444
rect 2832 9336 4476 9364
rect 2832 9324 2838 9336
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 4801 9367 4859 9373
rect 4801 9364 4813 9367
rect 4672 9336 4813 9364
rect 4672 9324 4678 9336
rect 4801 9333 4813 9336
rect 4847 9333 4859 9367
rect 4801 9327 4859 9333
rect 4982 9324 4988 9376
rect 5040 9364 5046 9376
rect 8662 9364 8668 9376
rect 5040 9336 8668 9364
rect 5040 9324 5046 9336
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 14642 9364 14648 9376
rect 12943 9336 14648 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 14737 9367 14795 9373
rect 14737 9333 14749 9367
rect 14783 9364 14795 9367
rect 14826 9364 14832 9376
rect 14783 9336 14832 9364
rect 14783 9333 14795 9336
rect 14737 9327 14795 9333
rect 14826 9324 14832 9336
rect 14884 9324 14890 9376
rect 14936 9364 14964 9472
rect 15197 9469 15209 9503
rect 15243 9500 15255 9503
rect 15654 9500 15660 9512
rect 15243 9472 15660 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 15654 9460 15660 9472
rect 15712 9460 15718 9512
rect 15102 9392 15108 9444
rect 15160 9432 15166 9444
rect 15764 9432 15792 9540
rect 15925 9537 15937 9540
rect 15971 9537 15983 9571
rect 15925 9531 15983 9537
rect 16025 9503 16083 9509
rect 16025 9469 16037 9503
rect 16071 9500 16083 9503
rect 16942 9500 16948 9512
rect 16071 9472 16948 9500
rect 16071 9469 16083 9472
rect 16025 9463 16083 9469
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17034 9460 17040 9512
rect 17092 9500 17098 9512
rect 17880 9509 17908 9608
rect 18138 9577 18144 9580
rect 18132 9568 18144 9577
rect 18099 9540 18144 9568
rect 18132 9531 18144 9540
rect 18138 9528 18144 9531
rect 18196 9528 18202 9580
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9537 19763 9571
rect 19705 9531 19763 9537
rect 17865 9503 17923 9509
rect 17865 9500 17877 9503
rect 17092 9472 17877 9500
rect 17092 9460 17098 9472
rect 17865 9469 17877 9472
rect 17911 9469 17923 9503
rect 17865 9463 17923 9469
rect 15160 9404 15792 9432
rect 15160 9392 15166 9404
rect 16206 9364 16212 9376
rect 14936 9336 16212 9364
rect 16206 9324 16212 9336
rect 16264 9364 16270 9376
rect 19720 9364 19748 9531
rect 20916 9500 20944 9608
rect 21910 9528 21916 9580
rect 21968 9568 21974 9580
rect 22077 9571 22135 9577
rect 22077 9568 22089 9571
rect 21968 9540 22089 9568
rect 21968 9528 21974 9540
rect 22077 9537 22089 9540
rect 22123 9537 22135 9571
rect 22077 9531 22135 9537
rect 21818 9500 21824 9512
rect 20916 9472 21824 9500
rect 21818 9460 21824 9472
rect 21876 9460 21882 9512
rect 16264 9336 19748 9364
rect 16264 9324 16270 9336
rect 22002 9324 22008 9376
rect 22060 9364 22066 9376
rect 23201 9367 23259 9373
rect 23201 9364 23213 9367
rect 22060 9336 23213 9364
rect 22060 9324 22066 9336
rect 23201 9333 23213 9336
rect 23247 9333 23259 9367
rect 23201 9327 23259 9333
rect 1104 9274 30820 9296
rect 1104 9222 5915 9274
rect 5967 9222 5979 9274
rect 6031 9222 6043 9274
rect 6095 9222 6107 9274
rect 6159 9222 6171 9274
rect 6223 9222 15846 9274
rect 15898 9222 15910 9274
rect 15962 9222 15974 9274
rect 16026 9222 16038 9274
rect 16090 9222 16102 9274
rect 16154 9222 25776 9274
rect 25828 9222 25840 9274
rect 25892 9222 25904 9274
rect 25956 9222 25968 9274
rect 26020 9222 26032 9274
rect 26084 9222 30820 9274
rect 1104 9200 30820 9222
rect 5169 9163 5227 9169
rect 5169 9160 5181 9163
rect 2884 9132 5181 9160
rect 2682 9024 2688 9036
rect 2643 8996 2688 9024
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 2314 8956 2320 8968
rect 2275 8928 2320 8956
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 2498 8956 2504 8968
rect 2459 8928 2504 8956
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 2884 8965 2912 9132
rect 5169 9129 5181 9132
rect 5215 9160 5227 9163
rect 5258 9160 5264 9172
rect 5215 9132 5264 9160
rect 5215 9129 5227 9132
rect 5169 9123 5227 9129
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 6822 9160 6828 9172
rect 6783 9132 6828 9160
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 9674 9160 9680 9172
rect 9635 9132 9680 9160
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10226 9160 10232 9172
rect 10187 9132 10232 9160
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 12912 9132 16620 9160
rect 3602 8984 3608 9036
rect 3660 9024 3666 9036
rect 9217 9027 9275 9033
rect 3660 8996 3924 9024
rect 3660 8984 3666 8996
rect 2869 8959 2927 8965
rect 2648 8928 2693 8956
rect 2648 8916 2654 8928
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 3896 8956 3924 8996
rect 8128 8996 9168 9024
rect 8128 8956 8156 8996
rect 3896 8928 8156 8956
rect 8205 8959 8263 8965
rect 3789 8919 3847 8925
rect 8205 8925 8217 8959
rect 8251 8956 8263 8959
rect 8294 8956 8300 8968
rect 8251 8928 8300 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 1486 8848 1492 8900
rect 1544 8888 1550 8900
rect 3804 8888 3832 8919
rect 8294 8916 8300 8928
rect 8352 8956 8358 8968
rect 8662 8956 8668 8968
rect 8352 8928 8668 8956
rect 8352 8916 8358 8928
rect 8662 8916 8668 8928
rect 8720 8916 8726 8968
rect 8938 8956 8944 8968
rect 8899 8928 8944 8956
rect 8938 8916 8944 8928
rect 8996 8916 9002 8968
rect 9140 8965 9168 8996
rect 9217 8993 9229 9027
rect 9263 9024 9275 9027
rect 9674 9024 9680 9036
rect 9263 8996 9680 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 10226 8984 10232 9036
rect 10284 9024 10290 9036
rect 10284 8996 11468 9024
rect 10284 8984 10290 8996
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8925 9367 8959
rect 9490 8956 9496 8968
rect 9451 8928 9496 8956
rect 9309 8919 9367 8925
rect 3878 8888 3884 8900
rect 1544 8860 3884 8888
rect 1544 8848 1550 8860
rect 3878 8848 3884 8860
rect 3936 8848 3942 8900
rect 4045 8891 4103 8897
rect 4045 8888 4057 8891
rect 3988 8860 4057 8888
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 1670 8820 1676 8832
rect 1627 8792 1676 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 3053 8823 3111 8829
rect 3053 8789 3065 8823
rect 3099 8820 3111 8823
rect 3988 8820 4016 8860
rect 4045 8857 4057 8860
rect 4091 8857 4103 8891
rect 4045 8851 4103 8857
rect 4338 8848 4344 8900
rect 4396 8888 4402 8900
rect 4982 8888 4988 8900
rect 4396 8860 4988 8888
rect 4396 8848 4402 8860
rect 4982 8848 4988 8860
rect 5040 8848 5046 8900
rect 5442 8848 5448 8900
rect 5500 8888 5506 8900
rect 5813 8891 5871 8897
rect 5813 8888 5825 8891
rect 5500 8860 5825 8888
rect 5500 8848 5506 8860
rect 5813 8857 5825 8860
rect 5859 8857 5871 8891
rect 5813 8851 5871 8857
rect 6362 8848 6368 8900
rect 6420 8888 6426 8900
rect 6638 8888 6644 8900
rect 6420 8860 6644 8888
rect 6420 8848 6426 8860
rect 6638 8848 6644 8860
rect 6696 8848 6702 8900
rect 7190 8848 7196 8900
rect 7248 8888 7254 8900
rect 7938 8891 7996 8897
rect 7938 8888 7950 8891
rect 7248 8860 7950 8888
rect 7248 8848 7254 8860
rect 7938 8857 7950 8860
rect 7984 8857 7996 8891
rect 7938 8851 7996 8857
rect 9214 8848 9220 8900
rect 9272 8888 9278 8900
rect 9324 8888 9352 8919
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 10134 8956 10140 8968
rect 10095 8928 10140 8956
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 11440 8965 11468 8996
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12713 9027 12771 9033
rect 12713 9024 12725 9027
rect 12492 8996 12725 9024
rect 12492 8984 12498 8996
rect 12713 8993 12725 8996
rect 12759 8993 12771 9027
rect 12713 8987 12771 8993
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10560 8928 10977 8956
rect 10560 8916 10566 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8925 11483 8959
rect 11606 8956 11612 8968
rect 11567 8928 11612 8956
rect 11425 8919 11483 8925
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 12912 8956 12940 9132
rect 16117 9095 16175 9101
rect 16117 9092 16129 9095
rect 15304 9064 16129 9092
rect 12406 8928 12940 8956
rect 12989 8959 13047 8965
rect 12406 8888 12434 8928
rect 12989 8925 13001 8959
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8956 14335 8959
rect 14366 8956 14372 8968
rect 14323 8928 14372 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 9272 8860 12434 8888
rect 9272 8848 9278 8860
rect 3099 8792 4016 8820
rect 5721 8823 5779 8829
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 5721 8789 5733 8823
rect 5767 8820 5779 8823
rect 6730 8820 6736 8832
rect 5767 8792 6736 8820
rect 5767 8789 5779 8792
rect 5721 8783 5779 8789
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7374 8820 7380 8832
rect 6972 8792 7380 8820
rect 6972 8780 6978 8792
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 10873 8823 10931 8829
rect 10873 8820 10885 8823
rect 10836 8792 10885 8820
rect 10836 8780 10842 8792
rect 10873 8789 10885 8792
rect 10919 8789 10931 8823
rect 11514 8820 11520 8832
rect 11475 8792 11520 8820
rect 10873 8783 10931 8789
rect 11514 8780 11520 8792
rect 11572 8780 11578 8832
rect 13004 8820 13032 8919
rect 14366 8916 14372 8928
rect 14424 8956 14430 8968
rect 15304 8958 15332 9064
rect 16117 9061 16129 9064
rect 16163 9061 16175 9095
rect 16592 9092 16620 9132
rect 16666 9120 16672 9172
rect 16724 9160 16730 9172
rect 19061 9163 19119 9169
rect 19061 9160 19073 9163
rect 16724 9132 19073 9160
rect 16724 9120 16730 9132
rect 19061 9129 19073 9132
rect 19107 9129 19119 9163
rect 19061 9123 19119 9129
rect 19613 9163 19671 9169
rect 19613 9129 19625 9163
rect 19659 9160 19671 9163
rect 20162 9160 20168 9172
rect 19659 9132 20168 9160
rect 19659 9129 19671 9132
rect 19613 9123 19671 9129
rect 20162 9120 20168 9132
rect 20220 9120 20226 9172
rect 20257 9163 20315 9169
rect 20257 9129 20269 9163
rect 20303 9160 20315 9163
rect 20346 9160 20352 9172
rect 20303 9132 20352 9160
rect 20303 9129 20315 9132
rect 20257 9123 20315 9129
rect 20346 9120 20352 9132
rect 20404 9120 20410 9172
rect 21910 9160 21916 9172
rect 21871 9132 21916 9160
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 17770 9092 17776 9104
rect 16592 9064 17776 9092
rect 16117 9055 16175 9061
rect 17770 9052 17776 9064
rect 17828 9052 17834 9104
rect 17862 9052 17868 9104
rect 17920 9092 17926 9104
rect 22002 9092 22008 9104
rect 17920 9064 22008 9092
rect 17920 9052 17926 9064
rect 19242 9024 19248 9036
rect 17972 8996 19248 9024
rect 17972 8968 18000 8996
rect 19242 8984 19248 8996
rect 19300 9024 19306 9036
rect 21453 9027 21511 9033
rect 19300 8996 21220 9024
rect 19300 8984 19306 8996
rect 15212 8956 15332 8958
rect 14424 8930 15332 8956
rect 14424 8928 15240 8930
rect 14424 8916 14430 8928
rect 15562 8916 15568 8968
rect 15620 8956 15626 8968
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 15620 8928 16313 8956
rect 15620 8916 15626 8928
rect 16301 8925 16313 8928
rect 16347 8956 16359 8959
rect 16945 8959 17003 8965
rect 16945 8956 16957 8959
rect 16347 8928 16957 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 16945 8925 16957 8928
rect 16991 8925 17003 8959
rect 16945 8919 17003 8925
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8956 17923 8959
rect 17954 8956 17960 8968
rect 17911 8928 17960 8956
rect 17911 8925 17923 8928
rect 17865 8919 17923 8925
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 18049 8959 18107 8965
rect 18049 8925 18061 8959
rect 18095 8925 18107 8959
rect 18049 8919 18107 8925
rect 18135 8959 18193 8965
rect 18135 8925 18147 8959
rect 18181 8925 18193 8959
rect 18135 8919 18193 8925
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18322 8956 18328 8968
rect 18279 8928 18328 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 14090 8848 14096 8900
rect 14148 8888 14154 8900
rect 14522 8891 14580 8897
rect 14522 8888 14534 8891
rect 14148 8860 14534 8888
rect 14148 8848 14154 8860
rect 14522 8857 14534 8860
rect 14568 8857 14580 8891
rect 14522 8851 14580 8857
rect 14642 8848 14648 8900
rect 14700 8888 14706 8900
rect 17678 8888 17684 8900
rect 14700 8860 17684 8888
rect 14700 8848 14706 8860
rect 15470 8820 15476 8832
rect 13004 8792 15476 8820
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 15672 8829 15700 8860
rect 17678 8848 17684 8860
rect 17736 8848 17742 8900
rect 15657 8823 15715 8829
rect 15657 8789 15669 8823
rect 15703 8789 15715 8823
rect 17034 8820 17040 8832
rect 16995 8792 17040 8820
rect 15657 8783 15715 8789
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 18064 8820 18092 8919
rect 18156 8888 18184 8919
rect 18322 8916 18328 8928
rect 18380 8916 18386 8968
rect 21192 8965 21220 8996
rect 21453 8993 21465 9027
rect 21499 9024 21511 9027
rect 21634 9024 21640 9036
rect 21499 8996 21640 9024
rect 21499 8993 21511 8996
rect 21453 8987 21511 8993
rect 21634 8984 21640 8996
rect 21692 8984 21698 9036
rect 18417 8959 18475 8965
rect 18417 8925 18429 8959
rect 18463 8925 18475 8959
rect 18417 8919 18475 8925
rect 19061 8959 19119 8965
rect 19061 8925 19073 8959
rect 19107 8956 19119 8959
rect 19521 8959 19579 8965
rect 19521 8956 19533 8959
rect 19107 8928 19533 8956
rect 19107 8925 19119 8928
rect 19061 8919 19119 8925
rect 19521 8925 19533 8928
rect 19567 8925 19579 8959
rect 19521 8919 19579 8925
rect 20165 8959 20223 8965
rect 20165 8925 20177 8959
rect 20211 8925 20223 8959
rect 20165 8919 20223 8925
rect 21177 8959 21235 8965
rect 21177 8925 21189 8959
rect 21223 8925 21235 8959
rect 21177 8919 21235 8925
rect 21361 8959 21419 8965
rect 21361 8925 21373 8959
rect 21407 8925 21419 8959
rect 21542 8956 21548 8968
rect 21503 8928 21548 8956
rect 21361 8919 21419 8925
rect 18156 8860 18276 8888
rect 18248 8832 18276 8860
rect 18432 8832 18460 8919
rect 19150 8848 19156 8900
rect 19208 8888 19214 8900
rect 20180 8888 20208 8919
rect 19208 8860 20208 8888
rect 19208 8848 19214 8860
rect 18138 8820 18144 8832
rect 18064 8792 18144 8820
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 18230 8780 18236 8832
rect 18288 8780 18294 8832
rect 18414 8780 18420 8832
rect 18472 8780 18478 8832
rect 18601 8823 18659 8829
rect 18601 8789 18613 8823
rect 18647 8820 18659 8823
rect 18782 8820 18788 8832
rect 18647 8792 18788 8820
rect 18647 8789 18659 8792
rect 18601 8783 18659 8789
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 21192 8820 21220 8919
rect 21376 8888 21404 8919
rect 21542 8916 21548 8928
rect 21600 8916 21606 8968
rect 21744 8965 21772 9064
rect 22002 9052 22008 9064
rect 22060 9052 22066 9104
rect 21729 8959 21787 8965
rect 21729 8925 21741 8959
rect 21775 8925 21787 8959
rect 21729 8919 21787 8925
rect 22002 8888 22008 8900
rect 21376 8860 22008 8888
rect 22002 8848 22008 8860
rect 22060 8848 22066 8900
rect 21542 8820 21548 8832
rect 21192 8792 21548 8820
rect 21542 8780 21548 8792
rect 21600 8780 21606 8832
rect 1104 8730 30820 8752
rect 1104 8678 10880 8730
rect 10932 8678 10944 8730
rect 10996 8678 11008 8730
rect 11060 8678 11072 8730
rect 11124 8678 11136 8730
rect 11188 8678 20811 8730
rect 20863 8678 20875 8730
rect 20927 8678 20939 8730
rect 20991 8678 21003 8730
rect 21055 8678 21067 8730
rect 21119 8678 30820 8730
rect 1104 8656 30820 8678
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 2832 8588 2877 8616
rect 2832 8576 2838 8588
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 5721 8619 5779 8625
rect 5721 8616 5733 8619
rect 4856 8588 5733 8616
rect 4856 8576 4862 8588
rect 5721 8585 5733 8588
rect 5767 8585 5779 8619
rect 5721 8579 5779 8585
rect 6638 8576 6644 8628
rect 6696 8616 6702 8628
rect 10229 8619 10287 8625
rect 6696 8588 8340 8616
rect 6696 8576 6702 8588
rect 2682 8508 2688 8560
rect 2740 8548 2746 8560
rect 3605 8551 3663 8557
rect 3605 8548 3617 8551
rect 2740 8520 3617 8548
rect 2740 8508 2746 8520
rect 3605 8517 3617 8520
rect 3651 8517 3663 8551
rect 5534 8548 5540 8560
rect 3605 8511 3663 8517
rect 4356 8520 5540 8548
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8480 1455 8483
rect 1486 8480 1492 8492
rect 1443 8452 1492 8480
rect 1443 8449 1455 8452
rect 1397 8443 1455 8449
rect 1486 8440 1492 8452
rect 1544 8440 1550 8492
rect 1664 8483 1722 8489
rect 1664 8449 1676 8483
rect 1710 8480 1722 8483
rect 2222 8480 2228 8492
rect 1710 8452 2228 8480
rect 1710 8449 1722 8452
rect 1664 8443 1722 8449
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 3786 8480 3792 8492
rect 3747 8452 3792 8480
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 4356 8489 4384 8520
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 6880 8520 7052 8548
rect 6880 8508 6886 8520
rect 4614 8489 4620 8492
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 3936 8452 4353 8480
rect 3936 8440 3942 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 4608 8480 4620 8489
rect 4575 8452 4620 8480
rect 4341 8443 4399 8449
rect 4608 8443 4620 8452
rect 4614 8440 4620 8443
rect 4672 8440 4678 8492
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 6457 8483 6515 8489
rect 6457 8480 6469 8483
rect 6328 8452 6469 8480
rect 6328 8440 6334 8452
rect 6457 8449 6469 8452
rect 6503 8449 6515 8483
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 6457 8443 6515 8449
rect 6559 8452 6653 8480
rect 3694 8236 3700 8288
rect 3752 8276 3758 8288
rect 6559 8276 6587 8452
rect 6641 8449 6653 8452
rect 6687 8480 6699 8483
rect 6914 8480 6920 8492
rect 6687 8452 6920 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 7024 8489 7052 8520
rect 7190 8508 7196 8560
rect 7248 8548 7254 8560
rect 7834 8548 7840 8560
rect 7248 8520 7293 8548
rect 7795 8520 7840 8548
rect 7248 8508 7254 8520
rect 7834 8508 7840 8520
rect 7892 8508 7898 8560
rect 8312 8548 8340 8588
rect 10229 8585 10241 8619
rect 10275 8616 10287 8619
rect 10318 8616 10324 8628
rect 10275 8588 10324 8616
rect 10275 8585 10287 8588
rect 10229 8579 10287 8585
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10597 8619 10655 8625
rect 10597 8585 10609 8619
rect 10643 8616 10655 8619
rect 11514 8616 11520 8628
rect 10643 8588 11520 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 14090 8616 14096 8628
rect 11716 8588 12434 8616
rect 14051 8588 14096 8616
rect 8312 8520 11192 8548
rect 7009 8483 7067 8489
rect 7009 8449 7021 8483
rect 7055 8449 7067 8483
rect 8312 8480 8340 8520
rect 8389 8483 8447 8489
rect 8389 8480 8401 8483
rect 8312 8452 8401 8480
rect 7009 8443 7067 8449
rect 8389 8449 8401 8452
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 8536 8452 8677 8480
rect 8536 8440 8542 8452
rect 8665 8449 8677 8452
rect 8711 8480 8723 8483
rect 8938 8480 8944 8492
rect 8711 8452 8944 8480
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 11164 8480 11192 8520
rect 11716 8480 11744 8588
rect 11790 8508 11796 8560
rect 11848 8548 11854 8560
rect 11977 8551 12035 8557
rect 11977 8548 11989 8551
rect 11848 8520 11989 8548
rect 11848 8508 11854 8520
rect 11977 8517 11989 8520
rect 12023 8517 12035 8551
rect 12406 8548 12434 8588
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 16850 8616 16856 8628
rect 14476 8588 16856 8616
rect 14476 8548 14504 8588
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 19610 8616 19616 8628
rect 18196 8588 19616 8616
rect 18196 8576 18202 8588
rect 19610 8576 19616 8588
rect 19668 8616 19674 8628
rect 19889 8619 19947 8625
rect 19889 8616 19901 8619
rect 19668 8588 19901 8616
rect 19668 8576 19674 8588
rect 19889 8585 19901 8588
rect 19935 8585 19947 8619
rect 22554 8616 22560 8628
rect 22515 8588 22560 8616
rect 19889 8579 19947 8585
rect 22554 8576 22560 8588
rect 22612 8576 22618 8628
rect 12406 8520 14504 8548
rect 11977 8511 12035 8517
rect 14550 8508 14556 8560
rect 14608 8548 14614 8560
rect 17034 8548 17040 8560
rect 14608 8520 17040 8548
rect 14608 8508 14614 8520
rect 11882 8480 11888 8492
rect 11164 8452 11744 8480
rect 11843 8452 11888 8480
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 13357 8483 13415 8489
rect 13357 8480 13369 8483
rect 13320 8452 13369 8480
rect 13320 8440 13326 8452
rect 13357 8449 13369 8452
rect 13403 8449 13415 8483
rect 13357 8443 13415 8449
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8480 13599 8483
rect 13814 8480 13820 8492
rect 13587 8452 13820 8480
rect 13587 8449 13599 8452
rect 13541 8443 13599 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8480 13967 8483
rect 14642 8480 14648 8492
rect 13955 8452 14648 8480
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 14826 8489 14832 8492
rect 14820 8480 14832 8489
rect 14787 8452 14832 8480
rect 14820 8443 14832 8452
rect 14826 8440 14832 8443
rect 14884 8440 14890 8492
rect 16684 8489 16712 8520
rect 17034 8508 17040 8520
rect 17092 8508 17098 8560
rect 21266 8508 21272 8560
rect 21324 8548 21330 8560
rect 21324 8520 22416 8548
rect 21324 8508 21330 8520
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 16925 8483 16983 8489
rect 16925 8480 16937 8483
rect 16816 8452 16937 8480
rect 16816 8440 16822 8452
rect 16925 8449 16937 8452
rect 16971 8449 16983 8483
rect 17052 8480 17080 8508
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 17052 8452 18521 8480
rect 16925 8443 16983 8449
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18782 8480 18788 8492
rect 18743 8452 18788 8480
rect 18509 8443 18567 8449
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 21542 8440 21548 8492
rect 21600 8480 21606 8492
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21600 8452 21833 8480
rect 21600 8440 21606 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 22005 8483 22063 8489
rect 22005 8449 22017 8483
rect 22051 8480 22063 8483
rect 22278 8480 22284 8492
rect 22051 8452 22284 8480
rect 22051 8449 22063 8452
rect 22005 8443 22063 8449
rect 22278 8440 22284 8452
rect 22336 8440 22342 8492
rect 22388 8489 22416 8520
rect 22373 8483 22431 8489
rect 22373 8449 22385 8483
rect 22419 8449 22431 8483
rect 22373 8443 22431 8449
rect 29638 8440 29644 8492
rect 29696 8480 29702 8492
rect 29825 8483 29883 8489
rect 29825 8480 29837 8483
rect 29696 8452 29837 8480
rect 29696 8440 29702 8452
rect 29825 8449 29837 8452
rect 29871 8449 29883 8483
rect 29825 8443 29883 8449
rect 6733 8415 6791 8421
rect 6733 8381 6745 8415
rect 6779 8381 6791 8415
rect 6733 8375 6791 8381
rect 6748 8344 6776 8375
rect 6822 8372 6828 8424
rect 6880 8412 6886 8424
rect 6880 8384 6925 8412
rect 6880 8372 6886 8384
rect 10134 8372 10140 8424
rect 10192 8412 10198 8424
rect 10318 8412 10324 8424
rect 10192 8384 10324 8412
rect 10192 8372 10198 8384
rect 10318 8372 10324 8384
rect 10376 8412 10382 8424
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 10376 8384 10701 8412
rect 10376 8372 10382 8384
rect 10689 8381 10701 8384
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 10873 8415 10931 8421
rect 10873 8381 10885 8415
rect 10919 8412 10931 8415
rect 12066 8412 12072 8424
rect 10919 8384 12072 8412
rect 10919 8381 10931 8384
rect 10873 8375 10931 8381
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 13633 8415 13691 8421
rect 13633 8381 13645 8415
rect 13679 8381 13691 8415
rect 13633 8375 13691 8381
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8412 13783 8415
rect 14458 8412 14464 8424
rect 13771 8384 14464 8412
rect 13771 8381 13783 8384
rect 13725 8375 13783 8381
rect 7650 8344 7656 8356
rect 6748 8316 6868 8344
rect 7611 8316 7656 8344
rect 6840 8288 6868 8316
rect 7650 8304 7656 8316
rect 7708 8304 7714 8356
rect 11330 8304 11336 8356
rect 11388 8344 11394 8356
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 11388 8316 11529 8344
rect 11388 8304 11394 8316
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 3752 8248 6587 8276
rect 3752 8236 3758 8248
rect 6822 8236 6828 8288
rect 6880 8236 6886 8288
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 10410 8276 10416 8288
rect 7064 8248 10416 8276
rect 7064 8236 7070 8248
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 10686 8236 10692 8288
rect 10744 8276 10750 8288
rect 10962 8276 10968 8288
rect 10744 8248 10968 8276
rect 10744 8236 10750 8248
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 13648 8276 13676 8375
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 14608 8384 14653 8412
rect 14608 8372 14614 8384
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 21450 8412 21456 8424
rect 17828 8384 21456 8412
rect 17828 8372 17834 8384
rect 21450 8372 21456 8384
rect 21508 8372 21514 8424
rect 21634 8372 21640 8424
rect 21692 8412 21698 8424
rect 21910 8412 21916 8424
rect 21692 8384 21916 8412
rect 21692 8372 21698 8384
rect 21910 8372 21916 8384
rect 21968 8412 21974 8424
rect 22097 8415 22155 8421
rect 22097 8412 22109 8415
rect 21968 8384 22109 8412
rect 21968 8372 21974 8384
rect 22097 8381 22109 8384
rect 22143 8381 22155 8415
rect 22097 8375 22155 8381
rect 22189 8415 22247 8421
rect 22189 8381 22201 8415
rect 22235 8381 22247 8415
rect 22189 8375 22247 8381
rect 15933 8347 15991 8353
rect 15933 8313 15945 8347
rect 15979 8344 15991 8347
rect 16206 8344 16212 8356
rect 15979 8316 16212 8344
rect 15979 8313 15991 8316
rect 15933 8307 15991 8313
rect 16206 8304 16212 8316
rect 16264 8304 16270 8356
rect 21468 8344 21496 8372
rect 22204 8344 22232 8375
rect 30006 8344 30012 8356
rect 21468 8316 22232 8344
rect 29967 8316 30012 8344
rect 30006 8304 30012 8316
rect 30064 8304 30070 8356
rect 15654 8276 15660 8288
rect 13648 8248 15660 8276
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 16482 8236 16488 8288
rect 16540 8276 16546 8288
rect 18049 8279 18107 8285
rect 18049 8276 18061 8279
rect 16540 8248 18061 8276
rect 16540 8236 16546 8248
rect 18049 8245 18061 8248
rect 18095 8276 18107 8279
rect 19150 8276 19156 8288
rect 18095 8248 19156 8276
rect 18095 8245 18107 8248
rect 18049 8239 18107 8245
rect 19150 8236 19156 8248
rect 19208 8236 19214 8288
rect 1104 8186 30820 8208
rect 1104 8134 5915 8186
rect 5967 8134 5979 8186
rect 6031 8134 6043 8186
rect 6095 8134 6107 8186
rect 6159 8134 6171 8186
rect 6223 8134 15846 8186
rect 15898 8134 15910 8186
rect 15962 8134 15974 8186
rect 16026 8134 16038 8186
rect 16090 8134 16102 8186
rect 16154 8134 25776 8186
rect 25828 8134 25840 8186
rect 25892 8134 25904 8186
rect 25956 8134 25968 8186
rect 26020 8134 26032 8186
rect 26084 8134 30820 8186
rect 1104 8112 30820 8134
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 2314 8072 2320 8084
rect 1636 8044 2320 8072
rect 1636 8032 1642 8044
rect 2314 8032 2320 8044
rect 2372 8072 2378 8084
rect 2639 8075 2697 8081
rect 2639 8072 2651 8075
rect 2372 8044 2651 8072
rect 2372 8032 2378 8044
rect 2639 8041 2651 8044
rect 2685 8041 2697 8075
rect 2639 8035 2697 8041
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8904 8044 9045 8072
rect 8904 8032 8910 8044
rect 9033 8041 9045 8044
rect 9079 8041 9091 8075
rect 9033 8035 9091 8041
rect 9401 8075 9459 8081
rect 9401 8041 9413 8075
rect 9447 8072 9459 8075
rect 10321 8075 10379 8081
rect 10321 8072 10333 8075
rect 9447 8044 10333 8072
rect 9447 8041 9459 8044
rect 9401 8035 9459 8041
rect 10321 8041 10333 8044
rect 10367 8072 10379 8075
rect 10781 8075 10839 8081
rect 10781 8072 10793 8075
rect 10367 8044 10793 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 10781 8041 10793 8044
rect 10827 8041 10839 8075
rect 10781 8035 10839 8041
rect 12529 8075 12587 8081
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 13354 8072 13360 8084
rect 12575 8044 13360 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 16393 8075 16451 8081
rect 16393 8041 16405 8075
rect 16439 8072 16451 8075
rect 16758 8072 16764 8084
rect 16439 8044 16764 8072
rect 16439 8041 16451 8044
rect 16393 8035 16451 8041
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 21085 8075 21143 8081
rect 21085 8041 21097 8075
rect 21131 8072 21143 8075
rect 21174 8072 21180 8084
rect 21131 8044 21180 8072
rect 21131 8041 21143 8044
rect 21085 8035 21143 8041
rect 21174 8032 21180 8044
rect 21232 8032 21238 8084
rect 21450 8032 21456 8084
rect 21508 8072 21514 8084
rect 21508 8044 22048 8072
rect 21508 8032 21514 8044
rect 8389 8007 8447 8013
rect 8389 7973 8401 8007
rect 8435 8004 8447 8007
rect 9214 8004 9220 8016
rect 8435 7976 9220 8004
rect 8435 7973 8447 7976
rect 8389 7967 8447 7973
rect 9214 7964 9220 7976
rect 9272 7964 9278 8016
rect 9582 7964 9588 8016
rect 9640 8004 9646 8016
rect 9861 8007 9919 8013
rect 9861 8004 9873 8007
rect 9640 7976 9873 8004
rect 9640 7964 9646 7976
rect 9861 7973 9873 7976
rect 9907 7973 9919 8007
rect 17954 8004 17960 8016
rect 9861 7967 9919 7973
rect 9968 7976 10824 8004
rect 2406 7936 2412 7948
rect 2367 7908 2412 7936
rect 2406 7896 2412 7908
rect 2464 7936 2470 7948
rect 9309 7939 9367 7945
rect 2464 7908 4384 7936
rect 2464 7896 2470 7908
rect 4356 7880 4384 7908
rect 9309 7905 9321 7939
rect 9355 7936 9367 7939
rect 9968 7936 9996 7976
rect 10796 7948 10824 7976
rect 10888 7976 17960 8004
rect 9355 7908 9996 7936
rect 10229 7939 10287 7945
rect 9355 7905 9367 7908
rect 9309 7899 9367 7905
rect 10229 7905 10241 7939
rect 10275 7936 10287 7939
rect 10502 7936 10508 7948
rect 10275 7908 10508 7936
rect 10275 7905 10287 7908
rect 10229 7899 10287 7905
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 10778 7896 10784 7948
rect 10836 7896 10842 7948
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3844 7840 3985 7868
rect 3844 7828 3850 7840
rect 3973 7837 3985 7840
rect 4019 7868 4031 7871
rect 4249 7871 4307 7877
rect 4019 7840 4108 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 1854 7732 1860 7744
rect 1627 7704 1860 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 4080 7732 4108 7840
rect 4249 7837 4261 7871
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4154 7760 4160 7812
rect 4212 7800 4218 7812
rect 4264 7800 4292 7831
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 5721 7871 5779 7877
rect 5721 7868 5733 7871
rect 4396 7840 5733 7868
rect 4396 7828 4402 7840
rect 5721 7837 5733 7840
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 5997 7871 6055 7877
rect 5997 7837 6009 7871
rect 6043 7868 6055 7871
rect 6270 7868 6276 7880
rect 6043 7840 6276 7868
rect 6043 7837 6055 7840
rect 5997 7831 6055 7837
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7868 10103 7871
rect 10134 7868 10140 7880
rect 10091 7840 10140 7868
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 4430 7800 4436 7812
rect 4212 7772 4436 7800
rect 4212 7760 4218 7772
rect 4430 7760 4436 7772
rect 4488 7760 4494 7812
rect 5442 7760 5448 7812
rect 5500 7800 5506 7812
rect 7101 7803 7159 7809
rect 7101 7800 7113 7803
rect 5500 7772 7113 7800
rect 5500 7760 5506 7772
rect 7101 7769 7113 7772
rect 7147 7769 7159 7803
rect 7101 7763 7159 7769
rect 7190 7760 7196 7812
rect 7248 7800 7254 7812
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 7248 7772 7297 7800
rect 7248 7760 7254 7772
rect 7285 7769 7297 7772
rect 7331 7800 7343 7803
rect 8205 7803 8263 7809
rect 8205 7800 8217 7803
rect 7331 7772 8217 7800
rect 7331 7769 7343 7772
rect 7285 7763 7343 7769
rect 8205 7769 8217 7772
rect 8251 7800 8263 7803
rect 9416 7800 9444 7831
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10321 7803 10379 7809
rect 10321 7800 10333 7803
rect 8251 7772 8800 7800
rect 9416 7772 10333 7800
rect 8251 7769 8263 7772
rect 8205 7763 8263 7769
rect 5460 7732 5488 7760
rect 4080 7704 5488 7732
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7650 7732 7656 7744
rect 6972 7704 7656 7732
rect 6972 7692 6978 7704
rect 7650 7692 7656 7704
rect 7708 7692 7714 7744
rect 8772 7732 8800 7772
rect 10321 7769 10333 7772
rect 10367 7800 10379 7803
rect 10686 7800 10692 7812
rect 10367 7772 10692 7800
rect 10367 7769 10379 7772
rect 10321 7763 10379 7769
rect 10686 7760 10692 7772
rect 10744 7760 10750 7812
rect 10888 7732 10916 7976
rect 17954 7964 17960 7976
rect 18012 7964 18018 8016
rect 21910 8004 21916 8016
rect 21836 7976 21916 8004
rect 11977 7939 12035 7945
rect 11977 7905 11989 7939
rect 12023 7936 12035 7939
rect 12066 7936 12072 7948
rect 12023 7908 12072 7936
rect 12023 7905 12035 7908
rect 11977 7899 12035 7905
rect 12066 7896 12072 7908
rect 12124 7936 12130 7948
rect 13170 7936 13176 7948
rect 12124 7908 13176 7936
rect 12124 7896 12130 7908
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 21836 7945 21864 7976
rect 21910 7964 21916 7976
rect 21968 7964 21974 8016
rect 15933 7939 15991 7945
rect 15933 7936 15945 7939
rect 15620 7908 15945 7936
rect 15620 7896 15626 7908
rect 15933 7905 15945 7908
rect 15979 7905 15991 7939
rect 15933 7899 15991 7905
rect 21821 7939 21879 7945
rect 21821 7905 21833 7939
rect 21867 7905 21879 7939
rect 21821 7899 21879 7905
rect 10962 7828 10968 7880
rect 11020 7868 11026 7880
rect 11790 7868 11796 7880
rect 11020 7840 11796 7868
rect 11020 7828 11026 7840
rect 11790 7828 11796 7840
rect 11848 7868 11854 7880
rect 11848 7840 12112 7868
rect 11848 7828 11854 7840
rect 11149 7803 11207 7809
rect 11149 7769 11161 7803
rect 11195 7800 11207 7803
rect 11330 7800 11336 7812
rect 11195 7772 11336 7800
rect 11195 7769 11207 7772
rect 11149 7763 11207 7769
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 12084 7809 12112 7840
rect 12342 7828 12348 7880
rect 12400 7868 12406 7880
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 12400 7840 13001 7868
rect 12400 7828 12406 7840
rect 12989 7837 13001 7840
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7868 13323 7871
rect 13354 7868 13360 7880
rect 13311 7840 13360 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 12069 7803 12127 7809
rect 12069 7769 12081 7803
rect 12115 7769 12127 7803
rect 12069 7763 12127 7769
rect 12526 7760 12532 7812
rect 12584 7800 12590 7812
rect 13096 7800 13124 7831
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 15657 7871 15715 7877
rect 15657 7868 15669 7871
rect 15528 7840 15669 7868
rect 15528 7828 15534 7840
rect 15657 7837 15669 7840
rect 15703 7837 15715 7871
rect 15657 7831 15715 7837
rect 15746 7828 15752 7880
rect 15804 7868 15810 7880
rect 15841 7871 15899 7877
rect 15841 7868 15853 7871
rect 15804 7840 15853 7868
rect 15804 7828 15810 7840
rect 15841 7837 15853 7840
rect 15887 7837 15899 7871
rect 16022 7868 16028 7880
rect 15983 7840 16028 7868
rect 15841 7831 15899 7837
rect 16022 7828 16028 7840
rect 16080 7828 16086 7880
rect 16209 7871 16267 7877
rect 16209 7837 16221 7871
rect 16255 7868 16267 7871
rect 16482 7868 16488 7880
rect 16255 7840 16488 7868
rect 16255 7837 16267 7840
rect 16209 7831 16267 7837
rect 16482 7828 16488 7840
rect 16540 7828 16546 7880
rect 16850 7828 16856 7880
rect 16908 7868 16914 7880
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 16908 7840 17049 7868
rect 16908 7828 16914 7840
rect 17037 7837 17049 7840
rect 17083 7868 17095 7871
rect 17681 7871 17739 7877
rect 17681 7868 17693 7871
rect 17083 7840 17693 7868
rect 17083 7837 17095 7840
rect 17037 7831 17095 7837
rect 17681 7837 17693 7840
rect 17727 7837 17739 7871
rect 17681 7831 17739 7837
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7868 18015 7871
rect 18046 7868 18052 7880
rect 18003 7840 18052 7868
rect 18003 7837 18015 7840
rect 17957 7831 18015 7837
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7868 19763 7871
rect 19794 7868 19800 7880
rect 19751 7840 19800 7868
rect 19751 7837 19763 7840
rect 19705 7831 19763 7837
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 21542 7868 21548 7880
rect 21503 7840 21548 7868
rect 21542 7828 21548 7840
rect 21600 7828 21606 7880
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7837 21787 7871
rect 21729 7831 21787 7837
rect 21913 7871 21971 7877
rect 21913 7837 21925 7871
rect 21959 7868 21971 7871
rect 22020 7868 22048 8044
rect 21959 7840 22048 7868
rect 21959 7837 21971 7840
rect 21913 7831 21971 7837
rect 12584 7772 13124 7800
rect 17221 7803 17279 7809
rect 12584 7760 12590 7772
rect 17221 7769 17233 7803
rect 17267 7800 17279 7803
rect 17494 7800 17500 7812
rect 17267 7772 17500 7800
rect 17267 7769 17279 7772
rect 17221 7763 17279 7769
rect 17494 7760 17500 7772
rect 17552 7760 17558 7812
rect 19972 7803 20030 7809
rect 19972 7769 19984 7803
rect 20018 7800 20030 7803
rect 20070 7800 20076 7812
rect 20018 7772 20076 7800
rect 20018 7769 20030 7772
rect 19972 7763 20030 7769
rect 20070 7760 20076 7772
rect 20128 7760 20134 7812
rect 8772 7704 10916 7732
rect 12158 7692 12164 7744
rect 12216 7732 12222 7744
rect 13446 7732 13452 7744
rect 12216 7704 12261 7732
rect 13407 7704 13452 7732
rect 12216 7692 12222 7704
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 14918 7692 14924 7744
rect 14976 7732 14982 7744
rect 15286 7732 15292 7744
rect 14976 7704 15292 7732
rect 14976 7692 14982 7704
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 21744 7732 21772 7831
rect 22094 7828 22100 7880
rect 22152 7868 22158 7880
rect 22152 7840 22197 7868
rect 22152 7828 22158 7840
rect 22094 7732 22100 7744
rect 21744 7704 22100 7732
rect 22094 7692 22100 7704
rect 22152 7692 22158 7744
rect 22278 7732 22284 7744
rect 22239 7704 22284 7732
rect 22278 7692 22284 7704
rect 22336 7692 22342 7744
rect 1104 7642 30820 7664
rect 1104 7590 10880 7642
rect 10932 7590 10944 7642
rect 10996 7590 11008 7642
rect 11060 7590 11072 7642
rect 11124 7590 11136 7642
rect 11188 7590 20811 7642
rect 20863 7590 20875 7642
rect 20927 7590 20939 7642
rect 20991 7590 21003 7642
rect 21055 7590 21067 7642
rect 21119 7590 30820 7642
rect 1104 7568 30820 7590
rect 2222 7528 2228 7540
rect 2183 7500 2228 7528
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 6914 7488 6920 7540
rect 6972 7488 6978 7540
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 7374 7528 7380 7540
rect 7064 7500 7380 7528
rect 7064 7488 7070 7500
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 10137 7531 10195 7537
rect 10137 7528 10149 7531
rect 9824 7500 10149 7528
rect 9824 7488 9830 7500
rect 10137 7497 10149 7500
rect 10183 7497 10195 7531
rect 10137 7491 10195 7497
rect 11609 7531 11667 7537
rect 11609 7497 11621 7531
rect 11655 7528 11667 7531
rect 11882 7528 11888 7540
rect 11655 7500 11888 7528
rect 11655 7497 11667 7500
rect 11609 7491 11667 7497
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 13446 7528 13452 7540
rect 13407 7500 13452 7528
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 13817 7531 13875 7537
rect 13817 7497 13829 7531
rect 13863 7528 13875 7531
rect 14274 7528 14280 7540
rect 13863 7500 14280 7528
rect 13863 7497 13875 7500
rect 13817 7491 13875 7497
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 22186 7488 22192 7540
rect 22244 7528 22250 7540
rect 23201 7531 23259 7537
rect 23201 7528 23213 7531
rect 22244 7500 23213 7528
rect 22244 7488 22250 7500
rect 23201 7497 23213 7500
rect 23247 7497 23259 7531
rect 23201 7491 23259 7497
rect 1578 7460 1584 7472
rect 1504 7432 1584 7460
rect 1504 7401 1532 7432
rect 1578 7420 1584 7432
rect 1636 7420 1642 7472
rect 2590 7460 2596 7472
rect 1780 7432 2596 7460
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7361 1547 7395
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1489 7355 1547 7361
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 1780 7401 1808 7432
rect 2590 7420 2596 7432
rect 2648 7420 2654 7472
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 5534 7460 5540 7472
rect 4304 7432 4568 7460
rect 5495 7432 5540 7460
rect 4304 7420 4310 7432
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7361 1823 7395
rect 1765 7355 1823 7361
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 2774 7392 2780 7404
rect 2087 7364 2780 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 3510 7392 3516 7404
rect 3471 7364 3516 7392
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7392 3847 7395
rect 4338 7392 4344 7404
rect 3835 7364 4344 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 4338 7352 4344 7364
rect 4396 7352 4402 7404
rect 4540 7401 4568 7432
rect 5534 7420 5540 7432
rect 5592 7420 5598 7472
rect 5721 7463 5779 7469
rect 5721 7429 5733 7463
rect 5767 7460 5779 7463
rect 6932 7460 6960 7488
rect 5767 7432 6960 7460
rect 5767 7429 5779 7432
rect 5721 7423 5779 7429
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 6328 7364 6745 7392
rect 6328 7352 6334 7364
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 6917 7395 6975 7401
rect 6917 7361 6929 7395
rect 6963 7392 6975 7395
rect 7024 7392 7052 7488
rect 9674 7460 9680 7472
rect 8772 7432 9680 7460
rect 7282 7392 7288 7404
rect 6963 7364 7052 7392
rect 7243 7364 7288 7392
rect 6963 7361 6975 7364
rect 6917 7355 6975 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 8478 7392 8484 7404
rect 8439 7364 8484 7392
rect 8478 7352 8484 7364
rect 8536 7352 8542 7404
rect 8570 7352 8576 7404
rect 8628 7392 8634 7404
rect 8772 7401 8800 7432
rect 9674 7420 9680 7432
rect 9732 7420 9738 7472
rect 14369 7463 14427 7469
rect 14369 7460 14381 7463
rect 11716 7432 14381 7460
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 8628 7364 8677 7392
rect 8628 7352 8634 7364
rect 8665 7361 8677 7364
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 10226 7392 10232 7404
rect 9079 7364 10232 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 10318 7352 10324 7404
rect 10376 7392 10382 7404
rect 10597 7395 10655 7401
rect 10376 7364 10421 7392
rect 10376 7352 10382 7364
rect 10597 7361 10609 7395
rect 10643 7392 10655 7395
rect 10686 7392 10692 7404
rect 10643 7364 10692 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 10778 7352 10784 7404
rect 10836 7392 10842 7404
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 10836 7364 11529 7392
rect 10836 7352 10842 7364
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 11716 7401 11744 7432
rect 14369 7429 14381 7432
rect 14415 7429 14427 7463
rect 18138 7460 18144 7472
rect 14369 7423 14427 7429
rect 14936 7432 18144 7460
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11664 7364 11713 7392
rect 11664 7352 11670 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7392 12219 7395
rect 12342 7392 12348 7404
rect 12207 7364 12348 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 12492 7364 12537 7392
rect 12492 7352 12498 7364
rect 13906 7352 13912 7404
rect 13964 7392 13970 7404
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13964 7364 14289 7392
rect 13964 7352 13970 7364
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14458 7392 14464 7404
rect 14419 7364 14464 7392
rect 14277 7355 14335 7361
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 1857 7327 1915 7333
rect 1857 7293 1869 7327
rect 1903 7324 1915 7327
rect 2682 7324 2688 7336
rect 1903 7296 2688 7324
rect 1903 7293 1915 7296
rect 1857 7287 1915 7293
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7324 4307 7327
rect 5258 7324 5264 7336
rect 4295 7296 5264 7324
rect 4295 7293 4307 7296
rect 4249 7287 4307 7293
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 7009 7327 7067 7333
rect 7009 7324 7021 7327
rect 6880 7296 7021 7324
rect 6880 7284 6886 7296
rect 7009 7293 7021 7296
rect 7055 7293 7067 7327
rect 7009 7287 7067 7293
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7190 7324 7196 7336
rect 7147 7296 7196 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7024 7256 7052 7287
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 8849 7327 8907 7333
rect 8849 7293 8861 7327
rect 8895 7324 8907 7327
rect 9214 7324 9220 7336
rect 8895 7296 9220 7324
rect 8895 7293 8907 7296
rect 8849 7287 8907 7293
rect 9214 7284 9220 7296
rect 9272 7284 9278 7336
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7324 10563 7327
rect 11330 7324 11336 7336
rect 10551 7296 11336 7324
rect 10551 7293 10563 7296
rect 10505 7287 10563 7293
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7324 12311 7327
rect 12526 7324 12532 7336
rect 12299 7296 12532 7324
rect 12299 7293 12311 7296
rect 12253 7287 12311 7293
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 13170 7324 13176 7336
rect 13131 7296 13176 7324
rect 13170 7284 13176 7296
rect 13228 7284 13234 7336
rect 13354 7324 13360 7336
rect 13315 7296 13360 7324
rect 13354 7284 13360 7296
rect 13412 7284 13418 7336
rect 14936 7256 14964 7432
rect 18138 7420 18144 7432
rect 18196 7460 18202 7472
rect 18414 7460 18420 7472
rect 18196 7432 18420 7460
rect 18196 7420 18202 7432
rect 18414 7420 18420 7432
rect 18472 7420 18478 7472
rect 22088 7463 22146 7469
rect 22088 7429 22100 7463
rect 22134 7460 22146 7463
rect 22278 7460 22284 7472
rect 22134 7432 22284 7460
rect 22134 7429 22146 7432
rect 22088 7423 22146 7429
rect 22278 7420 22284 7432
rect 22336 7420 22342 7472
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7392 15347 7395
rect 15378 7392 15384 7404
rect 15335 7364 15384 7392
rect 15335 7361 15347 7364
rect 15289 7355 15347 7361
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 15488 7324 15516 7355
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 15841 7395 15899 7401
rect 15620 7364 15665 7392
rect 15620 7352 15626 7364
rect 15841 7361 15853 7395
rect 15887 7392 15899 7395
rect 16666 7392 16672 7404
rect 15887 7364 16672 7392
rect 15887 7361 15899 7364
rect 15841 7355 15899 7361
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 17954 7392 17960 7404
rect 17915 7364 17960 7392
rect 17954 7352 17960 7364
rect 18012 7392 18018 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18012 7364 18613 7392
rect 18012 7352 18018 7364
rect 18601 7361 18613 7364
rect 18647 7392 18659 7395
rect 20901 7395 20959 7401
rect 20901 7392 20913 7395
rect 18647 7364 20913 7392
rect 18647 7361 18659 7364
rect 18601 7355 18659 7361
rect 20901 7361 20913 7364
rect 20947 7361 20959 7395
rect 29822 7392 29828 7404
rect 29783 7364 29828 7392
rect 20901 7355 20959 7361
rect 29822 7352 29828 7364
rect 29880 7352 29886 7404
rect 15068 7296 15516 7324
rect 15657 7327 15715 7333
rect 15068 7284 15074 7296
rect 15657 7293 15669 7327
rect 15703 7324 15715 7327
rect 16022 7324 16028 7336
rect 15703 7296 16028 7324
rect 15703 7293 15715 7296
rect 15657 7287 15715 7293
rect 7024 7228 14964 7256
rect 7469 7191 7527 7197
rect 7469 7157 7481 7191
rect 7515 7188 7527 7191
rect 8110 7188 8116 7200
rect 7515 7160 8116 7188
rect 7515 7157 7527 7160
rect 7469 7151 7527 7157
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 9214 7188 9220 7200
rect 9175 7160 9220 7188
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 10502 7188 10508 7200
rect 10463 7160 10508 7188
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 12618 7188 12624 7200
rect 12579 7160 12624 7188
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 15672 7188 15700 7287
rect 16022 7284 16028 7296
rect 16080 7324 16086 7336
rect 16942 7324 16948 7336
rect 16080 7296 16948 7324
rect 16080 7284 16086 7296
rect 16942 7284 16948 7296
rect 17000 7324 17006 7336
rect 17681 7327 17739 7333
rect 17681 7324 17693 7327
rect 17000 7296 17693 7324
rect 17000 7284 17006 7296
rect 17681 7293 17693 7296
rect 17727 7293 17739 7327
rect 19426 7324 19432 7336
rect 19387 7296 19432 7324
rect 17681 7287 17739 7293
rect 19426 7284 19432 7296
rect 19484 7284 19490 7336
rect 19610 7284 19616 7336
rect 19668 7324 19674 7336
rect 19705 7327 19763 7333
rect 19705 7324 19717 7327
rect 19668 7296 19717 7324
rect 19668 7284 19674 7296
rect 19705 7293 19717 7296
rect 19751 7324 19763 7327
rect 20622 7324 20628 7336
rect 19751 7296 20628 7324
rect 19751 7293 19763 7296
rect 19705 7287 19763 7293
rect 20622 7284 20628 7296
rect 20680 7324 20686 7336
rect 21634 7324 21640 7336
rect 20680 7296 21640 7324
rect 20680 7284 20686 7296
rect 21634 7284 21640 7296
rect 21692 7284 21698 7336
rect 21818 7324 21824 7336
rect 21779 7296 21824 7324
rect 21818 7284 21824 7296
rect 21876 7284 21882 7336
rect 15436 7160 15700 7188
rect 15436 7148 15442 7160
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 16025 7191 16083 7197
rect 16025 7188 16037 7191
rect 15804 7160 16037 7188
rect 15804 7148 15810 7160
rect 16025 7157 16037 7160
rect 16071 7157 16083 7191
rect 16025 7151 16083 7157
rect 18322 7148 18328 7200
rect 18380 7188 18386 7200
rect 18509 7191 18567 7197
rect 18509 7188 18521 7191
rect 18380 7160 18521 7188
rect 18380 7148 18386 7160
rect 18509 7157 18521 7160
rect 18555 7157 18567 7191
rect 18509 7151 18567 7157
rect 20809 7191 20867 7197
rect 20809 7157 20821 7191
rect 20855 7188 20867 7191
rect 21266 7188 21272 7200
rect 20855 7160 21272 7188
rect 20855 7157 20867 7160
rect 20809 7151 20867 7157
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 30006 7188 30012 7200
rect 29967 7160 30012 7188
rect 30006 7148 30012 7160
rect 30064 7148 30070 7200
rect 1104 7098 30820 7120
rect 1104 7046 5915 7098
rect 5967 7046 5979 7098
rect 6031 7046 6043 7098
rect 6095 7046 6107 7098
rect 6159 7046 6171 7098
rect 6223 7046 15846 7098
rect 15898 7046 15910 7098
rect 15962 7046 15974 7098
rect 16026 7046 16038 7098
rect 16090 7046 16102 7098
rect 16154 7046 25776 7098
rect 25828 7046 25840 7098
rect 25892 7046 25904 7098
rect 25956 7046 25968 7098
rect 26020 7046 26032 7098
rect 26084 7046 30820 7098
rect 1104 7024 30820 7046
rect 4154 6944 4160 6996
rect 4212 6944 4218 6996
rect 7006 6984 7012 6996
rect 6919 6956 7012 6984
rect 7006 6944 7012 6956
rect 7064 6984 7070 6996
rect 7282 6984 7288 6996
rect 7064 6956 7288 6984
rect 7064 6944 7070 6956
rect 7282 6944 7288 6956
rect 7340 6944 7346 6996
rect 9306 6944 9312 6996
rect 9364 6984 9370 6996
rect 9364 6956 9904 6984
rect 9364 6944 9370 6956
rect 3786 6916 3792 6928
rect 2056 6888 3792 6916
rect 2056 6857 2084 6888
rect 3786 6876 3792 6888
rect 3844 6916 3850 6928
rect 4172 6916 4200 6944
rect 9876 6916 9904 6956
rect 10226 6944 10232 6996
rect 10284 6984 10290 6996
rect 10321 6987 10379 6993
rect 10321 6984 10333 6987
rect 10284 6956 10333 6984
rect 10284 6944 10290 6956
rect 10321 6953 10333 6956
rect 10367 6953 10379 6987
rect 18322 6984 18328 6996
rect 10321 6947 10379 6953
rect 12406 6956 18328 6984
rect 12406 6916 12434 6956
rect 18322 6944 18328 6956
rect 18380 6944 18386 6996
rect 20070 6984 20076 6996
rect 20031 6956 20076 6984
rect 20070 6944 20076 6956
rect 20128 6944 20134 6996
rect 29822 6944 29828 6996
rect 29880 6984 29886 6996
rect 29917 6987 29975 6993
rect 29917 6984 29929 6987
rect 29880 6956 29929 6984
rect 29880 6944 29886 6956
rect 29917 6953 29929 6956
rect 29963 6953 29975 6987
rect 29917 6947 29975 6953
rect 3844 6888 4200 6916
rect 3844 6876 3850 6888
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6817 2099 6851
rect 4062 6848 4068 6860
rect 4023 6820 4068 6848
rect 2041 6811 2099 6817
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4172 6857 4200 6888
rect 5736 6888 6684 6916
rect 9876 6888 12434 6916
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6817 4215 6851
rect 4157 6811 4215 6817
rect 5169 6851 5227 6857
rect 5169 6817 5181 6851
rect 5215 6848 5227 6851
rect 5442 6848 5448 6860
rect 5215 6820 5448 6848
rect 5215 6817 5227 6820
rect 5169 6811 5227 6817
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 1673 6783 1731 6789
rect 1673 6780 1685 6783
rect 1636 6752 1685 6780
rect 1636 6740 1642 6752
rect 1673 6749 1685 6752
rect 1719 6749 1731 6783
rect 1854 6780 1860 6792
rect 1815 6752 1860 6780
rect 1673 6743 1731 6749
rect 1854 6740 1860 6752
rect 1912 6740 1918 6792
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 1949 6743 2007 6749
rect 1964 6712 1992 6743
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 3510 6740 3516 6792
rect 3568 6780 3574 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3568 6752 3801 6780
rect 3568 6740 3574 6752
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3936 6752 3985 6780
rect 3936 6740 3942 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 4338 6780 4344 6792
rect 4299 6752 4344 6780
rect 3973 6743 4031 6749
rect 4338 6740 4344 6752
rect 4396 6740 4402 6792
rect 5258 6780 5264 6792
rect 5171 6752 5264 6780
rect 5258 6740 5264 6752
rect 5316 6780 5322 6792
rect 5736 6780 5764 6888
rect 6089 6851 6147 6857
rect 5828 6820 6040 6848
rect 5828 6789 5856 6820
rect 5316 6752 5764 6780
rect 5813 6783 5871 6789
rect 5316 6740 5322 6752
rect 5813 6749 5825 6783
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 2590 6712 2596 6724
rect 1964 6684 2596 6712
rect 2590 6672 2596 6684
rect 2648 6712 2654 6724
rect 3145 6715 3203 6721
rect 2648 6684 2774 6712
rect 2648 6672 2654 6684
rect 2406 6644 2412 6656
rect 2367 6616 2412 6644
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 2746 6644 2774 6684
rect 3145 6681 3157 6715
rect 3191 6712 3203 6715
rect 5276 6712 5304 6740
rect 3191 6684 5304 6712
rect 3191 6681 3203 6684
rect 3145 6675 3203 6681
rect 3050 6644 3056 6656
rect 2746 6616 3056 6644
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 4522 6644 4528 6656
rect 4483 6616 4528 6644
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 5920 6644 5948 6743
rect 6012 6712 6040 6820
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 6546 6848 6552 6860
rect 6135 6820 6552 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 6656 6848 6684 6888
rect 15470 6876 15476 6928
rect 15528 6916 15534 6928
rect 16206 6916 16212 6928
rect 15528 6888 16212 6916
rect 15528 6876 15534 6888
rect 16206 6876 16212 6888
rect 16264 6916 16270 6928
rect 18138 6916 18144 6928
rect 16264 6888 16528 6916
rect 18099 6888 18144 6916
rect 16264 6876 16270 6888
rect 6656 6820 7052 6848
rect 6178 6780 6184 6792
rect 6139 6752 6184 6780
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6454 6780 6460 6792
rect 6415 6752 6460 6780
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 6914 6712 6920 6724
rect 6012 6684 6920 6712
rect 6914 6672 6920 6684
rect 6972 6672 6978 6724
rect 7024 6712 7052 6820
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 12124 6820 12265 6848
rect 12124 6808 12130 6820
rect 12253 6817 12265 6820
rect 12299 6848 12311 6851
rect 12710 6848 12716 6860
rect 12299 6820 12716 6848
rect 12299 6817 12311 6820
rect 12253 6811 12311 6817
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 14829 6851 14887 6857
rect 14829 6817 14841 6851
rect 14875 6848 14887 6851
rect 15562 6848 15568 6860
rect 14875 6820 15568 6848
rect 14875 6817 14887 6820
rect 14829 6811 14887 6817
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 15948 6820 16436 6848
rect 8110 6740 8116 6792
rect 8168 6789 8174 6792
rect 8168 6780 8180 6789
rect 8389 6783 8447 6789
rect 8168 6752 8213 6780
rect 8168 6743 8180 6752
rect 8389 6749 8401 6783
rect 8435 6780 8447 6783
rect 8662 6780 8668 6792
rect 8435 6752 8668 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 8168 6740 8174 6743
rect 8662 6740 8668 6752
rect 8720 6780 8726 6792
rect 9214 6789 9220 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8720 6752 8953 6780
rect 8720 6740 8726 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 9208 6780 9220 6789
rect 9175 6752 9220 6780
rect 8941 6743 8999 6749
rect 9208 6743 9220 6752
rect 9214 6740 9220 6743
rect 9272 6740 9278 6792
rect 12529 6783 12587 6789
rect 12529 6749 12541 6783
rect 12575 6780 12587 6783
rect 12618 6780 12624 6792
rect 12575 6752 12624 6780
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 15948 6780 15976 6820
rect 14599 6752 15976 6780
rect 16025 6783 16083 6789
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 16025 6749 16037 6783
rect 16071 6749 16083 6783
rect 16025 6743 16083 6749
rect 10965 6715 11023 6721
rect 10965 6712 10977 6715
rect 7024 6684 10977 6712
rect 10965 6681 10977 6684
rect 11011 6681 11023 6715
rect 14568 6712 14596 6743
rect 10965 6675 11023 6681
rect 11164 6684 14596 6712
rect 6822 6644 6828 6656
rect 5920 6616 6828 6644
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 10468 6616 10885 6644
rect 10468 6604 10474 6616
rect 10873 6613 10885 6616
rect 10919 6644 10931 6647
rect 11164 6644 11192 6684
rect 14826 6672 14832 6724
rect 14884 6712 14890 6724
rect 16040 6712 16068 6743
rect 14884 6684 16068 6712
rect 16408 6712 16436 6820
rect 16500 6780 16528 6888
rect 18138 6876 18144 6888
rect 18196 6876 18202 6928
rect 16942 6848 16948 6860
rect 16903 6820 16948 6848
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 19610 6848 19616 6860
rect 19571 6820 19616 6848
rect 19610 6808 19616 6820
rect 19668 6808 19674 6860
rect 19794 6808 19800 6860
rect 19852 6848 19858 6860
rect 20533 6851 20591 6857
rect 20533 6848 20545 6851
rect 19852 6820 20545 6848
rect 19852 6808 19858 6820
rect 20533 6817 20545 6820
rect 20579 6817 20591 6851
rect 20533 6811 20591 6817
rect 16577 6783 16635 6789
rect 16577 6780 16589 6783
rect 16500 6752 16589 6780
rect 16577 6749 16589 6752
rect 16623 6749 16635 6783
rect 16758 6780 16764 6792
rect 16719 6752 16764 6780
rect 16577 6743 16635 6749
rect 16758 6740 16764 6752
rect 16816 6740 16822 6792
rect 16850 6740 16856 6792
rect 16908 6780 16914 6792
rect 17129 6783 17187 6789
rect 16908 6752 16953 6780
rect 16908 6740 16914 6752
rect 17129 6749 17141 6783
rect 17175 6780 17187 6783
rect 17402 6780 17408 6792
rect 17175 6752 17408 6780
rect 17175 6749 17187 6752
rect 17129 6743 17187 6749
rect 17402 6740 17408 6752
rect 17460 6740 17466 6792
rect 17494 6740 17500 6792
rect 17552 6780 17558 6792
rect 19337 6783 19395 6789
rect 19337 6780 19349 6783
rect 17552 6752 19349 6780
rect 17552 6740 17558 6752
rect 19337 6749 19349 6752
rect 19383 6749 19395 6783
rect 19518 6780 19524 6792
rect 19479 6752 19524 6780
rect 19337 6743 19395 6749
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6780 19763 6783
rect 19889 6783 19947 6789
rect 19751 6752 19840 6780
rect 19751 6749 19763 6752
rect 19705 6743 19763 6749
rect 17957 6715 18015 6721
rect 17957 6712 17969 6715
rect 16408 6684 17969 6712
rect 14884 6672 14890 6684
rect 17957 6681 17969 6684
rect 18003 6712 18015 6715
rect 19426 6712 19432 6724
rect 18003 6684 19432 6712
rect 18003 6681 18015 6684
rect 17957 6675 18015 6681
rect 19426 6672 19432 6684
rect 19484 6672 19490 6724
rect 10919 6616 11192 6644
rect 10919 6613 10931 6616
rect 10873 6607 10931 6613
rect 12066 6604 12072 6656
rect 12124 6644 12130 6656
rect 12250 6644 12256 6656
rect 12124 6616 12256 6644
rect 12124 6604 12130 6616
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 12802 6644 12808 6656
rect 12492 6616 12808 6644
rect 12492 6604 12498 6616
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 12897 6647 12955 6653
rect 12897 6613 12909 6647
rect 12943 6644 12955 6647
rect 13538 6644 13544 6656
rect 12943 6616 13544 6644
rect 12943 6613 12955 6616
rect 12897 6607 12955 6613
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 13630 6604 13636 6656
rect 13688 6644 13694 6656
rect 15286 6644 15292 6656
rect 13688 6616 15292 6644
rect 13688 6604 13694 6616
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 15470 6604 15476 6656
rect 15528 6644 15534 6656
rect 15841 6647 15899 6653
rect 15841 6644 15853 6647
rect 15528 6616 15853 6644
rect 15528 6604 15534 6616
rect 15841 6613 15853 6616
rect 15887 6613 15899 6647
rect 17310 6644 17316 6656
rect 17271 6616 17316 6644
rect 15841 6607 15899 6613
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 19812 6644 19840 6752
rect 19889 6749 19901 6783
rect 19935 6780 19947 6783
rect 21082 6780 21088 6792
rect 19935 6752 21088 6780
rect 19935 6749 19947 6752
rect 19889 6743 19947 6749
rect 21082 6740 21088 6752
rect 21140 6740 21146 6792
rect 29638 6740 29644 6792
rect 29696 6780 29702 6792
rect 29917 6783 29975 6789
rect 29917 6780 29929 6783
rect 29696 6752 29929 6780
rect 29696 6740 29702 6752
rect 29917 6749 29929 6752
rect 29963 6749 29975 6783
rect 30098 6780 30104 6792
rect 30059 6752 30104 6780
rect 29917 6743 29975 6749
rect 30098 6740 30104 6752
rect 30156 6740 30162 6792
rect 20800 6715 20858 6721
rect 20800 6681 20812 6715
rect 20846 6712 20858 6715
rect 21174 6712 21180 6724
rect 20846 6684 21180 6712
rect 20846 6681 20858 6684
rect 20800 6675 20858 6681
rect 21174 6672 21180 6684
rect 21232 6672 21238 6724
rect 21266 6644 21272 6656
rect 19812 6616 21272 6644
rect 21266 6604 21272 6616
rect 21324 6604 21330 6656
rect 21726 6604 21732 6656
rect 21784 6644 21790 6656
rect 21913 6647 21971 6653
rect 21913 6644 21925 6647
rect 21784 6616 21925 6644
rect 21784 6604 21790 6616
rect 21913 6613 21925 6616
rect 21959 6613 21971 6647
rect 21913 6607 21971 6613
rect 1104 6554 30820 6576
rect 1104 6502 10880 6554
rect 10932 6502 10944 6554
rect 10996 6502 11008 6554
rect 11060 6502 11072 6554
rect 11124 6502 11136 6554
rect 11188 6502 20811 6554
rect 20863 6502 20875 6554
rect 20927 6502 20939 6554
rect 20991 6502 21003 6554
rect 21055 6502 21067 6554
rect 21119 6502 30820 6554
rect 1104 6480 30820 6502
rect 2222 6400 2228 6452
rect 2280 6440 2286 6452
rect 2961 6443 3019 6449
rect 2961 6440 2973 6443
rect 2280 6412 2973 6440
rect 2280 6400 2286 6412
rect 2961 6409 2973 6412
rect 3007 6440 3019 6443
rect 3007 6412 4108 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 1486 6332 1492 6384
rect 1544 6372 1550 6384
rect 1544 6344 4016 6372
rect 1544 6332 1550 6344
rect 1596 6313 1624 6344
rect 3988 6316 4016 6344
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 1848 6307 1906 6313
rect 1627 6276 1661 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 1848 6273 1860 6307
rect 1894 6304 1906 6307
rect 2406 6304 2412 6316
rect 1894 6276 2412 6304
rect 1894 6273 1906 6276
rect 1848 6267 1906 6273
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 3970 6304 3976 6316
rect 3883 6276 3976 6304
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4080 6304 4108 6412
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 5353 6443 5411 6449
rect 5353 6440 5365 6443
rect 4396 6412 5365 6440
rect 4396 6400 4402 6412
rect 5353 6409 5365 6412
rect 5399 6440 5411 6443
rect 6914 6440 6920 6452
rect 5399 6412 6592 6440
rect 5399 6409 5411 6412
rect 5353 6403 5411 6409
rect 4240 6375 4298 6381
rect 4240 6341 4252 6375
rect 4286 6372 4298 6375
rect 4522 6372 4528 6384
rect 4286 6344 4528 6372
rect 4286 6341 4298 6344
rect 4240 6335 4298 6341
rect 4522 6332 4528 6344
rect 4580 6332 4586 6384
rect 6564 6381 6592 6412
rect 6656 6412 6920 6440
rect 6549 6375 6607 6381
rect 6549 6341 6561 6375
rect 6595 6341 6607 6375
rect 6656 6372 6684 6412
rect 6914 6400 6920 6412
rect 6972 6440 6978 6452
rect 7742 6440 7748 6452
rect 6972 6412 7748 6440
rect 6972 6400 6978 6412
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 11885 6443 11943 6449
rect 11885 6409 11897 6443
rect 11931 6440 11943 6443
rect 12158 6440 12164 6452
rect 11931 6412 12164 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 12250 6400 12256 6452
rect 12308 6440 12314 6452
rect 12308 6412 15056 6440
rect 12308 6400 12314 6412
rect 6779 6375 6837 6381
rect 6779 6372 6791 6375
rect 6656 6344 6791 6372
rect 6549 6335 6607 6341
rect 6779 6341 6791 6344
rect 6825 6341 6837 6375
rect 6779 6335 6837 6341
rect 7650 6332 7656 6384
rect 7708 6372 7714 6384
rect 8573 6375 8631 6381
rect 8573 6372 8585 6375
rect 7708 6344 8585 6372
rect 7708 6332 7714 6344
rect 8573 6341 8585 6344
rect 8619 6341 8631 6375
rect 8573 6335 8631 6341
rect 10962 6332 10968 6384
rect 11020 6372 11026 6384
rect 13630 6372 13636 6384
rect 11020 6344 13636 6372
rect 11020 6332 11026 6344
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 6178 6304 6184 6316
rect 4080 6276 6184 6304
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 6454 6313 6460 6316
rect 6452 6304 6460 6313
rect 6415 6276 6460 6304
rect 6452 6267 6460 6276
rect 6454 6264 6460 6267
rect 6512 6264 6518 6316
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 7006 6304 7012 6316
rect 6687 6294 6776 6304
rect 6932 6294 7012 6304
rect 6687 6276 7012 6294
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 6748 6266 6960 6276
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7341 6307 7399 6313
rect 7341 6273 7353 6307
rect 7387 6273 7399 6307
rect 7341 6267 7399 6273
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 6472 6236 6500 6264
rect 7356 6236 7384 6267
rect 6472 6208 7384 6236
rect 7484 6168 7512 6267
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7616 6276 7661 6304
rect 7616 6264 7622 6276
rect 7742 6264 7748 6316
rect 7800 6304 7806 6316
rect 7800 6276 7845 6304
rect 7800 6264 7806 6276
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 10045 6307 10103 6313
rect 10045 6304 10057 6307
rect 9732 6276 10057 6304
rect 9732 6264 9738 6276
rect 10045 6273 10057 6276
rect 10091 6273 10103 6307
rect 10045 6267 10103 6273
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6304 10379 6307
rect 10410 6304 10416 6316
rect 10367 6276 10416 6304
rect 10367 6273 10379 6276
rect 10321 6267 10379 6273
rect 10410 6264 10416 6276
rect 10468 6264 10474 6316
rect 11790 6264 11796 6316
rect 11848 6304 11854 6316
rect 12069 6307 12127 6313
rect 12069 6304 12081 6307
rect 11848 6276 12081 6304
rect 11848 6264 11854 6276
rect 12069 6273 12081 6276
rect 12115 6273 12127 6307
rect 12342 6304 12348 6316
rect 12303 6276 12348 6304
rect 12069 6267 12127 6273
rect 4908 6140 7512 6168
rect 7745 6171 7803 6177
rect 3234 6060 3240 6112
rect 3292 6100 3298 6112
rect 4908 6100 4936 6140
rect 7745 6137 7757 6171
rect 7791 6168 7803 6171
rect 7926 6168 7932 6180
rect 7791 6140 7932 6168
rect 7791 6137 7803 6140
rect 7745 6131 7803 6137
rect 7926 6128 7932 6140
rect 7984 6128 7990 6180
rect 12084 6168 12112 6267
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 14366 6304 14372 6316
rect 14327 6276 14372 6304
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 14642 6313 14648 6316
rect 14636 6267 14648 6313
rect 14700 6304 14706 6316
rect 14700 6276 14736 6304
rect 15028 6302 15056 6412
rect 15194 6400 15200 6452
rect 15252 6440 15258 6452
rect 15749 6443 15807 6449
rect 15749 6440 15761 6443
rect 15252 6412 15761 6440
rect 15252 6400 15258 6412
rect 15749 6409 15761 6412
rect 15795 6409 15807 6443
rect 15749 6403 15807 6409
rect 16669 6443 16727 6449
rect 16669 6409 16681 6443
rect 16715 6440 16727 6443
rect 17402 6440 17408 6452
rect 16715 6412 17408 6440
rect 16715 6409 16727 6412
rect 16669 6403 16727 6409
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 18046 6400 18052 6452
rect 18104 6440 18110 6452
rect 18509 6443 18567 6449
rect 18509 6440 18521 6443
rect 18104 6412 18521 6440
rect 18104 6400 18110 6412
rect 18509 6409 18521 6412
rect 18555 6440 18567 6443
rect 18874 6440 18880 6452
rect 18555 6412 18880 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 21085 6443 21143 6449
rect 19300 6412 20392 6440
rect 19300 6400 19306 6412
rect 15102 6332 15108 6384
rect 15160 6372 15166 6384
rect 19334 6372 19340 6384
rect 15160 6344 19340 6372
rect 15160 6332 15166 6344
rect 16298 6304 16304 6316
rect 15212 6302 16304 6304
rect 15028 6276 16304 6302
rect 14642 6264 14648 6267
rect 14700 6264 14706 6276
rect 15028 6274 15240 6276
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 18064 6313 18092 6344
rect 19334 6332 19340 6344
rect 19392 6372 19398 6384
rect 19794 6372 19800 6384
rect 19392 6344 19800 6372
rect 19392 6332 19398 6344
rect 19794 6332 19800 6344
rect 19852 6372 19858 6384
rect 19852 6344 19932 6372
rect 19852 6332 19858 6344
rect 17782 6307 17840 6313
rect 17782 6304 17794 6307
rect 17368 6276 17794 6304
rect 17368 6264 17374 6276
rect 17782 6273 17794 6276
rect 17828 6273 17840 6307
rect 17782 6267 17840 6273
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6273 18107 6307
rect 18049 6267 18107 6273
rect 18230 6264 18236 6316
rect 18288 6304 18294 6316
rect 19904 6313 19932 6344
rect 20364 6313 20392 6412
rect 21085 6409 21097 6443
rect 21131 6440 21143 6443
rect 21174 6440 21180 6452
rect 21131 6412 21180 6440
rect 21131 6409 21143 6412
rect 21085 6403 21143 6409
rect 21174 6400 21180 6412
rect 21232 6400 21238 6452
rect 19622 6307 19680 6313
rect 19622 6304 19634 6307
rect 18288 6276 19634 6304
rect 18288 6264 18294 6276
rect 19622 6273 19634 6276
rect 19668 6273 19680 6307
rect 19622 6267 19680 6273
rect 19889 6307 19947 6313
rect 19889 6273 19901 6307
rect 19935 6273 19947 6307
rect 19889 6267 19947 6273
rect 20349 6307 20407 6313
rect 20349 6273 20361 6307
rect 20395 6273 20407 6307
rect 20530 6304 20536 6316
rect 20491 6276 20536 6304
rect 20349 6267 20407 6273
rect 20530 6264 20536 6276
rect 20588 6264 20594 6316
rect 20622 6264 20628 6316
rect 20680 6304 20686 6316
rect 20901 6307 20959 6313
rect 20680 6276 20725 6304
rect 20680 6264 20686 6276
rect 20901 6273 20913 6307
rect 20947 6304 20959 6307
rect 21726 6304 21732 6316
rect 20947 6276 21732 6304
rect 20947 6273 20959 6276
rect 20901 6267 20959 6273
rect 21726 6264 21732 6276
rect 21784 6264 21790 6316
rect 13633 6239 13691 6245
rect 13633 6205 13645 6239
rect 13679 6236 13691 6239
rect 13722 6236 13728 6248
rect 13679 6208 13728 6236
rect 13679 6205 13691 6208
rect 13633 6199 13691 6205
rect 12618 6168 12624 6180
rect 12084 6140 12624 6168
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 13648 6168 13676 6199
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 13906 6236 13912 6248
rect 13867 6208 13912 6236
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 20438 6196 20444 6248
rect 20496 6236 20502 6248
rect 20717 6239 20775 6245
rect 20717 6236 20729 6239
rect 20496 6208 20729 6236
rect 20496 6196 20502 6208
rect 20717 6205 20729 6208
rect 20763 6236 20775 6239
rect 21266 6236 21272 6248
rect 20763 6208 21272 6236
rect 20763 6205 20775 6208
rect 20717 6199 20775 6205
rect 21266 6196 21272 6208
rect 21324 6196 21330 6248
rect 13004 6140 13676 6168
rect 3292 6072 4936 6100
rect 3292 6060 3298 6072
rect 6362 6060 6368 6112
rect 6420 6100 6426 6112
rect 6825 6103 6883 6109
rect 6825 6100 6837 6103
rect 6420 6072 6837 6100
rect 6420 6060 6426 6072
rect 6825 6069 6837 6072
rect 6871 6069 6883 6103
rect 8662 6100 8668 6112
rect 8623 6072 8668 6100
rect 6825 6063 6883 6069
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 12253 6103 12311 6109
rect 12253 6069 12265 6103
rect 12299 6100 12311 6103
rect 12434 6100 12440 6112
rect 12299 6072 12440 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 12434 6060 12440 6072
rect 12492 6100 12498 6112
rect 13004 6100 13032 6140
rect 12492 6072 13032 6100
rect 12492 6060 12498 6072
rect 13262 6060 13268 6112
rect 13320 6100 13326 6112
rect 30098 6100 30104 6112
rect 13320 6072 30104 6100
rect 13320 6060 13326 6072
rect 30098 6060 30104 6072
rect 30156 6060 30162 6112
rect 1104 6010 30820 6032
rect 1104 5958 5915 6010
rect 5967 5958 5979 6010
rect 6031 5958 6043 6010
rect 6095 5958 6107 6010
rect 6159 5958 6171 6010
rect 6223 5958 15846 6010
rect 15898 5958 15910 6010
rect 15962 5958 15974 6010
rect 16026 5958 16038 6010
rect 16090 5958 16102 6010
rect 16154 5958 25776 6010
rect 25828 5958 25840 6010
rect 25892 5958 25904 6010
rect 25956 5958 25968 6010
rect 26020 5958 26032 6010
rect 26084 5958 30820 6010
rect 1104 5936 30820 5958
rect 3234 5896 3240 5908
rect 3195 5868 3240 5896
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 5537 5899 5595 5905
rect 5537 5865 5549 5899
rect 5583 5896 5595 5899
rect 5718 5896 5724 5908
rect 5583 5868 5724 5896
rect 5583 5865 5595 5868
rect 5537 5859 5595 5865
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 13173 5899 13231 5905
rect 13173 5896 13185 5899
rect 11388 5868 13185 5896
rect 11388 5856 11394 5868
rect 13173 5865 13185 5868
rect 13219 5865 13231 5899
rect 13173 5859 13231 5865
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 13541 5899 13599 5905
rect 13541 5896 13553 5899
rect 13412 5868 13553 5896
rect 13412 5856 13418 5868
rect 13541 5865 13553 5868
rect 13587 5896 13599 5899
rect 15013 5899 15071 5905
rect 15013 5896 15025 5899
rect 13587 5868 15025 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 15013 5865 15025 5868
rect 15059 5865 15071 5899
rect 15013 5859 15071 5865
rect 16666 5856 16672 5908
rect 16724 5896 16730 5908
rect 17037 5899 17095 5905
rect 17037 5896 17049 5899
rect 16724 5868 17049 5896
rect 16724 5856 16730 5868
rect 17037 5865 17049 5868
rect 17083 5865 17095 5899
rect 18230 5896 18236 5908
rect 18191 5868 18236 5896
rect 17037 5859 17095 5865
rect 18230 5856 18236 5868
rect 18288 5856 18294 5908
rect 19702 5856 19708 5908
rect 19760 5896 19766 5908
rect 20625 5899 20683 5905
rect 20625 5896 20637 5899
rect 19760 5868 20637 5896
rect 19760 5856 19766 5868
rect 20625 5865 20637 5868
rect 20671 5865 20683 5899
rect 20625 5859 20683 5865
rect 29454 5856 29460 5908
rect 29512 5896 29518 5908
rect 29822 5896 29828 5908
rect 29512 5868 29828 5896
rect 29512 5856 29518 5868
rect 29822 5856 29828 5868
rect 29880 5856 29886 5908
rect 6730 5828 6736 5840
rect 6564 5800 6736 5828
rect 1486 5720 1492 5772
rect 1544 5760 1550 5772
rect 1857 5763 1915 5769
rect 1857 5760 1869 5763
rect 1544 5732 1869 5760
rect 1544 5720 1550 5732
rect 1857 5729 1869 5732
rect 1903 5729 1915 5763
rect 1857 5723 1915 5729
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 6564 5769 6592 5800
rect 6730 5788 6736 5800
rect 6788 5788 6794 5840
rect 11974 5828 11980 5840
rect 11935 5800 11980 5828
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 12342 5788 12348 5840
rect 12400 5828 12406 5840
rect 12400 5800 14136 5828
rect 12400 5788 12406 5800
rect 4157 5763 4215 5769
rect 4157 5760 4169 5763
rect 4028 5732 4169 5760
rect 4028 5720 4034 5732
rect 4157 5729 4169 5732
rect 4203 5729 4215 5763
rect 4157 5723 4215 5729
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5729 6607 5763
rect 12250 5760 12256 5772
rect 11546 5732 12256 5760
rect 6549 5723 6607 5729
rect 12250 5720 12256 5732
rect 12308 5720 12314 5772
rect 12621 5763 12679 5769
rect 12621 5729 12633 5763
rect 12667 5760 12679 5763
rect 12710 5760 12716 5772
rect 12667 5732 12716 5760
rect 12667 5729 12679 5732
rect 12621 5723 12679 5729
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 14108 5769 14136 5800
rect 14366 5788 14372 5840
rect 14424 5788 14430 5840
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5729 14151 5763
rect 14384 5760 14412 5788
rect 15102 5760 15108 5772
rect 14384 5732 15108 5760
rect 14093 5723 14151 5729
rect 15102 5720 15108 5732
rect 15160 5760 15166 5772
rect 15657 5763 15715 5769
rect 15657 5760 15669 5763
rect 15160 5732 15669 5760
rect 15160 5720 15166 5732
rect 15657 5729 15669 5732
rect 15703 5729 15715 5763
rect 15657 5723 15715 5729
rect 16942 5720 16948 5772
rect 17000 5760 17006 5772
rect 17865 5763 17923 5769
rect 17865 5760 17877 5763
rect 17000 5732 17877 5760
rect 17000 5720 17006 5732
rect 17865 5729 17877 5732
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 19245 5763 19303 5769
rect 19245 5729 19257 5763
rect 19291 5760 19303 5763
rect 19426 5760 19432 5772
rect 19291 5732 19432 5760
rect 19291 5729 19303 5732
rect 19245 5723 19303 5729
rect 19426 5720 19432 5732
rect 19484 5720 19490 5772
rect 6270 5692 6276 5704
rect 6231 5664 6276 5692
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5661 6515 5695
rect 6457 5655 6515 5661
rect 2124 5627 2182 5633
rect 2124 5593 2136 5627
rect 2170 5624 2182 5627
rect 2682 5624 2688 5636
rect 2170 5596 2688 5624
rect 2170 5593 2182 5596
rect 2124 5587 2182 5593
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 4424 5627 4482 5633
rect 4424 5593 4436 5627
rect 4470 5624 4482 5627
rect 4706 5624 4712 5636
rect 4470 5596 4712 5624
rect 4470 5593 4482 5596
rect 4424 5587 4482 5593
rect 4706 5584 4712 5596
rect 4764 5584 4770 5636
rect 6362 5584 6368 5636
rect 6420 5624 6426 5636
rect 6472 5624 6500 5655
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 6822 5692 6828 5704
rect 6696 5664 6741 5692
rect 6783 5664 6828 5692
rect 6696 5652 6702 5664
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 13262 5692 13268 5704
rect 10060 5664 13268 5692
rect 8386 5624 8392 5636
rect 6420 5596 8392 5624
rect 6420 5584 6426 5596
rect 8386 5584 8392 5596
rect 8444 5584 8450 5636
rect 7006 5556 7012 5568
rect 6967 5528 7012 5556
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 10060 5565 10088 5664
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 13357 5695 13415 5701
rect 13357 5661 13369 5695
rect 13403 5661 13415 5695
rect 13357 5655 13415 5661
rect 10226 5624 10232 5636
rect 10187 5596 10232 5624
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 10594 5624 10600 5636
rect 10555 5596 10600 5624
rect 10594 5584 10600 5596
rect 10652 5584 10658 5636
rect 10962 5624 10968 5636
rect 10923 5596 10968 5624
rect 10962 5584 10968 5596
rect 11020 5584 11026 5636
rect 11057 5627 11115 5633
rect 11057 5593 11069 5627
rect 11103 5624 11115 5627
rect 11422 5624 11428 5636
rect 11103 5596 11428 5624
rect 11103 5593 11115 5596
rect 11057 5587 11115 5593
rect 11422 5584 11428 5596
rect 11480 5584 11486 5636
rect 11790 5584 11796 5636
rect 11848 5624 11854 5636
rect 12437 5627 12495 5633
rect 12437 5624 12449 5627
rect 11848 5596 12449 5624
rect 11848 5584 11854 5596
rect 12437 5593 12449 5596
rect 12483 5593 12495 5627
rect 12437 5587 12495 5593
rect 12802 5584 12808 5636
rect 12860 5624 12866 5636
rect 13372 5624 13400 5655
rect 13446 5652 13452 5704
rect 13504 5692 13510 5704
rect 13541 5695 13599 5701
rect 13541 5692 13553 5695
rect 13504 5664 13553 5692
rect 13504 5652 13510 5664
rect 13541 5661 13553 5664
rect 13587 5661 13599 5695
rect 13541 5655 13599 5661
rect 12860 5596 13400 5624
rect 13556 5624 13584 5655
rect 13722 5652 13728 5704
rect 13780 5692 13786 5704
rect 14185 5695 14243 5701
rect 14185 5692 14197 5695
rect 13780 5664 14197 5692
rect 13780 5652 13786 5664
rect 14185 5661 14197 5664
rect 14231 5661 14243 5695
rect 14369 5695 14427 5701
rect 14369 5692 14381 5695
rect 14185 5655 14243 5661
rect 14292 5664 14381 5692
rect 14292 5624 14320 5664
rect 14369 5661 14381 5664
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 15197 5695 15255 5701
rect 15197 5661 15209 5695
rect 15243 5661 15255 5695
rect 15197 5655 15255 5661
rect 15212 5624 15240 5655
rect 15746 5652 15752 5704
rect 15804 5692 15810 5704
rect 15913 5695 15971 5701
rect 15913 5692 15925 5695
rect 15804 5664 15925 5692
rect 15804 5652 15810 5664
rect 15913 5661 15925 5664
rect 15959 5661 15971 5695
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 15913 5655 15971 5661
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 17678 5692 17684 5704
rect 17639 5664 17684 5692
rect 17678 5652 17684 5664
rect 17736 5652 17742 5704
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5661 17831 5695
rect 18046 5692 18052 5704
rect 18007 5664 18052 5692
rect 17773 5655 17831 5661
rect 13556 5596 14320 5624
rect 14384 5596 15240 5624
rect 12860 5584 12866 5596
rect 10045 5559 10103 5565
rect 10045 5525 10057 5559
rect 10091 5525 10103 5559
rect 10045 5519 10103 5525
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 10836 5528 11345 5556
rect 10836 5516 10842 5528
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 12342 5556 12348 5568
rect 12303 5528 12348 5556
rect 11333 5519 11391 5525
rect 12342 5516 12348 5528
rect 12400 5516 12406 5568
rect 13262 5516 13268 5568
rect 13320 5556 13326 5568
rect 14384 5556 14412 5596
rect 16850 5584 16856 5636
rect 16908 5624 16914 5636
rect 17788 5624 17816 5655
rect 18046 5652 18052 5664
rect 18104 5652 18110 5704
rect 19521 5695 19579 5701
rect 19521 5661 19533 5695
rect 19567 5661 19579 5695
rect 20714 5692 20720 5704
rect 20675 5664 20720 5692
rect 19521 5655 19579 5661
rect 18230 5624 18236 5636
rect 16908 5596 18236 5624
rect 16908 5584 16914 5596
rect 18230 5584 18236 5596
rect 18288 5624 18294 5636
rect 19536 5624 19564 5655
rect 20714 5652 20720 5664
rect 20772 5652 20778 5704
rect 29730 5652 29736 5704
rect 29788 5692 29794 5704
rect 29825 5695 29883 5701
rect 29825 5692 29837 5695
rect 29788 5664 29837 5692
rect 29788 5652 29794 5664
rect 29825 5661 29837 5664
rect 29871 5661 29883 5695
rect 29825 5655 29883 5661
rect 19702 5624 19708 5636
rect 18288 5596 19708 5624
rect 18288 5584 18294 5596
rect 19702 5584 19708 5596
rect 19760 5584 19766 5636
rect 14550 5556 14556 5568
rect 13320 5528 14412 5556
rect 14511 5528 14556 5556
rect 13320 5516 13326 5528
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 1104 5466 30820 5488
rect 1104 5414 10880 5466
rect 10932 5414 10944 5466
rect 10996 5414 11008 5466
rect 11060 5414 11072 5466
rect 11124 5414 11136 5466
rect 11188 5414 20811 5466
rect 20863 5414 20875 5466
rect 20927 5414 20939 5466
rect 20991 5414 21003 5466
rect 21055 5414 21067 5466
rect 21119 5414 30820 5466
rect 1104 5392 30820 5414
rect 2682 5352 2688 5364
rect 2643 5324 2688 5352
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 3234 5352 3240 5364
rect 2884 5324 3240 5352
rect 2884 5225 2912 5324
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 4154 5312 4160 5364
rect 4212 5312 4218 5364
rect 4706 5352 4712 5364
rect 4667 5324 4712 5352
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 6641 5355 6699 5361
rect 6641 5321 6653 5355
rect 6687 5352 6699 5355
rect 6822 5352 6828 5364
rect 6687 5324 6828 5352
rect 6687 5321 6699 5324
rect 6641 5315 6699 5321
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 11609 5355 11667 5361
rect 11609 5321 11621 5355
rect 11655 5352 11667 5355
rect 12342 5352 12348 5364
rect 11655 5324 12348 5352
rect 11655 5321 11667 5324
rect 11609 5315 11667 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12986 5352 12992 5364
rect 12947 5324 12992 5352
rect 12986 5312 12992 5324
rect 13044 5312 13050 5364
rect 13357 5355 13415 5361
rect 13357 5321 13369 5355
rect 13403 5352 13415 5355
rect 14550 5352 14556 5364
rect 13403 5324 14556 5352
rect 13403 5321 13415 5324
rect 13357 5315 13415 5321
rect 14550 5312 14556 5324
rect 14608 5312 14614 5364
rect 14642 5312 14648 5364
rect 14700 5352 14706 5364
rect 15105 5355 15163 5361
rect 15105 5352 15117 5355
rect 14700 5324 15117 5352
rect 14700 5312 14706 5324
rect 15105 5321 15117 5324
rect 15151 5321 15163 5355
rect 15105 5315 15163 5321
rect 19889 5355 19947 5361
rect 19889 5321 19901 5355
rect 19935 5352 19947 5355
rect 20622 5352 20628 5364
rect 19935 5324 20628 5352
rect 19935 5321 19947 5324
rect 19889 5315 19947 5321
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 30006 5352 30012 5364
rect 29967 5324 30012 5352
rect 30006 5312 30012 5324
rect 30064 5312 30070 5364
rect 3050 5244 3056 5296
rect 3108 5284 3114 5296
rect 3881 5287 3939 5293
rect 3881 5284 3893 5287
rect 3108 5256 3188 5284
rect 3108 5244 3114 5256
rect 3160 5225 3188 5256
rect 3252 5256 3893 5284
rect 3252 5225 3280 5256
rect 3881 5253 3893 5256
rect 3927 5253 3939 5287
rect 4172 5284 4200 5312
rect 4172 5256 5396 5284
rect 3881 5247 3939 5253
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5185 2927 5219
rect 2869 5179 2927 5185
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5216 3479 5219
rect 3510 5216 3516 5228
rect 3467 5188 3516 5216
rect 3467 5185 3479 5188
rect 3421 5179 3479 5185
rect 3510 5176 3516 5188
rect 3568 5216 3574 5228
rect 3970 5216 3976 5228
rect 3568 5188 3976 5216
rect 3568 5176 3574 5188
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4154 5216 4160 5228
rect 4115 5188 4160 5216
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 4246 5176 4252 5228
rect 4304 5216 4310 5228
rect 5368 5225 5396 5256
rect 7006 5244 7012 5296
rect 7064 5284 7070 5296
rect 7754 5287 7812 5293
rect 7754 5284 7766 5287
rect 7064 5256 7766 5284
rect 7064 5244 7070 5256
rect 7754 5253 7766 5256
rect 7800 5253 7812 5287
rect 9398 5284 9404 5296
rect 7754 5247 7812 5253
rect 7852 5256 9404 5284
rect 4525 5219 4583 5225
rect 4304 5188 4349 5216
rect 4304 5176 4310 5188
rect 4525 5185 4537 5219
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 5353 5219 5411 5225
rect 5353 5185 5365 5219
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5148 1731 5151
rect 3053 5151 3111 5157
rect 1719 5120 2774 5148
rect 1719 5117 1731 5120
rect 1673 5111 1731 5117
rect 2746 5012 2774 5120
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3786 5148 3792 5160
rect 3099 5120 3792 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 3786 5108 3792 5120
rect 3844 5148 3850 5160
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 3844 5120 4353 5148
rect 3844 5108 3850 5120
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4540 5148 4568 5179
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 7852 5216 7880 5256
rect 9398 5244 9404 5256
rect 9456 5244 9462 5296
rect 21024 5287 21082 5293
rect 21024 5253 21036 5287
rect 21070 5284 21082 5287
rect 21174 5284 21180 5296
rect 21070 5256 21180 5284
rect 21070 5253 21082 5256
rect 21024 5247 21082 5253
rect 21174 5244 21180 5256
rect 21232 5244 21238 5296
rect 6512 5188 7880 5216
rect 6512 5176 6518 5188
rect 8386 5176 8392 5228
rect 8444 5216 8450 5228
rect 8737 5219 8795 5225
rect 8737 5216 8749 5219
rect 8444 5188 8749 5216
rect 8444 5176 8450 5188
rect 8737 5185 8749 5188
rect 8783 5185 8795 5219
rect 8737 5179 8795 5185
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5216 10839 5219
rect 11330 5216 11336 5228
rect 10827 5188 11336 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 11790 5216 11796 5228
rect 11751 5188 11796 5216
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12023 5188 12434 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12406 5160 12434 5188
rect 12710 5176 12716 5228
rect 12768 5216 12774 5228
rect 13078 5216 13084 5228
rect 12768 5188 13084 5216
rect 12768 5176 12774 5188
rect 13078 5176 13084 5188
rect 13136 5216 13142 5228
rect 14366 5216 14372 5228
rect 13136 5188 13584 5216
rect 14327 5188 14372 5216
rect 13136 5176 13142 5188
rect 5718 5148 5724 5160
rect 4540 5120 5724 5148
rect 4341 5111 4399 5117
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5148 8079 5151
rect 8481 5151 8539 5157
rect 8481 5148 8493 5151
rect 8067 5120 8493 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 8481 5117 8493 5120
rect 8527 5117 8539 5151
rect 8481 5111 8539 5117
rect 12069 5151 12127 5157
rect 12069 5117 12081 5151
rect 12115 5148 12127 5151
rect 12250 5148 12256 5160
rect 12115 5120 12256 5148
rect 12115 5117 12127 5120
rect 12069 5111 12127 5117
rect 3881 5083 3939 5089
rect 3881 5049 3893 5083
rect 3927 5080 3939 5083
rect 5169 5083 5227 5089
rect 5169 5080 5181 5083
rect 3927 5052 5181 5080
rect 3927 5049 3939 5052
rect 3881 5043 3939 5049
rect 5169 5049 5181 5052
rect 5215 5049 5227 5083
rect 5169 5043 5227 5049
rect 4062 5012 4068 5024
rect 2746 4984 4068 5012
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 8018 5012 8024 5024
rect 4212 4984 8024 5012
rect 4212 4972 4218 4984
rect 8018 4972 8024 4984
rect 8076 4972 8082 5024
rect 8496 5012 8524 5111
rect 12250 5108 12256 5120
rect 12308 5108 12314 5160
rect 12406 5120 12440 5160
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 13446 5148 13452 5160
rect 13359 5120 13452 5148
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 13556 5157 13584 5188
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 15194 5176 15200 5228
rect 15252 5216 15258 5228
rect 15289 5219 15347 5225
rect 15289 5216 15301 5219
rect 15252 5188 15301 5216
rect 15252 5176 15258 5188
rect 15289 5185 15301 5188
rect 15335 5185 15347 5219
rect 15289 5179 15347 5185
rect 15378 5176 15384 5228
rect 15436 5216 15442 5228
rect 15473 5219 15531 5225
rect 15473 5216 15485 5219
rect 15436 5188 15485 5216
rect 15436 5176 15442 5188
rect 15473 5185 15485 5188
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 15841 5219 15899 5225
rect 15841 5185 15853 5219
rect 15887 5216 15899 5219
rect 16206 5216 16212 5228
rect 15887 5188 16212 5216
rect 15887 5185 15899 5188
rect 15841 5179 15899 5185
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5117 13599 5151
rect 15562 5148 15568 5160
rect 15523 5120 15568 5148
rect 13541 5111 13599 5117
rect 15562 5108 15568 5120
rect 15620 5108 15626 5160
rect 15672 5148 15700 5179
rect 16206 5176 16212 5188
rect 16264 5176 16270 5228
rect 17310 5216 17316 5228
rect 17271 5188 17316 5216
rect 17310 5176 17316 5188
rect 17368 5176 17374 5228
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5216 18383 5219
rect 19242 5216 19248 5228
rect 18371 5188 19248 5216
rect 18371 5185 18383 5188
rect 18325 5179 18383 5185
rect 19242 5176 19248 5188
rect 19300 5176 19306 5228
rect 19610 5176 19616 5228
rect 19668 5216 19674 5228
rect 21269 5219 21327 5225
rect 21269 5216 21281 5219
rect 19668 5188 21281 5216
rect 19668 5176 19674 5188
rect 21269 5185 21281 5188
rect 21315 5216 21327 5219
rect 21818 5216 21824 5228
rect 21315 5188 21824 5216
rect 21315 5185 21327 5188
rect 21269 5179 21327 5185
rect 21818 5176 21824 5188
rect 21876 5176 21882 5228
rect 29822 5216 29828 5228
rect 29783 5188 29828 5216
rect 29822 5176 29828 5188
rect 29880 5176 29886 5228
rect 16666 5148 16672 5160
rect 15672 5120 16672 5148
rect 16666 5108 16672 5120
rect 16724 5108 16730 5160
rect 17589 5151 17647 5157
rect 17589 5117 17601 5151
rect 17635 5148 17647 5151
rect 17954 5148 17960 5160
rect 17635 5120 17960 5148
rect 17635 5117 17647 5120
rect 17589 5111 17647 5117
rect 17954 5108 17960 5120
rect 18012 5148 18018 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 18012 5120 18061 5148
rect 18012 5108 18018 5120
rect 18049 5117 18061 5120
rect 18095 5148 18107 5151
rect 18782 5148 18788 5160
rect 18095 5120 18788 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 18782 5108 18788 5120
rect 18840 5108 18846 5160
rect 10965 5083 11023 5089
rect 10965 5049 10977 5083
rect 11011 5080 11023 5083
rect 13464 5080 13492 5108
rect 11011 5052 13492 5080
rect 11011 5049 11023 5052
rect 10965 5043 11023 5049
rect 13906 5040 13912 5092
rect 13964 5080 13970 5092
rect 14185 5083 14243 5089
rect 14185 5080 14197 5083
rect 13964 5052 14197 5080
rect 13964 5040 13970 5052
rect 14185 5049 14197 5052
rect 14231 5080 14243 5083
rect 17497 5083 17555 5089
rect 17497 5080 17509 5083
rect 14231 5052 17509 5080
rect 14231 5049 14243 5052
rect 14185 5043 14243 5049
rect 17497 5049 17509 5052
rect 17543 5080 17555 5083
rect 18141 5083 18199 5089
rect 18141 5080 18153 5083
rect 17543 5052 18153 5080
rect 17543 5049 17555 5052
rect 17497 5043 17555 5049
rect 18141 5049 18153 5052
rect 18187 5080 18199 5083
rect 18598 5080 18604 5092
rect 18187 5052 18604 5080
rect 18187 5049 18199 5052
rect 18141 5043 18199 5049
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 8662 5012 8668 5024
rect 8496 4984 8668 5012
rect 8662 4972 8668 4984
rect 8720 5012 8726 5024
rect 9398 5012 9404 5024
rect 8720 4984 9404 5012
rect 8720 4972 8726 4984
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 9858 5012 9864 5024
rect 9819 4984 9864 5012
rect 9858 4972 9864 4984
rect 9916 5012 9922 5024
rect 10594 5012 10600 5024
rect 9916 4984 10600 5012
rect 9916 4972 9922 4984
rect 10594 4972 10600 4984
rect 10652 4972 10658 5024
rect 17126 5012 17132 5024
rect 17087 4984 17132 5012
rect 17126 4972 17132 4984
rect 17184 4972 17190 5024
rect 18506 5012 18512 5024
rect 18467 4984 18512 5012
rect 18506 4972 18512 4984
rect 18564 4972 18570 5024
rect 1104 4922 30820 4944
rect 1104 4870 5915 4922
rect 5967 4870 5979 4922
rect 6031 4870 6043 4922
rect 6095 4870 6107 4922
rect 6159 4870 6171 4922
rect 6223 4870 15846 4922
rect 15898 4870 15910 4922
rect 15962 4870 15974 4922
rect 16026 4870 16038 4922
rect 16090 4870 16102 4922
rect 16154 4870 25776 4922
rect 25828 4870 25840 4922
rect 25892 4870 25904 4922
rect 25956 4870 25968 4922
rect 26020 4870 26032 4922
rect 26084 4870 30820 4922
rect 1104 4848 30820 4870
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 3878 4808 3884 4820
rect 2915 4780 3884 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 4982 4808 4988 4820
rect 4120 4780 4988 4808
rect 4120 4768 4126 4780
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 5810 4808 5816 4820
rect 5368 4780 5816 4808
rect 1210 4632 1216 4684
rect 1268 4672 1274 4684
rect 1397 4675 1455 4681
rect 1397 4672 1409 4675
rect 1268 4644 1409 4672
rect 1268 4632 1274 4644
rect 1397 4641 1409 4644
rect 1443 4641 1455 4675
rect 1397 4635 1455 4641
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4672 1731 4675
rect 4154 4672 4160 4684
rect 1719 4644 4160 4672
rect 1719 4641 1731 4644
rect 1673 4635 1731 4641
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 2774 4604 2780 4616
rect 2731 4576 2780 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 5368 4613 5396 4780
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 8386 4808 8392 4820
rect 8347 4780 8392 4808
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 10686 4768 10692 4820
rect 10744 4808 10750 4820
rect 11333 4811 11391 4817
rect 11333 4808 11345 4811
rect 10744 4780 11345 4808
rect 10744 4768 10750 4780
rect 11333 4777 11345 4780
rect 11379 4777 11391 4811
rect 11333 4771 11391 4777
rect 15010 4768 15016 4820
rect 15068 4808 15074 4820
rect 15105 4811 15163 4817
rect 15105 4808 15117 4811
rect 15068 4780 15117 4808
rect 15068 4768 15074 4780
rect 15105 4777 15117 4780
rect 15151 4777 15163 4811
rect 17954 4808 17960 4820
rect 15105 4771 15163 4777
rect 15488 4780 17960 4808
rect 5626 4700 5632 4752
rect 5684 4700 5690 4752
rect 6638 4700 6644 4752
rect 6696 4740 6702 4752
rect 8478 4740 8484 4752
rect 6696 4712 6776 4740
rect 6696 4700 6702 4712
rect 5537 4675 5595 4681
rect 5537 4641 5549 4675
rect 5583 4672 5595 4675
rect 5644 4672 5672 4700
rect 6748 4681 6776 4712
rect 7760 4712 8484 4740
rect 6733 4675 6791 4681
rect 6733 4672 6745 4675
rect 5583 4644 6745 4672
rect 5583 4641 5595 4644
rect 5537 4635 5595 4641
rect 6733 4641 6745 4644
rect 6779 4641 6791 4675
rect 7098 4672 7104 4684
rect 6733 4635 6791 4641
rect 6840 4644 7104 4672
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4604 5963 4607
rect 6270 4604 6276 4616
rect 5951 4576 6276 4604
rect 5951 4573 5963 4576
rect 5905 4567 5963 4573
rect 4522 4496 4528 4548
rect 4580 4536 4586 4548
rect 5644 4536 5672 4567
rect 4580 4508 5672 4536
rect 5736 4536 5764 4567
rect 6270 4564 6276 4576
rect 6328 4604 6334 4616
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 6328 4576 6377 4604
rect 6328 4564 6334 4576
rect 6365 4573 6377 4576
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 6178 4536 6184 4548
rect 5736 4508 6184 4536
rect 4580 4496 4586 4508
rect 6178 4496 6184 4508
rect 6236 4536 6242 4548
rect 6454 4536 6460 4548
rect 6236 4508 6460 4536
rect 6236 4496 6242 4508
rect 6454 4496 6460 4508
rect 6512 4496 6518 4548
rect 6564 4536 6592 4567
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 6696 4576 6741 4604
rect 6696 4564 6702 4576
rect 6840 4536 6868 4644
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7760 4672 7788 4712
rect 8478 4700 8484 4712
rect 8536 4700 8542 4752
rect 14458 4700 14464 4752
rect 14516 4740 14522 4752
rect 14645 4743 14703 4749
rect 14645 4740 14657 4743
rect 14516 4712 14657 4740
rect 14516 4700 14522 4712
rect 14645 4709 14657 4712
rect 14691 4740 14703 4743
rect 15488 4740 15516 4780
rect 17954 4768 17960 4780
rect 18012 4768 18018 4820
rect 19794 4808 19800 4820
rect 18156 4780 19334 4808
rect 17221 4743 17279 4749
rect 17221 4740 17233 4743
rect 14691 4712 15516 4740
rect 15580 4712 17233 4740
rect 14691 4709 14703 4712
rect 14645 4703 14703 4709
rect 7926 4672 7932 4684
rect 7668 4644 7788 4672
rect 7887 4644 7932 4672
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 7558 4604 7564 4616
rect 6963 4576 7564 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7558 4564 7564 4576
rect 7616 4564 7622 4616
rect 7668 4613 7696 4644
rect 7926 4632 7932 4644
rect 7984 4632 7990 4684
rect 9858 4672 9864 4684
rect 8220 4644 9864 4672
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4573 7711 4607
rect 7834 4604 7840 4616
rect 7795 4576 7840 4604
rect 7653 4567 7711 4573
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4604 8079 4607
rect 8110 4604 8116 4616
rect 8067 4576 8116 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8220 4613 8248 4644
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 10778 4672 10784 4684
rect 10612 4644 10784 4672
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 8478 4564 8484 4616
rect 8536 4604 8542 4616
rect 8846 4604 8852 4616
rect 8536 4576 8852 4604
rect 8536 4564 8542 4576
rect 8846 4564 8852 4576
rect 8904 4604 8910 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8904 4576 8953 4604
rect 8904 4564 8910 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 6564 4508 6868 4536
rect 5166 4468 5172 4480
rect 5127 4440 5172 4468
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 5718 4428 5724 4480
rect 5776 4468 5782 4480
rect 6564 4468 6592 4508
rect 8662 4496 8668 4548
rect 8720 4536 8726 4548
rect 9140 4536 9168 4567
rect 8720 4508 9168 4536
rect 9232 4536 9260 4567
rect 9306 4564 9312 4616
rect 9364 4604 9370 4616
rect 9493 4607 9551 4613
rect 9364 4576 9409 4604
rect 9364 4564 9370 4576
rect 9493 4573 9505 4607
rect 9539 4604 9551 4607
rect 10612 4604 10640 4644
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 13265 4675 13323 4681
rect 13265 4672 13277 4675
rect 12308 4644 13277 4672
rect 12308 4632 12314 4644
rect 13265 4641 13277 4644
rect 13311 4641 13323 4675
rect 13265 4635 13323 4641
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 15580 4672 15608 4712
rect 17221 4709 17233 4712
rect 17267 4709 17279 4743
rect 18156 4740 18184 4780
rect 17221 4703 17279 4709
rect 17972 4712 18184 4740
rect 15746 4672 15752 4684
rect 15160 4644 15608 4672
rect 15707 4644 15752 4672
rect 15160 4632 15166 4644
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 16850 4672 16856 4684
rect 16500 4644 16856 4672
rect 9539 4576 10640 4604
rect 9539 4573 9551 4576
rect 9493 4567 9551 4573
rect 10686 4564 10692 4616
rect 10744 4604 10750 4616
rect 10744 4576 10789 4604
rect 10744 4564 10750 4576
rect 13170 4564 13176 4616
rect 13228 4604 13234 4616
rect 16500 4613 16528 4644
rect 16850 4632 16856 4644
rect 16908 4632 16914 4684
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 13228 4576 13553 4604
rect 13228 4564 13234 4576
rect 13541 4573 13553 4576
rect 13587 4604 13599 4607
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 13587 4576 14473 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 14461 4573 14473 4576
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 16485 4607 16543 4613
rect 16485 4573 16497 4607
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 16669 4607 16727 4613
rect 16669 4573 16681 4607
rect 16715 4573 16727 4607
rect 16669 4567 16727 4573
rect 16761 4607 16819 4613
rect 16761 4573 16773 4607
rect 16807 4604 16819 4607
rect 17034 4604 17040 4616
rect 16807 4576 17040 4604
rect 16807 4573 16819 4576
rect 16761 4567 16819 4573
rect 9582 4536 9588 4548
rect 9232 4508 9588 4536
rect 8720 4496 8726 4508
rect 7098 4468 7104 4480
rect 5776 4440 6592 4468
rect 7059 4440 7104 4468
rect 5776 4428 5782 4440
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 7926 4428 7932 4480
rect 7984 4468 7990 4480
rect 9232 4468 9260 4508
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 11514 4536 11520 4548
rect 11475 4508 11520 4536
rect 11514 4496 11520 4508
rect 11572 4496 11578 4548
rect 11698 4536 11704 4548
rect 11659 4508 11704 4536
rect 11698 4496 11704 4508
rect 11756 4496 11762 4548
rect 15473 4539 15531 4545
rect 15473 4505 15485 4539
rect 15519 4536 15531 4539
rect 16574 4536 16580 4548
rect 15519 4508 16580 4536
rect 15519 4505 15531 4508
rect 15473 4499 15531 4505
rect 16574 4496 16580 4508
rect 16632 4496 16638 4548
rect 16684 4536 16712 4567
rect 17034 4564 17040 4576
rect 17092 4564 17098 4616
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4573 17463 4607
rect 17405 4567 17463 4573
rect 16942 4536 16948 4548
rect 16684 4508 16948 4536
rect 16942 4496 16948 4508
rect 17000 4496 17006 4548
rect 7984 4440 9260 4468
rect 9677 4471 9735 4477
rect 7984 4428 7990 4440
rect 9677 4437 9689 4471
rect 9723 4468 9735 4471
rect 9766 4468 9772 4480
rect 9723 4440 9772 4468
rect 9723 4437 9735 4440
rect 9677 4431 9735 4437
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 10781 4471 10839 4477
rect 10781 4437 10793 4471
rect 10827 4468 10839 4471
rect 11238 4468 11244 4480
rect 10827 4440 11244 4468
rect 10827 4437 10839 4440
rect 10781 4431 10839 4437
rect 11238 4428 11244 4440
rect 11296 4428 11302 4480
rect 15562 4468 15568 4480
rect 15523 4440 15568 4468
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 16298 4468 16304 4480
rect 16259 4440 16304 4468
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 16390 4428 16396 4480
rect 16448 4468 16454 4480
rect 17420 4468 17448 4567
rect 17494 4564 17500 4616
rect 17552 4604 17558 4616
rect 17972 4613 18000 4712
rect 18230 4632 18236 4684
rect 18288 4672 18294 4684
rect 19306 4672 19334 4780
rect 19536 4780 19800 4808
rect 19426 4672 19432 4684
rect 18288 4644 18333 4672
rect 19306 4644 19432 4672
rect 18288 4632 18294 4644
rect 19426 4632 19432 4644
rect 19484 4632 19490 4684
rect 17957 4607 18015 4613
rect 17957 4604 17969 4607
rect 17552 4576 17969 4604
rect 17552 4564 17558 4576
rect 17957 4573 17969 4576
rect 18003 4573 18015 4607
rect 18138 4604 18144 4616
rect 18196 4613 18202 4616
rect 18103 4576 18144 4604
rect 17957 4567 18015 4573
rect 18138 4564 18144 4576
rect 18196 4567 18203 4613
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4573 18383 4607
rect 18325 4567 18383 4573
rect 18509 4607 18567 4613
rect 18509 4573 18521 4607
rect 18555 4604 18567 4607
rect 19536 4604 19564 4780
rect 19794 4768 19800 4780
rect 19852 4808 19858 4820
rect 21358 4808 21364 4820
rect 19852 4780 21364 4808
rect 19852 4768 19858 4780
rect 21358 4768 21364 4780
rect 21416 4768 21422 4820
rect 19610 4632 19616 4684
rect 19668 4672 19674 4684
rect 19668 4644 19713 4672
rect 19668 4632 19674 4644
rect 30098 4604 30104 4616
rect 18555 4576 19564 4604
rect 30059 4576 30104 4604
rect 18555 4573 18567 4576
rect 18509 4567 18567 4573
rect 18196 4564 18202 4567
rect 18340 4536 18368 4567
rect 30098 4564 30104 4576
rect 30156 4564 30162 4616
rect 19880 4539 19938 4545
rect 18340 4508 18828 4536
rect 18690 4468 18696 4480
rect 16448 4440 17448 4468
rect 18651 4440 18696 4468
rect 16448 4428 16454 4440
rect 18690 4428 18696 4440
rect 18748 4428 18754 4480
rect 18800 4468 18828 4508
rect 19880 4505 19892 4539
rect 19926 4536 19938 4539
rect 20162 4536 20168 4548
rect 19926 4508 20168 4536
rect 19926 4505 19938 4508
rect 19880 4499 19938 4505
rect 20162 4496 20168 4508
rect 20220 4496 20226 4548
rect 20438 4468 20444 4480
rect 18800 4440 20444 4468
rect 20438 4428 20444 4440
rect 20496 4428 20502 4480
rect 20714 4428 20720 4480
rect 20772 4468 20778 4480
rect 20993 4471 21051 4477
rect 20993 4468 21005 4471
rect 20772 4440 21005 4468
rect 20772 4428 20778 4440
rect 20993 4437 21005 4440
rect 21039 4437 21051 4471
rect 29914 4468 29920 4480
rect 29875 4440 29920 4468
rect 20993 4431 21051 4437
rect 29914 4428 29920 4440
rect 29972 4428 29978 4480
rect 1104 4378 30820 4400
rect 1104 4326 10880 4378
rect 10932 4326 10944 4378
rect 10996 4326 11008 4378
rect 11060 4326 11072 4378
rect 11124 4326 11136 4378
rect 11188 4326 20811 4378
rect 20863 4326 20875 4378
rect 20927 4326 20939 4378
rect 20991 4326 21003 4378
rect 21055 4326 21067 4378
rect 21119 4326 30820 4378
rect 1104 4304 30820 4326
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 4522 4264 4528 4276
rect 4304 4236 4528 4264
rect 4304 4224 4310 4236
rect 4522 4224 4528 4236
rect 4580 4224 4586 4276
rect 7558 4224 7564 4276
rect 7616 4264 7622 4276
rect 7745 4267 7803 4273
rect 7745 4264 7757 4267
rect 7616 4236 7757 4264
rect 7616 4224 7622 4236
rect 7745 4233 7757 4236
rect 7791 4233 7803 4267
rect 7745 4227 7803 4233
rect 12437 4267 12495 4273
rect 12437 4233 12449 4267
rect 12483 4264 12495 4267
rect 12894 4264 12900 4276
rect 12483 4236 12900 4264
rect 12483 4233 12495 4236
rect 12437 4227 12495 4233
rect 12894 4224 12900 4236
rect 12952 4224 12958 4276
rect 13170 4264 13176 4276
rect 13131 4236 13176 4264
rect 13170 4224 13176 4236
rect 13228 4224 13234 4276
rect 14918 4224 14924 4276
rect 14976 4264 14982 4276
rect 15013 4267 15071 4273
rect 15013 4264 15025 4267
rect 14976 4236 15025 4264
rect 14976 4224 14982 4236
rect 15013 4233 15025 4236
rect 15059 4233 15071 4267
rect 16666 4264 16672 4276
rect 16627 4236 16672 4264
rect 15013 4227 15071 4233
rect 16666 4224 16672 4236
rect 16724 4224 16730 4276
rect 19794 4264 19800 4276
rect 19755 4236 19800 4264
rect 19794 4224 19800 4236
rect 19852 4224 19858 4276
rect 20438 4224 20444 4276
rect 20496 4224 20502 4276
rect 20993 4267 21051 4273
rect 20993 4233 21005 4267
rect 21039 4264 21051 4267
rect 21174 4264 21180 4276
rect 21039 4236 21180 4264
rect 21039 4233 21051 4236
rect 20993 4227 21051 4233
rect 21174 4224 21180 4236
rect 21232 4224 21238 4276
rect 1854 4196 1860 4208
rect 1815 4168 1860 4196
rect 1854 4156 1860 4168
rect 1912 4156 1918 4208
rect 2225 4199 2283 4205
rect 2225 4165 2237 4199
rect 2271 4196 2283 4199
rect 3694 4196 3700 4208
rect 2271 4168 3700 4196
rect 2271 4165 2283 4168
rect 2225 4159 2283 4165
rect 3694 4156 3700 4168
rect 3752 4156 3758 4208
rect 7466 4196 7472 4208
rect 4448 4168 7472 4196
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2774 4128 2780 4140
rect 2731 4100 2780 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 2590 4020 2596 4072
rect 2648 4060 2654 4072
rect 3436 4060 3464 4091
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4448 4137 4476 4168
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 9674 4196 9680 4208
rect 9140 4168 9680 4196
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 4028 4100 4261 4128
rect 4028 4088 4034 4100
rect 4249 4097 4261 4100
rect 4295 4097 4307 4131
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 4249 4091 4307 4097
rect 4350 4100 4445 4128
rect 4350 4060 4378 4100
rect 4433 4097 4445 4100
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 4801 4131 4859 4137
rect 4801 4097 4813 4131
rect 4847 4128 4859 4131
rect 4890 4128 4896 4140
rect 4847 4100 4896 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 5592 4100 6377 4128
rect 5592 4088 5598 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 6632 4131 6690 4137
rect 6632 4097 6644 4131
rect 6678 4128 6690 4131
rect 7098 4128 7104 4140
rect 6678 4100 7104 4128
rect 6678 4097 6690 4100
rect 6632 4091 6690 4097
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 8846 4128 8852 4140
rect 8807 4100 8852 4128
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 9030 4128 9036 4140
rect 8991 4100 9036 4128
rect 9030 4088 9036 4100
rect 9088 4088 9094 4140
rect 9140 4137 9168 4168
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 11882 4156 11888 4208
rect 11940 4196 11946 4208
rect 15378 4196 15384 4208
rect 11940 4168 12112 4196
rect 15339 4168 15384 4196
rect 11940 4156 11946 4168
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4128 9275 4131
rect 9306 4128 9312 4140
rect 9263 4100 9312 4128
rect 9263 4097 9275 4100
rect 9217 4091 9275 4097
rect 4522 4060 4528 4072
rect 2648 4032 3464 4060
rect 3528 4032 4378 4060
rect 4483 4032 4528 4060
rect 2648 4020 2654 4032
rect 2869 3995 2927 4001
rect 2869 3961 2881 3995
rect 2915 3992 2927 3995
rect 3528 3992 3556 4032
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 4617 4063 4675 4069
rect 4617 4029 4629 4063
rect 4663 4060 4675 4063
rect 5626 4060 5632 4072
rect 4663 4032 5632 4060
rect 4663 4029 4675 4032
rect 4617 4023 4675 4029
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 9232 4060 9260 4091
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 9490 4128 9496 4140
rect 9447 4100 9496 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 9640 4100 10149 4128
rect 9640 4088 9646 4100
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10226 4088 10232 4140
rect 10284 4128 10290 4140
rect 10781 4131 10839 4137
rect 10781 4128 10793 4131
rect 10284 4100 10793 4128
rect 10284 4088 10290 4100
rect 10781 4097 10793 4100
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 11054 4088 11060 4140
rect 11112 4128 11118 4140
rect 11974 4128 11980 4140
rect 11112 4100 11980 4128
rect 11112 4088 11118 4100
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 12084 4137 12112 4168
rect 15378 4156 15384 4168
rect 15436 4156 15442 4208
rect 17037 4199 17095 4205
rect 17037 4165 17049 4199
rect 17083 4196 17095 4199
rect 18414 4196 18420 4208
rect 17083 4168 18420 4196
rect 17083 4165 17095 4168
rect 17037 4159 17095 4165
rect 18414 4156 18420 4168
rect 18472 4156 18478 4208
rect 18690 4205 18696 4208
rect 18684 4196 18696 4205
rect 18651 4168 18696 4196
rect 18684 4159 18696 4168
rect 18690 4156 18696 4159
rect 18748 4156 18754 4208
rect 20456 4196 20484 4224
rect 20456 4168 20576 4196
rect 12069 4131 12127 4137
rect 12069 4097 12081 4131
rect 12115 4097 12127 4131
rect 12069 4091 12127 4097
rect 12250 4088 12256 4140
rect 12308 4128 12314 4140
rect 13173 4131 13231 4137
rect 12308 4100 13124 4128
rect 12308 4088 12314 4100
rect 8352 4032 9260 4060
rect 10873 4063 10931 4069
rect 8352 4020 8358 4032
rect 10873 4029 10885 4063
rect 10919 4060 10931 4063
rect 11606 4060 11612 4072
rect 10919 4032 11612 4060
rect 10919 4029 10931 4032
rect 10873 4023 10931 4029
rect 11606 4020 11612 4032
rect 11664 4060 11670 4072
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 11664 4032 12173 4060
rect 11664 4020 11670 4032
rect 12161 4029 12173 4032
rect 12207 4060 12219 4063
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12207 4032 12909 4060
rect 12207 4029 12219 4032
rect 12161 4023 12219 4029
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 13096 4060 13124 4100
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 13354 4128 13360 4140
rect 13219 4100 13360 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 14366 4128 14372 4140
rect 13832 4100 14372 4128
rect 13832 4060 13860 4100
rect 14366 4088 14372 4100
rect 14424 4128 14430 4140
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14424 4100 14565 4128
rect 14424 4088 14430 4100
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 14553 4091 14611 4097
rect 15194 4088 15200 4140
rect 15252 4128 15258 4140
rect 15470 4128 15476 4140
rect 15252 4100 15476 4128
rect 15252 4088 15258 4100
rect 15470 4088 15476 4100
rect 15528 4088 15534 4140
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 18322 4128 18328 4140
rect 17175 4100 18328 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 18322 4088 18328 4100
rect 18380 4088 18386 4140
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 20257 4131 20315 4137
rect 20257 4128 20269 4131
rect 19484 4100 20269 4128
rect 19484 4088 19490 4100
rect 20257 4097 20269 4100
rect 20303 4097 20315 4131
rect 20438 4128 20444 4140
rect 20399 4100 20444 4128
rect 20257 4091 20315 4097
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 20548 4128 20576 4168
rect 20622 4156 20628 4208
rect 20680 4196 20686 4208
rect 20680 4168 20852 4196
rect 20680 4156 20686 4168
rect 20824 4137 20852 4168
rect 20809 4131 20867 4137
rect 20548 4100 20668 4128
rect 13096 4032 13860 4060
rect 14277 4063 14335 4069
rect 12897 4023 12955 4029
rect 14277 4029 14289 4063
rect 14323 4060 14335 4063
rect 14458 4060 14464 4072
rect 14323 4032 14464 4060
rect 14323 4029 14335 4032
rect 14277 4023 14335 4029
rect 14458 4020 14464 4032
rect 14516 4060 14522 4072
rect 15657 4063 15715 4069
rect 14516 4032 15516 4060
rect 14516 4020 14522 4032
rect 2915 3964 3556 3992
rect 3605 3995 3663 4001
rect 2915 3961 2927 3964
rect 2869 3955 2927 3961
rect 3605 3961 3617 3995
rect 3651 3992 3663 3995
rect 10686 3992 10692 4004
rect 3651 3964 6408 3992
rect 3651 3961 3663 3964
rect 3605 3955 3663 3961
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5074 3884 5080 3936
rect 5132 3924 5138 3936
rect 6270 3924 6276 3936
rect 5132 3896 6276 3924
rect 5132 3884 5138 3896
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 6380 3924 6408 3964
rect 9232 3964 10692 3992
rect 9232 3924 9260 3964
rect 10686 3952 10692 3964
rect 10744 3952 10750 4004
rect 13081 3995 13139 4001
rect 13081 3992 13093 3995
rect 12406 3964 13093 3992
rect 12406 3936 12434 3964
rect 13081 3961 13093 3964
rect 13127 3961 13139 3995
rect 15488 3992 15516 4032
rect 15657 4029 15669 4063
rect 15703 4060 15715 4063
rect 15746 4060 15752 4072
rect 15703 4032 15752 4060
rect 15703 4029 15715 4032
rect 15657 4023 15715 4029
rect 15746 4020 15752 4032
rect 15804 4060 15810 4072
rect 17221 4063 17279 4069
rect 17221 4060 17233 4063
rect 15804 4032 17233 4060
rect 15804 4020 15810 4032
rect 17221 4029 17233 4032
rect 17267 4060 17279 4063
rect 17402 4060 17408 4072
rect 17267 4032 17408 4060
rect 17267 4029 17279 4032
rect 17221 4023 17279 4029
rect 17402 4020 17408 4032
rect 17460 4020 17466 4072
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4029 18475 4063
rect 18417 4023 18475 4029
rect 16942 3992 16948 4004
rect 15488 3964 16948 3992
rect 13081 3955 13139 3961
rect 16942 3952 16948 3964
rect 17000 3952 17006 4004
rect 6380 3896 9260 3924
rect 9585 3927 9643 3933
rect 9585 3893 9597 3927
rect 9631 3924 9643 3927
rect 9674 3924 9680 3936
rect 9631 3896 9680 3924
rect 9631 3893 9643 3896
rect 9585 3887 9643 3893
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 10229 3927 10287 3933
rect 10229 3893 10241 3927
rect 10275 3924 10287 3927
rect 11054 3924 11060 3936
rect 10275 3896 11060 3924
rect 10275 3893 10287 3896
rect 10229 3887 10287 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 11296 3896 12081 3924
rect 11296 3884 11302 3896
rect 12069 3893 12081 3896
rect 12115 3924 12127 3927
rect 12342 3924 12348 3936
rect 12115 3896 12348 3924
rect 12115 3893 12127 3896
rect 12069 3887 12127 3893
rect 12342 3884 12348 3896
rect 12400 3896 12434 3936
rect 12400 3884 12406 3896
rect 14090 3884 14096 3936
rect 14148 3924 14154 3936
rect 16390 3924 16396 3936
rect 14148 3896 16396 3924
rect 14148 3884 14154 3896
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 18432 3924 18460 4023
rect 19702 4020 19708 4072
rect 19760 4060 19766 4072
rect 20640 4069 20668 4100
rect 20809 4097 20821 4131
rect 20855 4097 20867 4131
rect 20809 4091 20867 4097
rect 28537 4131 28595 4137
rect 28537 4097 28549 4131
rect 28583 4097 28595 4131
rect 28537 4091 28595 4097
rect 29181 4131 29239 4137
rect 29181 4097 29193 4131
rect 29227 4097 29239 4131
rect 29181 4091 29239 4097
rect 20533 4063 20591 4069
rect 20533 4060 20545 4063
rect 19760 4032 20545 4060
rect 19760 4020 19766 4032
rect 20533 4029 20545 4032
rect 20579 4029 20591 4063
rect 20533 4023 20591 4029
rect 20625 4063 20683 4069
rect 20625 4029 20637 4063
rect 20671 4029 20683 4063
rect 20625 4023 20683 4029
rect 19518 3952 19524 4004
rect 19576 3992 19582 4004
rect 23566 3992 23572 4004
rect 19576 3964 23572 3992
rect 19576 3952 19582 3964
rect 23566 3952 23572 3964
rect 23624 3952 23630 4004
rect 28552 3992 28580 4091
rect 29196 4060 29224 4091
rect 29730 4088 29736 4140
rect 29788 4128 29794 4140
rect 29825 4131 29883 4137
rect 29825 4128 29837 4131
rect 29788 4100 29837 4128
rect 29788 4088 29794 4100
rect 29825 4097 29837 4100
rect 29871 4097 29883 4131
rect 29825 4091 29883 4097
rect 30834 4060 30840 4072
rect 29196 4032 30840 4060
rect 30834 4020 30840 4032
rect 30892 4020 30898 4072
rect 31570 3992 31576 4004
rect 28552 3964 31576 3992
rect 31570 3952 31576 3964
rect 31628 3952 31634 4004
rect 19334 3924 19340 3936
rect 18432 3896 19340 3924
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 20530 3884 20536 3936
rect 20588 3924 20594 3936
rect 22922 3924 22928 3936
rect 20588 3896 22928 3924
rect 20588 3884 20594 3896
rect 22922 3884 22928 3896
rect 22980 3884 22986 3936
rect 28718 3924 28724 3936
rect 28679 3896 28724 3924
rect 28718 3884 28724 3896
rect 28776 3884 28782 3936
rect 29365 3927 29423 3933
rect 29365 3893 29377 3927
rect 29411 3924 29423 3927
rect 29546 3924 29552 3936
rect 29411 3896 29552 3924
rect 29411 3893 29423 3896
rect 29365 3887 29423 3893
rect 29546 3884 29552 3896
rect 29604 3884 29610 3936
rect 30006 3924 30012 3936
rect 29967 3896 30012 3924
rect 30006 3884 30012 3896
rect 30064 3884 30070 3936
rect 1104 3834 30820 3856
rect 1104 3782 5915 3834
rect 5967 3782 5979 3834
rect 6031 3782 6043 3834
rect 6095 3782 6107 3834
rect 6159 3782 6171 3834
rect 6223 3782 15846 3834
rect 15898 3782 15910 3834
rect 15962 3782 15974 3834
rect 16026 3782 16038 3834
rect 16090 3782 16102 3834
rect 16154 3782 25776 3834
rect 25828 3782 25840 3834
rect 25892 3782 25904 3834
rect 25956 3782 25968 3834
rect 26020 3782 26032 3834
rect 26084 3782 30820 3834
rect 1104 3760 30820 3782
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 3973 3723 4031 3729
rect 2179 3692 2774 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 2746 3584 2774 3692
rect 3973 3689 3985 3723
rect 4019 3720 4031 3723
rect 10226 3720 10232 3732
rect 4019 3692 10232 3720
rect 4019 3689 4031 3692
rect 3973 3683 4031 3689
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 10836 3692 10885 3720
rect 10836 3680 10842 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 10873 3683 10931 3689
rect 11238 3680 11244 3732
rect 11296 3720 11302 3732
rect 11609 3723 11667 3729
rect 11609 3720 11621 3723
rect 11296 3692 11621 3720
rect 11296 3680 11302 3692
rect 11609 3689 11621 3692
rect 11655 3689 11667 3723
rect 15654 3720 15660 3732
rect 15615 3692 15660 3720
rect 11609 3683 11667 3689
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 16758 3680 16764 3732
rect 16816 3720 16822 3732
rect 16853 3723 16911 3729
rect 16853 3720 16865 3723
rect 16816 3692 16865 3720
rect 16816 3680 16822 3692
rect 16853 3689 16865 3692
rect 16899 3689 16911 3723
rect 16853 3683 16911 3689
rect 16942 3680 16948 3732
rect 17000 3720 17006 3732
rect 18141 3723 18199 3729
rect 18141 3720 18153 3723
rect 17000 3692 18153 3720
rect 17000 3680 17006 3692
rect 18141 3689 18153 3692
rect 18187 3689 18199 3723
rect 18141 3683 18199 3689
rect 18414 3680 18420 3732
rect 18472 3720 18478 3732
rect 18509 3723 18567 3729
rect 18509 3720 18521 3723
rect 18472 3692 18521 3720
rect 18472 3680 18478 3692
rect 18509 3689 18521 3692
rect 18555 3689 18567 3723
rect 20162 3720 20168 3732
rect 20123 3692 20168 3720
rect 18509 3683 18567 3689
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20714 3680 20720 3732
rect 20772 3720 20778 3732
rect 20809 3723 20867 3729
rect 20809 3720 20821 3723
rect 20772 3692 20821 3720
rect 20772 3680 20778 3692
rect 20809 3689 20821 3692
rect 20855 3689 20867 3723
rect 22281 3723 22339 3729
rect 22281 3720 22293 3723
rect 20809 3683 20867 3689
rect 20916 3692 22293 3720
rect 3053 3655 3111 3661
rect 3053 3621 3065 3655
rect 3099 3652 3111 3655
rect 5074 3652 5080 3664
rect 3099 3624 5080 3652
rect 3099 3621 3111 3624
rect 3053 3615 3111 3621
rect 5074 3612 5080 3624
rect 5132 3612 5138 3664
rect 13078 3652 13084 3664
rect 13039 3624 13084 3652
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 17034 3652 17040 3664
rect 15028 3624 17040 3652
rect 2746 3556 3096 3584
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 2958 3516 2964 3528
rect 1903 3488 2964 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 2774 3408 2780 3460
rect 2832 3448 2838 3460
rect 2832 3420 2877 3448
rect 2832 3408 2838 3420
rect 3068 3380 3096 3556
rect 11606 3544 11612 3596
rect 11664 3584 11670 3596
rect 11701 3587 11759 3593
rect 11701 3584 11713 3587
rect 11664 3556 11713 3584
rect 11664 3544 11670 3556
rect 11701 3553 11713 3556
rect 11747 3584 11759 3587
rect 11747 3556 12296 3584
rect 11747 3553 11759 3556
rect 11701 3547 11759 3553
rect 3418 3476 3424 3528
rect 3476 3516 3482 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3476 3488 3801 3516
rect 3476 3476 3482 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 5123 3488 5580 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5552 3460 5580 3488
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9766 3525 9772 3528
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 9456 3488 9505 3516
rect 9456 3476 9462 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9760 3516 9772 3525
rect 9727 3488 9772 3516
rect 9493 3479 9551 3485
rect 9760 3479 9772 3488
rect 9766 3476 9772 3479
rect 9824 3476 9830 3528
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11793 3519 11851 3525
rect 11793 3516 11805 3519
rect 11572 3488 11805 3516
rect 11572 3476 11578 3488
rect 11793 3485 11805 3488
rect 11839 3516 11851 3519
rect 11974 3516 11980 3528
rect 11839 3488 11980 3516
rect 11839 3485 11851 3488
rect 11793 3479 11851 3485
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12268 3525 12296 3556
rect 13170 3544 13176 3596
rect 13228 3584 13234 3596
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 13228 3556 14105 3584
rect 13228 3544 13234 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 15028 3528 15056 3624
rect 17034 3612 17040 3624
rect 17092 3652 17098 3664
rect 17092 3624 18092 3652
rect 17092 3612 17098 3624
rect 15746 3544 15752 3596
rect 15804 3584 15810 3596
rect 16209 3587 16267 3593
rect 16209 3584 16221 3587
rect 15804 3556 16221 3584
rect 15804 3544 15810 3556
rect 16209 3553 16221 3556
rect 16255 3553 16267 3587
rect 17310 3584 17316 3596
rect 17271 3556 17316 3584
rect 16209 3547 16267 3553
rect 17310 3544 17316 3556
rect 17368 3544 17374 3596
rect 17402 3544 17408 3596
rect 17460 3584 17466 3596
rect 17954 3584 17960 3596
rect 17460 3556 17960 3584
rect 17460 3544 17466 3556
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 18064 3593 18092 3624
rect 20438 3612 20444 3664
rect 20496 3652 20502 3664
rect 20916 3652 20944 3692
rect 22281 3689 22293 3692
rect 22327 3689 22339 3723
rect 22922 3720 22928 3732
rect 22883 3692 22928 3720
rect 22281 3683 22339 3689
rect 22922 3680 22928 3692
rect 22980 3680 22986 3732
rect 20496 3624 20944 3652
rect 20496 3612 20502 3624
rect 20990 3612 20996 3664
rect 21048 3652 21054 3664
rect 21818 3652 21824 3664
rect 21048 3624 21824 3652
rect 21048 3612 21054 3624
rect 21818 3612 21824 3624
rect 21876 3612 21882 3664
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3553 18107 3587
rect 19702 3584 19708 3596
rect 19663 3556 19708 3584
rect 18049 3547 18107 3553
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 19797 3587 19855 3593
rect 19797 3553 19809 3587
rect 19843 3584 19855 3587
rect 20346 3584 20352 3596
rect 19843 3556 20352 3584
rect 19843 3553 19855 3556
rect 19797 3547 19855 3553
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3485 12311 3519
rect 12253 3479 12311 3485
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 12713 3519 12771 3525
rect 12713 3516 12725 3519
rect 12400 3488 12725 3516
rect 12400 3476 12406 3488
rect 12713 3485 12725 3488
rect 12759 3485 12771 3519
rect 12713 3479 12771 3485
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3516 13139 3519
rect 14369 3519 14427 3525
rect 13127 3488 14044 3516
rect 13127 3485 13139 3488
rect 13081 3479 13139 3485
rect 13188 3460 13216 3488
rect 5166 3408 5172 3460
rect 5224 3448 5230 3460
rect 5322 3451 5380 3457
rect 5322 3448 5334 3451
rect 5224 3420 5334 3448
rect 5224 3408 5230 3420
rect 5322 3417 5334 3420
rect 5368 3417 5380 3451
rect 5322 3411 5380 3417
rect 5534 3408 5540 3460
rect 5592 3408 5598 3460
rect 11330 3408 11336 3460
rect 11388 3448 11394 3460
rect 12434 3448 12440 3460
rect 11388 3420 12440 3448
rect 11388 3408 11394 3420
rect 12434 3408 12440 3420
rect 12492 3408 12498 3460
rect 13170 3408 13176 3460
rect 13228 3408 13234 3460
rect 5718 3380 5724 3392
rect 3068 3352 5724 3380
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 6457 3383 6515 3389
rect 6457 3380 6469 3383
rect 5868 3352 6469 3380
rect 5868 3340 5874 3352
rect 6457 3349 6469 3352
rect 6503 3349 6515 3383
rect 6457 3343 6515 3349
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 11425 3383 11483 3389
rect 11425 3380 11437 3383
rect 9640 3352 11437 3380
rect 9640 3340 9646 3352
rect 11425 3349 11437 3352
rect 11471 3349 11483 3383
rect 14016 3380 14044 3488
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 15010 3516 15016 3528
rect 14415 3488 15016 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 15010 3476 15016 3488
rect 15068 3476 15074 3528
rect 16025 3519 16083 3525
rect 16025 3485 16037 3519
rect 16071 3516 16083 3519
rect 16298 3516 16304 3528
rect 16071 3488 16304 3516
rect 16071 3485 16083 3488
rect 16025 3479 16083 3485
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 17126 3476 17132 3528
rect 17184 3516 17190 3528
rect 17221 3519 17279 3525
rect 17221 3516 17233 3519
rect 17184 3488 17233 3516
rect 17184 3476 17190 3488
rect 17221 3485 17233 3488
rect 17267 3485 17279 3519
rect 18322 3516 18328 3528
rect 18283 3488 18328 3516
rect 17221 3479 17279 3485
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 19426 3516 19432 3528
rect 19387 3488 19432 3516
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3516 19671 3519
rect 19886 3516 19892 3528
rect 19659 3488 19892 3516
rect 19659 3485 19671 3488
rect 19613 3479 19671 3485
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 19981 3519 20039 3525
rect 19981 3485 19993 3519
rect 20027 3516 20039 3519
rect 20806 3516 20812 3528
rect 20027 3488 20812 3516
rect 20027 3485 20039 3488
rect 19981 3479 20039 3485
rect 20806 3476 20812 3488
rect 20864 3476 20870 3528
rect 20901 3519 20959 3525
rect 20901 3485 20913 3519
rect 20947 3485 20959 3519
rect 20901 3479 20959 3485
rect 16117 3451 16175 3457
rect 16117 3417 16129 3451
rect 16163 3448 16175 3451
rect 16666 3448 16672 3460
rect 16163 3420 16672 3448
rect 16163 3417 16175 3420
rect 16117 3411 16175 3417
rect 16666 3408 16672 3420
rect 16724 3448 16730 3460
rect 16850 3448 16856 3460
rect 16724 3420 16856 3448
rect 16724 3408 16730 3420
rect 16850 3408 16856 3420
rect 16908 3408 16914 3460
rect 20916 3448 20944 3479
rect 20990 3476 20996 3528
rect 21048 3516 21054 3528
rect 21048 3488 21093 3516
rect 21048 3476 21054 3488
rect 21174 3476 21180 3528
rect 21232 3516 21238 3528
rect 22465 3519 22523 3525
rect 22465 3516 22477 3519
rect 21232 3488 22477 3516
rect 21232 3476 21238 3488
rect 22465 3485 22477 3488
rect 22511 3485 22523 3519
rect 22465 3479 22523 3485
rect 22554 3476 22560 3528
rect 22612 3516 22618 3528
rect 23109 3519 23167 3525
rect 23109 3516 23121 3519
rect 22612 3488 23121 3516
rect 22612 3476 22618 3488
rect 23109 3485 23121 3488
rect 23155 3485 23167 3519
rect 23109 3479 23167 3485
rect 27798 3476 27804 3528
rect 27856 3516 27862 3528
rect 28077 3519 28135 3525
rect 28077 3516 28089 3519
rect 27856 3488 28089 3516
rect 27856 3476 27862 3488
rect 28077 3485 28089 3488
rect 28123 3485 28135 3519
rect 28077 3479 28135 3485
rect 28534 3476 28540 3528
rect 28592 3516 28598 3528
rect 28813 3519 28871 3525
rect 28813 3516 28825 3519
rect 28592 3488 28825 3516
rect 28592 3476 28598 3488
rect 28813 3485 28825 3488
rect 28859 3485 28871 3519
rect 28813 3479 28871 3485
rect 29270 3476 29276 3528
rect 29328 3516 29334 3528
rect 29733 3519 29791 3525
rect 29733 3516 29745 3519
rect 29328 3488 29745 3516
rect 29328 3476 29334 3488
rect 29733 3485 29745 3488
rect 29779 3485 29791 3519
rect 29733 3479 29791 3485
rect 21358 3448 21364 3460
rect 16960 3420 20760 3448
rect 20916 3420 21364 3448
rect 16960 3380 16988 3420
rect 14016 3352 16988 3380
rect 11425 3343 11483 3349
rect 17126 3340 17132 3392
rect 17184 3380 17190 3392
rect 20625 3383 20683 3389
rect 20625 3380 20637 3383
rect 17184 3352 20637 3380
rect 17184 3340 17190 3352
rect 20625 3349 20637 3352
rect 20671 3349 20683 3383
rect 20732 3380 20760 3420
rect 21358 3408 21364 3420
rect 21416 3408 21422 3460
rect 21453 3451 21511 3457
rect 21453 3417 21465 3451
rect 21499 3417 21511 3451
rect 21453 3411 21511 3417
rect 21637 3451 21695 3457
rect 21637 3417 21649 3451
rect 21683 3417 21695 3451
rect 21637 3411 21695 3417
rect 21468 3380 21496 3411
rect 20732 3352 21496 3380
rect 21652 3380 21680 3411
rect 21818 3408 21824 3460
rect 21876 3448 21882 3460
rect 22738 3448 22744 3460
rect 21876 3420 22744 3448
rect 21876 3408 21882 3420
rect 22738 3408 22744 3420
rect 22796 3408 22802 3460
rect 22462 3380 22468 3392
rect 21652 3352 22468 3380
rect 20625 3343 20683 3349
rect 22462 3340 22468 3352
rect 22520 3380 22526 3392
rect 25682 3380 25688 3392
rect 22520 3352 25688 3380
rect 22520 3340 22526 3352
rect 25682 3340 25688 3352
rect 25740 3340 25746 3392
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 27893 3383 27951 3389
rect 27893 3380 27905 3383
rect 27764 3352 27905 3380
rect 27764 3340 27770 3352
rect 27893 3349 27905 3352
rect 27939 3349 27951 3383
rect 27893 3343 27951 3349
rect 27982 3340 27988 3392
rect 28040 3380 28046 3392
rect 28629 3383 28687 3389
rect 28629 3380 28641 3383
rect 28040 3352 28641 3380
rect 28040 3340 28046 3352
rect 28629 3349 28641 3352
rect 28675 3349 28687 3383
rect 28629 3343 28687 3349
rect 29549 3383 29607 3389
rect 29549 3349 29561 3383
rect 29595 3380 29607 3383
rect 29914 3380 29920 3392
rect 29595 3352 29920 3380
rect 29595 3349 29607 3352
rect 29549 3343 29607 3349
rect 29914 3340 29920 3352
rect 29972 3340 29978 3392
rect 1104 3290 30820 3312
rect 1104 3238 10880 3290
rect 10932 3238 10944 3290
rect 10996 3238 11008 3290
rect 11060 3238 11072 3290
rect 11124 3238 11136 3290
rect 11188 3238 20811 3290
rect 20863 3238 20875 3290
rect 20927 3238 20939 3290
rect 20991 3238 21003 3290
rect 21055 3238 21067 3290
rect 21119 3238 30820 3290
rect 1104 3216 30820 3238
rect 4798 3176 4804 3188
rect 3896 3148 4804 3176
rect 1857 3111 1915 3117
rect 1857 3077 1869 3111
rect 1903 3108 1915 3111
rect 2866 3108 2872 3120
rect 1903 3080 2872 3108
rect 1903 3077 1915 3080
rect 1857 3071 1915 3077
rect 2866 3068 2872 3080
rect 2924 3068 2930 3120
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 2832 3012 2877 3040
rect 2832 3000 2838 3012
rect 2133 2907 2191 2913
rect 2133 2873 2145 2907
rect 2179 2904 2191 2907
rect 3896 2904 3924 3148
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 4890 3136 4896 3188
rect 4948 3176 4954 3188
rect 5353 3179 5411 3185
rect 5353 3176 5365 3179
rect 4948 3148 5365 3176
rect 4948 3136 4954 3148
rect 5353 3145 5365 3148
rect 5399 3145 5411 3179
rect 5353 3139 5411 3145
rect 7469 3179 7527 3185
rect 7469 3145 7481 3179
rect 7515 3176 7527 3179
rect 9030 3176 9036 3188
rect 7515 3148 9036 3176
rect 7515 3145 7527 3148
rect 7469 3139 7527 3145
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 9548 3148 10793 3176
rect 9548 3136 9554 3148
rect 10781 3145 10793 3148
rect 10827 3176 10839 3179
rect 11422 3176 11428 3188
rect 10827 3148 11428 3176
rect 10827 3145 10839 3148
rect 10781 3139 10839 3145
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 11517 3179 11575 3185
rect 11517 3145 11529 3179
rect 11563 3176 11575 3179
rect 11698 3176 11704 3188
rect 11563 3148 11704 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 13814 3176 13820 3188
rect 13775 3148 13820 3176
rect 13814 3136 13820 3148
rect 13872 3136 13878 3188
rect 17126 3176 17132 3188
rect 14016 3148 17132 3176
rect 5534 3108 5540 3120
rect 3988 3080 5540 3108
rect 3988 3049 4016 3080
rect 5534 3068 5540 3080
rect 5592 3068 5598 3120
rect 8294 3068 8300 3120
rect 8352 3108 8358 3120
rect 8352 3080 10456 3108
rect 8352 3068 8358 3080
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4240 3043 4298 3049
rect 4240 3009 4252 3043
rect 4286 3040 4298 3043
rect 4982 3040 4988 3052
rect 4286 3012 4988 3040
rect 4286 3009 4298 3012
rect 4240 3003 4298 3009
rect 4982 3000 4988 3012
rect 5040 3000 5046 3052
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 6512 3012 6561 3040
rect 6512 3000 6518 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 7248 3012 7297 3040
rect 7248 3000 7254 3012
rect 7285 3009 7297 3012
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7466 3000 7472 3052
rect 7524 3040 7530 3052
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 7524 3012 8401 3040
rect 7524 3000 7530 3012
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 8754 3040 8760 3052
rect 8619 3012 8760 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3040 8999 3043
rect 9122 3040 9128 3052
rect 8987 3012 9128 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 9398 3040 9404 3052
rect 9359 3012 9404 3040
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 9674 3049 9680 3052
rect 9668 3040 9680 3049
rect 9635 3012 9680 3040
rect 9668 3003 9680 3012
rect 9674 3000 9680 3003
rect 9732 3000 9738 3052
rect 2179 2876 3924 2904
rect 2179 2873 2191 2876
rect 2133 2867 2191 2873
rect 4982 2864 4988 2916
rect 5040 2904 5046 2916
rect 7374 2904 7380 2916
rect 5040 2876 7380 2904
rect 5040 2864 5046 2876
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 10428 2904 10456 3080
rect 11882 3068 11888 3120
rect 11940 3108 11946 3120
rect 12713 3111 12771 3117
rect 12713 3108 12725 3111
rect 11940 3080 12725 3108
rect 11940 3068 11946 3080
rect 12713 3077 12725 3080
rect 12759 3077 12771 3111
rect 12713 3071 12771 3077
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3040 11759 3043
rect 11790 3040 11796 3052
rect 11747 3012 11796 3040
rect 11747 3009 11759 3012
rect 11701 3003 11759 3009
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 12986 3040 12992 3052
rect 12023 3012 12992 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 13170 3040 13176 3052
rect 13131 3012 13176 3040
rect 13170 3000 13176 3012
rect 13228 3000 13234 3052
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3040 13323 3043
rect 13354 3040 13360 3052
rect 13311 3012 13360 3040
rect 13311 3009 13323 3012
rect 13265 3003 13323 3009
rect 13354 3000 13360 3012
rect 13412 3040 13418 3052
rect 14016 3040 14044 3148
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 17589 3179 17647 3185
rect 17589 3145 17601 3179
rect 17635 3176 17647 3179
rect 17678 3176 17684 3188
rect 17635 3148 17684 3176
rect 17635 3145 17647 3148
rect 17589 3139 17647 3145
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 17954 3136 17960 3188
rect 18012 3136 18018 3188
rect 18506 3136 18512 3188
rect 18564 3176 18570 3188
rect 19153 3179 19211 3185
rect 19153 3176 19165 3179
rect 18564 3148 19165 3176
rect 18564 3136 18570 3148
rect 19153 3145 19165 3148
rect 19199 3145 19211 3179
rect 19153 3139 19211 3145
rect 19242 3136 19248 3188
rect 19300 3176 19306 3188
rect 19300 3148 19345 3176
rect 19444 3148 20760 3176
rect 19300 3136 19306 3148
rect 14277 3111 14335 3117
rect 14277 3077 14289 3111
rect 14323 3108 14335 3111
rect 15102 3108 15108 3120
rect 14323 3080 15108 3108
rect 14323 3077 14335 3080
rect 14277 3071 14335 3077
rect 15102 3068 15108 3080
rect 15160 3068 15166 3120
rect 15473 3111 15531 3117
rect 15473 3077 15485 3111
rect 15519 3108 15531 3111
rect 15562 3108 15568 3120
rect 15519 3080 15568 3108
rect 15519 3077 15531 3080
rect 15473 3071 15531 3077
rect 15562 3068 15568 3080
rect 15620 3068 15626 3120
rect 16482 3108 16488 3120
rect 15948 3080 16488 3108
rect 14182 3040 14188 3052
rect 13412 3012 14044 3040
rect 14143 3012 14188 3040
rect 13412 3000 13418 3012
rect 14182 3000 14188 3012
rect 14240 3000 14246 3052
rect 15194 3040 15200 3052
rect 15155 3012 15200 3040
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 15746 3040 15752 3052
rect 15304 3012 15752 3040
rect 11885 2975 11943 2981
rect 11885 2941 11897 2975
rect 11931 2972 11943 2975
rect 11931 2944 12434 2972
rect 11931 2941 11943 2944
rect 11885 2935 11943 2941
rect 12406 2904 12434 2944
rect 13078 2932 13084 2984
rect 13136 2972 13142 2984
rect 14369 2975 14427 2981
rect 14369 2972 14381 2975
rect 13136 2944 14381 2972
rect 13136 2932 13142 2944
rect 14369 2941 14381 2944
rect 14415 2972 14427 2975
rect 15304 2972 15332 3012
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 15948 3049 15976 3080
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 16669 3111 16727 3117
rect 16669 3108 16681 3111
rect 16632 3080 16681 3108
rect 16632 3068 16638 3080
rect 16669 3077 16681 3080
rect 16715 3077 16727 3111
rect 17972 3108 18000 3136
rect 17972 3080 18184 3108
rect 16669 3071 16727 3077
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3009 15991 3043
rect 16883 3043 16941 3049
rect 16883 3040 16895 3043
rect 15933 3003 15991 3009
rect 16868 3009 16895 3040
rect 16929 3009 16941 3043
rect 16868 3003 16941 3009
rect 14415 2944 15332 2972
rect 15381 2975 15439 2981
rect 14415 2941 14427 2944
rect 14369 2935 14427 2941
rect 15381 2941 15393 2975
rect 15427 2972 15439 2975
rect 15427 2944 15516 2972
rect 15427 2941 15439 2944
rect 15381 2935 15439 2941
rect 15013 2907 15071 2913
rect 15013 2904 15025 2907
rect 10428 2876 11928 2904
rect 12406 2876 15025 2904
rect 3053 2839 3111 2845
rect 3053 2805 3065 2839
rect 3099 2836 3111 2839
rect 6362 2836 6368 2848
rect 3099 2808 6368 2836
rect 3099 2805 3111 2808
rect 3053 2799 3111 2805
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 6733 2839 6791 2845
rect 6733 2805 6745 2839
rect 6779 2836 6791 2839
rect 8662 2836 8668 2848
rect 6779 2808 8668 2836
rect 6779 2805 6791 2808
rect 6733 2799 6791 2805
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 9306 2796 9312 2848
rect 9364 2836 9370 2848
rect 11790 2836 11796 2848
rect 9364 2808 11796 2836
rect 9364 2796 9370 2808
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 11900 2845 11928 2876
rect 15013 2873 15025 2876
rect 15059 2873 15071 2907
rect 15013 2867 15071 2873
rect 15102 2864 15108 2916
rect 15160 2904 15166 2916
rect 15160 2876 15240 2904
rect 15160 2864 15166 2876
rect 11885 2839 11943 2845
rect 11885 2805 11897 2839
rect 11931 2805 11943 2839
rect 11885 2799 11943 2805
rect 14918 2796 14924 2848
rect 14976 2836 14982 2848
rect 15212 2845 15240 2876
rect 15197 2839 15255 2845
rect 15197 2836 15209 2839
rect 14976 2808 15209 2836
rect 14976 2796 14982 2808
rect 15197 2805 15209 2808
rect 15243 2805 15255 2839
rect 15488 2836 15516 2944
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 16868 2972 16896 3003
rect 17034 3000 17040 3052
rect 17092 3040 17098 3052
rect 17129 3043 17187 3049
rect 17129 3040 17141 3043
rect 17092 3012 17141 3040
rect 17092 3000 17098 3012
rect 17129 3009 17141 3012
rect 17175 3009 17187 3043
rect 17954 3040 17960 3052
rect 17915 3012 17960 3040
rect 17129 3003 17187 3009
rect 17954 3000 17960 3012
rect 18012 3000 18018 3052
rect 18046 2972 18052 2984
rect 15620 2944 16896 2972
rect 18007 2944 18052 2972
rect 15620 2932 15626 2944
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18156 2981 18184 3080
rect 18141 2975 18199 2981
rect 18141 2941 18153 2975
rect 18187 2972 18199 2975
rect 19337 2975 19395 2981
rect 19337 2972 19349 2975
rect 18187 2944 19349 2972
rect 18187 2941 18199 2944
rect 18141 2935 18199 2941
rect 19337 2941 19349 2944
rect 19383 2941 19395 2975
rect 19337 2935 19395 2941
rect 16117 2907 16175 2913
rect 16117 2873 16129 2907
rect 16163 2904 16175 2907
rect 16758 2904 16764 2916
rect 16163 2876 16764 2904
rect 16163 2873 16175 2876
rect 16117 2867 16175 2873
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 16942 2864 16948 2916
rect 17000 2904 17006 2916
rect 17037 2907 17095 2913
rect 17037 2904 17049 2907
rect 17000 2876 17049 2904
rect 17000 2864 17006 2876
rect 17037 2873 17049 2876
rect 17083 2873 17095 2907
rect 17037 2867 17095 2873
rect 17218 2864 17224 2916
rect 17276 2904 17282 2916
rect 19444 2904 19472 3148
rect 20530 3068 20536 3120
rect 20588 3108 20594 3120
rect 20732 3108 20760 3148
rect 21358 3136 21364 3188
rect 21416 3176 21422 3188
rect 21818 3176 21824 3188
rect 21416 3148 21824 3176
rect 21416 3136 21422 3148
rect 21818 3136 21824 3148
rect 21876 3136 21882 3188
rect 22922 3176 22928 3188
rect 22883 3148 22928 3176
rect 22922 3136 22928 3148
rect 22980 3136 22986 3188
rect 23566 3176 23572 3188
rect 23527 3148 23572 3176
rect 23566 3136 23572 3148
rect 23624 3136 23630 3188
rect 27249 3179 27307 3185
rect 27249 3145 27261 3179
rect 27295 3176 27307 3179
rect 29365 3179 29423 3185
rect 27295 3148 28212 3176
rect 27295 3145 27307 3148
rect 27249 3139 27307 3145
rect 21634 3108 21640 3120
rect 20588 3080 20668 3108
rect 20732 3080 21640 3108
rect 20588 3068 20594 3080
rect 20162 3040 20168 3052
rect 20123 3012 20168 3040
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 20438 3000 20444 3052
rect 20496 3040 20502 3052
rect 20640 3049 20668 3080
rect 21634 3068 21640 3080
rect 21692 3068 21698 3120
rect 21726 3068 21732 3120
rect 21784 3108 21790 3120
rect 27709 3111 27767 3117
rect 21784 3080 23796 3108
rect 21784 3068 21790 3080
rect 20625 3043 20683 3049
rect 20496 3012 20541 3040
rect 20496 3000 20502 3012
rect 20625 3009 20637 3043
rect 20671 3009 20683 3043
rect 22002 3040 22008 3052
rect 21963 3012 22008 3040
rect 20625 3003 20683 3009
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 22094 3000 22100 3052
rect 22152 3040 22158 3052
rect 22462 3040 22468 3052
rect 22152 3012 22197 3040
rect 22423 3012 22468 3040
rect 22152 3000 22158 3012
rect 22462 3000 22468 3012
rect 22520 3000 22526 3052
rect 23768 3049 23796 3080
rect 27709 3077 27721 3111
rect 27755 3108 27767 3111
rect 27982 3108 27988 3120
rect 27755 3080 27988 3108
rect 27755 3077 27767 3080
rect 27709 3071 27767 3077
rect 27982 3068 27988 3080
rect 28040 3068 28046 3120
rect 28184 3117 28212 3148
rect 29365 3145 29377 3179
rect 29411 3145 29423 3179
rect 29365 3139 29423 3145
rect 28169 3111 28227 3117
rect 28169 3077 28181 3111
rect 28215 3077 28227 3111
rect 28169 3071 28227 3077
rect 28353 3111 28411 3117
rect 28353 3077 28365 3111
rect 28399 3108 28411 3111
rect 29380 3108 29408 3139
rect 28399 3080 29408 3108
rect 28399 3077 28411 3080
rect 28353 3071 28411 3077
rect 23109 3043 23167 3049
rect 23109 3009 23121 3043
rect 23155 3009 23167 3043
rect 23109 3003 23167 3009
rect 23753 3043 23811 3049
rect 23753 3009 23765 3043
rect 23799 3009 23811 3043
rect 23753 3003 23811 3009
rect 23124 2972 23152 3003
rect 23934 3000 23940 3052
rect 23992 3040 23998 3052
rect 24397 3043 24455 3049
rect 24397 3040 24409 3043
rect 23992 3012 24409 3040
rect 23992 3000 23998 3012
rect 24397 3009 24409 3012
rect 24443 3009 24455 3043
rect 27430 3040 27436 3052
rect 27391 3012 27436 3040
rect 24397 3003 24455 3009
rect 27430 3000 27436 3012
rect 27488 3000 27494 3052
rect 28718 3000 28724 3052
rect 28776 3040 28782 3052
rect 29549 3043 29607 3049
rect 29549 3040 29561 3043
rect 28776 3012 29561 3040
rect 28776 3000 28782 3012
rect 29549 3009 29561 3012
rect 29595 3009 29607 3043
rect 29914 3040 29920 3052
rect 29875 3012 29920 3040
rect 29549 3003 29607 3009
rect 29914 3000 29920 3012
rect 29972 3000 29978 3052
rect 30006 3000 30012 3052
rect 30064 3040 30070 3052
rect 30064 3012 30109 3040
rect 30064 3000 30070 3012
rect 27614 2972 27620 2984
rect 20548 2944 23152 2972
rect 27575 2944 27620 2972
rect 17276 2876 19472 2904
rect 17276 2864 17282 2876
rect 20162 2864 20168 2916
rect 20220 2904 20226 2916
rect 20548 2904 20576 2944
rect 27614 2932 27620 2944
rect 27672 2932 27678 2984
rect 20220 2876 20576 2904
rect 20809 2907 20867 2913
rect 20220 2864 20226 2876
rect 20809 2873 20821 2907
rect 20855 2904 20867 2907
rect 22094 2904 22100 2916
rect 20855 2876 22100 2904
rect 20855 2873 20867 2876
rect 20809 2867 20867 2873
rect 22094 2864 22100 2876
rect 22152 2864 22158 2916
rect 22738 2864 22744 2916
rect 22796 2904 22802 2916
rect 28537 2907 28595 2913
rect 28537 2904 28549 2907
rect 22796 2876 28549 2904
rect 22796 2864 22802 2876
rect 28537 2873 28549 2876
rect 28583 2873 28595 2907
rect 28537 2867 28595 2873
rect 16666 2836 16672 2848
rect 15488 2808 16672 2836
rect 15197 2799 15255 2805
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 18138 2796 18144 2848
rect 18196 2836 18202 2848
rect 18785 2839 18843 2845
rect 18785 2836 18797 2839
rect 18196 2808 18797 2836
rect 18196 2796 18202 2808
rect 18785 2805 18797 2808
rect 18831 2805 18843 2839
rect 18785 2799 18843 2805
rect 19518 2796 19524 2848
rect 19576 2836 19582 2848
rect 20254 2836 20260 2848
rect 19576 2808 20260 2836
rect 19576 2796 19582 2808
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 22370 2836 22376 2848
rect 22331 2808 22376 2836
rect 22370 2796 22376 2808
rect 22428 2836 22434 2848
rect 24213 2839 24271 2845
rect 24213 2836 24225 2839
rect 22428 2808 24225 2836
rect 22428 2796 22434 2808
rect 24213 2805 24225 2808
rect 24259 2805 24271 2839
rect 27706 2836 27712 2848
rect 27667 2808 27712 2836
rect 24213 2799 24271 2805
rect 27706 2796 27712 2808
rect 27764 2796 27770 2848
rect 29546 2836 29552 2848
rect 29507 2808 29552 2836
rect 29546 2796 29552 2808
rect 29604 2796 29610 2848
rect 1104 2746 30820 2768
rect 1104 2694 5915 2746
rect 5967 2694 5979 2746
rect 6031 2694 6043 2746
rect 6095 2694 6107 2746
rect 6159 2694 6171 2746
rect 6223 2694 15846 2746
rect 15898 2694 15910 2746
rect 15962 2694 15974 2746
rect 16026 2694 16038 2746
rect 16090 2694 16102 2746
rect 16154 2694 25776 2746
rect 25828 2694 25840 2746
rect 25892 2694 25904 2746
rect 25956 2694 25968 2746
rect 26020 2694 26032 2746
rect 26084 2694 30820 2746
rect 1104 2672 30820 2694
rect 4430 2632 4436 2644
rect 4391 2604 4436 2632
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 7834 2632 7840 2644
rect 6595 2604 7840 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8205 2635 8263 2641
rect 8205 2601 8217 2635
rect 8251 2632 8263 2635
rect 8294 2632 8300 2644
rect 8251 2604 8300 2632
rect 8251 2601 8263 2604
rect 8205 2595 8263 2601
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 11698 2632 11704 2644
rect 9171 2604 11704 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 14093 2635 14151 2641
rect 14093 2601 14105 2635
rect 14139 2632 14151 2635
rect 14182 2632 14188 2644
rect 14139 2604 14188 2632
rect 14139 2601 14151 2604
rect 14093 2595 14151 2601
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 14458 2632 14464 2644
rect 14419 2604 14464 2632
rect 14458 2592 14464 2604
rect 14516 2632 14522 2644
rect 15105 2635 15163 2641
rect 15105 2632 15117 2635
rect 14516 2604 15117 2632
rect 14516 2592 14522 2604
rect 15105 2601 15117 2604
rect 15151 2601 15163 2635
rect 15105 2595 15163 2601
rect 15378 2592 15384 2644
rect 15436 2632 15442 2644
rect 15473 2635 15531 2641
rect 15473 2632 15485 2635
rect 15436 2604 15485 2632
rect 15436 2592 15442 2604
rect 15473 2601 15485 2604
rect 15519 2601 15531 2635
rect 15473 2595 15531 2601
rect 15562 2592 15568 2644
rect 15620 2632 15626 2644
rect 16117 2635 16175 2641
rect 16117 2632 16129 2635
rect 15620 2604 16129 2632
rect 15620 2592 15626 2604
rect 16117 2601 16129 2604
rect 16163 2601 16175 2635
rect 16666 2632 16672 2644
rect 16627 2604 16672 2632
rect 16117 2595 16175 2601
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 17773 2635 17831 2641
rect 17773 2601 17785 2635
rect 17819 2601 17831 2635
rect 17773 2595 17831 2601
rect 3053 2567 3111 2573
rect 3053 2533 3065 2567
rect 3099 2564 3111 2567
rect 7466 2564 7472 2576
rect 3099 2536 7472 2564
rect 3099 2533 3111 2536
rect 3053 2527 3111 2533
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 7561 2567 7619 2573
rect 7561 2533 7573 2567
rect 7607 2564 7619 2567
rect 12894 2564 12900 2576
rect 7607 2536 12900 2564
rect 7607 2533 7619 2536
rect 7561 2527 7619 2533
rect 12894 2524 12900 2536
rect 12952 2524 12958 2576
rect 12986 2524 12992 2576
rect 13044 2564 13050 2576
rect 17313 2567 17371 2573
rect 17313 2564 17325 2567
rect 13044 2536 17325 2564
rect 13044 2524 13050 2536
rect 17313 2533 17325 2536
rect 17359 2533 17371 2567
rect 17788 2564 17816 2595
rect 17954 2592 17960 2644
rect 18012 2632 18018 2644
rect 18233 2635 18291 2641
rect 18233 2632 18245 2635
rect 18012 2604 18245 2632
rect 18012 2592 18018 2604
rect 18233 2601 18245 2604
rect 18279 2601 18291 2635
rect 19245 2635 19303 2641
rect 19245 2632 19257 2635
rect 18233 2595 18291 2601
rect 18340 2604 19257 2632
rect 18340 2576 18368 2604
rect 19245 2601 19257 2604
rect 19291 2601 19303 2635
rect 20254 2632 20260 2644
rect 20215 2604 20260 2632
rect 19245 2595 19303 2601
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 20714 2632 20720 2644
rect 20675 2604 20720 2632
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 21634 2592 21640 2644
rect 21692 2632 21698 2644
rect 21821 2635 21879 2641
rect 21821 2632 21833 2635
rect 21692 2604 21833 2632
rect 21692 2592 21698 2604
rect 21821 2601 21833 2604
rect 21867 2601 21879 2635
rect 21821 2595 21879 2601
rect 22094 2592 22100 2644
rect 22152 2632 22158 2644
rect 22152 2604 22197 2632
rect 22152 2592 22158 2604
rect 22278 2592 22284 2644
rect 22336 2632 22342 2644
rect 24397 2635 24455 2641
rect 24397 2632 24409 2635
rect 22336 2604 24409 2632
rect 22336 2592 22342 2604
rect 24397 2601 24409 2604
rect 24443 2601 24455 2635
rect 25682 2632 25688 2644
rect 25643 2604 25688 2632
rect 24397 2595 24455 2601
rect 25682 2592 25688 2604
rect 25740 2592 25746 2644
rect 27157 2635 27215 2641
rect 27157 2601 27169 2635
rect 27203 2632 27215 2635
rect 27430 2632 27436 2644
rect 27203 2604 27436 2632
rect 27203 2601 27215 2604
rect 27157 2595 27215 2601
rect 27430 2592 27436 2604
rect 27488 2592 27494 2644
rect 27614 2632 27620 2644
rect 27575 2604 27620 2632
rect 27614 2592 27620 2604
rect 27672 2592 27678 2644
rect 18322 2564 18328 2576
rect 17788 2536 18328 2564
rect 17313 2527 17371 2533
rect 18322 2524 18328 2536
rect 18380 2524 18386 2576
rect 18598 2524 18604 2576
rect 18656 2564 18662 2576
rect 18656 2536 22876 2564
rect 18656 2524 18662 2536
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2496 2283 2499
rect 9306 2496 9312 2508
rect 2271 2468 4568 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 1854 2388 1860 2440
rect 1912 2428 1918 2440
rect 1949 2431 2007 2437
rect 1949 2428 1961 2431
rect 1912 2400 1961 2428
rect 1912 2388 1918 2400
rect 1949 2397 1961 2400
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 382 2320 388 2372
rect 440 2360 446 2372
rect 2884 2360 2912 2391
rect 4154 2360 4160 2372
rect 440 2332 2912 2360
rect 4115 2332 4160 2360
rect 440 2320 446 2332
rect 4154 2320 4160 2332
rect 4212 2320 4218 2372
rect 4540 2292 4568 2468
rect 7392 2468 9312 2496
rect 4890 2388 4896 2440
rect 4948 2428 4954 2440
rect 4985 2431 5043 2437
rect 4985 2428 4997 2431
rect 4948 2400 4997 2428
rect 4948 2388 4954 2400
rect 4985 2397 4997 2400
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 5276 2360 5304 2391
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 7392 2437 7420 2468
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 10318 2496 10324 2508
rect 9907 2468 10324 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 10502 2456 10508 2508
rect 10560 2496 10566 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 10560 2468 11805 2496
rect 10560 2456 10566 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 14553 2499 14611 2505
rect 14553 2465 14565 2499
rect 14599 2496 14611 2499
rect 15010 2496 15016 2508
rect 14599 2468 15016 2496
rect 14599 2465 14611 2468
rect 14553 2459 14611 2465
rect 15010 2456 15016 2468
rect 15068 2456 15074 2508
rect 16758 2456 16764 2508
rect 16816 2496 16822 2508
rect 16816 2468 16988 2496
rect 16816 2456 16822 2468
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5776 2400 6377 2428
rect 5776 2388 5782 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7984 2400 8033 2428
rect 7984 2388 7990 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8812 2400 8953 2428
rect 8812 2388 8818 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9490 2388 9496 2440
rect 9548 2428 9554 2440
rect 9585 2431 9643 2437
rect 9585 2428 9597 2431
rect 9548 2400 9597 2428
rect 9548 2388 9554 2400
rect 9585 2397 9597 2400
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 10284 2400 11529 2428
rect 10284 2388 10290 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 12805 2431 12863 2437
rect 12805 2397 12817 2431
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2428 14335 2431
rect 14918 2428 14924 2440
rect 14323 2400 14924 2428
rect 14323 2397 14335 2400
rect 14277 2391 14335 2397
rect 8386 2360 8392 2372
rect 5276 2332 8392 2360
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 11330 2320 11336 2372
rect 11388 2360 11394 2372
rect 12820 2360 12848 2391
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 15286 2428 15292 2440
rect 15247 2400 15292 2428
rect 15286 2388 15292 2400
rect 15344 2388 15350 2440
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 15933 2431 15991 2437
rect 15933 2428 15945 2431
rect 15620 2400 15945 2428
rect 15620 2388 15626 2400
rect 15933 2397 15945 2400
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 16390 2388 16396 2440
rect 16448 2428 16454 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16448 2400 16865 2428
rect 16448 2388 16454 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16960 2428 16988 2468
rect 17126 2456 17132 2508
rect 17184 2496 17190 2508
rect 20438 2496 20444 2508
rect 17184 2468 19472 2496
rect 20399 2468 20444 2496
rect 17184 2456 17190 2468
rect 17402 2428 17408 2440
rect 16960 2400 17408 2428
rect 16853 2391 16911 2397
rect 17402 2388 17408 2400
rect 17460 2428 17466 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17460 2400 17509 2428
rect 17460 2388 17466 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 17589 2431 17647 2437
rect 17589 2397 17601 2431
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2428 17831 2431
rect 18046 2428 18052 2440
rect 17819 2400 18052 2428
rect 17819 2397 17831 2400
rect 17773 2391 17831 2397
rect 11388 2332 12848 2360
rect 11388 2320 11394 2332
rect 8938 2292 8944 2304
rect 4540 2264 8944 2292
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 12618 2252 12624 2304
rect 12676 2292 12682 2304
rect 12989 2295 13047 2301
rect 12989 2292 13001 2295
rect 12676 2264 13001 2292
rect 12676 2252 12682 2264
rect 12989 2261 13001 2264
rect 13035 2261 13047 2295
rect 17604 2292 17632 2391
rect 18046 2388 18052 2400
rect 18104 2428 18110 2440
rect 18417 2431 18475 2437
rect 18417 2428 18429 2431
rect 18104 2400 18429 2428
rect 18104 2388 18110 2400
rect 18417 2397 18429 2400
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 18432 2360 18460 2391
rect 18506 2388 18512 2440
rect 18564 2428 18570 2440
rect 18601 2431 18659 2437
rect 18601 2428 18613 2431
rect 18564 2400 18613 2428
rect 18564 2388 18570 2400
rect 18601 2397 18613 2400
rect 18647 2397 18659 2431
rect 18601 2391 18659 2397
rect 18693 2431 18751 2437
rect 18693 2397 18705 2431
rect 18739 2428 18751 2431
rect 18782 2428 18788 2440
rect 18739 2400 18788 2428
rect 18739 2397 18751 2400
rect 18693 2391 18751 2397
rect 18782 2388 18788 2400
rect 18840 2388 18846 2440
rect 19444 2437 19472 2468
rect 20438 2456 20444 2468
rect 20496 2456 20502 2508
rect 22646 2496 22652 2508
rect 20640 2468 22652 2496
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2397 19487 2431
rect 20530 2428 20536 2440
rect 19429 2391 19487 2397
rect 19536 2400 20392 2428
rect 20491 2400 20536 2428
rect 19536 2360 19564 2400
rect 18432 2332 19564 2360
rect 20070 2320 20076 2372
rect 20128 2360 20134 2372
rect 20257 2363 20315 2369
rect 20257 2360 20269 2363
rect 20128 2332 20269 2360
rect 20128 2320 20134 2332
rect 20257 2329 20269 2332
rect 20303 2329 20315 2363
rect 20364 2360 20392 2400
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 20640 2360 20668 2468
rect 22646 2456 22652 2468
rect 22704 2456 22710 2508
rect 21818 2388 21824 2440
rect 21876 2428 21882 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21876 2400 22017 2428
rect 21876 2388 21882 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2428 22247 2431
rect 22738 2428 22744 2440
rect 22235 2400 22744 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 22738 2388 22744 2400
rect 22796 2388 22802 2440
rect 22848 2437 22876 2536
rect 23198 2456 23204 2508
rect 23256 2496 23262 2508
rect 23256 2468 24624 2496
rect 23256 2456 23262 2468
rect 24596 2437 24624 2468
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 24581 2431 24639 2437
rect 24581 2397 24593 2431
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 23492 2360 23520 2391
rect 24762 2388 24768 2440
rect 24820 2428 24826 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 24820 2400 25237 2428
rect 24820 2388 24826 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 25498 2388 25504 2440
rect 25556 2428 25562 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 25556 2400 25881 2428
rect 25556 2388 25562 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 26234 2388 26240 2440
rect 26292 2428 26298 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26292 2400 26985 2428
rect 26292 2388 26298 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27120 2400 27813 2428
rect 27120 2388 27126 2400
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 28718 2428 28724 2440
rect 28679 2400 28724 2428
rect 27801 2391 27859 2397
rect 28718 2388 28724 2400
rect 28776 2388 28782 2440
rect 29454 2388 29460 2440
rect 29512 2428 29518 2440
rect 29825 2431 29883 2437
rect 29825 2428 29837 2431
rect 29512 2400 29837 2428
rect 29512 2388 29518 2400
rect 29825 2397 29837 2400
rect 29871 2397 29883 2431
rect 29825 2391 29883 2397
rect 20364 2332 20668 2360
rect 20732 2332 23520 2360
rect 20257 2323 20315 2329
rect 19242 2292 19248 2304
rect 17604 2264 19248 2292
rect 12989 2255 13047 2261
rect 19242 2252 19248 2264
rect 19300 2252 19306 2304
rect 19426 2252 19432 2304
rect 19484 2292 19490 2304
rect 20732 2292 20760 2332
rect 22646 2292 22652 2304
rect 19484 2264 20760 2292
rect 22607 2264 22652 2292
rect 19484 2252 19490 2264
rect 22646 2252 22652 2264
rect 22704 2252 22710 2304
rect 23290 2292 23296 2304
rect 23251 2264 23296 2292
rect 23290 2252 23296 2264
rect 23348 2252 23354 2304
rect 25038 2292 25044 2304
rect 24999 2264 25044 2292
rect 25038 2252 25044 2264
rect 25096 2252 25102 2304
rect 28902 2292 28908 2304
rect 28863 2264 28908 2292
rect 28902 2252 28908 2264
rect 28960 2252 28966 2304
rect 30006 2292 30012 2304
rect 29967 2264 30012 2292
rect 30006 2252 30012 2264
rect 30064 2252 30070 2304
rect 1104 2202 30820 2224
rect 1104 2150 10880 2202
rect 10932 2150 10944 2202
rect 10996 2150 11008 2202
rect 11060 2150 11072 2202
rect 11124 2150 11136 2202
rect 11188 2150 20811 2202
rect 20863 2150 20875 2202
rect 20927 2150 20939 2202
rect 20991 2150 21003 2202
rect 21055 2150 21067 2202
rect 21119 2150 30820 2202
rect 1104 2128 30820 2150
rect 22002 2048 22008 2100
rect 22060 2088 22066 2100
rect 25038 2088 25044 2100
rect 22060 2060 25044 2088
rect 22060 2048 22066 2060
rect 25038 2048 25044 2060
rect 25096 2048 25102 2100
rect 19242 1980 19248 2032
rect 19300 2020 19306 2032
rect 23290 2020 23296 2032
rect 19300 1992 23296 2020
rect 19300 1980 19306 1992
rect 23290 1980 23296 1992
rect 23348 1980 23354 2032
<< via1 >>
rect 10880 45670 10932 45722
rect 10944 45670 10996 45722
rect 11008 45670 11060 45722
rect 11072 45670 11124 45722
rect 11136 45670 11188 45722
rect 20811 45670 20863 45722
rect 20875 45670 20927 45722
rect 20939 45670 20991 45722
rect 21003 45670 21055 45722
rect 21067 45670 21119 45722
rect 1400 45432 1452 45484
rect 2872 45432 2924 45484
rect 3056 45432 3108 45484
rect 3148 45475 3200 45484
rect 3148 45441 3157 45475
rect 3157 45441 3191 45475
rect 3191 45441 3200 45475
rect 3148 45432 3200 45441
rect 4804 45432 4856 45484
rect 30104 45475 30156 45484
rect 30104 45441 30113 45475
rect 30113 45441 30147 45475
rect 30147 45441 30156 45475
rect 30104 45432 30156 45441
rect 2228 45339 2280 45348
rect 2228 45305 2237 45339
rect 2237 45305 2271 45339
rect 2271 45305 2280 45339
rect 2228 45296 2280 45305
rect 2964 45339 3016 45348
rect 2964 45305 2973 45339
rect 2973 45305 3007 45339
rect 3007 45305 3016 45339
rect 2964 45296 3016 45305
rect 5264 45364 5316 45416
rect 2780 45228 2832 45280
rect 2872 45228 2924 45280
rect 29920 45271 29972 45280
rect 29920 45237 29929 45271
rect 29929 45237 29963 45271
rect 29963 45237 29972 45271
rect 29920 45228 29972 45237
rect 5915 45126 5967 45178
rect 5979 45126 6031 45178
rect 6043 45126 6095 45178
rect 6107 45126 6159 45178
rect 6171 45126 6223 45178
rect 15846 45126 15898 45178
rect 15910 45126 15962 45178
rect 15974 45126 16026 45178
rect 16038 45126 16090 45178
rect 16102 45126 16154 45178
rect 25776 45126 25828 45178
rect 25840 45126 25892 45178
rect 25904 45126 25956 45178
rect 25968 45126 26020 45178
rect 26032 45126 26084 45178
rect 3056 45024 3108 45076
rect 3148 45024 3200 45076
rect 5172 45024 5224 45076
rect 2872 44820 2924 44872
rect 5724 44888 5776 44940
rect 4528 44820 4580 44872
rect 1492 44727 1544 44736
rect 1492 44693 1501 44727
rect 1501 44693 1535 44727
rect 1535 44693 1544 44727
rect 1492 44684 1544 44693
rect 2872 44727 2924 44736
rect 2872 44693 2881 44727
rect 2881 44693 2915 44727
rect 2915 44693 2924 44727
rect 2872 44684 2924 44693
rect 5540 44820 5592 44872
rect 6552 44820 6604 44872
rect 8392 44820 8444 44872
rect 30196 44820 30248 44872
rect 7012 44752 7064 44804
rect 6276 44684 6328 44736
rect 7196 44684 7248 44736
rect 8944 44727 8996 44736
rect 8944 44693 8953 44727
rect 8953 44693 8987 44727
rect 8987 44693 8996 44727
rect 8944 44684 8996 44693
rect 29000 44684 29052 44736
rect 10880 44582 10932 44634
rect 10944 44582 10996 44634
rect 11008 44582 11060 44634
rect 11072 44582 11124 44634
rect 11136 44582 11188 44634
rect 20811 44582 20863 44634
rect 20875 44582 20927 44634
rect 20939 44582 20991 44634
rect 21003 44582 21055 44634
rect 21067 44582 21119 44634
rect 4804 44523 4856 44532
rect 4804 44489 4813 44523
rect 4813 44489 4847 44523
rect 4847 44489 4856 44523
rect 4804 44480 4856 44489
rect 5264 44523 5316 44532
rect 5264 44489 5273 44523
rect 5273 44489 5307 44523
rect 5307 44489 5316 44523
rect 5264 44480 5316 44489
rect 6552 44523 6604 44532
rect 6552 44489 6561 44523
rect 6561 44489 6595 44523
rect 6595 44489 6604 44523
rect 6552 44480 6604 44489
rect 7012 44523 7064 44532
rect 7012 44489 7021 44523
rect 7021 44489 7055 44523
rect 7055 44489 7064 44523
rect 7012 44480 7064 44489
rect 7564 44480 7616 44532
rect 2872 44412 2924 44464
rect 8760 44480 8812 44532
rect 10508 44480 10560 44532
rect 18144 44480 18196 44532
rect 2320 44387 2372 44396
rect 2320 44353 2329 44387
rect 2329 44353 2363 44387
rect 2363 44353 2372 44387
rect 2320 44344 2372 44353
rect 4252 44344 4304 44396
rect 3976 44276 4028 44328
rect 6368 44387 6420 44396
rect 6368 44353 6377 44387
rect 6377 44353 6411 44387
rect 6411 44353 6420 44387
rect 6368 44344 6420 44353
rect 7196 44387 7248 44396
rect 7196 44353 7205 44387
rect 7205 44353 7239 44387
rect 7239 44353 7248 44387
rect 7196 44344 7248 44353
rect 7564 44387 7616 44396
rect 7564 44353 7573 44387
rect 7573 44353 7607 44387
rect 7607 44353 7616 44387
rect 7564 44344 7616 44353
rect 7748 44387 7800 44396
rect 7748 44353 7757 44387
rect 7757 44353 7791 44387
rect 7791 44353 7800 44387
rect 7748 44344 7800 44353
rect 8300 44344 8352 44396
rect 7380 44319 7432 44328
rect 5540 44208 5592 44260
rect 7380 44285 7389 44319
rect 7389 44285 7423 44319
rect 7423 44285 7432 44319
rect 7380 44276 7432 44285
rect 7840 44276 7892 44328
rect 9128 44344 9180 44396
rect 8852 44208 8904 44260
rect 9956 44208 10008 44260
rect 18328 44387 18380 44396
rect 18328 44353 18337 44387
rect 18337 44353 18371 44387
rect 18371 44353 18380 44387
rect 18328 44344 18380 44353
rect 30104 44387 30156 44396
rect 30104 44353 30113 44387
rect 30113 44353 30147 44387
rect 30147 44353 30156 44387
rect 30104 44344 30156 44353
rect 29920 44276 29972 44328
rect 18052 44208 18104 44260
rect 1492 44183 1544 44192
rect 1492 44149 1501 44183
rect 1501 44149 1535 44183
rect 1535 44149 1544 44183
rect 1492 44140 1544 44149
rect 1952 44140 2004 44192
rect 2964 44140 3016 44192
rect 3424 44183 3476 44192
rect 3424 44149 3433 44183
rect 3433 44149 3467 44183
rect 3467 44149 3476 44183
rect 3424 44140 3476 44149
rect 5172 44140 5224 44192
rect 8300 44140 8352 44192
rect 8760 44140 8812 44192
rect 10232 44140 10284 44192
rect 17960 44140 18012 44192
rect 29920 44183 29972 44192
rect 29920 44149 29929 44183
rect 29929 44149 29963 44183
rect 29963 44149 29972 44183
rect 29920 44140 29972 44149
rect 5915 44038 5967 44090
rect 5979 44038 6031 44090
rect 6043 44038 6095 44090
rect 6107 44038 6159 44090
rect 6171 44038 6223 44090
rect 15846 44038 15898 44090
rect 15910 44038 15962 44090
rect 15974 44038 16026 44090
rect 16038 44038 16090 44090
rect 16102 44038 16154 44090
rect 25776 44038 25828 44090
rect 25840 44038 25892 44090
rect 25904 44038 25956 44090
rect 25968 44038 26020 44090
rect 26032 44038 26084 44090
rect 4528 43936 4580 43988
rect 3148 43868 3200 43920
rect 5172 43868 5224 43920
rect 6368 43936 6420 43988
rect 7748 43936 7800 43988
rect 18144 43979 18196 43988
rect 18144 43945 18153 43979
rect 18153 43945 18187 43979
rect 18187 43945 18196 43979
rect 18144 43936 18196 43945
rect 6276 43868 6328 43920
rect 7380 43800 7432 43852
rect 1860 43775 1912 43784
rect 1860 43741 1869 43775
rect 1869 43741 1903 43775
rect 1903 43741 1912 43775
rect 1860 43732 1912 43741
rect 2504 43732 2556 43784
rect 5080 43732 5132 43784
rect 5540 43732 5592 43784
rect 5908 43732 5960 43784
rect 6644 43732 6696 43784
rect 5632 43664 5684 43716
rect 7748 43664 7800 43716
rect 1584 43596 1636 43648
rect 3240 43596 3292 43648
rect 5356 43596 5408 43648
rect 7196 43596 7248 43648
rect 7288 43596 7340 43648
rect 7932 43775 7984 43784
rect 7932 43741 7941 43775
rect 7941 43741 7975 43775
rect 7975 43741 7984 43775
rect 8944 43843 8996 43852
rect 8944 43809 8953 43843
rect 8953 43809 8987 43843
rect 8987 43809 8996 43843
rect 8944 43800 8996 43809
rect 7932 43732 7984 43741
rect 18328 43775 18380 43784
rect 18328 43741 18337 43775
rect 18337 43741 18371 43775
rect 18371 43741 18380 43775
rect 18328 43732 18380 43741
rect 29000 43732 29052 43784
rect 10692 43664 10744 43716
rect 17960 43664 18012 43716
rect 10880 43494 10932 43546
rect 10944 43494 10996 43546
rect 11008 43494 11060 43546
rect 11072 43494 11124 43546
rect 11136 43494 11188 43546
rect 20811 43494 20863 43546
rect 20875 43494 20927 43546
rect 20939 43494 20991 43546
rect 21003 43494 21055 43546
rect 21067 43494 21119 43546
rect 7196 43392 7248 43444
rect 8852 43435 8904 43444
rect 8852 43401 8861 43435
rect 8861 43401 8895 43435
rect 8895 43401 8904 43435
rect 8852 43392 8904 43401
rect 18052 43392 18104 43444
rect 3424 43324 3476 43376
rect 9956 43367 10008 43376
rect 9956 43333 9974 43367
rect 9974 43333 10008 43367
rect 9956 43324 10008 43333
rect 2872 43256 2924 43308
rect 3884 43299 3936 43308
rect 3884 43265 3893 43299
rect 3893 43265 3927 43299
rect 3927 43265 3936 43299
rect 3884 43256 3936 43265
rect 4528 43299 4580 43308
rect 4528 43265 4537 43299
rect 4537 43265 4571 43299
rect 4571 43265 4580 43299
rect 4528 43256 4580 43265
rect 5080 43256 5132 43308
rect 5908 43256 5960 43308
rect 7012 43299 7064 43308
rect 7012 43265 7046 43299
rect 7046 43265 7064 43299
rect 10232 43299 10284 43308
rect 7012 43256 7064 43265
rect 10232 43265 10241 43299
rect 10241 43265 10275 43299
rect 10275 43265 10284 43299
rect 10232 43256 10284 43265
rect 18328 43299 18380 43308
rect 18328 43265 18337 43299
rect 18337 43265 18371 43299
rect 18371 43265 18380 43299
rect 18328 43256 18380 43265
rect 19064 43256 19116 43308
rect 6736 43231 6788 43240
rect 6736 43197 6745 43231
rect 6745 43197 6779 43231
rect 6779 43197 6788 43231
rect 6736 43188 6788 43197
rect 29920 43188 29972 43240
rect 1492 43095 1544 43104
rect 1492 43061 1501 43095
rect 1501 43061 1535 43095
rect 1535 43061 1544 43095
rect 1492 43052 1544 43061
rect 2780 43052 2832 43104
rect 3056 43052 3108 43104
rect 4344 43095 4396 43104
rect 4344 43061 4353 43095
rect 4353 43061 4387 43095
rect 4387 43061 4396 43095
rect 4344 43052 4396 43061
rect 5172 43095 5224 43104
rect 5172 43061 5181 43095
rect 5181 43061 5215 43095
rect 5215 43061 5224 43095
rect 5172 43052 5224 43061
rect 6920 43052 6972 43104
rect 5915 42950 5967 43002
rect 5979 42950 6031 43002
rect 6043 42950 6095 43002
rect 6107 42950 6159 43002
rect 6171 42950 6223 43002
rect 15846 42950 15898 43002
rect 15910 42950 15962 43002
rect 15974 42950 16026 43002
rect 16038 42950 16090 43002
rect 16102 42950 16154 43002
rect 25776 42950 25828 43002
rect 25840 42950 25892 43002
rect 25904 42950 25956 43002
rect 25968 42950 26020 43002
rect 26032 42950 26084 43002
rect 5172 42848 5224 42900
rect 7012 42891 7064 42900
rect 7012 42857 7021 42891
rect 7021 42857 7055 42891
rect 7055 42857 7064 42891
rect 7012 42848 7064 42857
rect 2964 42712 3016 42764
rect 2136 42687 2188 42696
rect 2136 42653 2145 42687
rect 2145 42653 2179 42687
rect 2179 42653 2188 42687
rect 2136 42644 2188 42653
rect 3056 42687 3108 42696
rect 3056 42653 3065 42687
rect 3065 42653 3099 42687
rect 3099 42653 3108 42687
rect 3056 42644 3108 42653
rect 1492 42551 1544 42560
rect 1492 42517 1501 42551
rect 1501 42517 1535 42551
rect 1535 42517 1544 42551
rect 1492 42508 1544 42517
rect 2596 42508 2648 42560
rect 5908 42644 5960 42696
rect 7196 42687 7248 42696
rect 7196 42653 7205 42687
rect 7205 42653 7239 42687
rect 7239 42653 7248 42687
rect 7196 42644 7248 42653
rect 7380 42687 7432 42696
rect 7380 42653 7389 42687
rect 7389 42653 7423 42687
rect 7423 42653 7432 42687
rect 7380 42644 7432 42653
rect 7840 42780 7892 42832
rect 7656 42644 7708 42696
rect 7748 42687 7800 42696
rect 7748 42653 7757 42687
rect 7757 42653 7791 42687
rect 7791 42653 7800 42687
rect 7748 42644 7800 42653
rect 8024 42644 8076 42696
rect 30104 42687 30156 42696
rect 30104 42653 30113 42687
rect 30113 42653 30147 42687
rect 30147 42653 30156 42687
rect 30104 42644 30156 42653
rect 4436 42619 4488 42628
rect 4436 42585 4470 42619
rect 4470 42585 4488 42619
rect 4436 42576 4488 42585
rect 5724 42576 5776 42628
rect 5816 42508 5868 42560
rect 10324 42576 10376 42628
rect 7932 42508 7984 42560
rect 8392 42551 8444 42560
rect 8392 42517 8401 42551
rect 8401 42517 8435 42551
rect 8435 42517 8444 42551
rect 8392 42508 8444 42517
rect 9128 42551 9180 42560
rect 9128 42517 9137 42551
rect 9137 42517 9171 42551
rect 9171 42517 9180 42551
rect 9128 42508 9180 42517
rect 29920 42551 29972 42560
rect 29920 42517 29929 42551
rect 29929 42517 29963 42551
rect 29963 42517 29972 42551
rect 29920 42508 29972 42517
rect 10880 42406 10932 42458
rect 10944 42406 10996 42458
rect 11008 42406 11060 42458
rect 11072 42406 11124 42458
rect 11136 42406 11188 42458
rect 20811 42406 20863 42458
rect 20875 42406 20927 42458
rect 20939 42406 20991 42458
rect 21003 42406 21055 42458
rect 21067 42406 21119 42458
rect 4252 42304 4304 42356
rect 6736 42347 6788 42356
rect 6736 42313 6745 42347
rect 6745 42313 6779 42347
rect 6779 42313 6788 42347
rect 6736 42304 6788 42313
rect 7380 42304 7432 42356
rect 7748 42304 7800 42356
rect 7932 42347 7984 42356
rect 7932 42313 7941 42347
rect 7941 42313 7975 42347
rect 7975 42313 7984 42347
rect 7932 42304 7984 42313
rect 4344 42236 4396 42288
rect 6552 42236 6604 42288
rect 2412 42168 2464 42220
rect 2780 42211 2832 42220
rect 2780 42177 2789 42211
rect 2789 42177 2823 42211
rect 2823 42177 2832 42211
rect 2780 42168 2832 42177
rect 3424 42168 3476 42220
rect 3516 42168 3568 42220
rect 5908 42168 5960 42220
rect 6276 42168 6328 42220
rect 6920 42211 6972 42220
rect 6920 42177 6929 42211
rect 6929 42177 6963 42211
rect 6963 42177 6972 42211
rect 6920 42168 6972 42177
rect 8116 42168 8168 42220
rect 5264 42100 5316 42152
rect 8300 42100 8352 42152
rect 9312 42143 9364 42152
rect 9312 42109 9321 42143
rect 9321 42109 9355 42143
rect 9355 42109 9364 42143
rect 9312 42100 9364 42109
rect 4068 42032 4120 42084
rect 1492 42007 1544 42016
rect 1492 41973 1501 42007
rect 1501 41973 1535 42007
rect 1535 41973 1544 42007
rect 1492 41964 1544 41973
rect 2044 41964 2096 42016
rect 3700 41964 3752 42016
rect 5356 41964 5408 42016
rect 5915 41862 5967 41914
rect 5979 41862 6031 41914
rect 6043 41862 6095 41914
rect 6107 41862 6159 41914
rect 6171 41862 6223 41914
rect 15846 41862 15898 41914
rect 15910 41862 15962 41914
rect 15974 41862 16026 41914
rect 16038 41862 16090 41914
rect 16102 41862 16154 41914
rect 25776 41862 25828 41914
rect 25840 41862 25892 41914
rect 25904 41862 25956 41914
rect 25968 41862 26020 41914
rect 26032 41862 26084 41914
rect 2872 41803 2924 41812
rect 2872 41769 2881 41803
rect 2881 41769 2915 41803
rect 2915 41769 2924 41803
rect 2872 41760 2924 41769
rect 4436 41803 4488 41812
rect 4436 41769 4445 41803
rect 4445 41769 4479 41803
rect 4479 41769 4488 41803
rect 4436 41760 4488 41769
rect 5632 41803 5684 41812
rect 5632 41769 5641 41803
rect 5641 41769 5675 41803
rect 5675 41769 5684 41803
rect 5632 41760 5684 41769
rect 8116 41803 8168 41812
rect 5356 41692 5408 41744
rect 8116 41769 8125 41803
rect 8125 41769 8159 41803
rect 8159 41769 8168 41803
rect 8116 41760 8168 41769
rect 9312 41760 9364 41812
rect 6276 41692 6328 41744
rect 4344 41624 4396 41676
rect 1768 41556 1820 41608
rect 2780 41556 2832 41608
rect 3884 41556 3936 41608
rect 4436 41556 4488 41608
rect 4712 41556 4764 41608
rect 5264 41624 5316 41676
rect 7012 41692 7064 41744
rect 7656 41692 7708 41744
rect 10232 41692 10284 41744
rect 5172 41599 5224 41608
rect 5172 41565 5181 41599
rect 5181 41565 5215 41599
rect 5215 41565 5224 41599
rect 5172 41556 5224 41565
rect 6644 41556 6696 41608
rect 5816 41531 5868 41540
rect 5816 41497 5825 41531
rect 5825 41497 5859 41531
rect 5859 41497 5868 41531
rect 5816 41488 5868 41497
rect 6368 41488 6420 41540
rect 1676 41463 1728 41472
rect 1676 41429 1685 41463
rect 1685 41429 1719 41463
rect 1719 41429 1728 41463
rect 1676 41420 1728 41429
rect 2964 41420 3016 41472
rect 7472 41420 7524 41472
rect 7748 41599 7800 41608
rect 7748 41565 7757 41599
rect 7757 41565 7791 41599
rect 7791 41565 7800 41599
rect 7932 41599 7984 41608
rect 7748 41556 7800 41565
rect 7932 41565 7941 41599
rect 7941 41565 7975 41599
rect 7975 41565 7984 41599
rect 7932 41556 7984 41565
rect 12992 41599 13044 41608
rect 12992 41565 13001 41599
rect 13001 41565 13035 41599
rect 13035 41565 13044 41599
rect 12992 41556 13044 41565
rect 15752 41556 15804 41608
rect 7840 41488 7892 41540
rect 10140 41488 10192 41540
rect 29920 41556 29972 41608
rect 12624 41420 12676 41472
rect 16304 41420 16356 41472
rect 22008 41488 22060 41540
rect 21916 41420 21968 41472
rect 10880 41318 10932 41370
rect 10944 41318 10996 41370
rect 11008 41318 11060 41370
rect 11072 41318 11124 41370
rect 11136 41318 11188 41370
rect 20811 41318 20863 41370
rect 20875 41318 20927 41370
rect 20939 41318 20991 41370
rect 21003 41318 21055 41370
rect 21067 41318 21119 41370
rect 2320 41216 2372 41268
rect 3424 41259 3476 41268
rect 3424 41225 3433 41259
rect 3433 41225 3467 41259
rect 3467 41225 3476 41259
rect 3424 41216 3476 41225
rect 3976 41216 4028 41268
rect 6552 41259 6604 41268
rect 6552 41225 6561 41259
rect 6561 41225 6595 41259
rect 6595 41225 6604 41259
rect 6552 41216 6604 41225
rect 21916 41259 21968 41268
rect 21916 41225 21925 41259
rect 21925 41225 21959 41259
rect 21959 41225 21968 41259
rect 21916 41216 21968 41225
rect 5172 41148 5224 41200
rect 6368 41148 6420 41200
rect 6920 41148 6972 41200
rect 7564 41148 7616 41200
rect 3700 41080 3752 41132
rect 3976 41123 4028 41132
rect 3976 41089 3985 41123
rect 3985 41089 4019 41123
rect 4019 41089 4028 41123
rect 3976 41080 4028 41089
rect 4436 41080 4488 41132
rect 5816 41080 5868 41132
rect 6644 41080 6696 41132
rect 6736 41080 6788 41132
rect 7840 41080 7892 41132
rect 14464 41080 14516 41132
rect 15568 41080 15620 41132
rect 3240 41012 3292 41064
rect 2964 40987 3016 40996
rect 2964 40953 2973 40987
rect 2973 40953 3007 40987
rect 3007 40953 3016 40987
rect 2964 40944 3016 40953
rect 4252 41012 4304 41064
rect 4160 40944 4212 40996
rect 4712 41012 4764 41064
rect 5448 41012 5500 41064
rect 6920 41012 6972 41064
rect 7932 41055 7984 41064
rect 7932 41021 7941 41055
rect 7941 41021 7975 41055
rect 7975 41021 7984 41055
rect 7932 41012 7984 41021
rect 12624 41055 12676 41064
rect 1492 40919 1544 40928
rect 1492 40885 1501 40919
rect 1501 40885 1535 40919
rect 1535 40885 1544 40919
rect 1492 40876 1544 40885
rect 5356 40944 5408 40996
rect 4804 40919 4856 40928
rect 4804 40885 4813 40919
rect 4813 40885 4847 40919
rect 4847 40885 4856 40919
rect 4804 40876 4856 40885
rect 5724 40944 5776 40996
rect 6276 40944 6328 40996
rect 6828 40944 6880 40996
rect 7196 40876 7248 40928
rect 12624 41021 12633 41055
rect 12633 41021 12667 41055
rect 12667 41021 12676 41055
rect 12624 41012 12676 41021
rect 12900 41012 12952 41064
rect 13544 41055 13596 41064
rect 13544 41021 13553 41055
rect 13553 41021 13587 41055
rect 13587 41021 13596 41055
rect 13544 41012 13596 41021
rect 13728 41012 13780 41064
rect 14004 41012 14056 41064
rect 14924 40944 14976 40996
rect 16304 41080 16356 41132
rect 17408 41123 17460 41132
rect 17408 41089 17417 41123
rect 17417 41089 17451 41123
rect 17451 41089 17460 41123
rect 17408 41080 17460 41089
rect 22008 41080 22060 41132
rect 30104 41123 30156 41132
rect 30104 41089 30113 41123
rect 30113 41089 30147 41123
rect 30147 41089 30156 41123
rect 30104 41080 30156 41089
rect 14740 40876 14792 40928
rect 16488 40876 16540 40928
rect 16672 40919 16724 40928
rect 16672 40885 16681 40919
rect 16681 40885 16715 40919
rect 16715 40885 16724 40919
rect 16672 40876 16724 40885
rect 17040 40876 17092 40928
rect 5915 40774 5967 40826
rect 5979 40774 6031 40826
rect 6043 40774 6095 40826
rect 6107 40774 6159 40826
rect 6171 40774 6223 40826
rect 15846 40774 15898 40826
rect 15910 40774 15962 40826
rect 15974 40774 16026 40826
rect 16038 40774 16090 40826
rect 16102 40774 16154 40826
rect 25776 40774 25828 40826
rect 25840 40774 25892 40826
rect 25904 40774 25956 40826
rect 25968 40774 26020 40826
rect 26032 40774 26084 40826
rect 3976 40672 4028 40724
rect 2228 40604 2280 40656
rect 4252 40579 4304 40588
rect 4252 40545 4261 40579
rect 4261 40545 4295 40579
rect 4295 40545 4304 40579
rect 4252 40536 4304 40545
rect 1952 40468 2004 40520
rect 2780 40468 2832 40520
rect 3976 40511 4028 40520
rect 3976 40477 3985 40511
rect 3985 40477 4019 40511
rect 4019 40477 4028 40511
rect 3976 40468 4028 40477
rect 4160 40511 4212 40520
rect 4160 40477 4169 40511
rect 4169 40477 4203 40511
rect 4203 40477 4212 40511
rect 4160 40468 4212 40477
rect 4436 40468 4488 40520
rect 4620 40468 4672 40520
rect 5080 40468 5132 40520
rect 6460 40604 6512 40656
rect 6736 40672 6788 40724
rect 6828 40672 6880 40724
rect 12992 40672 13044 40724
rect 17316 40672 17368 40724
rect 7288 40604 7340 40656
rect 7748 40536 7800 40588
rect 5448 40400 5500 40452
rect 1492 40375 1544 40384
rect 1492 40341 1501 40375
rect 1501 40341 1535 40375
rect 1535 40341 1544 40375
rect 1492 40332 1544 40341
rect 3056 40332 3108 40384
rect 3792 40375 3844 40384
rect 3792 40341 3801 40375
rect 3801 40341 3835 40375
rect 3835 40341 3844 40375
rect 3792 40332 3844 40341
rect 6552 40468 6604 40520
rect 6920 40468 6972 40520
rect 8576 40468 8628 40520
rect 9772 40511 9824 40520
rect 9772 40477 9781 40511
rect 9781 40477 9815 40511
rect 9815 40477 9824 40511
rect 9772 40468 9824 40477
rect 13544 40536 13596 40588
rect 16856 40604 16908 40656
rect 14740 40579 14792 40588
rect 14740 40545 14749 40579
rect 14749 40545 14783 40579
rect 14783 40545 14792 40579
rect 14740 40536 14792 40545
rect 16672 40536 16724 40588
rect 16764 40579 16816 40588
rect 16764 40545 16773 40579
rect 16773 40545 16807 40579
rect 16807 40545 16816 40579
rect 17040 40579 17092 40588
rect 16764 40536 16816 40545
rect 17040 40545 17049 40579
rect 17049 40545 17083 40579
rect 17083 40545 17092 40579
rect 17040 40536 17092 40545
rect 17500 40536 17552 40588
rect 12992 40511 13044 40520
rect 12992 40477 13001 40511
rect 13001 40477 13035 40511
rect 13035 40477 13044 40511
rect 12992 40468 13044 40477
rect 16304 40511 16356 40520
rect 16304 40477 16313 40511
rect 16313 40477 16347 40511
rect 16347 40477 16356 40511
rect 16304 40468 16356 40477
rect 17316 40511 17368 40520
rect 17316 40477 17325 40511
rect 17325 40477 17359 40511
rect 17359 40477 17368 40511
rect 17316 40468 17368 40477
rect 18604 40511 18656 40520
rect 18604 40477 18613 40511
rect 18613 40477 18647 40511
rect 18647 40477 18656 40511
rect 18604 40468 18656 40477
rect 6736 40400 6788 40452
rect 8944 40332 8996 40384
rect 9128 40375 9180 40384
rect 9128 40341 9137 40375
rect 9137 40341 9171 40375
rect 9171 40341 9180 40375
rect 9128 40332 9180 40341
rect 13820 40332 13872 40384
rect 14832 40375 14884 40384
rect 14832 40341 14841 40375
rect 14841 40341 14875 40375
rect 14875 40341 14884 40375
rect 14832 40332 14884 40341
rect 19800 40400 19852 40452
rect 17960 40375 18012 40384
rect 17960 40341 17969 40375
rect 17969 40341 18003 40375
rect 18003 40341 18012 40375
rect 17960 40332 18012 40341
rect 18420 40375 18472 40384
rect 18420 40341 18429 40375
rect 18429 40341 18463 40375
rect 18463 40341 18472 40375
rect 18420 40332 18472 40341
rect 10880 40230 10932 40282
rect 10944 40230 10996 40282
rect 11008 40230 11060 40282
rect 11072 40230 11124 40282
rect 11136 40230 11188 40282
rect 20811 40230 20863 40282
rect 20875 40230 20927 40282
rect 20939 40230 20991 40282
rect 21003 40230 21055 40282
rect 21067 40230 21119 40282
rect 3976 40128 4028 40180
rect 4804 40128 4856 40180
rect 3792 40060 3844 40112
rect 7288 40060 7340 40112
rect 7932 40128 7984 40180
rect 8576 40171 8628 40180
rect 8576 40137 8585 40171
rect 8585 40137 8619 40171
rect 8619 40137 8628 40171
rect 8576 40128 8628 40137
rect 2964 39992 3016 40044
rect 5724 39992 5776 40044
rect 6736 39992 6788 40044
rect 7196 39992 7248 40044
rect 7380 39992 7432 40044
rect 8024 40060 8076 40112
rect 14832 40128 14884 40180
rect 16580 40128 16632 40180
rect 15568 40103 15620 40112
rect 15568 40069 15577 40103
rect 15577 40069 15611 40103
rect 15611 40069 15620 40103
rect 15568 40060 15620 40069
rect 16488 40060 16540 40112
rect 17408 40128 17460 40180
rect 18420 40128 18472 40180
rect 17960 40103 18012 40112
rect 12624 39992 12676 40044
rect 12900 39992 12952 40044
rect 15660 39992 15712 40044
rect 17960 40069 17969 40103
rect 17969 40069 18003 40103
rect 18003 40069 18012 40103
rect 17960 40060 18012 40069
rect 18052 40060 18104 40112
rect 19800 40103 19852 40112
rect 19800 40069 19809 40103
rect 19809 40069 19843 40103
rect 19843 40069 19852 40103
rect 19800 40060 19852 40069
rect 18696 40035 18748 40044
rect 18696 40001 18705 40035
rect 18705 40001 18739 40035
rect 18739 40001 18748 40035
rect 18696 39992 18748 40001
rect 2872 39967 2924 39976
rect 2872 39933 2881 39967
rect 2881 39933 2915 39967
rect 2915 39933 2924 39967
rect 2872 39924 2924 39933
rect 13544 39924 13596 39976
rect 13820 39967 13872 39976
rect 13820 39933 13854 39967
rect 13854 39933 13872 39967
rect 13820 39924 13872 39933
rect 14004 39967 14056 39976
rect 14004 39933 14013 39967
rect 14013 39933 14047 39967
rect 14047 39933 14056 39967
rect 14004 39924 14056 39933
rect 16212 39924 16264 39976
rect 16764 39924 16816 39976
rect 18880 39924 18932 39976
rect 4528 39856 4580 39908
rect 2228 39831 2280 39840
rect 2228 39797 2237 39831
rect 2237 39797 2271 39831
rect 2271 39797 2280 39831
rect 2228 39788 2280 39797
rect 3516 39788 3568 39840
rect 4344 39788 4396 39840
rect 4896 39788 4948 39840
rect 5356 39788 5408 39840
rect 6920 39831 6972 39840
rect 6920 39797 6929 39831
rect 6929 39797 6963 39831
rect 6963 39797 6972 39831
rect 6920 39788 6972 39797
rect 9680 39831 9732 39840
rect 9680 39797 9689 39831
rect 9689 39797 9723 39831
rect 9723 39797 9732 39831
rect 9680 39788 9732 39797
rect 15752 39856 15804 39908
rect 15660 39788 15712 39840
rect 19432 39788 19484 39840
rect 20076 39788 20128 39840
rect 5915 39686 5967 39738
rect 5979 39686 6031 39738
rect 6043 39686 6095 39738
rect 6107 39686 6159 39738
rect 6171 39686 6223 39738
rect 15846 39686 15898 39738
rect 15910 39686 15962 39738
rect 15974 39686 16026 39738
rect 16038 39686 16090 39738
rect 16102 39686 16154 39738
rect 25776 39686 25828 39738
rect 25840 39686 25892 39738
rect 25904 39686 25956 39738
rect 25968 39686 26020 39738
rect 26032 39686 26084 39738
rect 2872 39627 2924 39636
rect 2872 39593 2881 39627
rect 2881 39593 2915 39627
rect 2915 39593 2924 39627
rect 2872 39584 2924 39593
rect 5816 39627 5868 39636
rect 5816 39593 5825 39627
rect 5825 39593 5859 39627
rect 5859 39593 5868 39627
rect 5816 39584 5868 39593
rect 6644 39584 6696 39636
rect 4528 39516 4580 39568
rect 7012 39516 7064 39568
rect 8024 39584 8076 39636
rect 8852 39516 8904 39568
rect 1584 39380 1636 39432
rect 4068 39448 4120 39500
rect 6368 39448 6420 39500
rect 9680 39584 9732 39636
rect 12992 39627 13044 39636
rect 12992 39593 13001 39627
rect 13001 39593 13035 39627
rect 13035 39593 13044 39627
rect 12992 39584 13044 39593
rect 15660 39584 15712 39636
rect 18604 39584 18656 39636
rect 22284 39516 22336 39568
rect 3056 39423 3108 39432
rect 3056 39389 3065 39423
rect 3065 39389 3099 39423
rect 3099 39389 3108 39423
rect 3056 39380 3108 39389
rect 3792 39423 3844 39432
rect 3792 39389 3801 39423
rect 3801 39389 3835 39423
rect 3835 39389 3844 39423
rect 3792 39380 3844 39389
rect 1492 39287 1544 39296
rect 1492 39253 1501 39287
rect 1501 39253 1535 39287
rect 1535 39253 1544 39287
rect 1492 39244 1544 39253
rect 2228 39287 2280 39296
rect 2228 39253 2237 39287
rect 2237 39253 2271 39287
rect 2271 39253 2280 39287
rect 2228 39244 2280 39253
rect 3976 39287 4028 39296
rect 3976 39253 3985 39287
rect 3985 39253 4019 39287
rect 4019 39253 4028 39287
rect 3976 39244 4028 39253
rect 4712 39287 4764 39296
rect 4712 39253 4721 39287
rect 4721 39253 4755 39287
rect 4755 39253 4764 39287
rect 4712 39244 4764 39253
rect 5816 39380 5868 39432
rect 6460 39423 6512 39432
rect 6460 39389 6469 39423
rect 6469 39389 6503 39423
rect 6503 39389 6512 39423
rect 6460 39380 6512 39389
rect 6644 39423 6696 39432
rect 6644 39389 6653 39423
rect 6653 39389 6687 39423
rect 6687 39389 6696 39423
rect 6644 39380 6696 39389
rect 6736 39423 6788 39432
rect 6736 39389 6745 39423
rect 6745 39389 6779 39423
rect 6779 39389 6788 39423
rect 6736 39380 6788 39389
rect 6920 39380 6972 39432
rect 14280 39448 14332 39500
rect 15016 39448 15068 39500
rect 15384 39448 15436 39500
rect 16856 39448 16908 39500
rect 12900 39380 12952 39432
rect 14832 39423 14884 39432
rect 14832 39389 14841 39423
rect 14841 39389 14875 39423
rect 14875 39389 14884 39423
rect 14832 39380 14884 39389
rect 15568 39423 15620 39432
rect 15568 39389 15577 39423
rect 15577 39389 15611 39423
rect 15611 39389 15620 39423
rect 15844 39423 15896 39432
rect 15568 39380 15620 39389
rect 15844 39389 15853 39423
rect 15853 39389 15887 39423
rect 15887 39389 15896 39423
rect 15844 39380 15896 39389
rect 17960 39380 18012 39432
rect 19432 39423 19484 39432
rect 19432 39389 19441 39423
rect 19441 39389 19475 39423
rect 19475 39389 19484 39423
rect 19432 39380 19484 39389
rect 30104 39423 30156 39432
rect 9680 39355 9732 39364
rect 9680 39321 9714 39355
rect 9714 39321 9732 39355
rect 9680 39312 9732 39321
rect 14096 39312 14148 39364
rect 14464 39312 14516 39364
rect 18052 39312 18104 39364
rect 18880 39312 18932 39364
rect 20260 39355 20312 39364
rect 20260 39321 20269 39355
rect 20269 39321 20303 39355
rect 20303 39321 20312 39355
rect 20260 39312 20312 39321
rect 22008 39312 22060 39364
rect 6828 39244 6880 39296
rect 7196 39287 7248 39296
rect 7196 39253 7205 39287
rect 7205 39253 7239 39287
rect 7239 39253 7248 39287
rect 7196 39244 7248 39253
rect 10784 39287 10836 39296
rect 10784 39253 10793 39287
rect 10793 39253 10827 39287
rect 10827 39253 10836 39287
rect 10784 39244 10836 39253
rect 15016 39244 15068 39296
rect 15568 39244 15620 39296
rect 16120 39244 16172 39296
rect 18696 39244 18748 39296
rect 19156 39244 19208 39296
rect 19800 39244 19852 39296
rect 21548 39287 21600 39296
rect 21548 39253 21557 39287
rect 21557 39253 21591 39287
rect 21591 39253 21600 39287
rect 21548 39244 21600 39253
rect 30104 39389 30113 39423
rect 30113 39389 30147 39423
rect 30147 39389 30156 39423
rect 30104 39380 30156 39389
rect 10880 39142 10932 39194
rect 10944 39142 10996 39194
rect 11008 39142 11060 39194
rect 11072 39142 11124 39194
rect 11136 39142 11188 39194
rect 20811 39142 20863 39194
rect 20875 39142 20927 39194
rect 20939 39142 20991 39194
rect 21003 39142 21055 39194
rect 21067 39142 21119 39194
rect 2504 39040 2556 39092
rect 6368 39040 6420 39092
rect 13544 39083 13596 39092
rect 13544 39049 13553 39083
rect 13553 39049 13587 39083
rect 13587 39049 13596 39083
rect 13544 39040 13596 39049
rect 15292 39040 15344 39092
rect 16120 39083 16172 39092
rect 16120 39049 16129 39083
rect 16129 39049 16163 39083
rect 16163 39049 16172 39083
rect 16120 39040 16172 39049
rect 19156 39083 19208 39092
rect 19156 39049 19165 39083
rect 19165 39049 19199 39083
rect 19199 39049 19208 39083
rect 19156 39040 19208 39049
rect 20260 39083 20312 39092
rect 20260 39049 20269 39083
rect 20269 39049 20303 39083
rect 20303 39049 20312 39083
rect 20260 39040 20312 39049
rect 3148 38904 3200 38956
rect 4712 38972 4764 39024
rect 4160 38904 4212 38956
rect 4436 38947 4488 38956
rect 4436 38913 4445 38947
rect 4445 38913 4479 38947
rect 4479 38913 4488 38947
rect 4436 38904 4488 38913
rect 4620 38947 4672 38956
rect 4620 38913 4629 38947
rect 4629 38913 4663 38947
rect 4663 38913 4672 38947
rect 4620 38904 4672 38913
rect 5816 38947 5868 38956
rect 5816 38913 5825 38947
rect 5825 38913 5859 38947
rect 5859 38913 5868 38947
rect 5816 38904 5868 38913
rect 7196 38972 7248 39024
rect 13820 39015 13872 39024
rect 13820 38981 13829 39015
rect 13829 38981 13863 39015
rect 13863 38981 13872 39015
rect 13820 38972 13872 38981
rect 18696 38972 18748 39024
rect 9128 38904 9180 38956
rect 9496 38947 9548 38956
rect 9496 38913 9530 38947
rect 9530 38913 9548 38947
rect 9496 38904 9548 38913
rect 12624 38904 12676 38956
rect 14280 38947 14332 38956
rect 14280 38913 14289 38947
rect 14289 38913 14323 38947
rect 14323 38913 14332 38947
rect 14280 38904 14332 38913
rect 15292 38947 15344 38956
rect 15292 38913 15326 38947
rect 15326 38913 15344 38947
rect 20076 38947 20128 38956
rect 15292 38904 15344 38913
rect 20076 38913 20085 38947
rect 20085 38913 20119 38947
rect 20119 38913 20128 38947
rect 20076 38904 20128 38913
rect 2964 38836 3016 38888
rect 4252 38879 4304 38888
rect 4252 38845 4261 38879
rect 4261 38845 4295 38879
rect 4295 38845 4304 38879
rect 4252 38836 4304 38845
rect 4344 38879 4396 38888
rect 4344 38845 4353 38879
rect 4353 38845 4387 38879
rect 4387 38845 4396 38879
rect 4344 38836 4396 38845
rect 14004 38836 14056 38888
rect 14832 38836 14884 38888
rect 15200 38879 15252 38888
rect 2872 38768 2924 38820
rect 4988 38768 5040 38820
rect 15200 38845 15209 38879
rect 15209 38845 15243 38879
rect 15243 38845 15252 38879
rect 15200 38836 15252 38845
rect 15844 38836 15896 38888
rect 16212 38836 16264 38888
rect 18880 38879 18932 38888
rect 18880 38845 18889 38879
rect 18889 38845 18923 38879
rect 18923 38845 18932 38879
rect 18880 38836 18932 38845
rect 1952 38700 2004 38752
rect 2320 38700 2372 38752
rect 3056 38743 3108 38752
rect 3056 38709 3065 38743
rect 3065 38709 3099 38743
rect 3099 38709 3108 38743
rect 3056 38700 3108 38709
rect 4252 38700 4304 38752
rect 5724 38743 5776 38752
rect 5724 38709 5733 38743
rect 5733 38709 5767 38743
rect 5767 38709 5776 38743
rect 5724 38700 5776 38709
rect 6460 38700 6512 38752
rect 7012 38700 7064 38752
rect 9220 38700 9272 38752
rect 14924 38700 14976 38752
rect 20260 38700 20312 38752
rect 5915 38598 5967 38650
rect 5979 38598 6031 38650
rect 6043 38598 6095 38650
rect 6107 38598 6159 38650
rect 6171 38598 6223 38650
rect 15846 38598 15898 38650
rect 15910 38598 15962 38650
rect 15974 38598 16026 38650
rect 16038 38598 16090 38650
rect 16102 38598 16154 38650
rect 25776 38598 25828 38650
rect 25840 38598 25892 38650
rect 25904 38598 25956 38650
rect 25968 38598 26020 38650
rect 26032 38598 26084 38650
rect 1952 38496 2004 38548
rect 2136 38496 2188 38548
rect 4160 38496 4212 38548
rect 2964 38428 3016 38480
rect 2872 38403 2924 38412
rect 2872 38369 2881 38403
rect 2881 38369 2915 38403
rect 2915 38369 2924 38403
rect 2872 38360 2924 38369
rect 2688 38335 2740 38344
rect 2688 38301 2697 38335
rect 2697 38301 2731 38335
rect 2731 38301 2740 38335
rect 2688 38292 2740 38301
rect 3976 38403 4028 38412
rect 3976 38369 3985 38403
rect 3985 38369 4019 38403
rect 4019 38369 4028 38403
rect 3976 38360 4028 38369
rect 4988 38360 5040 38412
rect 3148 38292 3200 38344
rect 4068 38292 4120 38344
rect 4252 38335 4304 38344
rect 4252 38301 4286 38335
rect 4286 38301 4304 38335
rect 4252 38292 4304 38301
rect 5816 38335 5868 38344
rect 5816 38301 5825 38335
rect 5825 38301 5859 38335
rect 5859 38301 5868 38335
rect 9312 38496 9364 38548
rect 9404 38496 9456 38548
rect 7012 38428 7064 38480
rect 6920 38360 6972 38412
rect 7288 38335 7340 38344
rect 5816 38292 5868 38301
rect 7288 38301 7297 38335
rect 7297 38301 7331 38335
rect 7331 38301 7340 38335
rect 7288 38292 7340 38301
rect 7380 38292 7432 38344
rect 7656 38335 7708 38344
rect 7656 38301 7665 38335
rect 7665 38301 7699 38335
rect 7699 38301 7708 38335
rect 7656 38292 7708 38301
rect 2504 38199 2556 38208
rect 2504 38165 2513 38199
rect 2513 38165 2547 38199
rect 2547 38165 2556 38199
rect 2504 38156 2556 38165
rect 4344 38156 4396 38208
rect 7104 38199 7156 38208
rect 7104 38165 7113 38199
rect 7113 38165 7147 38199
rect 7147 38165 7156 38199
rect 7104 38156 7156 38165
rect 8760 38360 8812 38412
rect 8668 38224 8720 38276
rect 9036 38292 9088 38344
rect 9312 38335 9364 38344
rect 9312 38301 9321 38335
rect 9321 38301 9355 38335
rect 9355 38301 9364 38335
rect 9312 38292 9364 38301
rect 10784 38428 10836 38480
rect 12900 38496 12952 38548
rect 14832 38496 14884 38548
rect 17408 38539 17460 38548
rect 17408 38505 17417 38539
rect 17417 38505 17451 38539
rect 17451 38505 17460 38539
rect 17408 38496 17460 38505
rect 19432 38496 19484 38548
rect 9588 38360 9640 38412
rect 9680 38335 9732 38344
rect 9680 38301 9689 38335
rect 9689 38301 9723 38335
rect 9723 38301 9732 38335
rect 9680 38292 9732 38301
rect 10600 38292 10652 38344
rect 12716 38292 12768 38344
rect 13176 38335 13228 38344
rect 13176 38301 13185 38335
rect 13185 38301 13219 38335
rect 13219 38301 13228 38335
rect 13176 38292 13228 38301
rect 17592 38335 17644 38344
rect 17592 38301 17601 38335
rect 17601 38301 17635 38335
rect 17635 38301 17644 38335
rect 17592 38292 17644 38301
rect 18420 38335 18472 38344
rect 18420 38301 18429 38335
rect 18429 38301 18463 38335
rect 18463 38301 18472 38335
rect 18420 38292 18472 38301
rect 30104 38335 30156 38344
rect 30104 38301 30113 38335
rect 30113 38301 30147 38335
rect 30147 38301 30156 38335
rect 30104 38292 30156 38301
rect 8852 38156 8904 38208
rect 9588 38156 9640 38208
rect 9956 38156 10008 38208
rect 12532 38156 12584 38208
rect 21548 38224 21600 38276
rect 17316 38156 17368 38208
rect 18972 38156 19024 38208
rect 29920 38199 29972 38208
rect 29920 38165 29929 38199
rect 29929 38165 29963 38199
rect 29963 38165 29972 38199
rect 29920 38156 29972 38165
rect 10880 38054 10932 38106
rect 10944 38054 10996 38106
rect 11008 38054 11060 38106
rect 11072 38054 11124 38106
rect 11136 38054 11188 38106
rect 20811 38054 20863 38106
rect 20875 38054 20927 38106
rect 20939 38054 20991 38106
rect 21003 38054 21055 38106
rect 21067 38054 21119 38106
rect 1860 37952 1912 38004
rect 2688 37952 2740 38004
rect 3148 37952 3200 38004
rect 3700 37952 3752 38004
rect 7472 37952 7524 38004
rect 2504 37884 2556 37936
rect 6368 37884 6420 37936
rect 6552 37884 6604 37936
rect 9496 37952 9548 38004
rect 12716 37995 12768 38004
rect 12716 37961 12725 37995
rect 12725 37961 12759 37995
rect 12759 37961 12768 37995
rect 12716 37952 12768 37961
rect 15108 37952 15160 38004
rect 17316 37952 17368 38004
rect 4344 37816 4396 37868
rect 5724 37816 5776 37868
rect 8024 37859 8076 37868
rect 2964 37748 3016 37800
rect 4436 37791 4488 37800
rect 4436 37757 4445 37791
rect 4445 37757 4479 37791
rect 4479 37757 4488 37791
rect 4436 37748 4488 37757
rect 6368 37791 6420 37800
rect 6368 37757 6377 37791
rect 6377 37757 6411 37791
rect 6411 37757 6420 37791
rect 6368 37748 6420 37757
rect 8024 37825 8033 37859
rect 8033 37825 8067 37859
rect 8067 37825 8076 37859
rect 8024 37816 8076 37825
rect 8300 37816 8352 37868
rect 8668 37859 8720 37868
rect 8668 37825 8677 37859
rect 8677 37825 8711 37859
rect 8711 37825 8720 37859
rect 8668 37816 8720 37825
rect 8852 37859 8904 37868
rect 8852 37825 8861 37859
rect 8861 37825 8895 37859
rect 8895 37825 8904 37859
rect 8852 37816 8904 37825
rect 9220 37859 9272 37868
rect 9220 37825 9229 37859
rect 9229 37825 9263 37859
rect 9263 37825 9272 37859
rect 9956 37859 10008 37868
rect 9220 37816 9272 37825
rect 4620 37680 4672 37732
rect 8484 37748 8536 37800
rect 8760 37748 8812 37800
rect 9128 37748 9180 37800
rect 9312 37748 9364 37800
rect 9956 37825 9965 37859
rect 9965 37825 9999 37859
rect 9999 37825 10008 37859
rect 9956 37816 10008 37825
rect 10048 37816 10100 37868
rect 10600 37859 10652 37868
rect 10600 37825 10609 37859
rect 10609 37825 10643 37859
rect 10643 37825 10652 37859
rect 10600 37816 10652 37825
rect 1952 37612 2004 37664
rect 4160 37612 4212 37664
rect 5448 37612 5500 37664
rect 12532 37884 12584 37936
rect 17408 37884 17460 37936
rect 18052 37884 18104 37936
rect 12624 37816 12676 37868
rect 13084 37859 13136 37868
rect 13084 37825 13093 37859
rect 13093 37825 13127 37859
rect 13127 37825 13136 37859
rect 13084 37816 13136 37825
rect 14004 37859 14056 37868
rect 14004 37825 14013 37859
rect 14013 37825 14047 37859
rect 14047 37825 14056 37859
rect 14004 37816 14056 37825
rect 14924 37859 14976 37868
rect 14924 37825 14933 37859
rect 14933 37825 14967 37859
rect 14967 37825 14976 37859
rect 14924 37816 14976 37825
rect 17868 37859 17920 37868
rect 17868 37825 17877 37859
rect 17877 37825 17911 37859
rect 17911 37825 17920 37859
rect 17868 37816 17920 37825
rect 18420 37884 18472 37936
rect 20720 37884 20772 37936
rect 18972 37859 19024 37868
rect 18972 37825 18981 37859
rect 18981 37825 19015 37859
rect 19015 37825 19024 37859
rect 18972 37816 19024 37825
rect 19248 37859 19300 37868
rect 19248 37825 19282 37859
rect 19282 37825 19300 37859
rect 19248 37816 19300 37825
rect 22008 37816 22060 37868
rect 14280 37791 14332 37800
rect 14280 37757 14289 37791
rect 14289 37757 14323 37791
rect 14323 37757 14332 37791
rect 14280 37748 14332 37757
rect 29920 37748 29972 37800
rect 17592 37680 17644 37732
rect 9312 37612 9364 37664
rect 10876 37612 10928 37664
rect 11520 37655 11572 37664
rect 11520 37621 11529 37655
rect 11529 37621 11563 37655
rect 11563 37621 11572 37655
rect 11520 37612 11572 37621
rect 12716 37612 12768 37664
rect 14188 37655 14240 37664
rect 14188 37621 14197 37655
rect 14197 37621 14231 37655
rect 14231 37621 14240 37655
rect 14188 37612 14240 37621
rect 17960 37612 18012 37664
rect 19340 37612 19392 37664
rect 20352 37655 20404 37664
rect 20352 37621 20361 37655
rect 20361 37621 20395 37655
rect 20395 37621 20404 37655
rect 20352 37612 20404 37621
rect 5915 37510 5967 37562
rect 5979 37510 6031 37562
rect 6043 37510 6095 37562
rect 6107 37510 6159 37562
rect 6171 37510 6223 37562
rect 15846 37510 15898 37562
rect 15910 37510 15962 37562
rect 15974 37510 16026 37562
rect 16038 37510 16090 37562
rect 16102 37510 16154 37562
rect 25776 37510 25828 37562
rect 25840 37510 25892 37562
rect 25904 37510 25956 37562
rect 25968 37510 26020 37562
rect 26032 37510 26084 37562
rect 1952 37408 2004 37460
rect 7288 37408 7340 37460
rect 7196 37340 7248 37392
rect 13176 37408 13228 37460
rect 14188 37408 14240 37460
rect 15108 37408 15160 37460
rect 16304 37408 16356 37460
rect 13084 37340 13136 37392
rect 2320 37204 2372 37256
rect 5448 37272 5500 37324
rect 10876 37315 10928 37324
rect 10876 37281 10885 37315
rect 10885 37281 10919 37315
rect 10919 37281 10928 37315
rect 10876 37272 10928 37281
rect 12624 37272 12676 37324
rect 2596 37204 2648 37256
rect 2964 37204 3016 37256
rect 3976 37247 4028 37256
rect 3976 37213 3985 37247
rect 3985 37213 4019 37247
rect 4019 37213 4028 37247
rect 3976 37204 4028 37213
rect 4988 37204 5040 37256
rect 7104 37204 7156 37256
rect 9680 37204 9732 37256
rect 9772 37204 9824 37256
rect 12716 37247 12768 37256
rect 12716 37213 12725 37247
rect 12725 37213 12759 37247
rect 12759 37213 12768 37247
rect 12716 37204 12768 37213
rect 14096 37247 14148 37256
rect 14096 37213 14105 37247
rect 14105 37213 14139 37247
rect 14139 37213 14148 37247
rect 14096 37204 14148 37213
rect 15200 37272 15252 37324
rect 15568 37315 15620 37324
rect 15568 37281 15577 37315
rect 15577 37281 15611 37315
rect 15611 37281 15620 37315
rect 15568 37272 15620 37281
rect 16304 37272 16356 37324
rect 17868 37315 17920 37324
rect 15108 37247 15160 37256
rect 9036 37136 9088 37188
rect 11244 37136 11296 37188
rect 13084 37136 13136 37188
rect 15108 37213 15117 37247
rect 15117 37213 15151 37247
rect 15151 37213 15160 37247
rect 15108 37204 15160 37213
rect 16120 37247 16172 37256
rect 16120 37213 16129 37247
rect 16129 37213 16163 37247
rect 16163 37213 16172 37247
rect 16120 37204 16172 37213
rect 14556 37136 14608 37188
rect 17868 37281 17877 37315
rect 17877 37281 17911 37315
rect 17911 37281 17920 37315
rect 17868 37272 17920 37281
rect 17960 37247 18012 37256
rect 17960 37213 17969 37247
rect 17969 37213 18003 37247
rect 18003 37213 18012 37247
rect 17960 37204 18012 37213
rect 19340 37204 19392 37256
rect 19984 37204 20036 37256
rect 20352 37204 20404 37256
rect 2412 37111 2464 37120
rect 2412 37077 2421 37111
rect 2421 37077 2455 37111
rect 2455 37077 2464 37111
rect 2412 37068 2464 37077
rect 2872 37068 2924 37120
rect 3056 37111 3108 37120
rect 3056 37077 3065 37111
rect 3065 37077 3099 37111
rect 3099 37077 3108 37111
rect 3056 37068 3108 37077
rect 3792 37111 3844 37120
rect 3792 37077 3801 37111
rect 3801 37077 3835 37111
rect 3835 37077 3844 37111
rect 3792 37068 3844 37077
rect 3884 37068 3936 37120
rect 8576 37068 8628 37120
rect 8760 37068 8812 37120
rect 11428 37068 11480 37120
rect 15292 37068 15344 37120
rect 16212 37068 16264 37120
rect 20076 37136 20128 37188
rect 16764 37111 16816 37120
rect 16764 37077 16773 37111
rect 16773 37077 16807 37111
rect 16807 37077 16816 37111
rect 16764 37068 16816 37077
rect 18144 37068 18196 37120
rect 18420 37068 18472 37120
rect 20352 37111 20404 37120
rect 20352 37077 20361 37111
rect 20361 37077 20395 37111
rect 20395 37077 20404 37111
rect 20352 37068 20404 37077
rect 10880 36966 10932 37018
rect 10944 36966 10996 37018
rect 11008 36966 11060 37018
rect 11072 36966 11124 37018
rect 11136 36966 11188 37018
rect 20811 36966 20863 37018
rect 20875 36966 20927 37018
rect 20939 36966 20991 37018
rect 21003 36966 21055 37018
rect 21067 36966 21119 37018
rect 1400 36864 1452 36916
rect 2596 36864 2648 36916
rect 4436 36864 4488 36916
rect 4988 36907 5040 36916
rect 4988 36873 4997 36907
rect 4997 36873 5031 36907
rect 5031 36873 5040 36907
rect 4988 36864 5040 36873
rect 6828 36864 6880 36916
rect 6736 36796 6788 36848
rect 9036 36864 9088 36916
rect 9864 36864 9916 36916
rect 10324 36864 10376 36916
rect 2044 36728 2096 36780
rect 2780 36728 2832 36780
rect 2412 36592 2464 36644
rect 4160 36728 4212 36780
rect 5172 36728 5224 36780
rect 5632 36771 5684 36780
rect 5632 36737 5641 36771
rect 5641 36737 5675 36771
rect 5675 36737 5684 36771
rect 5632 36728 5684 36737
rect 4896 36660 4948 36712
rect 7196 36728 7248 36780
rect 8300 36728 8352 36780
rect 8392 36771 8444 36780
rect 8392 36737 8401 36771
rect 8401 36737 8435 36771
rect 8435 36737 8444 36771
rect 8760 36771 8812 36780
rect 8392 36728 8444 36737
rect 8760 36737 8769 36771
rect 8769 36737 8803 36771
rect 8803 36737 8812 36771
rect 8760 36728 8812 36737
rect 9680 36796 9732 36848
rect 10416 36771 10468 36780
rect 8484 36703 8536 36712
rect 1400 36524 1452 36576
rect 2320 36567 2372 36576
rect 2320 36533 2329 36567
rect 2329 36533 2363 36567
rect 2363 36533 2372 36567
rect 2320 36524 2372 36533
rect 3976 36592 4028 36644
rect 8484 36669 8493 36703
rect 8493 36669 8527 36703
rect 8527 36669 8536 36703
rect 8484 36660 8536 36669
rect 9036 36660 9088 36712
rect 10416 36737 10425 36771
rect 10425 36737 10459 36771
rect 10459 36737 10468 36771
rect 10416 36728 10468 36737
rect 10508 36771 10560 36780
rect 10508 36737 10517 36771
rect 10517 36737 10551 36771
rect 10551 36737 10560 36771
rect 13084 36796 13136 36848
rect 10508 36728 10560 36737
rect 11520 36771 11572 36780
rect 11520 36737 11529 36771
rect 11529 36737 11563 36771
rect 11563 36737 11572 36771
rect 11520 36728 11572 36737
rect 10324 36660 10376 36712
rect 10692 36660 10744 36712
rect 13268 36728 13320 36780
rect 7656 36592 7708 36644
rect 8392 36592 8444 36644
rect 6644 36524 6696 36576
rect 9220 36524 9272 36576
rect 9588 36524 9640 36576
rect 9956 36524 10008 36576
rect 11888 36524 11940 36576
rect 15108 36864 15160 36916
rect 16764 36864 16816 36916
rect 17868 36864 17920 36916
rect 14188 36771 14240 36780
rect 14188 36737 14197 36771
rect 14197 36737 14231 36771
rect 14231 36737 14240 36771
rect 14188 36728 14240 36737
rect 14556 36771 14608 36780
rect 14556 36737 14565 36771
rect 14565 36737 14599 36771
rect 14599 36737 14608 36771
rect 14556 36728 14608 36737
rect 14832 36728 14884 36780
rect 19064 36796 19116 36848
rect 20444 36796 20496 36848
rect 14096 36660 14148 36712
rect 14648 36660 14700 36712
rect 15292 36703 15344 36712
rect 15292 36669 15301 36703
rect 15301 36669 15335 36703
rect 15335 36669 15344 36703
rect 15292 36660 15344 36669
rect 18420 36728 18472 36780
rect 18604 36771 18656 36780
rect 18604 36737 18638 36771
rect 18638 36737 18656 36771
rect 20536 36771 20588 36780
rect 18604 36728 18656 36737
rect 20536 36737 20545 36771
rect 20545 36737 20579 36771
rect 20579 36737 20588 36771
rect 20536 36728 20588 36737
rect 14372 36592 14424 36644
rect 15200 36524 15252 36576
rect 16764 36660 16816 36712
rect 17040 36703 17092 36712
rect 17040 36669 17049 36703
rect 17049 36669 17083 36703
rect 17083 36669 17092 36703
rect 17040 36660 17092 36669
rect 20628 36703 20680 36712
rect 20628 36669 20637 36703
rect 20637 36669 20671 36703
rect 20671 36669 20680 36703
rect 20628 36660 20680 36669
rect 21364 36728 21416 36780
rect 22008 36728 22060 36780
rect 30104 36771 30156 36780
rect 30104 36737 30113 36771
rect 30113 36737 30147 36771
rect 30147 36737 30156 36771
rect 30104 36728 30156 36737
rect 19984 36592 20036 36644
rect 19800 36524 19852 36576
rect 20812 36524 20864 36576
rect 5915 36422 5967 36474
rect 5979 36422 6031 36474
rect 6043 36422 6095 36474
rect 6107 36422 6159 36474
rect 6171 36422 6223 36474
rect 15846 36422 15898 36474
rect 15910 36422 15962 36474
rect 15974 36422 16026 36474
rect 16038 36422 16090 36474
rect 16102 36422 16154 36474
rect 25776 36422 25828 36474
rect 25840 36422 25892 36474
rect 25904 36422 25956 36474
rect 25968 36422 26020 36474
rect 26032 36422 26084 36474
rect 5172 36363 5224 36372
rect 5172 36329 5181 36363
rect 5181 36329 5215 36363
rect 5215 36329 5224 36363
rect 5172 36320 5224 36329
rect 7196 36363 7248 36372
rect 7196 36329 7205 36363
rect 7205 36329 7239 36363
rect 7239 36329 7248 36363
rect 7196 36320 7248 36329
rect 9772 36363 9824 36372
rect 9772 36329 9781 36363
rect 9781 36329 9815 36363
rect 9815 36329 9824 36363
rect 9772 36320 9824 36329
rect 10416 36320 10468 36372
rect 1676 36159 1728 36168
rect 1676 36125 1685 36159
rect 1685 36125 1719 36159
rect 1719 36125 1728 36159
rect 1676 36116 1728 36125
rect 9680 36252 9732 36304
rect 4252 36116 4304 36168
rect 5540 36184 5592 36236
rect 6460 36184 6512 36236
rect 6644 36227 6696 36236
rect 6644 36193 6653 36227
rect 6653 36193 6687 36227
rect 6687 36193 6696 36227
rect 6644 36184 6696 36193
rect 6736 36184 6788 36236
rect 10048 36184 10100 36236
rect 8024 36159 8076 36168
rect 3516 36048 3568 36100
rect 5448 36048 5500 36100
rect 8024 36125 8033 36159
rect 8033 36125 8067 36159
rect 8067 36125 8076 36159
rect 8024 36116 8076 36125
rect 9128 36159 9180 36168
rect 9128 36125 9137 36159
rect 9137 36125 9171 36159
rect 9171 36125 9180 36159
rect 9128 36116 9180 36125
rect 9312 36116 9364 36168
rect 10324 36159 10376 36168
rect 10324 36125 10333 36159
rect 10333 36125 10367 36159
rect 10367 36125 10376 36159
rect 10324 36116 10376 36125
rect 10600 36320 10652 36372
rect 10692 36320 10744 36372
rect 11244 36320 11296 36372
rect 11336 36320 11388 36372
rect 11520 36295 11572 36304
rect 11520 36261 11529 36295
rect 11529 36261 11563 36295
rect 11563 36261 11572 36295
rect 11520 36252 11572 36261
rect 14004 36320 14056 36372
rect 15200 36252 15252 36304
rect 17040 36320 17092 36372
rect 18604 36363 18656 36372
rect 18604 36329 18613 36363
rect 18613 36329 18647 36363
rect 18647 36329 18656 36363
rect 18604 36320 18656 36329
rect 20628 36320 20680 36372
rect 15108 36227 15160 36236
rect 15108 36193 15117 36227
rect 15117 36193 15151 36227
rect 15151 36193 15160 36227
rect 15108 36184 15160 36193
rect 11428 36116 11480 36168
rect 11704 36159 11756 36168
rect 11704 36125 11713 36159
rect 11713 36125 11747 36159
rect 11747 36125 11756 36159
rect 11704 36116 11756 36125
rect 14188 36116 14240 36168
rect 14280 36159 14332 36168
rect 14280 36125 14289 36159
rect 14289 36125 14323 36159
rect 14323 36125 14332 36159
rect 14280 36116 14332 36125
rect 15016 36116 15068 36168
rect 19616 36252 19668 36304
rect 16304 36184 16356 36236
rect 16120 36159 16172 36168
rect 16120 36125 16129 36159
rect 16129 36125 16163 36159
rect 16163 36125 16172 36159
rect 16120 36116 16172 36125
rect 1492 36023 1544 36032
rect 1492 35989 1501 36023
rect 1501 35989 1535 36023
rect 1535 35989 1544 36023
rect 1492 35980 1544 35989
rect 2228 35980 2280 36032
rect 2964 36023 3016 36032
rect 2964 35989 2973 36023
rect 2973 35989 3007 36023
rect 3007 35989 3016 36023
rect 2964 35980 3016 35989
rect 5080 35980 5132 36032
rect 7472 35980 7524 36032
rect 8392 35980 8444 36032
rect 8944 36023 8996 36032
rect 8944 35989 8953 36023
rect 8953 35989 8987 36023
rect 8987 35989 8996 36023
rect 8944 35980 8996 35989
rect 9036 35980 9088 36032
rect 11336 35980 11388 36032
rect 13268 35980 13320 36032
rect 20812 36184 20864 36236
rect 21364 36227 21416 36236
rect 21364 36193 21373 36227
rect 21373 36193 21407 36227
rect 21407 36193 21416 36227
rect 21364 36184 21416 36193
rect 18236 36116 18288 36168
rect 18604 36159 18656 36168
rect 18052 36048 18104 36100
rect 18604 36125 18613 36159
rect 18613 36125 18647 36159
rect 18647 36125 18656 36159
rect 18604 36116 18656 36125
rect 19892 36116 19944 36168
rect 20076 36159 20128 36168
rect 20076 36125 20085 36159
rect 20085 36125 20119 36159
rect 20119 36125 20128 36159
rect 20076 36116 20128 36125
rect 20352 36159 20404 36168
rect 20352 36125 20361 36159
rect 20361 36125 20395 36159
rect 20395 36125 20404 36159
rect 20352 36116 20404 36125
rect 21548 36116 21600 36168
rect 17224 35980 17276 36032
rect 19984 35980 20036 36032
rect 10880 35878 10932 35930
rect 10944 35878 10996 35930
rect 11008 35878 11060 35930
rect 11072 35878 11124 35930
rect 11136 35878 11188 35930
rect 20811 35878 20863 35930
rect 20875 35878 20927 35930
rect 20939 35878 20991 35930
rect 21003 35878 21055 35930
rect 21067 35878 21119 35930
rect 8024 35776 8076 35828
rect 9128 35776 9180 35828
rect 11704 35776 11756 35828
rect 18236 35819 18288 35828
rect 18236 35785 18245 35819
rect 18245 35785 18279 35819
rect 18279 35785 18288 35819
rect 18236 35776 18288 35785
rect 18604 35776 18656 35828
rect 19156 35819 19208 35828
rect 19156 35785 19165 35819
rect 19165 35785 19199 35819
rect 19199 35785 19208 35819
rect 19156 35776 19208 35785
rect 20444 35776 20496 35828
rect 1860 35683 1912 35692
rect 1860 35649 1869 35683
rect 1869 35649 1903 35683
rect 1903 35649 1912 35683
rect 1860 35640 1912 35649
rect 2412 35640 2464 35692
rect 2964 35640 3016 35692
rect 3424 35683 3476 35692
rect 3424 35649 3458 35683
rect 3458 35649 3476 35683
rect 3424 35640 3476 35649
rect 4436 35640 4488 35692
rect 9680 35708 9732 35760
rect 6276 35640 6328 35692
rect 6736 35640 6788 35692
rect 7564 35640 7616 35692
rect 10416 35708 10468 35760
rect 20536 35708 20588 35760
rect 10048 35640 10100 35692
rect 10784 35683 10836 35692
rect 10784 35649 10793 35683
rect 10793 35649 10827 35683
rect 10827 35649 10836 35683
rect 10784 35640 10836 35649
rect 11520 35683 11572 35692
rect 11520 35649 11529 35683
rect 11529 35649 11563 35683
rect 11563 35649 11572 35683
rect 11520 35640 11572 35649
rect 16396 35640 16448 35692
rect 8760 35572 8812 35624
rect 10232 35572 10284 35624
rect 10324 35572 10376 35624
rect 10692 35504 10744 35556
rect 14464 35572 14516 35624
rect 16764 35615 16816 35624
rect 16764 35581 16773 35615
rect 16773 35581 16807 35615
rect 16807 35581 16816 35615
rect 16764 35572 16816 35581
rect 16856 35572 16908 35624
rect 17132 35504 17184 35556
rect 17960 35640 18012 35692
rect 18972 35640 19024 35692
rect 19800 35640 19852 35692
rect 20168 35640 20220 35692
rect 20352 35640 20404 35692
rect 21548 35640 21600 35692
rect 19524 35572 19576 35624
rect 2228 35479 2280 35488
rect 2228 35445 2237 35479
rect 2237 35445 2271 35479
rect 2271 35445 2280 35479
rect 2228 35436 2280 35445
rect 3792 35436 3844 35488
rect 4896 35436 4948 35488
rect 5540 35436 5592 35488
rect 9220 35479 9272 35488
rect 9220 35445 9229 35479
rect 9229 35445 9263 35479
rect 9263 35445 9272 35479
rect 9220 35436 9272 35445
rect 10600 35479 10652 35488
rect 10600 35445 10609 35479
rect 10609 35445 10643 35479
rect 10643 35445 10652 35479
rect 10600 35436 10652 35445
rect 17316 35436 17368 35488
rect 17408 35479 17460 35488
rect 17408 35445 17417 35479
rect 17417 35445 17451 35479
rect 17451 35445 17460 35479
rect 17408 35436 17460 35445
rect 19432 35436 19484 35488
rect 20628 35436 20680 35488
rect 5915 35334 5967 35386
rect 5979 35334 6031 35386
rect 6043 35334 6095 35386
rect 6107 35334 6159 35386
rect 6171 35334 6223 35386
rect 15846 35334 15898 35386
rect 15910 35334 15962 35386
rect 15974 35334 16026 35386
rect 16038 35334 16090 35386
rect 16102 35334 16154 35386
rect 25776 35334 25828 35386
rect 25840 35334 25892 35386
rect 25904 35334 25956 35386
rect 25968 35334 26020 35386
rect 26032 35334 26084 35386
rect 2228 35275 2280 35284
rect 2228 35241 2237 35275
rect 2237 35241 2271 35275
rect 2271 35241 2280 35275
rect 2228 35232 2280 35241
rect 4436 35275 4488 35284
rect 4436 35241 4445 35275
rect 4445 35241 4479 35275
rect 4479 35241 4488 35275
rect 4436 35232 4488 35241
rect 1860 35207 1912 35216
rect 1860 35173 1869 35207
rect 1869 35173 1903 35207
rect 1903 35173 1912 35207
rect 1860 35164 1912 35173
rect 8668 35232 8720 35284
rect 10048 35232 10100 35284
rect 10784 35275 10836 35284
rect 10784 35241 10793 35275
rect 10793 35241 10827 35275
rect 10827 35241 10836 35275
rect 10784 35232 10836 35241
rect 8852 35164 8904 35216
rect 4896 35139 4948 35148
rect 4252 35071 4304 35080
rect 4252 35037 4261 35071
rect 4261 35037 4295 35071
rect 4295 35037 4304 35071
rect 4252 35028 4304 35037
rect 4896 35105 4905 35139
rect 4905 35105 4939 35139
rect 4939 35105 4948 35139
rect 4896 35096 4948 35105
rect 8392 35139 8444 35148
rect 8392 35105 8401 35139
rect 8401 35105 8435 35139
rect 8435 35105 8444 35139
rect 8392 35096 8444 35105
rect 8944 35139 8996 35148
rect 8944 35105 8953 35139
rect 8953 35105 8987 35139
rect 8987 35105 8996 35139
rect 8944 35096 8996 35105
rect 12440 35232 12492 35284
rect 13084 35275 13136 35284
rect 13084 35241 13093 35275
rect 13093 35241 13127 35275
rect 13127 35241 13136 35275
rect 13084 35232 13136 35241
rect 15568 35232 15620 35284
rect 16396 35275 16448 35284
rect 16396 35241 16405 35275
rect 16405 35241 16439 35275
rect 16439 35241 16448 35275
rect 16396 35232 16448 35241
rect 20352 35232 20404 35284
rect 20168 35164 20220 35216
rect 13728 35096 13780 35148
rect 15292 35096 15344 35148
rect 17316 35139 17368 35148
rect 17316 35105 17325 35139
rect 17325 35105 17359 35139
rect 17359 35105 17368 35139
rect 17316 35096 17368 35105
rect 20444 35096 20496 35148
rect 20628 35096 20680 35148
rect 6368 35028 6420 35080
rect 9220 35071 9272 35080
rect 9220 35037 9254 35071
rect 9254 35037 9272 35071
rect 9220 35028 9272 35037
rect 9956 35028 10008 35080
rect 14372 35028 14424 35080
rect 14648 35028 14700 35080
rect 15476 35071 15528 35080
rect 15476 35037 15485 35071
rect 15485 35037 15519 35071
rect 15519 35037 15528 35071
rect 15752 35071 15804 35080
rect 15476 35028 15528 35037
rect 15752 35037 15761 35071
rect 15761 35037 15795 35071
rect 15795 35037 15804 35071
rect 15752 35028 15804 35037
rect 20168 35028 20220 35080
rect 3792 34960 3844 35012
rect 4712 34960 4764 35012
rect 7656 34960 7708 35012
rect 12072 34960 12124 35012
rect 2964 34935 3016 34944
rect 2964 34901 2973 34935
rect 2973 34901 3007 34935
rect 3007 34901 3016 34935
rect 2964 34892 3016 34901
rect 4896 34892 4948 34944
rect 7012 34935 7064 34944
rect 7012 34901 7021 34935
rect 7021 34901 7055 34935
rect 7055 34901 7064 34935
rect 7012 34892 7064 34901
rect 9680 34892 9732 34944
rect 10508 34892 10560 34944
rect 18236 34960 18288 35012
rect 15476 34892 15528 34944
rect 19708 34935 19760 34944
rect 19708 34901 19717 34935
rect 19717 34901 19751 34935
rect 19751 34901 19760 34935
rect 19708 34892 19760 34901
rect 20076 34935 20128 34944
rect 20076 34901 20085 34935
rect 20085 34901 20119 34935
rect 20119 34901 20128 34935
rect 20076 34892 20128 34901
rect 10880 34790 10932 34842
rect 10944 34790 10996 34842
rect 11008 34790 11060 34842
rect 11072 34790 11124 34842
rect 11136 34790 11188 34842
rect 20811 34790 20863 34842
rect 20875 34790 20927 34842
rect 20939 34790 20991 34842
rect 21003 34790 21055 34842
rect 21067 34790 21119 34842
rect 1768 34688 1820 34740
rect 3424 34688 3476 34740
rect 4712 34731 4764 34740
rect 4712 34697 4721 34731
rect 4721 34697 4755 34731
rect 4755 34697 4764 34731
rect 4712 34688 4764 34697
rect 7656 34688 7708 34740
rect 10324 34688 10376 34740
rect 16856 34688 16908 34740
rect 17040 34688 17092 34740
rect 17224 34688 17276 34740
rect 17408 34731 17460 34740
rect 17408 34697 17417 34731
rect 17417 34697 17451 34731
rect 17451 34697 17460 34731
rect 18236 34731 18288 34740
rect 17408 34688 17460 34697
rect 18236 34697 18245 34731
rect 18245 34697 18279 34731
rect 18279 34697 18288 34731
rect 18236 34688 18288 34697
rect 6920 34620 6972 34672
rect 2412 34595 2464 34604
rect 2412 34561 2421 34595
rect 2421 34561 2455 34595
rect 2455 34561 2464 34595
rect 2412 34552 2464 34561
rect 2872 34595 2924 34604
rect 2872 34561 2881 34595
rect 2881 34561 2915 34595
rect 2915 34561 2924 34595
rect 2872 34552 2924 34561
rect 3792 34552 3844 34604
rect 4068 34595 4120 34604
rect 4068 34561 4077 34595
rect 4077 34561 4111 34595
rect 4111 34561 4120 34595
rect 4068 34552 4120 34561
rect 4344 34552 4396 34604
rect 4896 34595 4948 34604
rect 4896 34561 4905 34595
rect 4905 34561 4939 34595
rect 4939 34561 4948 34595
rect 4896 34552 4948 34561
rect 5080 34595 5132 34604
rect 5080 34561 5089 34595
rect 5089 34561 5123 34595
rect 5123 34561 5132 34595
rect 5080 34552 5132 34561
rect 5264 34595 5316 34604
rect 5264 34561 5273 34595
rect 5273 34561 5307 34595
rect 5307 34561 5316 34595
rect 5264 34552 5316 34561
rect 5724 34552 5776 34604
rect 7012 34552 7064 34604
rect 8208 34552 8260 34604
rect 8668 34552 8720 34604
rect 9772 34620 9824 34672
rect 10232 34595 10284 34604
rect 10232 34561 10241 34595
rect 10241 34561 10275 34595
rect 10275 34561 10284 34595
rect 10232 34552 10284 34561
rect 10416 34595 10468 34604
rect 10416 34561 10425 34595
rect 10425 34561 10459 34595
rect 10459 34561 10468 34595
rect 10416 34552 10468 34561
rect 10692 34552 10744 34604
rect 11244 34552 11296 34604
rect 11520 34552 11572 34604
rect 12440 34620 12492 34672
rect 13728 34620 13780 34672
rect 14096 34552 14148 34604
rect 15292 34595 15344 34604
rect 15292 34561 15326 34595
rect 15326 34561 15344 34595
rect 15292 34552 15344 34561
rect 18052 34552 18104 34604
rect 19156 34688 19208 34740
rect 19524 34620 19576 34672
rect 19708 34552 19760 34604
rect 19800 34552 19852 34604
rect 19984 34552 20036 34604
rect 30104 34595 30156 34604
rect 30104 34561 30113 34595
rect 30113 34561 30147 34595
rect 30147 34561 30156 34595
rect 30104 34552 30156 34561
rect 7288 34484 7340 34536
rect 4068 34416 4120 34468
rect 8024 34527 8076 34536
rect 8024 34493 8033 34527
rect 8033 34493 8067 34527
rect 8067 34493 8076 34527
rect 8944 34527 8996 34536
rect 8024 34484 8076 34493
rect 8944 34493 8953 34527
rect 8953 34493 8987 34527
rect 8987 34493 8996 34527
rect 8944 34484 8996 34493
rect 9680 34484 9732 34536
rect 14648 34484 14700 34536
rect 15660 34484 15712 34536
rect 17592 34527 17644 34536
rect 17592 34493 17601 34527
rect 17601 34493 17635 34527
rect 17635 34493 17644 34527
rect 17592 34484 17644 34493
rect 19432 34527 19484 34536
rect 19432 34493 19441 34527
rect 19441 34493 19475 34527
rect 19475 34493 19484 34527
rect 19432 34484 19484 34493
rect 20260 34484 20312 34536
rect 29828 34527 29880 34536
rect 29828 34493 29837 34527
rect 29837 34493 29871 34527
rect 29871 34493 29880 34527
rect 29828 34484 29880 34493
rect 2228 34348 2280 34400
rect 3056 34391 3108 34400
rect 3056 34357 3065 34391
rect 3065 34357 3099 34391
rect 3099 34357 3108 34391
rect 3056 34348 3108 34357
rect 3976 34348 4028 34400
rect 5080 34348 5132 34400
rect 6460 34391 6512 34400
rect 6460 34357 6469 34391
rect 6469 34357 6503 34391
rect 6503 34357 6512 34391
rect 6460 34348 6512 34357
rect 7380 34348 7432 34400
rect 10876 34348 10928 34400
rect 14464 34348 14516 34400
rect 15016 34416 15068 34468
rect 19340 34416 19392 34468
rect 19984 34416 20036 34468
rect 20444 34348 20496 34400
rect 5915 34246 5967 34298
rect 5979 34246 6031 34298
rect 6043 34246 6095 34298
rect 6107 34246 6159 34298
rect 6171 34246 6223 34298
rect 15846 34246 15898 34298
rect 15910 34246 15962 34298
rect 15974 34246 16026 34298
rect 16038 34246 16090 34298
rect 16102 34246 16154 34298
rect 25776 34246 25828 34298
rect 25840 34246 25892 34298
rect 25904 34246 25956 34298
rect 25968 34246 26020 34298
rect 26032 34246 26084 34298
rect 2228 34187 2280 34196
rect 2228 34153 2237 34187
rect 2237 34153 2271 34187
rect 2271 34153 2280 34187
rect 2228 34144 2280 34153
rect 6276 34144 6328 34196
rect 7564 34187 7616 34196
rect 7564 34153 7573 34187
rect 7573 34153 7607 34187
rect 7607 34153 7616 34187
rect 7564 34144 7616 34153
rect 7656 34144 7708 34196
rect 20720 34144 20772 34196
rect 2412 34076 2464 34128
rect 4804 34076 4856 34128
rect 5356 34076 5408 34128
rect 9680 34076 9732 34128
rect 10140 34076 10192 34128
rect 12532 34076 12584 34128
rect 14096 34119 14148 34128
rect 3056 34008 3108 34060
rect 3884 33940 3936 33992
rect 8300 34008 8352 34060
rect 9772 34051 9824 34060
rect 9772 34017 9781 34051
rect 9781 34017 9815 34051
rect 9815 34017 9824 34051
rect 9772 34008 9824 34017
rect 10600 34051 10652 34060
rect 10600 34017 10609 34051
rect 10609 34017 10643 34051
rect 10643 34017 10652 34051
rect 10600 34008 10652 34017
rect 2780 33804 2832 33856
rect 2964 33847 3016 33856
rect 2964 33813 2973 33847
rect 2973 33813 3007 33847
rect 3007 33813 3016 33847
rect 2964 33804 3016 33813
rect 3608 33872 3660 33924
rect 7656 33940 7708 33992
rect 8208 33983 8260 33992
rect 8208 33949 8217 33983
rect 8217 33949 8251 33983
rect 8251 33949 8260 33983
rect 8208 33940 8260 33949
rect 9680 33940 9732 33992
rect 8392 33872 8444 33924
rect 10692 33940 10744 33992
rect 10876 33983 10928 33992
rect 10876 33949 10910 33983
rect 10910 33949 10928 33983
rect 10876 33940 10928 33949
rect 13452 34008 13504 34060
rect 14096 34085 14105 34119
rect 14105 34085 14139 34119
rect 14139 34085 14148 34119
rect 14096 34076 14148 34085
rect 14372 34076 14424 34128
rect 15016 34076 15068 34128
rect 12532 33983 12584 33992
rect 12532 33949 12542 33983
rect 12542 33949 12576 33983
rect 12576 33949 12584 33983
rect 12532 33940 12584 33949
rect 12992 33940 13044 33992
rect 19432 34076 19484 34128
rect 20444 34119 20496 34128
rect 20444 34085 20453 34119
rect 20453 34085 20487 34119
rect 20487 34085 20496 34119
rect 20444 34076 20496 34085
rect 10416 33872 10468 33924
rect 12716 33915 12768 33924
rect 12716 33881 12725 33915
rect 12725 33881 12759 33915
rect 12759 33881 12768 33915
rect 12716 33872 12768 33881
rect 12808 33915 12860 33924
rect 12808 33881 12817 33915
rect 12817 33881 12851 33915
rect 12851 33881 12860 33915
rect 14372 33915 14424 33924
rect 12808 33872 12860 33881
rect 14372 33881 14381 33915
rect 14381 33881 14415 33915
rect 14415 33881 14424 33915
rect 14372 33872 14424 33881
rect 14464 33915 14516 33924
rect 14464 33881 14473 33915
rect 14473 33881 14507 33915
rect 14507 33881 14516 33915
rect 14464 33872 14516 33881
rect 3792 33804 3844 33856
rect 6552 33804 6604 33856
rect 8484 33804 8536 33856
rect 8944 33804 8996 33856
rect 9404 33847 9456 33856
rect 9404 33813 9413 33847
rect 9413 33813 9447 33847
rect 9447 33813 9456 33847
rect 9404 33804 9456 33813
rect 11244 33804 11296 33856
rect 13176 33804 13228 33856
rect 13452 33804 13504 33856
rect 17408 33940 17460 33992
rect 18512 33983 18564 33992
rect 18512 33949 18521 33983
rect 18521 33949 18555 33983
rect 18555 33949 18564 33983
rect 18512 33940 18564 33949
rect 19892 33940 19944 33992
rect 20628 33983 20680 33992
rect 20628 33949 20637 33983
rect 20637 33949 20671 33983
rect 20671 33949 20680 33983
rect 20628 33940 20680 33949
rect 18880 33872 18932 33924
rect 21640 33940 21692 33992
rect 16948 33804 17000 33856
rect 19340 33804 19392 33856
rect 21180 33872 21232 33924
rect 20720 33847 20772 33856
rect 20720 33813 20729 33847
rect 20729 33813 20763 33847
rect 20763 33813 20772 33847
rect 20720 33804 20772 33813
rect 21272 33804 21324 33856
rect 22652 33804 22704 33856
rect 10880 33702 10932 33754
rect 10944 33702 10996 33754
rect 11008 33702 11060 33754
rect 11072 33702 11124 33754
rect 11136 33702 11188 33754
rect 20811 33702 20863 33754
rect 20875 33702 20927 33754
rect 20939 33702 20991 33754
rect 21003 33702 21055 33754
rect 21067 33702 21119 33754
rect 2872 33600 2924 33652
rect 3608 33643 3660 33652
rect 3608 33609 3617 33643
rect 3617 33609 3651 33643
rect 3651 33609 3660 33643
rect 3608 33600 3660 33609
rect 5632 33600 5684 33652
rect 7656 33600 7708 33652
rect 7840 33600 7892 33652
rect 8760 33600 8812 33652
rect 2044 33464 2096 33516
rect 3148 33507 3200 33516
rect 3148 33473 3157 33507
rect 3157 33473 3191 33507
rect 3191 33473 3200 33507
rect 3148 33464 3200 33473
rect 3792 33507 3844 33516
rect 3792 33473 3801 33507
rect 3801 33473 3835 33507
rect 3835 33473 3844 33507
rect 3792 33464 3844 33473
rect 4068 33507 4120 33516
rect 4068 33473 4077 33507
rect 4077 33473 4111 33507
rect 4111 33473 4120 33507
rect 4068 33464 4120 33473
rect 4804 33532 4856 33584
rect 7564 33532 7616 33584
rect 4344 33507 4396 33516
rect 4344 33473 4353 33507
rect 4353 33473 4387 33507
rect 4387 33473 4396 33507
rect 4344 33464 4396 33473
rect 6276 33464 6328 33516
rect 6552 33507 6604 33516
rect 6552 33473 6561 33507
rect 6561 33473 6595 33507
rect 6595 33473 6604 33507
rect 6552 33464 6604 33473
rect 7748 33507 7800 33516
rect 7748 33473 7757 33507
rect 7757 33473 7791 33507
rect 7791 33473 7800 33507
rect 7748 33464 7800 33473
rect 7840 33464 7892 33516
rect 3976 33439 4028 33448
rect 3976 33405 3985 33439
rect 3985 33405 4019 33439
rect 4019 33405 4028 33439
rect 3976 33396 4028 33405
rect 8668 33464 8720 33516
rect 1492 33303 1544 33312
rect 1492 33269 1501 33303
rect 1501 33269 1535 33303
rect 1535 33269 1544 33303
rect 1492 33260 1544 33269
rect 2136 33303 2188 33312
rect 2136 33269 2145 33303
rect 2145 33269 2179 33303
rect 2179 33269 2188 33303
rect 2136 33260 2188 33269
rect 3148 33328 3200 33380
rect 4252 33328 4304 33380
rect 8208 33396 8260 33448
rect 10692 33600 10744 33652
rect 12716 33600 12768 33652
rect 14924 33600 14976 33652
rect 9496 33532 9548 33584
rect 14372 33532 14424 33584
rect 15568 33532 15620 33584
rect 16396 33532 16448 33584
rect 17316 33575 17368 33584
rect 17316 33541 17325 33575
rect 17325 33541 17359 33575
rect 17359 33541 17368 33575
rect 17316 33532 17368 33541
rect 18328 33575 18380 33584
rect 18328 33541 18337 33575
rect 18337 33541 18371 33575
rect 18371 33541 18380 33575
rect 18328 33532 18380 33541
rect 19892 33600 19944 33652
rect 20720 33643 20772 33652
rect 20720 33609 20729 33643
rect 20729 33609 20763 33643
rect 20763 33609 20772 33643
rect 20720 33600 20772 33609
rect 8484 33328 8536 33380
rect 4160 33260 4212 33312
rect 7104 33260 7156 33312
rect 10416 33464 10468 33516
rect 10692 33464 10744 33516
rect 12348 33464 12400 33516
rect 12808 33464 12860 33516
rect 13176 33507 13228 33516
rect 13176 33473 13210 33507
rect 13210 33473 13228 33507
rect 13176 33464 13228 33473
rect 13452 33464 13504 33516
rect 15292 33507 15344 33516
rect 11520 33439 11572 33448
rect 11520 33405 11529 33439
rect 11529 33405 11563 33439
rect 11563 33405 11572 33439
rect 11520 33396 11572 33405
rect 12440 33396 12492 33448
rect 12900 33439 12952 33448
rect 12900 33405 12909 33439
rect 12909 33405 12943 33439
rect 12943 33405 12952 33439
rect 12900 33396 12952 33405
rect 15292 33473 15301 33507
rect 15301 33473 15335 33507
rect 15335 33473 15344 33507
rect 15292 33464 15344 33473
rect 15476 33507 15528 33516
rect 15476 33473 15490 33507
rect 15490 33473 15524 33507
rect 15524 33473 15528 33507
rect 15476 33464 15528 33473
rect 17960 33464 18012 33516
rect 19340 33464 19392 33516
rect 20168 33464 20220 33516
rect 20812 33575 20864 33584
rect 20812 33541 20839 33575
rect 20839 33541 20864 33575
rect 21272 33600 21324 33652
rect 20812 33532 20864 33541
rect 21180 33532 21232 33584
rect 21456 33464 21508 33516
rect 21824 33507 21876 33516
rect 21824 33473 21833 33507
rect 21833 33473 21867 33507
rect 21867 33473 21876 33507
rect 21824 33464 21876 33473
rect 22652 33507 22704 33516
rect 22652 33473 22661 33507
rect 22661 33473 22695 33507
rect 22695 33473 22704 33507
rect 22652 33464 22704 33473
rect 30104 33464 30156 33516
rect 9312 33260 9364 33312
rect 29828 33328 29880 33380
rect 15660 33303 15712 33312
rect 15660 33269 15669 33303
rect 15669 33269 15703 33303
rect 15703 33269 15712 33303
rect 15660 33260 15712 33269
rect 18696 33260 18748 33312
rect 19800 33303 19852 33312
rect 19800 33269 19809 33303
rect 19809 33269 19843 33303
rect 19843 33269 19852 33303
rect 19800 33260 19852 33269
rect 22376 33260 22428 33312
rect 30012 33303 30064 33312
rect 30012 33269 30021 33303
rect 30021 33269 30055 33303
rect 30055 33269 30064 33303
rect 30012 33260 30064 33269
rect 5915 33158 5967 33210
rect 5979 33158 6031 33210
rect 6043 33158 6095 33210
rect 6107 33158 6159 33210
rect 6171 33158 6223 33210
rect 15846 33158 15898 33210
rect 15910 33158 15962 33210
rect 15974 33158 16026 33210
rect 16038 33158 16090 33210
rect 16102 33158 16154 33210
rect 25776 33158 25828 33210
rect 25840 33158 25892 33210
rect 25904 33158 25956 33210
rect 25968 33158 26020 33210
rect 26032 33158 26084 33210
rect 2228 33099 2280 33108
rect 2228 33065 2237 33099
rect 2237 33065 2271 33099
rect 2271 33065 2280 33099
rect 2228 33056 2280 33065
rect 5724 33099 5776 33108
rect 5724 33065 5733 33099
rect 5733 33065 5767 33099
rect 5767 33065 5776 33099
rect 5724 33056 5776 33065
rect 7932 33056 7984 33108
rect 9220 33056 9272 33108
rect 9680 33056 9732 33108
rect 10324 33056 10376 33108
rect 12072 33099 12124 33108
rect 12072 33065 12081 33099
rect 12081 33065 12115 33099
rect 12115 33065 12124 33099
rect 12072 33056 12124 33065
rect 2136 32988 2188 33040
rect 10416 32988 10468 33040
rect 19064 33056 19116 33108
rect 19156 33056 19208 33108
rect 19800 33099 19852 33108
rect 19800 33065 19809 33099
rect 19809 33065 19843 33099
rect 19843 33065 19852 33099
rect 19800 33056 19852 33065
rect 20444 33056 20496 33108
rect 20536 33056 20588 33108
rect 16396 33031 16448 33040
rect 16396 32997 16405 33031
rect 16405 32997 16439 33031
rect 16439 32997 16448 33031
rect 16396 32988 16448 32997
rect 7932 32963 7984 32972
rect 7932 32929 7941 32963
rect 7941 32929 7975 32963
rect 7975 32929 7984 32963
rect 7932 32920 7984 32929
rect 8484 32920 8536 32972
rect 9312 32963 9364 32972
rect 9312 32929 9321 32963
rect 9321 32929 9355 32963
rect 9355 32929 9364 32963
rect 9312 32920 9364 32929
rect 10784 32920 10836 32972
rect 12992 32920 13044 32972
rect 15016 32963 15068 32972
rect 15016 32929 15025 32963
rect 15025 32929 15059 32963
rect 15059 32929 15068 32963
rect 15016 32920 15068 32929
rect 16948 32963 17000 32972
rect 16948 32929 16957 32963
rect 16957 32929 16991 32963
rect 16991 32929 17000 32963
rect 16948 32920 17000 32929
rect 19892 32920 19944 32972
rect 21824 33056 21876 33108
rect 3148 32852 3200 32904
rect 3332 32852 3384 32904
rect 7564 32852 7616 32904
rect 2412 32759 2464 32768
rect 2412 32725 2421 32759
rect 2421 32725 2455 32759
rect 2455 32725 2464 32759
rect 2412 32716 2464 32725
rect 3148 32716 3200 32768
rect 3884 32784 3936 32836
rect 5632 32784 5684 32836
rect 8116 32852 8168 32904
rect 9220 32852 9272 32904
rect 9404 32852 9456 32904
rect 11796 32895 11848 32904
rect 8668 32784 8720 32836
rect 11796 32861 11805 32895
rect 11805 32861 11839 32895
rect 11839 32861 11848 32895
rect 11796 32852 11848 32861
rect 11888 32895 11940 32904
rect 11888 32861 11897 32895
rect 11897 32861 11931 32895
rect 11931 32861 11940 32895
rect 11888 32852 11940 32861
rect 12072 32895 12124 32904
rect 12072 32861 12081 32895
rect 12081 32861 12115 32895
rect 12115 32861 12124 32895
rect 12072 32852 12124 32861
rect 15660 32852 15712 32904
rect 19432 32852 19484 32904
rect 19616 32895 19668 32904
rect 19616 32861 19625 32895
rect 19625 32861 19659 32895
rect 19659 32861 19668 32895
rect 19616 32852 19668 32861
rect 20168 32852 20220 32904
rect 12532 32784 12584 32836
rect 12992 32784 13044 32836
rect 17868 32784 17920 32836
rect 20628 32784 20680 32836
rect 21916 32784 21968 32836
rect 5172 32759 5224 32768
rect 5172 32725 5181 32759
rect 5181 32725 5215 32759
rect 5215 32725 5224 32759
rect 5172 32716 5224 32725
rect 6828 32759 6880 32768
rect 6828 32725 6837 32759
rect 6837 32725 6871 32759
rect 6871 32725 6880 32759
rect 6828 32716 6880 32725
rect 8760 32716 8812 32768
rect 18328 32759 18380 32768
rect 18328 32725 18337 32759
rect 18337 32725 18371 32759
rect 18371 32725 18380 32759
rect 18328 32716 18380 32725
rect 18420 32716 18472 32768
rect 20536 32716 20588 32768
rect 20720 32716 20772 32768
rect 21364 32716 21416 32768
rect 22192 32759 22244 32768
rect 22192 32725 22219 32759
rect 22219 32725 22244 32759
rect 22192 32716 22244 32725
rect 10880 32614 10932 32666
rect 10944 32614 10996 32666
rect 11008 32614 11060 32666
rect 11072 32614 11124 32666
rect 11136 32614 11188 32666
rect 20811 32614 20863 32666
rect 20875 32614 20927 32666
rect 20939 32614 20991 32666
rect 21003 32614 21055 32666
rect 21067 32614 21119 32666
rect 3332 32555 3384 32564
rect 3332 32521 3341 32555
rect 3341 32521 3375 32555
rect 3375 32521 3384 32555
rect 3332 32512 3384 32521
rect 3884 32512 3936 32564
rect 7748 32512 7800 32564
rect 8116 32512 8168 32564
rect 9220 32512 9272 32564
rect 15476 32555 15528 32564
rect 2780 32376 2832 32428
rect 3148 32419 3200 32428
rect 3148 32385 3157 32419
rect 3157 32385 3191 32419
rect 3191 32385 3200 32419
rect 3148 32376 3200 32385
rect 5172 32444 5224 32496
rect 7104 32487 7156 32496
rect 7104 32453 7138 32487
rect 7138 32453 7156 32487
rect 7104 32444 7156 32453
rect 4252 32419 4304 32428
rect 4252 32385 4261 32419
rect 4261 32385 4295 32419
rect 4295 32385 4304 32419
rect 4252 32376 4304 32385
rect 2964 32308 3016 32360
rect 4068 32308 4120 32360
rect 4436 32376 4488 32428
rect 5632 32376 5684 32428
rect 9956 32444 10008 32496
rect 8760 32376 8812 32428
rect 4528 32240 4580 32292
rect 6368 32308 6420 32360
rect 8668 32351 8720 32360
rect 8668 32317 8677 32351
rect 8677 32317 8711 32351
rect 8711 32317 8720 32351
rect 8668 32308 8720 32317
rect 6644 32240 6696 32292
rect 1492 32215 1544 32224
rect 1492 32181 1501 32215
rect 1501 32181 1535 32215
rect 1535 32181 1544 32215
rect 1492 32172 1544 32181
rect 2228 32215 2280 32224
rect 2228 32181 2237 32215
rect 2237 32181 2271 32215
rect 2271 32181 2280 32215
rect 2228 32172 2280 32181
rect 6736 32172 6788 32224
rect 10416 32240 10468 32292
rect 9772 32172 9824 32224
rect 15476 32521 15485 32555
rect 15485 32521 15519 32555
rect 15519 32521 15528 32555
rect 15476 32512 15528 32521
rect 17868 32555 17920 32564
rect 17868 32521 17877 32555
rect 17877 32521 17911 32555
rect 17911 32521 17920 32555
rect 17868 32512 17920 32521
rect 19248 32555 19300 32564
rect 19248 32521 19257 32555
rect 19257 32521 19291 32555
rect 19291 32521 19300 32555
rect 19248 32512 19300 32521
rect 19708 32512 19760 32564
rect 11520 32444 11572 32496
rect 12072 32444 12124 32496
rect 12532 32444 12584 32496
rect 13912 32444 13964 32496
rect 10876 32419 10928 32428
rect 10876 32385 10885 32419
rect 10885 32385 10919 32419
rect 10919 32385 10928 32419
rect 10876 32376 10928 32385
rect 12256 32376 12308 32428
rect 12900 32376 12952 32428
rect 15292 32376 15344 32428
rect 17132 32419 17184 32428
rect 17132 32385 17141 32419
rect 17141 32385 17175 32419
rect 17175 32385 17184 32419
rect 17132 32376 17184 32385
rect 17316 32419 17368 32428
rect 17316 32385 17325 32419
rect 17325 32385 17359 32419
rect 17359 32385 17368 32419
rect 17316 32376 17368 32385
rect 18328 32376 18380 32428
rect 18604 32444 18656 32496
rect 11336 32308 11388 32360
rect 17408 32351 17460 32360
rect 17408 32317 17417 32351
rect 17417 32317 17451 32351
rect 17451 32317 17460 32351
rect 17408 32308 17460 32317
rect 18420 32308 18472 32360
rect 17776 32240 17828 32292
rect 12164 32172 12216 32224
rect 14648 32172 14700 32224
rect 14740 32172 14792 32224
rect 18880 32419 18932 32428
rect 18880 32385 18889 32419
rect 18889 32385 18923 32419
rect 18923 32385 18932 32419
rect 18880 32376 18932 32385
rect 19800 32444 19852 32496
rect 20260 32512 20312 32564
rect 20628 32444 20680 32496
rect 19616 32376 19668 32428
rect 20444 32376 20496 32428
rect 21364 32444 21416 32496
rect 21640 32512 21692 32564
rect 22192 32487 22244 32496
rect 22192 32453 22201 32487
rect 22201 32453 22235 32487
rect 22235 32453 22244 32487
rect 22192 32444 22244 32453
rect 21272 32419 21324 32428
rect 21272 32385 21281 32419
rect 21281 32385 21315 32419
rect 21315 32385 21324 32419
rect 21272 32376 21324 32385
rect 19156 32308 19208 32360
rect 18696 32240 18748 32292
rect 20720 32308 20772 32360
rect 21180 32308 21232 32360
rect 20536 32240 20588 32292
rect 19892 32172 19944 32224
rect 20904 32172 20956 32224
rect 21916 32172 21968 32224
rect 5915 32070 5967 32122
rect 5979 32070 6031 32122
rect 6043 32070 6095 32122
rect 6107 32070 6159 32122
rect 6171 32070 6223 32122
rect 15846 32070 15898 32122
rect 15910 32070 15962 32122
rect 15974 32070 16026 32122
rect 16038 32070 16090 32122
rect 16102 32070 16154 32122
rect 25776 32070 25828 32122
rect 25840 32070 25892 32122
rect 25904 32070 25956 32122
rect 25968 32070 26020 32122
rect 26032 32070 26084 32122
rect 2320 32011 2372 32020
rect 2320 31977 2329 32011
rect 2329 31977 2363 32011
rect 2363 31977 2372 32011
rect 2320 31968 2372 31977
rect 2964 32011 3016 32020
rect 2964 31977 2973 32011
rect 2973 31977 3007 32011
rect 3007 31977 3016 32011
rect 2964 31968 3016 31977
rect 6368 32011 6420 32020
rect 6368 31977 6377 32011
rect 6377 31977 6411 32011
rect 6411 31977 6420 32011
rect 6368 31968 6420 31977
rect 8668 31968 8720 32020
rect 9680 32011 9732 32020
rect 9680 31977 9689 32011
rect 9689 31977 9723 32011
rect 9723 31977 9732 32011
rect 9680 31968 9732 31977
rect 10140 31968 10192 32020
rect 10876 31968 10928 32020
rect 18512 32011 18564 32020
rect 18512 31977 18521 32011
rect 18521 31977 18555 32011
rect 18555 31977 18564 32011
rect 18512 31968 18564 31977
rect 19064 31968 19116 32020
rect 2136 31900 2188 31952
rect 3792 31900 3844 31952
rect 4068 31943 4120 31952
rect 4068 31909 4077 31943
rect 4077 31909 4111 31943
rect 4111 31909 4120 31943
rect 4068 31900 4120 31909
rect 2964 31832 3016 31884
rect 5632 31875 5684 31884
rect 5632 31841 5641 31875
rect 5641 31841 5675 31875
rect 5675 31841 5684 31875
rect 5632 31832 5684 31841
rect 9864 31900 9916 31952
rect 11152 31900 11204 31952
rect 11244 31900 11296 31952
rect 12624 31943 12676 31952
rect 12624 31909 12633 31943
rect 12633 31909 12667 31943
rect 12667 31909 12676 31943
rect 12624 31900 12676 31909
rect 12900 31900 12952 31952
rect 17408 31900 17460 31952
rect 3148 31807 3200 31816
rect 3148 31773 3157 31807
rect 3157 31773 3191 31807
rect 3191 31773 3200 31807
rect 3148 31764 3200 31773
rect 4528 31764 4580 31816
rect 5172 31764 5224 31816
rect 6460 31764 6512 31816
rect 6828 31807 6880 31816
rect 4804 31696 4856 31748
rect 6828 31773 6837 31807
rect 6837 31773 6871 31807
rect 6871 31773 6880 31807
rect 6828 31764 6880 31773
rect 7564 31764 7616 31816
rect 9128 31832 9180 31884
rect 8852 31764 8904 31816
rect 10048 31764 10100 31816
rect 11336 31764 11388 31816
rect 18420 31875 18472 31884
rect 11888 31696 11940 31748
rect 18420 31841 18429 31875
rect 18429 31841 18463 31875
rect 18463 31841 18472 31875
rect 18420 31832 18472 31841
rect 19984 31832 20036 31884
rect 20720 31832 20772 31884
rect 20904 31875 20956 31884
rect 20904 31841 20913 31875
rect 20913 31841 20947 31875
rect 20947 31841 20956 31875
rect 20904 31832 20956 31841
rect 21272 31832 21324 31884
rect 15476 31764 15528 31816
rect 18696 31807 18748 31816
rect 18696 31773 18705 31807
rect 18705 31773 18739 31807
rect 18739 31773 18748 31807
rect 18696 31764 18748 31773
rect 20628 31807 20680 31816
rect 20628 31773 20637 31807
rect 20637 31773 20671 31807
rect 20671 31773 20680 31807
rect 20628 31764 20680 31773
rect 13820 31696 13872 31748
rect 20444 31696 20496 31748
rect 21916 31764 21968 31816
rect 29828 31807 29880 31816
rect 29828 31773 29837 31807
rect 29837 31773 29871 31807
rect 29871 31773 29880 31807
rect 29828 31764 29880 31773
rect 21088 31696 21140 31748
rect 4160 31628 4212 31680
rect 7104 31628 7156 31680
rect 9772 31628 9824 31680
rect 15384 31628 15436 31680
rect 30012 31671 30064 31680
rect 30012 31637 30021 31671
rect 30021 31637 30055 31671
rect 30055 31637 30064 31671
rect 30012 31628 30064 31637
rect 10880 31526 10932 31578
rect 10944 31526 10996 31578
rect 11008 31526 11060 31578
rect 11072 31526 11124 31578
rect 11136 31526 11188 31578
rect 20811 31526 20863 31578
rect 20875 31526 20927 31578
rect 20939 31526 20991 31578
rect 21003 31526 21055 31578
rect 21067 31526 21119 31578
rect 3148 31424 3200 31476
rect 8392 31424 8444 31476
rect 12532 31424 12584 31476
rect 12900 31424 12952 31476
rect 13452 31424 13504 31476
rect 13820 31424 13872 31476
rect 15292 31424 15344 31476
rect 17040 31424 17092 31476
rect 18328 31424 18380 31476
rect 21916 31467 21968 31476
rect 2136 31288 2188 31340
rect 3700 31356 3752 31408
rect 3792 31331 3844 31340
rect 3516 31152 3568 31204
rect 3792 31297 3801 31331
rect 3801 31297 3835 31331
rect 3835 31297 3844 31331
rect 3792 31288 3844 31297
rect 4252 31356 4304 31408
rect 4436 31288 4488 31340
rect 6552 31331 6604 31340
rect 6552 31297 6561 31331
rect 6561 31297 6595 31331
rect 6595 31297 6604 31331
rect 6552 31288 6604 31297
rect 6736 31331 6788 31340
rect 6736 31297 6745 31331
rect 6745 31297 6779 31331
rect 6779 31297 6788 31331
rect 6736 31288 6788 31297
rect 7840 31356 7892 31408
rect 7104 31331 7156 31340
rect 7104 31297 7113 31331
rect 7113 31297 7147 31331
rect 7147 31297 7156 31331
rect 7104 31288 7156 31297
rect 7288 31288 7340 31340
rect 8300 31288 8352 31340
rect 9036 31331 9088 31340
rect 6828 31263 6880 31272
rect 6828 31229 6837 31263
rect 6837 31229 6871 31263
rect 6871 31229 6880 31263
rect 6828 31220 6880 31229
rect 5080 31152 5132 31204
rect 6920 31152 6972 31204
rect 9036 31297 9045 31331
rect 9045 31297 9079 31331
rect 9079 31297 9088 31331
rect 9036 31288 9088 31297
rect 10324 31288 10376 31340
rect 10508 31288 10560 31340
rect 12716 31356 12768 31408
rect 10232 31220 10284 31272
rect 12440 31331 12492 31340
rect 12440 31297 12449 31331
rect 12449 31297 12483 31331
rect 12483 31297 12492 31331
rect 12900 31331 12952 31340
rect 12440 31288 12492 31297
rect 12900 31297 12909 31331
rect 12909 31297 12943 31331
rect 12943 31297 12952 31331
rect 12900 31288 12952 31297
rect 12992 31331 13044 31340
rect 12992 31297 13002 31331
rect 13002 31297 13036 31331
rect 13036 31297 13044 31331
rect 12992 31288 13044 31297
rect 13084 31220 13136 31272
rect 13268 31331 13320 31340
rect 13268 31297 13277 31331
rect 13277 31297 13311 31331
rect 13311 31297 13320 31331
rect 13268 31288 13320 31297
rect 15568 31288 15620 31340
rect 15016 31220 15068 31272
rect 15384 31220 15436 31272
rect 17224 31288 17276 31340
rect 18420 31356 18472 31408
rect 21916 31433 21925 31467
rect 21925 31433 21959 31467
rect 21959 31433 21968 31467
rect 21916 31424 21968 31433
rect 19984 31356 20036 31408
rect 20168 31288 20220 31340
rect 21640 31288 21692 31340
rect 17132 31263 17184 31272
rect 2320 31127 2372 31136
rect 2320 31093 2329 31127
rect 2329 31093 2363 31127
rect 2363 31093 2372 31127
rect 2320 31084 2372 31093
rect 3424 31127 3476 31136
rect 3424 31093 3433 31127
rect 3433 31093 3467 31127
rect 3467 31093 3476 31127
rect 3424 31084 3476 31093
rect 4252 31084 4304 31136
rect 6368 31127 6420 31136
rect 6368 31093 6377 31127
rect 6377 31093 6411 31127
rect 6411 31093 6420 31127
rect 6368 31084 6420 31093
rect 7564 31127 7616 31136
rect 7564 31093 7573 31127
rect 7573 31093 7607 31127
rect 7607 31093 7616 31127
rect 7564 31084 7616 31093
rect 8852 31127 8904 31136
rect 8852 31093 8861 31127
rect 8861 31093 8895 31127
rect 8895 31093 8904 31127
rect 8852 31084 8904 31093
rect 9680 31084 9732 31136
rect 10048 31084 10100 31136
rect 14740 31152 14792 31204
rect 17132 31229 17141 31263
rect 17141 31229 17175 31263
rect 17175 31229 17184 31263
rect 17132 31220 17184 31229
rect 19708 31152 19760 31204
rect 20444 31152 20496 31204
rect 10692 31084 10744 31136
rect 15384 31084 15436 31136
rect 17868 31084 17920 31136
rect 20536 31084 20588 31136
rect 5915 30982 5967 31034
rect 5979 30982 6031 31034
rect 6043 30982 6095 31034
rect 6107 30982 6159 31034
rect 6171 30982 6223 31034
rect 15846 30982 15898 31034
rect 15910 30982 15962 31034
rect 15974 30982 16026 31034
rect 16038 30982 16090 31034
rect 16102 30982 16154 31034
rect 25776 30982 25828 31034
rect 25840 30982 25892 31034
rect 25904 30982 25956 31034
rect 25968 30982 26020 31034
rect 26032 30982 26084 31034
rect 2320 30923 2372 30932
rect 2320 30889 2329 30923
rect 2329 30889 2363 30923
rect 2363 30889 2372 30923
rect 2320 30880 2372 30889
rect 2688 30880 2740 30932
rect 8852 30880 8904 30932
rect 11888 30923 11940 30932
rect 11888 30889 11897 30923
rect 11897 30889 11931 30923
rect 11931 30889 11940 30923
rect 11888 30880 11940 30889
rect 29828 30880 29880 30932
rect 2136 30812 2188 30864
rect 3516 30744 3568 30796
rect 3056 30676 3108 30728
rect 4528 30676 4580 30728
rect 5080 30744 5132 30796
rect 10324 30812 10376 30864
rect 13268 30812 13320 30864
rect 20720 30812 20772 30864
rect 10600 30744 10652 30796
rect 4712 30676 4764 30728
rect 4804 30719 4856 30728
rect 4804 30685 4813 30719
rect 4813 30685 4847 30719
rect 4847 30685 4856 30719
rect 4804 30676 4856 30685
rect 5172 30719 5224 30728
rect 5172 30685 5181 30719
rect 5181 30685 5215 30719
rect 5215 30685 5224 30719
rect 5172 30676 5224 30685
rect 6368 30676 6420 30728
rect 7932 30676 7984 30728
rect 8116 30676 8168 30728
rect 9220 30676 9272 30728
rect 10048 30719 10100 30728
rect 10048 30685 10057 30719
rect 10057 30685 10091 30719
rect 10091 30685 10100 30719
rect 10048 30676 10100 30685
rect 10692 30719 10744 30728
rect 10692 30685 10701 30719
rect 10701 30685 10735 30719
rect 10735 30685 10744 30719
rect 10692 30676 10744 30685
rect 11888 30744 11940 30796
rect 12808 30744 12860 30796
rect 17132 30744 17184 30796
rect 17500 30744 17552 30796
rect 17960 30787 18012 30796
rect 17960 30753 17969 30787
rect 17969 30753 18003 30787
rect 18003 30753 18012 30787
rect 17960 30744 18012 30753
rect 11428 30719 11480 30728
rect 11428 30685 11437 30719
rect 11437 30685 11471 30719
rect 11471 30685 11480 30719
rect 11428 30676 11480 30685
rect 12624 30676 12676 30728
rect 12992 30676 13044 30728
rect 14188 30676 14240 30728
rect 17040 30676 17092 30728
rect 17868 30719 17920 30728
rect 17868 30685 17877 30719
rect 17877 30685 17911 30719
rect 17911 30685 17920 30719
rect 17868 30676 17920 30685
rect 19248 30744 19300 30796
rect 20260 30787 20312 30796
rect 20260 30753 20269 30787
rect 20269 30753 20303 30787
rect 20303 30753 20312 30787
rect 20260 30744 20312 30753
rect 20536 30787 20588 30796
rect 20536 30753 20545 30787
rect 20545 30753 20579 30787
rect 20579 30753 20588 30787
rect 20536 30744 20588 30753
rect 2504 30583 2556 30592
rect 2504 30549 2513 30583
rect 2513 30549 2547 30583
rect 2547 30549 2556 30583
rect 2504 30540 2556 30549
rect 3148 30583 3200 30592
rect 3148 30549 3157 30583
rect 3157 30549 3191 30583
rect 3191 30549 3200 30583
rect 3148 30540 3200 30549
rect 4160 30540 4212 30592
rect 14740 30608 14792 30660
rect 29552 30676 29604 30728
rect 30104 30719 30156 30728
rect 30104 30685 30113 30719
rect 30113 30685 30147 30719
rect 30147 30685 30156 30719
rect 30104 30676 30156 30685
rect 21180 30651 21232 30660
rect 6552 30540 6604 30592
rect 7932 30583 7984 30592
rect 7932 30549 7941 30583
rect 7941 30549 7975 30583
rect 7975 30549 7984 30583
rect 7932 30540 7984 30549
rect 8576 30540 8628 30592
rect 9220 30540 9272 30592
rect 10508 30583 10560 30592
rect 10508 30549 10517 30583
rect 10517 30549 10551 30583
rect 10551 30549 10560 30583
rect 10508 30540 10560 30549
rect 11520 30540 11572 30592
rect 15660 30583 15712 30592
rect 15660 30549 15669 30583
rect 15669 30549 15703 30583
rect 15703 30549 15712 30583
rect 15660 30540 15712 30549
rect 17224 30540 17276 30592
rect 21180 30617 21189 30651
rect 21189 30617 21223 30651
rect 21223 30617 21232 30651
rect 21180 30608 21232 30617
rect 21640 30608 21692 30660
rect 19432 30540 19484 30592
rect 10880 30438 10932 30490
rect 10944 30438 10996 30490
rect 11008 30438 11060 30490
rect 11072 30438 11124 30490
rect 11136 30438 11188 30490
rect 20811 30438 20863 30490
rect 20875 30438 20927 30490
rect 20939 30438 20991 30490
rect 21003 30438 21055 30490
rect 21067 30438 21119 30490
rect 4252 30379 4304 30388
rect 3424 30268 3476 30320
rect 4252 30345 4261 30379
rect 4261 30345 4295 30379
rect 4295 30345 4304 30379
rect 4252 30336 4304 30345
rect 4528 30336 4580 30388
rect 4804 30268 4856 30320
rect 2136 30200 2188 30252
rect 4620 30200 4672 30252
rect 5448 30268 5500 30320
rect 5356 30243 5408 30252
rect 5356 30209 5365 30243
rect 5365 30209 5399 30243
rect 5399 30209 5408 30243
rect 5356 30200 5408 30209
rect 6828 30243 6880 30252
rect 2872 30175 2924 30184
rect 2872 30141 2881 30175
rect 2881 30141 2915 30175
rect 2915 30141 2924 30175
rect 2872 30132 2924 30141
rect 5080 30132 5132 30184
rect 6828 30209 6837 30243
rect 6837 30209 6871 30243
rect 6871 30209 6880 30243
rect 6828 30200 6880 30209
rect 8024 30268 8076 30320
rect 10876 30268 10928 30320
rect 7104 30243 7156 30252
rect 7104 30209 7113 30243
rect 7113 30209 7147 30243
rect 7147 30209 7156 30243
rect 7104 30200 7156 30209
rect 7932 30243 7984 30252
rect 7932 30209 7941 30243
rect 7941 30209 7975 30243
rect 7975 30209 7984 30243
rect 7932 30200 7984 30209
rect 8576 30243 8628 30252
rect 8576 30209 8585 30243
rect 8585 30209 8619 30243
rect 8619 30209 8628 30243
rect 8576 30200 8628 30209
rect 9128 30243 9180 30252
rect 9128 30209 9137 30243
rect 9137 30209 9171 30243
rect 9171 30209 9180 30243
rect 9128 30200 9180 30209
rect 10416 30200 10468 30252
rect 11520 30243 11572 30252
rect 11520 30209 11529 30243
rect 11529 30209 11563 30243
rect 11563 30209 11572 30243
rect 11520 30200 11572 30209
rect 12992 30336 13044 30388
rect 14740 30379 14792 30388
rect 14740 30345 14749 30379
rect 14749 30345 14783 30379
rect 14783 30345 14792 30379
rect 14740 30336 14792 30345
rect 19524 30336 19576 30388
rect 20076 30336 20128 30388
rect 12256 30311 12308 30320
rect 12256 30277 12265 30311
rect 12265 30277 12299 30311
rect 12299 30277 12308 30311
rect 12256 30268 12308 30277
rect 12440 30268 12492 30320
rect 12164 30200 12216 30252
rect 13084 30243 13136 30252
rect 13084 30209 13093 30243
rect 13093 30209 13127 30243
rect 13127 30209 13136 30243
rect 13084 30200 13136 30209
rect 13360 30268 13412 30320
rect 15476 30311 15528 30320
rect 15476 30277 15485 30311
rect 15485 30277 15519 30311
rect 15519 30277 15528 30311
rect 15476 30268 15528 30277
rect 19340 30268 19392 30320
rect 20536 30268 20588 30320
rect 14096 30243 14148 30252
rect 14096 30209 14105 30243
rect 14105 30209 14139 30243
rect 14139 30209 14148 30243
rect 14096 30200 14148 30209
rect 6736 30175 6788 30184
rect 6736 30141 6745 30175
rect 6745 30141 6779 30175
rect 6779 30141 6788 30175
rect 6736 30132 6788 30141
rect 10600 30132 10652 30184
rect 10692 30132 10744 30184
rect 11888 30175 11940 30184
rect 11888 30141 11897 30175
rect 11897 30141 11931 30175
rect 11931 30141 11940 30175
rect 12808 30175 12860 30184
rect 11888 30132 11940 30141
rect 12808 30141 12817 30175
rect 12817 30141 12851 30175
rect 12851 30141 12860 30175
rect 12808 30132 12860 30141
rect 13452 30132 13504 30184
rect 2688 30064 2740 30116
rect 4896 30064 4948 30116
rect 5356 30064 5408 30116
rect 14464 30243 14516 30252
rect 14464 30209 14473 30243
rect 14473 30209 14507 30243
rect 14507 30209 14516 30243
rect 14464 30200 14516 30209
rect 14648 30200 14700 30252
rect 15660 30064 15712 30116
rect 16856 30200 16908 30252
rect 17868 30243 17920 30252
rect 17868 30209 17877 30243
rect 17877 30209 17911 30243
rect 17911 30209 17920 30243
rect 17868 30200 17920 30209
rect 19156 30243 19208 30252
rect 17132 30175 17184 30184
rect 17132 30141 17141 30175
rect 17141 30141 17175 30175
rect 17175 30141 17184 30175
rect 17132 30132 17184 30141
rect 17500 30132 17552 30184
rect 19156 30209 19165 30243
rect 19165 30209 19199 30243
rect 19199 30209 19208 30243
rect 19156 30200 19208 30209
rect 20720 30200 20772 30252
rect 22928 30243 22980 30252
rect 22928 30209 22937 30243
rect 22937 30209 22971 30243
rect 22971 30209 22980 30243
rect 22928 30200 22980 30209
rect 30104 30268 30156 30320
rect 20260 30132 20312 30184
rect 17040 30064 17092 30116
rect 18236 30064 18288 30116
rect 20168 30107 20220 30116
rect 20168 30073 20177 30107
rect 20177 30073 20211 30107
rect 20211 30073 20220 30107
rect 20168 30064 20220 30073
rect 30012 30107 30064 30116
rect 30012 30073 30021 30107
rect 30021 30073 30055 30107
rect 30055 30073 30064 30107
rect 30012 30064 30064 30073
rect 2320 29996 2372 30048
rect 6368 30039 6420 30048
rect 6368 30005 6377 30039
rect 6377 30005 6411 30039
rect 6411 30005 6420 30039
rect 6368 29996 6420 30005
rect 7288 29996 7340 30048
rect 7840 29996 7892 30048
rect 9312 30039 9364 30048
rect 9312 30005 9321 30039
rect 9321 30005 9355 30039
rect 9355 30005 9364 30039
rect 9312 29996 9364 30005
rect 9680 29996 9732 30048
rect 10232 29996 10284 30048
rect 15200 29996 15252 30048
rect 18052 30039 18104 30048
rect 18052 30005 18061 30039
rect 18061 30005 18095 30039
rect 18095 30005 18104 30039
rect 18052 29996 18104 30005
rect 21272 29996 21324 30048
rect 22652 29996 22704 30048
rect 5915 29894 5967 29946
rect 5979 29894 6031 29946
rect 6043 29894 6095 29946
rect 6107 29894 6159 29946
rect 6171 29894 6223 29946
rect 15846 29894 15898 29946
rect 15910 29894 15962 29946
rect 15974 29894 16026 29946
rect 16038 29894 16090 29946
rect 16102 29894 16154 29946
rect 25776 29894 25828 29946
rect 25840 29894 25892 29946
rect 25904 29894 25956 29946
rect 25968 29894 26020 29946
rect 26032 29894 26084 29946
rect 1492 29835 1544 29844
rect 1492 29801 1501 29835
rect 1501 29801 1535 29835
rect 1535 29801 1544 29835
rect 1492 29792 1544 29801
rect 2872 29792 2924 29844
rect 4804 29792 4856 29844
rect 11704 29792 11756 29844
rect 12348 29792 12400 29844
rect 13636 29792 13688 29844
rect 17132 29792 17184 29844
rect 17224 29792 17276 29844
rect 20076 29792 20128 29844
rect 11796 29767 11848 29776
rect 2320 29631 2372 29640
rect 2320 29597 2329 29631
rect 2329 29597 2363 29631
rect 2363 29597 2372 29631
rect 2320 29588 2372 29597
rect 11796 29733 11805 29767
rect 11805 29733 11839 29767
rect 11839 29733 11848 29767
rect 11796 29724 11848 29733
rect 12164 29724 12216 29776
rect 19156 29724 19208 29776
rect 21916 29767 21968 29776
rect 12716 29656 12768 29708
rect 17408 29656 17460 29708
rect 17500 29656 17552 29708
rect 18052 29699 18104 29708
rect 18052 29665 18061 29699
rect 18061 29665 18095 29699
rect 18095 29665 18104 29699
rect 18052 29656 18104 29665
rect 18144 29656 18196 29708
rect 19432 29699 19484 29708
rect 19432 29665 19441 29699
rect 19441 29665 19475 29699
rect 19475 29665 19484 29699
rect 19432 29656 19484 29665
rect 4620 29631 4672 29640
rect 4620 29597 4629 29631
rect 4629 29597 4663 29631
rect 4663 29597 4672 29631
rect 4620 29588 4672 29597
rect 5816 29588 5868 29640
rect 7472 29588 7524 29640
rect 11336 29588 11388 29640
rect 11612 29631 11664 29640
rect 11612 29597 11621 29631
rect 11621 29597 11655 29631
rect 11655 29597 11664 29631
rect 11612 29588 11664 29597
rect 14188 29631 14240 29640
rect 14188 29597 14197 29631
rect 14197 29597 14231 29631
rect 14231 29597 14240 29631
rect 14188 29588 14240 29597
rect 15292 29588 15344 29640
rect 16764 29631 16816 29640
rect 16764 29597 16773 29631
rect 16773 29597 16807 29631
rect 16807 29597 16816 29631
rect 16764 29588 16816 29597
rect 16948 29631 17000 29640
rect 16948 29597 16957 29631
rect 16957 29597 16991 29631
rect 16991 29597 17000 29631
rect 17132 29631 17184 29640
rect 16948 29588 17000 29597
rect 17132 29597 17141 29631
rect 17141 29597 17175 29631
rect 17175 29597 17184 29631
rect 17132 29588 17184 29597
rect 18512 29588 18564 29640
rect 21916 29733 21925 29767
rect 21925 29733 21959 29767
rect 21959 29733 21968 29767
rect 21916 29724 21968 29733
rect 21548 29656 21600 29708
rect 22376 29699 22428 29708
rect 22376 29665 22385 29699
rect 22385 29665 22419 29699
rect 22419 29665 22428 29699
rect 22376 29656 22428 29665
rect 6368 29520 6420 29572
rect 6552 29520 6604 29572
rect 9772 29520 9824 29572
rect 14004 29520 14056 29572
rect 19432 29520 19484 29572
rect 19984 29588 20036 29640
rect 20260 29520 20312 29572
rect 21456 29588 21508 29640
rect 22652 29631 22704 29640
rect 22652 29597 22686 29631
rect 22686 29597 22704 29631
rect 22652 29588 22704 29597
rect 21640 29520 21692 29572
rect 4436 29495 4488 29504
rect 4436 29461 4445 29495
rect 4445 29461 4479 29495
rect 4479 29461 4488 29495
rect 4436 29452 4488 29461
rect 6920 29452 6972 29504
rect 7656 29495 7708 29504
rect 7656 29461 7665 29495
rect 7665 29461 7699 29495
rect 7699 29461 7708 29495
rect 7656 29452 7708 29461
rect 18420 29452 18472 29504
rect 19340 29495 19392 29504
rect 19340 29461 19349 29495
rect 19349 29461 19383 29495
rect 19383 29461 19392 29495
rect 19340 29452 19392 29461
rect 21824 29452 21876 29504
rect 29736 29452 29788 29504
rect 10880 29350 10932 29402
rect 10944 29350 10996 29402
rect 11008 29350 11060 29402
rect 11072 29350 11124 29402
rect 11136 29350 11188 29402
rect 20811 29350 20863 29402
rect 20875 29350 20927 29402
rect 20939 29350 20991 29402
rect 21003 29350 21055 29402
rect 21067 29350 21119 29402
rect 2780 29291 2832 29300
rect 2780 29257 2789 29291
rect 2789 29257 2823 29291
rect 2823 29257 2832 29291
rect 2780 29248 2832 29257
rect 4712 29248 4764 29300
rect 5816 29291 5868 29300
rect 5816 29257 5825 29291
rect 5825 29257 5859 29291
rect 5859 29257 5868 29291
rect 5816 29248 5868 29257
rect 10508 29248 10560 29300
rect 11612 29248 11664 29300
rect 4160 29180 4212 29232
rect 9680 29180 9732 29232
rect 11060 29180 11112 29232
rect 1676 29155 1728 29164
rect 1676 29121 1685 29155
rect 1685 29121 1719 29155
rect 1719 29121 1728 29155
rect 1676 29112 1728 29121
rect 2504 29112 2556 29164
rect 2964 29155 3016 29164
rect 2964 29121 2973 29155
rect 2973 29121 3007 29155
rect 3007 29121 3016 29155
rect 2964 29112 3016 29121
rect 5632 29155 5684 29164
rect 5632 29121 5641 29155
rect 5641 29121 5675 29155
rect 5675 29121 5684 29155
rect 5632 29112 5684 29121
rect 8484 29112 8536 29164
rect 11796 29112 11848 29164
rect 12808 29248 12860 29300
rect 14004 29291 14056 29300
rect 12716 29180 12768 29232
rect 3792 29087 3844 29096
rect 3792 29053 3801 29087
rect 3801 29053 3835 29087
rect 3835 29053 3844 29087
rect 3792 29044 3844 29053
rect 7380 29087 7432 29096
rect 7380 29053 7389 29087
rect 7389 29053 7423 29087
rect 7423 29053 7432 29087
rect 7380 29044 7432 29053
rect 7748 29044 7800 29096
rect 13636 29223 13688 29232
rect 13636 29189 13645 29223
rect 13645 29189 13679 29223
rect 13679 29189 13688 29223
rect 13636 29180 13688 29189
rect 14004 29257 14013 29291
rect 14013 29257 14047 29291
rect 14047 29257 14056 29291
rect 14004 29248 14056 29257
rect 14096 29180 14148 29232
rect 15568 29180 15620 29232
rect 16948 29248 17000 29300
rect 17040 29248 17092 29300
rect 18236 29248 18288 29300
rect 18696 29248 18748 29300
rect 21548 29248 21600 29300
rect 21732 29248 21784 29300
rect 19984 29180 20036 29232
rect 13452 29155 13504 29164
rect 13452 29121 13462 29155
rect 13462 29121 13496 29155
rect 13496 29121 13504 29155
rect 13728 29155 13780 29164
rect 13452 29112 13504 29121
rect 13728 29121 13737 29155
rect 13737 29121 13771 29155
rect 13771 29121 13780 29155
rect 13728 29112 13780 29121
rect 14648 29112 14700 29164
rect 17040 29155 17092 29164
rect 14832 29044 14884 29096
rect 17040 29121 17049 29155
rect 17049 29121 17083 29155
rect 17083 29121 17092 29155
rect 17040 29112 17092 29121
rect 18144 29112 18196 29164
rect 18788 29155 18840 29164
rect 18236 29044 18288 29096
rect 18788 29121 18797 29155
rect 18797 29121 18831 29155
rect 18831 29121 18840 29155
rect 18788 29112 18840 29121
rect 19432 29155 19484 29164
rect 19432 29121 19441 29155
rect 19441 29121 19475 29155
rect 19475 29121 19484 29155
rect 19432 29112 19484 29121
rect 19800 29112 19852 29164
rect 21272 29112 21324 29164
rect 21456 29180 21508 29232
rect 29368 29112 29420 29164
rect 20444 29044 20496 29096
rect 1492 29019 1544 29028
rect 1492 28985 1501 29019
rect 1501 28985 1535 29019
rect 1535 28985 1544 29019
rect 1492 28976 1544 28985
rect 3056 28976 3108 29028
rect 6828 28976 6880 29028
rect 12348 28976 12400 29028
rect 14188 28976 14240 29028
rect 15660 28976 15712 29028
rect 22008 29044 22060 29096
rect 7012 28908 7064 28960
rect 18328 28908 18380 28960
rect 19616 28908 19668 28960
rect 5915 28806 5967 28858
rect 5979 28806 6031 28858
rect 6043 28806 6095 28858
rect 6107 28806 6159 28858
rect 6171 28806 6223 28858
rect 15846 28806 15898 28858
rect 15910 28806 15962 28858
rect 15974 28806 16026 28858
rect 16038 28806 16090 28858
rect 16102 28806 16154 28858
rect 25776 28806 25828 28858
rect 25840 28806 25892 28858
rect 25904 28806 25956 28858
rect 25968 28806 26020 28858
rect 26032 28806 26084 28858
rect 1676 28704 1728 28756
rect 3792 28747 3844 28756
rect 3792 28713 3801 28747
rect 3801 28713 3835 28747
rect 3835 28713 3844 28747
rect 3792 28704 3844 28713
rect 5632 28704 5684 28756
rect 7380 28704 7432 28756
rect 11428 28704 11480 28756
rect 12256 28704 12308 28756
rect 15292 28704 15344 28756
rect 15660 28747 15712 28756
rect 15660 28713 15669 28747
rect 15669 28713 15703 28747
rect 15703 28713 15712 28747
rect 15660 28704 15712 28713
rect 17224 28704 17276 28756
rect 12900 28636 12952 28688
rect 7748 28568 7800 28620
rect 11888 28568 11940 28620
rect 12532 28568 12584 28620
rect 4436 28500 4488 28552
rect 4620 28543 4672 28552
rect 4620 28509 4629 28543
rect 4629 28509 4663 28543
rect 4663 28509 4672 28543
rect 4620 28500 4672 28509
rect 6460 28500 6512 28552
rect 7656 28500 7708 28552
rect 9312 28543 9364 28552
rect 1492 28407 1544 28416
rect 1492 28373 1501 28407
rect 1501 28373 1535 28407
rect 1535 28373 1544 28407
rect 1492 28364 1544 28373
rect 3148 28432 3200 28484
rect 9312 28509 9321 28543
rect 9321 28509 9355 28543
rect 9355 28509 9364 28543
rect 9312 28500 9364 28509
rect 10324 28543 10376 28552
rect 10324 28509 10333 28543
rect 10333 28509 10367 28543
rect 10367 28509 10376 28543
rect 10324 28500 10376 28509
rect 10784 28500 10836 28552
rect 11060 28543 11112 28552
rect 11060 28509 11069 28543
rect 11069 28509 11103 28543
rect 11103 28509 11112 28543
rect 11060 28500 11112 28509
rect 11796 28543 11848 28552
rect 11796 28509 11805 28543
rect 11805 28509 11839 28543
rect 11839 28509 11848 28543
rect 11796 28500 11848 28509
rect 11980 28500 12032 28552
rect 13452 28568 13504 28620
rect 19432 28636 19484 28688
rect 14096 28568 14148 28620
rect 17868 28568 17920 28620
rect 13544 28500 13596 28552
rect 15200 28500 15252 28552
rect 15476 28500 15528 28552
rect 16948 28543 17000 28552
rect 16948 28509 16957 28543
rect 16957 28509 16991 28543
rect 16991 28509 17000 28543
rect 16948 28500 17000 28509
rect 17500 28500 17552 28552
rect 18052 28543 18104 28552
rect 18052 28509 18061 28543
rect 18061 28509 18095 28543
rect 18095 28509 18104 28543
rect 18052 28500 18104 28509
rect 9496 28432 9548 28484
rect 12164 28432 12216 28484
rect 14096 28432 14148 28484
rect 14832 28475 14884 28484
rect 14832 28441 14841 28475
rect 14841 28441 14875 28475
rect 14875 28441 14884 28475
rect 14832 28432 14884 28441
rect 18328 28543 18380 28552
rect 18328 28509 18337 28543
rect 18337 28509 18371 28543
rect 18371 28509 18380 28543
rect 18328 28500 18380 28509
rect 18604 28500 18656 28552
rect 21180 28704 21232 28756
rect 21548 28704 21600 28756
rect 22928 28704 22980 28756
rect 22008 28636 22060 28688
rect 21824 28611 21876 28620
rect 21824 28577 21833 28611
rect 21833 28577 21867 28611
rect 21867 28577 21876 28611
rect 21824 28568 21876 28577
rect 21916 28568 21968 28620
rect 7012 28364 7064 28416
rect 7104 28407 7156 28416
rect 7104 28373 7113 28407
rect 7113 28373 7147 28407
rect 7147 28373 7156 28407
rect 7104 28364 7156 28373
rect 8668 28364 8720 28416
rect 8944 28407 8996 28416
rect 8944 28373 8953 28407
rect 8953 28373 8987 28407
rect 8987 28373 8996 28407
rect 8944 28364 8996 28373
rect 9404 28407 9456 28416
rect 9404 28373 9413 28407
rect 9413 28373 9447 28407
rect 9447 28373 9456 28407
rect 9404 28364 9456 28373
rect 10232 28407 10284 28416
rect 10232 28373 10241 28407
rect 10241 28373 10275 28407
rect 10275 28373 10284 28407
rect 10232 28364 10284 28373
rect 13176 28364 13228 28416
rect 18236 28364 18288 28416
rect 18512 28364 18564 28416
rect 20628 28543 20680 28552
rect 20628 28509 20637 28543
rect 20637 28509 20671 28543
rect 20671 28509 20680 28543
rect 20628 28500 20680 28509
rect 22560 28500 22612 28552
rect 29828 28543 29880 28552
rect 29828 28509 29837 28543
rect 29837 28509 29871 28543
rect 29871 28509 29880 28543
rect 29828 28500 29880 28509
rect 20720 28432 20772 28484
rect 21916 28432 21968 28484
rect 21824 28364 21876 28416
rect 22192 28407 22244 28416
rect 22192 28373 22201 28407
rect 22201 28373 22235 28407
rect 22235 28373 22244 28407
rect 30012 28407 30064 28416
rect 22192 28364 22244 28373
rect 30012 28373 30021 28407
rect 30021 28373 30055 28407
rect 30055 28373 30064 28407
rect 30012 28364 30064 28373
rect 10880 28262 10932 28314
rect 10944 28262 10996 28314
rect 11008 28262 11060 28314
rect 11072 28262 11124 28314
rect 11136 28262 11188 28314
rect 20811 28262 20863 28314
rect 20875 28262 20927 28314
rect 20939 28262 20991 28314
rect 21003 28262 21055 28314
rect 21067 28262 21119 28314
rect 2044 28160 2096 28212
rect 7104 28160 7156 28212
rect 9404 28160 9456 28212
rect 2412 28024 2464 28076
rect 3332 28024 3384 28076
rect 8944 28092 8996 28144
rect 10048 28160 10100 28212
rect 14096 28160 14148 28212
rect 17132 28160 17184 28212
rect 18604 28203 18656 28212
rect 18604 28169 18613 28203
rect 18613 28169 18647 28203
rect 18647 28169 18656 28203
rect 18604 28160 18656 28169
rect 18788 28160 18840 28212
rect 20628 28160 20680 28212
rect 21916 28203 21968 28212
rect 21916 28169 21925 28203
rect 21925 28169 21959 28203
rect 21959 28169 21968 28203
rect 21916 28160 21968 28169
rect 22192 28160 22244 28212
rect 29460 28160 29512 28212
rect 29828 28160 29880 28212
rect 3148 27956 3200 28008
rect 8668 28067 8720 28076
rect 8668 28033 8677 28067
rect 8677 28033 8711 28067
rect 8711 28033 8720 28067
rect 8668 28024 8720 28033
rect 8760 28067 8812 28076
rect 8760 28033 8769 28067
rect 8769 28033 8803 28067
rect 8803 28033 8812 28067
rect 11336 28092 11388 28144
rect 12532 28092 12584 28144
rect 8760 28024 8812 28033
rect 9864 28067 9916 28076
rect 9864 28033 9898 28067
rect 9898 28033 9916 28067
rect 9864 28024 9916 28033
rect 10324 28024 10376 28076
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 12624 28024 12676 28076
rect 14188 28092 14240 28144
rect 13176 28067 13228 28076
rect 13176 28033 13210 28067
rect 13210 28033 13228 28067
rect 13176 28024 13228 28033
rect 13544 28024 13596 28076
rect 14464 28024 14516 28076
rect 14832 28024 14884 28076
rect 16672 28067 16724 28076
rect 11796 27956 11848 28008
rect 12532 27956 12584 28008
rect 14372 27956 14424 28008
rect 16672 28033 16681 28067
rect 16681 28033 16715 28067
rect 16715 28033 16724 28067
rect 16672 28024 16724 28033
rect 16856 28067 16908 28076
rect 16856 28033 16865 28067
rect 16865 28033 16899 28067
rect 16899 28033 16908 28067
rect 16856 28024 16908 28033
rect 17868 28067 17920 28076
rect 17868 28033 17877 28067
rect 17877 28033 17911 28067
rect 17911 28033 17920 28067
rect 17868 28024 17920 28033
rect 18052 28067 18104 28076
rect 18052 28033 18061 28067
rect 18061 28033 18095 28067
rect 18095 28033 18104 28067
rect 18052 28024 18104 28033
rect 18880 28092 18932 28144
rect 18420 28067 18472 28076
rect 18420 28033 18429 28067
rect 18429 28033 18463 28067
rect 18463 28033 18472 28067
rect 18420 28024 18472 28033
rect 18512 28024 18564 28076
rect 20444 28067 20496 28076
rect 20444 28033 20453 28067
rect 20453 28033 20487 28067
rect 20487 28033 20496 28067
rect 20444 28024 20496 28033
rect 20628 28024 20680 28076
rect 21456 28024 21508 28076
rect 21824 28067 21876 28076
rect 21824 28033 21833 28067
rect 21833 28033 21867 28067
rect 21867 28033 21876 28067
rect 21824 28024 21876 28033
rect 29644 28024 29696 28076
rect 30104 28067 30156 28076
rect 30104 28033 30113 28067
rect 30113 28033 30147 28067
rect 30147 28033 30156 28067
rect 30104 28024 30156 28033
rect 17960 27956 18012 28008
rect 19524 27999 19576 28008
rect 19524 27965 19533 27999
rect 19533 27965 19567 27999
rect 19567 27965 19576 27999
rect 19524 27956 19576 27965
rect 12072 27888 12124 27940
rect 18604 27888 18656 27940
rect 20536 27931 20588 27940
rect 20536 27897 20545 27931
rect 20545 27897 20579 27931
rect 20579 27897 20588 27931
rect 20536 27888 20588 27897
rect 21180 27888 21232 27940
rect 1492 27863 1544 27872
rect 1492 27829 1501 27863
rect 1501 27829 1535 27863
rect 1535 27829 1544 27863
rect 1492 27820 1544 27829
rect 2780 27820 2832 27872
rect 3608 27820 3660 27872
rect 7196 27820 7248 27872
rect 7932 27820 7984 27872
rect 9496 27820 9548 27872
rect 15568 27863 15620 27872
rect 15568 27829 15577 27863
rect 15577 27829 15611 27863
rect 15611 27829 15620 27863
rect 15568 27820 15620 27829
rect 16672 27820 16724 27872
rect 19432 27820 19484 27872
rect 5915 27718 5967 27770
rect 5979 27718 6031 27770
rect 6043 27718 6095 27770
rect 6107 27718 6159 27770
rect 6171 27718 6223 27770
rect 15846 27718 15898 27770
rect 15910 27718 15962 27770
rect 15974 27718 16026 27770
rect 16038 27718 16090 27770
rect 16102 27718 16154 27770
rect 25776 27718 25828 27770
rect 25840 27718 25892 27770
rect 25904 27718 25956 27770
rect 25968 27718 26020 27770
rect 26032 27718 26084 27770
rect 3332 27616 3384 27668
rect 9128 27616 9180 27668
rect 5816 27591 5868 27600
rect 5816 27557 5825 27591
rect 5825 27557 5859 27591
rect 5859 27557 5868 27591
rect 5816 27548 5868 27557
rect 7472 27548 7524 27600
rect 3148 27412 3200 27464
rect 1676 27276 1728 27328
rect 4620 27344 4672 27396
rect 5724 27455 5776 27464
rect 5724 27421 5733 27455
rect 5733 27421 5767 27455
rect 5767 27421 5776 27455
rect 5724 27412 5776 27421
rect 6368 27412 6420 27464
rect 7380 27455 7432 27464
rect 7380 27421 7389 27455
rect 7389 27421 7423 27455
rect 7423 27421 7432 27455
rect 7380 27412 7432 27421
rect 8760 27548 8812 27600
rect 9036 27548 9088 27600
rect 8208 27480 8260 27532
rect 9312 27548 9364 27600
rect 9496 27616 9548 27668
rect 10784 27616 10836 27668
rect 9680 27591 9732 27600
rect 9680 27557 9689 27591
rect 9689 27557 9723 27591
rect 9723 27557 9732 27591
rect 9680 27548 9732 27557
rect 11980 27616 12032 27668
rect 16856 27616 16908 27668
rect 18052 27616 18104 27668
rect 19616 27616 19668 27668
rect 19800 27616 19852 27668
rect 19984 27616 20036 27668
rect 20536 27616 20588 27668
rect 19524 27548 19576 27600
rect 20076 27591 20128 27600
rect 20076 27557 20085 27591
rect 20085 27557 20119 27591
rect 20119 27557 20128 27591
rect 20076 27548 20128 27557
rect 10324 27480 10376 27532
rect 11336 27523 11388 27532
rect 8392 27455 8444 27464
rect 8392 27421 8401 27455
rect 8401 27421 8435 27455
rect 8435 27421 8444 27455
rect 8392 27412 8444 27421
rect 8852 27412 8904 27464
rect 9128 27455 9180 27464
rect 9128 27421 9141 27455
rect 9141 27421 9175 27455
rect 9175 27421 9180 27455
rect 9128 27412 9180 27421
rect 6000 27344 6052 27396
rect 9312 27421 9321 27442
rect 9321 27421 9355 27442
rect 9355 27421 9364 27442
rect 9312 27390 9364 27421
rect 10232 27412 10284 27464
rect 6828 27276 6880 27328
rect 7104 27276 7156 27328
rect 10508 27344 10560 27396
rect 9588 27276 9640 27328
rect 11336 27489 11345 27523
rect 11345 27489 11379 27523
rect 11379 27489 11388 27523
rect 11336 27480 11388 27489
rect 14096 27480 14148 27532
rect 10784 27455 10836 27464
rect 10784 27421 10793 27455
rect 10793 27421 10827 27455
rect 10827 27421 10836 27455
rect 10784 27412 10836 27421
rect 10876 27455 10928 27464
rect 10876 27421 10885 27455
rect 10885 27421 10919 27455
rect 10919 27421 10928 27455
rect 14372 27455 14424 27464
rect 10876 27412 10928 27421
rect 14372 27421 14381 27455
rect 14381 27421 14415 27455
rect 14415 27421 14424 27455
rect 14372 27412 14424 27421
rect 15292 27455 15344 27464
rect 11428 27344 11480 27396
rect 15292 27421 15301 27455
rect 15301 27421 15335 27455
rect 15335 27421 15344 27455
rect 15292 27412 15344 27421
rect 10784 27276 10836 27328
rect 14740 27344 14792 27396
rect 17500 27480 17552 27532
rect 18604 27480 18656 27532
rect 17224 27412 17276 27464
rect 18420 27412 18472 27464
rect 17592 27344 17644 27396
rect 19800 27480 19852 27532
rect 19432 27412 19484 27464
rect 20260 27455 20312 27464
rect 20260 27421 20269 27455
rect 20269 27421 20303 27455
rect 20303 27421 20312 27455
rect 20260 27412 20312 27421
rect 21364 27455 21416 27464
rect 21364 27421 21373 27455
rect 21373 27421 21407 27455
rect 21407 27421 21416 27455
rect 21364 27412 21416 27421
rect 21640 27455 21692 27464
rect 21640 27421 21649 27455
rect 21649 27421 21683 27455
rect 21683 27421 21692 27455
rect 21640 27412 21692 27421
rect 29920 27412 29972 27464
rect 16488 27319 16540 27328
rect 16488 27285 16497 27319
rect 16497 27285 16531 27319
rect 16531 27285 16540 27319
rect 16488 27276 16540 27285
rect 18604 27276 18656 27328
rect 30012 27319 30064 27328
rect 30012 27285 30021 27319
rect 30021 27285 30055 27319
rect 30055 27285 30064 27319
rect 30012 27276 30064 27285
rect 10880 27174 10932 27226
rect 10944 27174 10996 27226
rect 11008 27174 11060 27226
rect 11072 27174 11124 27226
rect 11136 27174 11188 27226
rect 20811 27174 20863 27226
rect 20875 27174 20927 27226
rect 20939 27174 20991 27226
rect 21003 27174 21055 27226
rect 21067 27174 21119 27226
rect 6552 27072 6604 27124
rect 8576 27072 8628 27124
rect 10324 27072 10376 27124
rect 11428 27072 11480 27124
rect 11796 27072 11848 27124
rect 13728 27072 13780 27124
rect 17040 27072 17092 27124
rect 17224 27115 17276 27124
rect 17224 27081 17233 27115
rect 17233 27081 17267 27115
rect 17267 27081 17276 27115
rect 17224 27072 17276 27081
rect 18144 27115 18196 27124
rect 18144 27081 18153 27115
rect 18153 27081 18187 27115
rect 18187 27081 18196 27115
rect 18144 27072 18196 27081
rect 21364 27072 21416 27124
rect 21824 27072 21876 27124
rect 29920 27115 29972 27124
rect 29920 27081 29929 27115
rect 29929 27081 29963 27115
rect 29963 27081 29972 27115
rect 29920 27072 29972 27081
rect 7472 27004 7524 27056
rect 8024 27004 8076 27056
rect 13360 27004 13412 27056
rect 1676 26979 1728 26988
rect 1676 26945 1685 26979
rect 1685 26945 1719 26979
rect 1719 26945 1728 26979
rect 1676 26936 1728 26945
rect 5540 26979 5592 26988
rect 5540 26945 5558 26979
rect 5558 26945 5592 26979
rect 5540 26936 5592 26945
rect 7012 26936 7064 26988
rect 7104 26979 7156 26988
rect 7104 26945 7113 26979
rect 7113 26945 7147 26979
rect 7147 26945 7156 26979
rect 7104 26936 7156 26945
rect 8300 26936 8352 26988
rect 6828 26868 6880 26920
rect 1492 26843 1544 26852
rect 1492 26809 1501 26843
rect 1501 26809 1535 26843
rect 1535 26809 1544 26843
rect 1492 26800 1544 26809
rect 7932 26868 7984 26920
rect 8392 26800 8444 26852
rect 8944 26936 8996 26988
rect 9220 26979 9272 26988
rect 9220 26945 9230 26979
rect 9230 26945 9264 26979
rect 9264 26945 9272 26979
rect 9404 26979 9456 26988
rect 9220 26936 9272 26945
rect 9404 26945 9413 26979
rect 9413 26945 9447 26979
rect 9447 26945 9456 26979
rect 9404 26936 9456 26945
rect 8668 26868 8720 26920
rect 9588 26979 9640 26988
rect 9588 26945 9602 26979
rect 9602 26945 9636 26979
rect 9636 26945 9640 26979
rect 10232 26979 10284 26988
rect 9588 26936 9640 26945
rect 10232 26945 10241 26979
rect 10241 26945 10275 26979
rect 10275 26945 10284 26979
rect 10232 26936 10284 26945
rect 10324 26936 10376 26988
rect 10508 26979 10560 26988
rect 10508 26945 10517 26979
rect 10517 26945 10551 26979
rect 10551 26945 10560 26979
rect 10784 26979 10836 26988
rect 10508 26936 10560 26945
rect 10784 26945 10793 26979
rect 10793 26945 10827 26979
rect 10827 26945 10836 26979
rect 10784 26936 10836 26945
rect 12624 26979 12676 26988
rect 12624 26945 12633 26979
rect 12633 26945 12667 26979
rect 12667 26945 12676 26979
rect 12624 26936 12676 26945
rect 12716 26936 12768 26988
rect 14004 26936 14056 26988
rect 14372 26936 14424 26988
rect 14924 26979 14976 26988
rect 14924 26945 14933 26979
rect 14933 26945 14967 26979
rect 14967 26945 14976 26979
rect 14924 26936 14976 26945
rect 15568 27004 15620 27056
rect 21088 27004 21140 27056
rect 12348 26868 12400 26920
rect 14740 26911 14792 26920
rect 14740 26877 14749 26911
rect 14749 26877 14783 26911
rect 14783 26877 14792 26911
rect 14740 26868 14792 26877
rect 15108 26868 15160 26920
rect 18328 26936 18380 26988
rect 17316 26911 17368 26920
rect 17316 26877 17325 26911
rect 17325 26877 17359 26911
rect 17359 26877 17368 26911
rect 17316 26868 17368 26877
rect 17500 26911 17552 26920
rect 17500 26877 17509 26911
rect 17509 26877 17543 26911
rect 17543 26877 17552 26911
rect 17500 26868 17552 26877
rect 18604 26911 18656 26920
rect 18604 26877 18613 26911
rect 18613 26877 18647 26911
rect 18647 26877 18656 26911
rect 18604 26868 18656 26877
rect 18696 26911 18748 26920
rect 18696 26877 18705 26911
rect 18705 26877 18739 26911
rect 18739 26877 18748 26911
rect 20260 26936 20312 26988
rect 21916 26936 21968 26988
rect 22100 26979 22152 26988
rect 22100 26945 22134 26979
rect 22134 26945 22152 26979
rect 30104 26979 30156 26988
rect 22100 26936 22152 26945
rect 30104 26945 30113 26979
rect 30113 26945 30147 26979
rect 30147 26945 30156 26979
rect 30104 26936 30156 26945
rect 18696 26868 18748 26877
rect 20628 26868 20680 26920
rect 12440 26800 12492 26852
rect 20260 26800 20312 26852
rect 20536 26800 20588 26852
rect 21732 26868 21784 26920
rect 4896 26732 4948 26784
rect 7472 26732 7524 26784
rect 9312 26732 9364 26784
rect 9864 26732 9916 26784
rect 14004 26775 14056 26784
rect 14004 26741 14013 26775
rect 14013 26741 14047 26775
rect 14047 26741 14056 26775
rect 14004 26732 14056 26741
rect 16304 26732 16356 26784
rect 19432 26732 19484 26784
rect 21180 26732 21232 26784
rect 21548 26732 21600 26784
rect 22008 26732 22060 26784
rect 5915 26630 5967 26682
rect 5979 26630 6031 26682
rect 6043 26630 6095 26682
rect 6107 26630 6159 26682
rect 6171 26630 6223 26682
rect 15846 26630 15898 26682
rect 15910 26630 15962 26682
rect 15974 26630 16026 26682
rect 16038 26630 16090 26682
rect 16102 26630 16154 26682
rect 25776 26630 25828 26682
rect 25840 26630 25892 26682
rect 25904 26630 25956 26682
rect 25968 26630 26020 26682
rect 26032 26630 26084 26682
rect 2872 26324 2924 26376
rect 3148 26324 3200 26376
rect 8300 26571 8352 26580
rect 8300 26537 8309 26571
rect 8309 26537 8343 26571
rect 8343 26537 8352 26571
rect 8300 26528 8352 26537
rect 9772 26528 9824 26580
rect 10324 26528 10376 26580
rect 12072 26528 12124 26580
rect 12716 26528 12768 26580
rect 14740 26528 14792 26580
rect 14924 26528 14976 26580
rect 16488 26571 16540 26580
rect 3792 26503 3844 26512
rect 3792 26469 3801 26503
rect 3801 26469 3835 26503
rect 3835 26469 3844 26503
rect 3792 26460 3844 26469
rect 5908 26392 5960 26444
rect 5264 26324 5316 26376
rect 5356 26324 5408 26376
rect 7472 26435 7524 26444
rect 7472 26401 7481 26435
rect 7481 26401 7515 26435
rect 7515 26401 7524 26435
rect 7472 26392 7524 26401
rect 7656 26435 7708 26444
rect 7656 26401 7665 26435
rect 7665 26401 7699 26435
rect 7699 26401 7708 26435
rect 7656 26392 7708 26401
rect 6092 26367 6144 26376
rect 6092 26333 6137 26367
rect 6137 26333 6144 26367
rect 6092 26324 6144 26333
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6276 26324 6328 26333
rect 7840 26324 7892 26376
rect 8300 26324 8352 26376
rect 8576 26324 8628 26376
rect 8944 26324 8996 26376
rect 9220 26367 9272 26376
rect 9220 26333 9227 26367
rect 9227 26333 9272 26367
rect 9220 26324 9272 26333
rect 11704 26460 11756 26512
rect 9496 26367 9548 26376
rect 9496 26333 9510 26367
rect 9510 26333 9544 26367
rect 9544 26333 9548 26367
rect 9496 26324 9548 26333
rect 9680 26324 9732 26376
rect 10600 26324 10652 26376
rect 10784 26324 10836 26376
rect 11704 26324 11756 26376
rect 12072 26367 12124 26376
rect 12072 26333 12081 26367
rect 12081 26333 12115 26367
rect 12115 26333 12124 26367
rect 12072 26324 12124 26333
rect 14004 26392 14056 26444
rect 8116 26256 8168 26308
rect 9404 26299 9456 26308
rect 9404 26265 9413 26299
rect 9413 26265 9447 26299
rect 9447 26265 9456 26299
rect 9404 26256 9456 26265
rect 9588 26256 9640 26308
rect 1492 26231 1544 26240
rect 1492 26197 1501 26231
rect 1501 26197 1535 26231
rect 1535 26197 1544 26231
rect 1492 26188 1544 26197
rect 2964 26188 3016 26240
rect 4712 26188 4764 26240
rect 5356 26188 5408 26240
rect 5816 26188 5868 26240
rect 9772 26188 9824 26240
rect 10140 26256 10192 26308
rect 11796 26188 11848 26240
rect 14096 26324 14148 26376
rect 16488 26537 16497 26571
rect 16497 26537 16531 26571
rect 16531 26537 16540 26571
rect 16488 26528 16540 26537
rect 17868 26528 17920 26580
rect 19524 26528 19576 26580
rect 20444 26528 20496 26580
rect 19892 26460 19944 26512
rect 20720 26460 20772 26512
rect 21180 26392 21232 26444
rect 21732 26435 21784 26444
rect 21732 26401 21741 26435
rect 21741 26401 21775 26435
rect 21775 26401 21784 26435
rect 21732 26392 21784 26401
rect 16304 26367 16356 26376
rect 14924 26256 14976 26308
rect 15108 26256 15160 26308
rect 16304 26333 16313 26367
rect 16313 26333 16347 26367
rect 16347 26333 16356 26367
rect 16304 26324 16356 26333
rect 16764 26324 16816 26376
rect 18236 26367 18288 26376
rect 18236 26333 18245 26367
rect 18245 26333 18279 26367
rect 18279 26333 18288 26367
rect 18236 26324 18288 26333
rect 19432 26324 19484 26376
rect 19708 26324 19760 26376
rect 19892 26367 19944 26376
rect 19892 26333 19901 26367
rect 19901 26333 19935 26367
rect 19935 26333 19944 26367
rect 20536 26367 20588 26376
rect 19892 26324 19944 26333
rect 20536 26333 20545 26367
rect 20545 26333 20579 26367
rect 20579 26333 20588 26367
rect 20536 26324 20588 26333
rect 20628 26324 20680 26376
rect 21088 26367 21140 26376
rect 17592 26299 17644 26308
rect 17592 26265 17601 26299
rect 17601 26265 17635 26299
rect 17635 26265 17644 26299
rect 17592 26256 17644 26265
rect 17960 26256 18012 26308
rect 21088 26333 21097 26367
rect 21097 26333 21131 26367
rect 21131 26333 21140 26367
rect 21088 26324 21140 26333
rect 21364 26324 21416 26376
rect 12348 26188 12400 26240
rect 14556 26231 14608 26240
rect 14556 26197 14565 26231
rect 14565 26197 14599 26231
rect 14599 26197 14608 26231
rect 14556 26188 14608 26197
rect 15752 26231 15804 26240
rect 15752 26197 15761 26231
rect 15761 26197 15795 26231
rect 15795 26197 15804 26231
rect 15752 26188 15804 26197
rect 18052 26188 18104 26240
rect 18236 26188 18288 26240
rect 20720 26188 20772 26240
rect 22192 26188 22244 26240
rect 10880 26086 10932 26138
rect 10944 26086 10996 26138
rect 11008 26086 11060 26138
rect 11072 26086 11124 26138
rect 11136 26086 11188 26138
rect 20811 26086 20863 26138
rect 20875 26086 20927 26138
rect 20939 26086 20991 26138
rect 21003 26086 21055 26138
rect 21067 26086 21119 26138
rect 2872 25984 2924 26036
rect 5540 25984 5592 26036
rect 4896 25959 4948 25968
rect 4896 25925 4905 25959
rect 4905 25925 4939 25959
rect 4939 25925 4948 25959
rect 4896 25916 4948 25925
rect 2964 25848 3016 25900
rect 3148 25891 3200 25900
rect 3148 25857 3157 25891
rect 3157 25857 3191 25891
rect 3191 25857 3200 25891
rect 3148 25848 3200 25857
rect 4712 25891 4764 25900
rect 4712 25857 4716 25891
rect 4716 25857 4750 25891
rect 4750 25857 4764 25891
rect 4712 25848 4764 25857
rect 4804 25891 4856 25900
rect 4804 25857 4813 25891
rect 4813 25857 4847 25891
rect 4847 25857 4856 25891
rect 5080 25891 5132 25900
rect 4804 25848 4856 25857
rect 5080 25857 5088 25891
rect 5088 25857 5122 25891
rect 5122 25857 5132 25891
rect 5080 25848 5132 25857
rect 6276 25984 6328 26036
rect 6828 25984 6880 26036
rect 5816 25891 5868 25900
rect 5816 25857 5825 25891
rect 5825 25857 5859 25891
rect 5859 25857 5868 25891
rect 5816 25848 5868 25857
rect 5908 25848 5960 25900
rect 6736 25891 6788 25900
rect 6736 25857 6745 25891
rect 6745 25857 6779 25891
rect 6779 25857 6788 25891
rect 6736 25848 6788 25857
rect 7012 25916 7064 25968
rect 8024 25916 8076 25968
rect 9128 25916 9180 25968
rect 7380 25848 7432 25900
rect 8576 25848 8628 25900
rect 9772 25984 9824 26036
rect 10324 25984 10376 26036
rect 15752 25984 15804 26036
rect 17592 26027 17644 26036
rect 17592 25993 17601 26027
rect 17601 25993 17635 26027
rect 17635 25993 17644 26027
rect 17592 25984 17644 25993
rect 19892 25984 19944 26036
rect 21916 26027 21968 26036
rect 13360 25959 13412 25968
rect 13360 25925 13369 25959
rect 13369 25925 13403 25959
rect 13403 25925 13412 25959
rect 13360 25916 13412 25925
rect 18604 25916 18656 25968
rect 19524 25916 19576 25968
rect 19800 25916 19852 25968
rect 8760 25823 8812 25832
rect 5724 25712 5776 25764
rect 8760 25789 8769 25823
rect 8769 25789 8803 25823
rect 8803 25789 8812 25823
rect 8760 25780 8812 25789
rect 9588 25848 9640 25900
rect 9772 25891 9824 25900
rect 9772 25857 9806 25891
rect 9806 25857 9824 25891
rect 9772 25848 9824 25857
rect 11704 25848 11756 25900
rect 1492 25687 1544 25696
rect 1492 25653 1501 25687
rect 1501 25653 1535 25687
rect 1535 25653 1544 25687
rect 1492 25644 1544 25653
rect 6276 25644 6328 25696
rect 11428 25780 11480 25832
rect 12256 25891 12308 25900
rect 12256 25857 12265 25891
rect 12265 25857 12299 25891
rect 12299 25857 12308 25891
rect 12256 25848 12308 25857
rect 12900 25848 12952 25900
rect 16488 25848 16540 25900
rect 17040 25848 17092 25900
rect 18420 25848 18472 25900
rect 18972 25848 19024 25900
rect 12348 25823 12400 25832
rect 12348 25789 12357 25823
rect 12357 25789 12391 25823
rect 12391 25789 12400 25823
rect 12348 25780 12400 25789
rect 16856 25780 16908 25832
rect 18052 25823 18104 25832
rect 18052 25789 18061 25823
rect 18061 25789 18095 25823
rect 18095 25789 18104 25823
rect 18052 25780 18104 25789
rect 11888 25712 11940 25764
rect 17500 25712 17552 25764
rect 19524 25780 19576 25832
rect 20536 25891 20588 25900
rect 19800 25823 19852 25832
rect 19800 25789 19809 25823
rect 19809 25789 19843 25823
rect 19843 25789 19852 25823
rect 19800 25780 19852 25789
rect 20536 25857 20545 25891
rect 20545 25857 20579 25891
rect 20579 25857 20588 25891
rect 20536 25848 20588 25857
rect 21364 25916 21416 25968
rect 20812 25891 20864 25900
rect 20812 25857 20821 25891
rect 20821 25857 20855 25891
rect 20855 25857 20864 25891
rect 21088 25891 21140 25900
rect 20812 25848 20864 25857
rect 21088 25857 21097 25891
rect 21097 25857 21131 25891
rect 21131 25857 21140 25891
rect 21088 25848 21140 25857
rect 21916 25993 21925 26027
rect 21925 25993 21959 26027
rect 21959 25993 21968 26027
rect 21916 25984 21968 25993
rect 22008 25891 22060 25900
rect 22008 25857 22017 25891
rect 22017 25857 22051 25891
rect 22051 25857 22060 25891
rect 22008 25848 22060 25857
rect 29184 25848 29236 25900
rect 20812 25712 20864 25764
rect 22100 25780 22152 25832
rect 14004 25644 14056 25696
rect 16212 25644 16264 25696
rect 17684 25644 17736 25696
rect 19616 25687 19668 25696
rect 19616 25653 19625 25687
rect 19625 25653 19659 25687
rect 19659 25653 19668 25687
rect 19616 25644 19668 25653
rect 19984 25644 20036 25696
rect 20628 25644 20680 25696
rect 30012 25687 30064 25696
rect 30012 25653 30021 25687
rect 30021 25653 30055 25687
rect 30055 25653 30064 25687
rect 30012 25644 30064 25653
rect 5915 25542 5967 25594
rect 5979 25542 6031 25594
rect 6043 25542 6095 25594
rect 6107 25542 6159 25594
rect 6171 25542 6223 25594
rect 15846 25542 15898 25594
rect 15910 25542 15962 25594
rect 15974 25542 16026 25594
rect 16038 25542 16090 25594
rect 16102 25542 16154 25594
rect 25776 25542 25828 25594
rect 25840 25542 25892 25594
rect 25904 25542 25956 25594
rect 25968 25542 26020 25594
rect 26032 25542 26084 25594
rect 4160 25372 4212 25424
rect 7472 25347 7524 25356
rect 7472 25313 7481 25347
rect 7481 25313 7515 25347
rect 7515 25313 7524 25347
rect 7472 25304 7524 25313
rect 7656 25304 7708 25356
rect 7748 25304 7800 25356
rect 8392 25304 8444 25356
rect 6276 25279 6328 25288
rect 6276 25245 6285 25279
rect 6285 25245 6319 25279
rect 6319 25245 6328 25279
rect 6276 25236 6328 25245
rect 7840 25236 7892 25288
rect 8760 25236 8812 25288
rect 6552 25168 6604 25220
rect 7288 25211 7340 25220
rect 7288 25177 7297 25211
rect 7297 25177 7331 25211
rect 7331 25177 7340 25211
rect 7288 25168 7340 25177
rect 5632 25143 5684 25152
rect 5632 25109 5641 25143
rect 5641 25109 5675 25143
rect 5675 25109 5684 25143
rect 5632 25100 5684 25109
rect 7380 25143 7432 25152
rect 7380 25109 7389 25143
rect 7389 25109 7423 25143
rect 7423 25109 7432 25143
rect 7380 25100 7432 25109
rect 8944 25100 8996 25152
rect 9312 25279 9364 25288
rect 9312 25245 9321 25279
rect 9321 25245 9355 25279
rect 9355 25245 9364 25279
rect 9864 25440 9916 25492
rect 10416 25440 10468 25492
rect 18052 25440 18104 25492
rect 19708 25483 19760 25492
rect 19708 25449 19717 25483
rect 19717 25449 19751 25483
rect 19751 25449 19760 25483
rect 19708 25440 19760 25449
rect 20628 25483 20680 25492
rect 20628 25449 20637 25483
rect 20637 25449 20671 25483
rect 20671 25449 20680 25483
rect 20628 25440 20680 25449
rect 21180 25440 21232 25492
rect 12624 25415 12676 25424
rect 12624 25381 12633 25415
rect 12633 25381 12667 25415
rect 12667 25381 12676 25415
rect 12624 25372 12676 25381
rect 9312 25236 9364 25245
rect 9680 25279 9732 25288
rect 9680 25245 9689 25279
rect 9689 25245 9723 25279
rect 9723 25245 9732 25279
rect 9680 25236 9732 25245
rect 10508 25236 10560 25288
rect 12716 25236 12768 25288
rect 14280 25372 14332 25424
rect 21732 25372 21784 25424
rect 16212 25236 16264 25288
rect 11796 25168 11848 25220
rect 11888 25168 11940 25220
rect 16672 25304 16724 25356
rect 16856 25347 16908 25356
rect 16856 25313 16865 25347
rect 16865 25313 16899 25347
rect 16899 25313 16908 25347
rect 16856 25304 16908 25313
rect 19984 25304 20036 25356
rect 20536 25347 20588 25356
rect 20536 25313 20545 25347
rect 20545 25313 20579 25347
rect 20579 25313 20588 25347
rect 20536 25304 20588 25313
rect 16580 25236 16632 25288
rect 19524 25279 19576 25288
rect 19524 25245 19533 25279
rect 19533 25245 19567 25279
rect 19567 25245 19576 25279
rect 19524 25236 19576 25245
rect 16488 25168 16540 25220
rect 18420 25168 18472 25220
rect 19432 25168 19484 25220
rect 19708 25236 19760 25288
rect 20720 25279 20772 25288
rect 20720 25245 20729 25279
rect 20729 25245 20763 25279
rect 20763 25245 20772 25279
rect 21824 25304 21876 25356
rect 20720 25236 20772 25245
rect 22192 25236 22244 25288
rect 20076 25168 20128 25220
rect 21548 25168 21600 25220
rect 22100 25168 22152 25220
rect 11244 25100 11296 25152
rect 15752 25143 15804 25152
rect 15752 25109 15761 25143
rect 15761 25109 15795 25143
rect 15795 25109 15804 25143
rect 15752 25100 15804 25109
rect 17224 25100 17276 25152
rect 18052 25100 18104 25152
rect 10880 24998 10932 25050
rect 10944 24998 10996 25050
rect 11008 24998 11060 25050
rect 11072 24998 11124 25050
rect 11136 24998 11188 25050
rect 20811 24998 20863 25050
rect 20875 24998 20927 25050
rect 20939 24998 20991 25050
rect 21003 24998 21055 25050
rect 21067 24998 21119 25050
rect 7380 24896 7432 24948
rect 7656 24896 7708 24948
rect 8116 24896 8168 24948
rect 9772 24896 9824 24948
rect 11796 24896 11848 24948
rect 12900 24939 12952 24948
rect 12900 24905 12909 24939
rect 12909 24905 12943 24939
rect 12943 24905 12952 24939
rect 12900 24896 12952 24905
rect 17684 24939 17736 24948
rect 17684 24905 17693 24939
rect 17693 24905 17727 24939
rect 17727 24905 17736 24939
rect 17684 24896 17736 24905
rect 19616 24896 19668 24948
rect 22192 24939 22244 24948
rect 22192 24905 22201 24939
rect 22201 24905 22235 24939
rect 22235 24905 22244 24939
rect 22192 24896 22244 24905
rect 3148 24803 3200 24812
rect 3148 24769 3157 24803
rect 3157 24769 3191 24803
rect 3191 24769 3200 24803
rect 3148 24760 3200 24769
rect 4160 24760 4212 24812
rect 5540 24803 5592 24812
rect 5540 24769 5558 24803
rect 5558 24769 5592 24803
rect 5540 24760 5592 24769
rect 5724 24760 5776 24812
rect 7104 24803 7156 24812
rect 7104 24769 7113 24803
rect 7113 24769 7147 24803
rect 7147 24769 7156 24803
rect 7104 24760 7156 24769
rect 7196 24692 7248 24744
rect 8116 24803 8168 24812
rect 8116 24769 8125 24803
rect 8125 24769 8159 24803
rect 8159 24769 8168 24803
rect 8116 24760 8168 24769
rect 9588 24828 9640 24880
rect 15108 24828 15160 24880
rect 8576 24760 8628 24812
rect 8760 24760 8812 24812
rect 9036 24803 9088 24812
rect 9036 24769 9045 24803
rect 9045 24769 9079 24803
rect 9079 24769 9088 24803
rect 9036 24760 9088 24769
rect 9220 24803 9272 24812
rect 9220 24769 9227 24803
rect 9227 24769 9272 24803
rect 9220 24760 9272 24769
rect 9496 24803 9548 24812
rect 9496 24769 9510 24803
rect 9510 24769 9544 24803
rect 9544 24769 9548 24803
rect 10416 24803 10468 24812
rect 9496 24760 9548 24769
rect 10416 24769 10425 24803
rect 10425 24769 10459 24803
rect 10459 24769 10468 24803
rect 10416 24760 10468 24769
rect 10508 24803 10560 24812
rect 10508 24769 10517 24803
rect 10517 24769 10551 24803
rect 10551 24769 10560 24803
rect 10508 24760 10560 24769
rect 10784 24760 10836 24812
rect 11612 24760 11664 24812
rect 10324 24692 10376 24744
rect 1492 24667 1544 24676
rect 1492 24633 1501 24667
rect 1501 24633 1535 24667
rect 1535 24633 1544 24667
rect 1492 24624 1544 24633
rect 10692 24624 10744 24676
rect 5816 24556 5868 24608
rect 7472 24556 7524 24608
rect 12624 24760 12676 24812
rect 14004 24803 14056 24812
rect 14004 24769 14022 24803
rect 14022 24769 14056 24803
rect 14280 24803 14332 24812
rect 14004 24760 14056 24769
rect 14280 24769 14289 24803
rect 14289 24769 14323 24803
rect 14323 24769 14332 24803
rect 14280 24760 14332 24769
rect 14372 24760 14424 24812
rect 14832 24760 14884 24812
rect 22008 24828 22060 24880
rect 16764 24760 16816 24812
rect 18880 24803 18932 24812
rect 11980 24692 12032 24744
rect 12072 24624 12124 24676
rect 13084 24692 13136 24744
rect 15476 24692 15528 24744
rect 16212 24692 16264 24744
rect 18880 24769 18889 24803
rect 18889 24769 18923 24803
rect 18923 24769 18932 24803
rect 18880 24760 18932 24769
rect 19156 24692 19208 24744
rect 19892 24760 19944 24812
rect 20628 24760 20680 24812
rect 20720 24692 20772 24744
rect 16396 24624 16448 24676
rect 17684 24624 17736 24676
rect 21456 24692 21508 24744
rect 21916 24692 21968 24744
rect 22744 24624 22796 24676
rect 15292 24556 15344 24608
rect 16580 24556 16632 24608
rect 17776 24556 17828 24608
rect 18604 24556 18656 24608
rect 19984 24556 20036 24608
rect 21088 24556 21140 24608
rect 23756 24556 23808 24608
rect 5915 24454 5967 24506
rect 5979 24454 6031 24506
rect 6043 24454 6095 24506
rect 6107 24454 6159 24506
rect 6171 24454 6223 24506
rect 15846 24454 15898 24506
rect 15910 24454 15962 24506
rect 15974 24454 16026 24506
rect 16038 24454 16090 24506
rect 16102 24454 16154 24506
rect 25776 24454 25828 24506
rect 25840 24454 25892 24506
rect 25904 24454 25956 24506
rect 25968 24454 26020 24506
rect 26032 24454 26084 24506
rect 4436 24352 4488 24404
rect 4712 24352 4764 24404
rect 5540 24352 5592 24404
rect 7104 24352 7156 24404
rect 8576 24352 8628 24404
rect 9680 24352 9732 24404
rect 6092 24284 6144 24336
rect 3148 24216 3200 24268
rect 3792 24191 3844 24200
rect 1492 24055 1544 24064
rect 1492 24021 1501 24055
rect 1501 24021 1535 24055
rect 1535 24021 1544 24055
rect 1492 24012 1544 24021
rect 3792 24157 3801 24191
rect 3801 24157 3835 24191
rect 3835 24157 3844 24191
rect 3792 24148 3844 24157
rect 6184 24259 6236 24268
rect 6184 24225 6193 24259
rect 6193 24225 6227 24259
rect 6227 24225 6236 24259
rect 6184 24216 6236 24225
rect 5172 24148 5224 24200
rect 5816 24148 5868 24200
rect 6092 24191 6144 24200
rect 6092 24157 6101 24191
rect 6101 24157 6135 24191
rect 6135 24157 6144 24191
rect 6092 24148 6144 24157
rect 6736 24216 6788 24268
rect 7380 24216 7432 24268
rect 8208 24216 8260 24268
rect 6552 24148 6604 24200
rect 7564 24148 7616 24200
rect 7656 24148 7708 24200
rect 8944 24191 8996 24200
rect 4068 24123 4120 24132
rect 4068 24089 4102 24123
rect 4102 24089 4120 24123
rect 4068 24080 4120 24089
rect 4344 24012 4396 24064
rect 6276 24012 6328 24064
rect 7196 24080 7248 24132
rect 7932 24080 7984 24132
rect 8944 24157 8953 24191
rect 8953 24157 8987 24191
rect 8987 24157 8996 24191
rect 8944 24148 8996 24157
rect 9128 24148 9180 24200
rect 9864 24148 9916 24200
rect 10140 24191 10192 24200
rect 10140 24157 10149 24191
rect 10149 24157 10183 24191
rect 10183 24157 10192 24191
rect 10140 24148 10192 24157
rect 19708 24352 19760 24404
rect 19800 24352 19852 24404
rect 11244 24284 11296 24336
rect 12256 24284 12308 24336
rect 14372 24284 14424 24336
rect 8576 24080 8628 24132
rect 9772 24080 9824 24132
rect 7380 24055 7432 24064
rect 7380 24021 7389 24055
rect 7389 24021 7423 24055
rect 7423 24021 7432 24055
rect 7380 24012 7432 24021
rect 9128 24012 9180 24064
rect 9312 24012 9364 24064
rect 11244 24148 11296 24200
rect 11428 24148 11480 24200
rect 11520 24148 11572 24200
rect 11704 24148 11756 24200
rect 10692 24080 10744 24132
rect 12348 24148 12400 24200
rect 13084 24191 13136 24200
rect 13084 24157 13093 24191
rect 13093 24157 13127 24191
rect 13127 24157 13136 24191
rect 13084 24148 13136 24157
rect 13544 24148 13596 24200
rect 14556 24148 14608 24200
rect 15016 24216 15068 24268
rect 15108 24191 15160 24200
rect 15108 24157 15117 24191
rect 15117 24157 15151 24191
rect 15151 24157 15160 24191
rect 15108 24148 15160 24157
rect 16580 24284 16632 24336
rect 16764 24216 16816 24268
rect 17776 24259 17828 24268
rect 17776 24225 17785 24259
rect 17785 24225 17819 24259
rect 17819 24225 17828 24259
rect 17776 24216 17828 24225
rect 19340 24284 19392 24336
rect 21916 24284 21968 24336
rect 19984 24216 20036 24268
rect 15292 24191 15344 24200
rect 15292 24157 15306 24191
rect 15306 24157 15340 24191
rect 15340 24157 15344 24191
rect 15292 24148 15344 24157
rect 15752 24148 15804 24200
rect 16120 24148 16172 24200
rect 16580 24191 16632 24200
rect 15384 24080 15436 24132
rect 16580 24157 16589 24191
rect 16589 24157 16623 24191
rect 16623 24157 16632 24191
rect 16580 24148 16632 24157
rect 17132 24148 17184 24200
rect 18788 24148 18840 24200
rect 19156 24148 19208 24200
rect 19616 24148 19668 24200
rect 20536 24216 20588 24268
rect 21088 24259 21140 24268
rect 21088 24225 21097 24259
rect 21097 24225 21131 24259
rect 21131 24225 21140 24259
rect 21088 24216 21140 24225
rect 20628 24148 20680 24200
rect 21272 24148 21324 24200
rect 19432 24080 19484 24132
rect 20536 24080 20588 24132
rect 22008 24123 22060 24132
rect 12624 24055 12676 24064
rect 12624 24021 12633 24055
rect 12633 24021 12667 24055
rect 12667 24021 12676 24055
rect 12624 24012 12676 24021
rect 14740 24012 14792 24064
rect 16672 24012 16724 24064
rect 18788 24012 18840 24064
rect 19340 24055 19392 24064
rect 19340 24021 19349 24055
rect 19349 24021 19383 24055
rect 19383 24021 19392 24055
rect 19340 24012 19392 24021
rect 19708 24012 19760 24064
rect 20628 24012 20680 24064
rect 21364 24055 21416 24064
rect 21364 24021 21373 24055
rect 21373 24021 21407 24055
rect 21407 24021 21416 24055
rect 21364 24012 21416 24021
rect 22008 24089 22017 24123
rect 22017 24089 22051 24123
rect 22051 24089 22060 24123
rect 22008 24080 22060 24089
rect 22100 24080 22152 24132
rect 22928 24148 22980 24200
rect 23756 24191 23808 24200
rect 23756 24157 23765 24191
rect 23765 24157 23799 24191
rect 23799 24157 23808 24191
rect 23756 24148 23808 24157
rect 29920 24148 29972 24200
rect 22376 24055 22428 24064
rect 22376 24021 22385 24055
rect 22385 24021 22419 24055
rect 22419 24021 22428 24055
rect 22376 24012 22428 24021
rect 23112 24012 23164 24064
rect 30012 24055 30064 24064
rect 30012 24021 30021 24055
rect 30021 24021 30055 24055
rect 30055 24021 30064 24055
rect 30012 24012 30064 24021
rect 10880 23910 10932 23962
rect 10944 23910 10996 23962
rect 11008 23910 11060 23962
rect 11072 23910 11124 23962
rect 11136 23910 11188 23962
rect 20811 23910 20863 23962
rect 20875 23910 20927 23962
rect 20939 23910 20991 23962
rect 21003 23910 21055 23962
rect 21067 23910 21119 23962
rect 4068 23808 4120 23860
rect 3792 23740 3844 23792
rect 4252 23672 4304 23724
rect 1400 23647 1452 23656
rect 1400 23613 1409 23647
rect 1409 23613 1443 23647
rect 1443 23613 1452 23647
rect 1400 23604 1452 23613
rect 2136 23604 2188 23656
rect 4344 23647 4396 23656
rect 4344 23613 4353 23647
rect 4353 23613 4387 23647
rect 4387 23613 4396 23647
rect 4344 23604 4396 23613
rect 4896 23672 4948 23724
rect 6552 23808 6604 23860
rect 6736 23808 6788 23860
rect 6276 23740 6328 23792
rect 6368 23715 6420 23724
rect 6368 23681 6377 23715
rect 6377 23681 6411 23715
rect 6411 23681 6420 23715
rect 6368 23672 6420 23681
rect 6920 23740 6972 23792
rect 7012 23740 7064 23792
rect 10600 23808 10652 23860
rect 14372 23808 14424 23860
rect 14832 23808 14884 23860
rect 15292 23808 15344 23860
rect 16120 23851 16172 23860
rect 16120 23817 16129 23851
rect 16129 23817 16163 23851
rect 16163 23817 16172 23851
rect 16120 23808 16172 23817
rect 18604 23851 18656 23860
rect 18604 23817 18613 23851
rect 18613 23817 18647 23851
rect 18647 23817 18656 23851
rect 18604 23808 18656 23817
rect 19708 23808 19760 23860
rect 29920 23851 29972 23860
rect 29920 23817 29929 23851
rect 29929 23817 29963 23851
rect 29963 23817 29972 23851
rect 29920 23808 29972 23817
rect 9128 23740 9180 23792
rect 10508 23740 10560 23792
rect 11888 23740 11940 23792
rect 7104 23536 7156 23588
rect 4804 23468 4856 23520
rect 5080 23468 5132 23520
rect 7012 23468 7064 23520
rect 7196 23511 7248 23520
rect 7196 23477 7205 23511
rect 7205 23477 7239 23511
rect 7239 23477 7248 23511
rect 7196 23468 7248 23477
rect 8024 23468 8076 23520
rect 8760 23672 8812 23724
rect 9036 23715 9088 23724
rect 9036 23681 9045 23715
rect 9045 23681 9079 23715
rect 9079 23681 9088 23715
rect 9036 23672 9088 23681
rect 8944 23604 8996 23656
rect 10876 23672 10928 23724
rect 11428 23672 11480 23724
rect 9496 23604 9548 23656
rect 10600 23604 10652 23656
rect 11796 23715 11848 23724
rect 11796 23681 11805 23715
rect 11805 23681 11839 23715
rect 11839 23681 11848 23715
rect 12256 23740 12308 23792
rect 12624 23740 12676 23792
rect 14556 23783 14608 23792
rect 14556 23749 14565 23783
rect 14565 23749 14599 23783
rect 14599 23749 14608 23783
rect 14556 23740 14608 23749
rect 16488 23740 16540 23792
rect 17408 23740 17460 23792
rect 11796 23672 11848 23681
rect 12716 23715 12768 23724
rect 12256 23604 12308 23656
rect 12716 23681 12725 23715
rect 12725 23681 12759 23715
rect 12759 23681 12768 23715
rect 12716 23672 12768 23681
rect 13544 23672 13596 23724
rect 16672 23715 16724 23724
rect 16672 23681 16681 23715
rect 16681 23681 16715 23715
rect 16715 23681 16724 23715
rect 16672 23672 16724 23681
rect 17040 23672 17092 23724
rect 18512 23715 18564 23724
rect 18512 23681 18521 23715
rect 18521 23681 18555 23715
rect 18555 23681 18564 23715
rect 18512 23672 18564 23681
rect 19800 23672 19852 23724
rect 19892 23672 19944 23724
rect 20260 23672 20312 23724
rect 20533 23715 20585 23724
rect 20533 23681 20542 23715
rect 20542 23681 20576 23715
rect 20576 23681 20585 23715
rect 20533 23672 20585 23681
rect 15108 23604 15160 23656
rect 15660 23647 15712 23656
rect 15660 23613 15669 23647
rect 15669 23613 15703 23647
rect 15703 23613 15712 23647
rect 15660 23604 15712 23613
rect 17224 23647 17276 23656
rect 17224 23613 17233 23647
rect 17233 23613 17267 23647
rect 17267 23613 17276 23647
rect 17224 23604 17276 23613
rect 17408 23647 17460 23656
rect 17408 23613 17417 23647
rect 17417 23613 17451 23647
rect 17451 23613 17460 23647
rect 17408 23604 17460 23613
rect 18604 23604 18656 23656
rect 19524 23604 19576 23656
rect 19616 23604 19668 23656
rect 8484 23536 8536 23588
rect 9220 23536 9272 23588
rect 16856 23536 16908 23588
rect 20260 23536 20312 23588
rect 22376 23672 22428 23724
rect 30104 23715 30156 23724
rect 22468 23647 22520 23656
rect 22468 23613 22477 23647
rect 22477 23613 22511 23647
rect 22511 23613 22520 23647
rect 22468 23604 22520 23613
rect 22376 23536 22428 23588
rect 30104 23681 30113 23715
rect 30113 23681 30147 23715
rect 30147 23681 30156 23715
rect 30104 23672 30156 23681
rect 8392 23468 8444 23520
rect 9036 23468 9088 23520
rect 9588 23468 9640 23520
rect 9864 23468 9916 23520
rect 10784 23468 10836 23520
rect 12532 23468 12584 23520
rect 16304 23468 16356 23520
rect 16948 23468 17000 23520
rect 17224 23468 17276 23520
rect 18144 23511 18196 23520
rect 18144 23477 18153 23511
rect 18153 23477 18187 23511
rect 18187 23477 18196 23511
rect 18144 23468 18196 23477
rect 20168 23511 20220 23520
rect 20168 23477 20177 23511
rect 20177 23477 20211 23511
rect 20211 23477 20220 23511
rect 20168 23468 20220 23477
rect 20720 23468 20772 23520
rect 21548 23468 21600 23520
rect 22928 23468 22980 23520
rect 5915 23366 5967 23418
rect 5979 23366 6031 23418
rect 6043 23366 6095 23418
rect 6107 23366 6159 23418
rect 6171 23366 6223 23418
rect 15846 23366 15898 23418
rect 15910 23366 15962 23418
rect 15974 23366 16026 23418
rect 16038 23366 16090 23418
rect 16102 23366 16154 23418
rect 25776 23366 25828 23418
rect 25840 23366 25892 23418
rect 25904 23366 25956 23418
rect 25968 23366 26020 23418
rect 26032 23366 26084 23418
rect 7380 23264 7432 23316
rect 8392 23264 8444 23316
rect 8944 23264 8996 23316
rect 10876 23264 10928 23316
rect 13544 23307 13596 23316
rect 13544 23273 13553 23307
rect 13553 23273 13587 23307
rect 13587 23273 13596 23307
rect 13544 23264 13596 23273
rect 15384 23264 15436 23316
rect 17408 23264 17460 23316
rect 18512 23264 18564 23316
rect 20168 23264 20220 23316
rect 21180 23264 21232 23316
rect 6552 23196 6604 23248
rect 7472 23196 7524 23248
rect 4436 23128 4488 23180
rect 4804 23128 4856 23180
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 4896 23103 4948 23112
rect 1584 22967 1636 22976
rect 1584 22933 1593 22967
rect 1593 22933 1627 22967
rect 1627 22933 1636 22967
rect 1584 22924 1636 22933
rect 4160 22967 4212 22976
rect 4160 22933 4169 22967
rect 4169 22933 4203 22967
rect 4203 22933 4212 22967
rect 4160 22924 4212 22933
rect 4528 22924 4580 22976
rect 4896 23069 4905 23103
rect 4905 23069 4939 23103
rect 4939 23069 4948 23103
rect 4896 23060 4948 23069
rect 7380 23103 7432 23112
rect 7380 23069 7389 23103
rect 7389 23069 7423 23103
rect 7423 23069 7432 23103
rect 7380 23060 7432 23069
rect 7748 23196 7800 23248
rect 8208 23196 8260 23248
rect 15016 23196 15068 23248
rect 18052 23196 18104 23248
rect 19156 23196 19208 23248
rect 22560 23264 22612 23316
rect 7656 23171 7708 23180
rect 7656 23137 7665 23171
rect 7665 23137 7699 23171
rect 7699 23137 7708 23171
rect 7656 23128 7708 23137
rect 5632 23035 5684 23044
rect 5632 23001 5666 23035
rect 5666 23001 5684 23035
rect 5632 22992 5684 23001
rect 5724 22992 5776 23044
rect 5540 22924 5592 22976
rect 7012 22924 7064 22976
rect 8392 23060 8444 23112
rect 8484 23060 8536 23112
rect 9036 23060 9088 23112
rect 9864 23060 9916 23112
rect 11520 23060 11572 23112
rect 14740 23103 14792 23112
rect 14740 23069 14749 23103
rect 14749 23069 14783 23103
rect 14783 23069 14792 23103
rect 14740 23060 14792 23069
rect 14832 23103 14884 23112
rect 14832 23069 14841 23103
rect 14841 23069 14875 23103
rect 14875 23069 14884 23103
rect 14832 23060 14884 23069
rect 15016 23103 15068 23112
rect 15016 23069 15025 23103
rect 15025 23069 15059 23103
rect 15059 23069 15068 23103
rect 16764 23128 16816 23180
rect 18696 23128 18748 23180
rect 15016 23060 15068 23069
rect 16396 23060 16448 23112
rect 18052 23060 18104 23112
rect 12532 22992 12584 23044
rect 17408 22992 17460 23044
rect 19156 23060 19208 23112
rect 19524 23103 19576 23112
rect 19524 23069 19533 23103
rect 19533 23069 19567 23103
rect 19567 23069 19576 23103
rect 19524 23060 19576 23069
rect 18420 22992 18472 23044
rect 18604 22992 18656 23044
rect 20628 23060 20680 23112
rect 21364 23060 21416 23112
rect 22468 23060 22520 23112
rect 22928 23103 22980 23112
rect 22928 23069 22937 23103
rect 22937 23069 22971 23103
rect 22971 23069 22980 23103
rect 22928 23060 22980 23069
rect 23112 23103 23164 23112
rect 23112 23069 23121 23103
rect 23121 23069 23155 23103
rect 23155 23069 23164 23103
rect 23112 23060 23164 23069
rect 22744 23035 22796 23044
rect 22744 23001 22753 23035
rect 22753 23001 22787 23035
rect 22787 23001 22796 23035
rect 22744 22992 22796 23001
rect 16948 22924 17000 22976
rect 18880 22924 18932 22976
rect 10880 22822 10932 22874
rect 10944 22822 10996 22874
rect 11008 22822 11060 22874
rect 11072 22822 11124 22874
rect 11136 22822 11188 22874
rect 20811 22822 20863 22874
rect 20875 22822 20927 22874
rect 20939 22822 20991 22874
rect 21003 22822 21055 22874
rect 21067 22822 21119 22874
rect 4528 22720 4580 22772
rect 4160 22652 4212 22704
rect 5632 22720 5684 22772
rect 6276 22652 6328 22704
rect 2044 22627 2096 22636
rect 2044 22593 2053 22627
rect 2053 22593 2087 22627
rect 2087 22593 2096 22627
rect 2044 22584 2096 22593
rect 2780 22584 2832 22636
rect 3792 22584 3844 22636
rect 6552 22627 6604 22636
rect 6552 22593 6561 22627
rect 6561 22593 6595 22627
rect 6595 22593 6604 22627
rect 6552 22584 6604 22593
rect 7104 22720 7156 22772
rect 8116 22720 8168 22772
rect 9128 22763 9180 22772
rect 9128 22729 9137 22763
rect 9137 22729 9171 22763
rect 9171 22729 9180 22763
rect 9128 22720 9180 22729
rect 10416 22720 10468 22772
rect 11428 22720 11480 22772
rect 12072 22720 12124 22772
rect 7012 22584 7064 22636
rect 8300 22652 8352 22704
rect 9036 22652 9088 22704
rect 11152 22652 11204 22704
rect 11336 22652 11388 22704
rect 8024 22627 8076 22636
rect 8024 22593 8058 22627
rect 8058 22593 8076 22627
rect 8024 22584 8076 22593
rect 9128 22584 9180 22636
rect 9404 22584 9456 22636
rect 9956 22584 10008 22636
rect 10416 22584 10468 22636
rect 10692 22627 10744 22636
rect 10692 22593 10710 22627
rect 10710 22593 10744 22627
rect 10692 22584 10744 22593
rect 10876 22584 10928 22636
rect 11428 22584 11480 22636
rect 11888 22652 11940 22704
rect 12808 22720 12860 22772
rect 15660 22720 15712 22772
rect 16580 22720 16632 22772
rect 17408 22720 17460 22772
rect 20352 22720 20404 22772
rect 22468 22720 22520 22772
rect 12532 22652 12584 22704
rect 16396 22652 16448 22704
rect 19892 22652 19944 22704
rect 20996 22695 21048 22704
rect 20996 22661 21005 22695
rect 21005 22661 21039 22695
rect 21039 22661 21048 22695
rect 20996 22652 21048 22661
rect 12716 22627 12768 22636
rect 2872 22516 2924 22568
rect 6368 22516 6420 22568
rect 12716 22593 12725 22627
rect 12725 22593 12759 22627
rect 12759 22593 12768 22627
rect 12716 22584 12768 22593
rect 3976 22448 4028 22500
rect 6552 22448 6604 22500
rect 1952 22380 2004 22432
rect 4252 22380 4304 22432
rect 5816 22380 5868 22432
rect 12164 22516 12216 22568
rect 11520 22448 11572 22500
rect 12256 22423 12308 22432
rect 12256 22389 12265 22423
rect 12265 22389 12299 22423
rect 12299 22389 12308 22423
rect 12256 22380 12308 22389
rect 13728 22380 13780 22432
rect 16488 22584 16540 22636
rect 16764 22584 16816 22636
rect 19708 22584 19760 22636
rect 21180 22627 21232 22636
rect 21180 22593 21189 22627
rect 21189 22593 21223 22627
rect 21223 22593 21232 22627
rect 21180 22584 21232 22593
rect 23020 22584 23072 22636
rect 30196 22584 30248 22636
rect 15568 22516 15620 22568
rect 16396 22516 16448 22568
rect 15016 22448 15068 22500
rect 16212 22448 16264 22500
rect 16488 22448 16540 22500
rect 16856 22448 16908 22500
rect 15108 22380 15160 22432
rect 16672 22380 16724 22432
rect 18052 22516 18104 22568
rect 18880 22516 18932 22568
rect 22376 22516 22428 22568
rect 30104 22516 30156 22568
rect 19524 22448 19576 22500
rect 19432 22380 19484 22432
rect 19616 22423 19668 22432
rect 19616 22389 19625 22423
rect 19625 22389 19659 22423
rect 19659 22389 19668 22423
rect 19616 22380 19668 22389
rect 30012 22423 30064 22432
rect 30012 22389 30021 22423
rect 30021 22389 30055 22423
rect 30055 22389 30064 22423
rect 30012 22380 30064 22389
rect 5915 22278 5967 22330
rect 5979 22278 6031 22330
rect 6043 22278 6095 22330
rect 6107 22278 6159 22330
rect 6171 22278 6223 22330
rect 15846 22278 15898 22330
rect 15910 22278 15962 22330
rect 15974 22278 16026 22330
rect 16038 22278 16090 22330
rect 16102 22278 16154 22330
rect 25776 22278 25828 22330
rect 25840 22278 25892 22330
rect 25904 22278 25956 22330
rect 25968 22278 26020 22330
rect 26032 22278 26084 22330
rect 10692 22176 10744 22228
rect 8208 22108 8260 22160
rect 9404 22108 9456 22160
rect 4804 22040 4856 22092
rect 5724 22040 5776 22092
rect 8944 22083 8996 22092
rect 8944 22049 8953 22083
rect 8953 22049 8987 22083
rect 8987 22049 8996 22083
rect 8944 22040 8996 22049
rect 9496 22040 9548 22092
rect 11888 22083 11940 22092
rect 11888 22049 11897 22083
rect 11897 22049 11931 22083
rect 11931 22049 11940 22083
rect 11888 22040 11940 22049
rect 12532 22040 12584 22092
rect 1676 21972 1728 22024
rect 3700 21972 3752 22024
rect 5540 22015 5592 22024
rect 5540 21981 5549 22015
rect 5549 21981 5583 22015
rect 5583 21981 5592 22015
rect 5540 21972 5592 21981
rect 7196 21972 7248 22024
rect 9588 21972 9640 22024
rect 10324 21972 10376 22024
rect 10784 22015 10836 22024
rect 2412 21904 2464 21956
rect 6736 21904 6788 21956
rect 8300 21947 8352 21956
rect 8300 21913 8309 21947
rect 8309 21913 8343 21947
rect 8343 21913 8352 21947
rect 8300 21904 8352 21913
rect 9220 21904 9272 21956
rect 10784 21981 10793 22015
rect 10793 21981 10827 22015
rect 10827 21981 10836 22015
rect 10784 21972 10836 21981
rect 11244 21972 11296 22024
rect 11612 22015 11664 22024
rect 11612 21981 11621 22015
rect 11621 21981 11655 22015
rect 11655 21981 11664 22015
rect 11612 21972 11664 21981
rect 11980 22015 12032 22024
rect 2964 21836 3016 21888
rect 7012 21836 7064 21888
rect 7840 21836 7892 21888
rect 11980 21981 11989 22015
rect 11989 21981 12023 22015
rect 12023 21981 12032 22015
rect 11980 21972 12032 21981
rect 13728 21972 13780 22024
rect 15200 21972 15252 22024
rect 15384 22108 15436 22160
rect 17040 22176 17092 22228
rect 18696 22176 18748 22228
rect 19064 22176 19116 22228
rect 21456 22176 21508 22228
rect 19432 22108 19484 22160
rect 15660 22083 15712 22092
rect 15660 22049 15669 22083
rect 15669 22049 15703 22083
rect 15703 22049 15712 22083
rect 15660 22040 15712 22049
rect 18144 22083 18196 22092
rect 18144 22049 18153 22083
rect 18153 22049 18187 22083
rect 18187 22049 18196 22083
rect 18144 22040 18196 22049
rect 15752 22015 15804 22024
rect 15752 21981 15766 22015
rect 15766 21981 15800 22015
rect 15800 21981 15804 22015
rect 15752 21972 15804 21981
rect 16488 21972 16540 22024
rect 16672 22015 16724 22024
rect 16672 21981 16681 22015
rect 16681 21981 16715 22015
rect 16715 21981 16724 22015
rect 16672 21972 16724 21981
rect 16856 22015 16908 22024
rect 16856 21981 16865 22015
rect 16865 21981 16899 22015
rect 16899 21981 16908 22015
rect 16856 21972 16908 21981
rect 17040 21972 17092 22024
rect 15568 21947 15620 21956
rect 15568 21913 15577 21947
rect 15577 21913 15611 21947
rect 15611 21913 15620 21947
rect 15568 21904 15620 21913
rect 15844 21904 15896 21956
rect 17316 21972 17368 22024
rect 17684 21972 17736 22024
rect 18052 21972 18104 22024
rect 19340 22040 19392 22092
rect 20996 22040 21048 22092
rect 22008 22040 22060 22092
rect 22376 22083 22428 22092
rect 22376 22049 22385 22083
rect 22385 22049 22419 22083
rect 22419 22049 22428 22083
rect 22376 22040 22428 22049
rect 20444 21972 20496 22024
rect 21640 21972 21692 22024
rect 22468 21972 22520 22024
rect 18052 21879 18104 21888
rect 18052 21845 18061 21879
rect 18061 21845 18095 21879
rect 18095 21845 18104 21879
rect 18052 21836 18104 21845
rect 18144 21836 18196 21888
rect 19064 21836 19116 21888
rect 21180 21904 21232 21956
rect 23020 21904 23072 21956
rect 21824 21879 21876 21888
rect 21824 21845 21833 21879
rect 21833 21845 21867 21879
rect 21867 21845 21876 21879
rect 21824 21836 21876 21845
rect 10880 21734 10932 21786
rect 10944 21734 10996 21786
rect 11008 21734 11060 21786
rect 11072 21734 11124 21786
rect 11136 21734 11188 21786
rect 20811 21734 20863 21786
rect 20875 21734 20927 21786
rect 20939 21734 20991 21786
rect 21003 21734 21055 21786
rect 21067 21734 21119 21786
rect 4436 21632 4488 21684
rect 7380 21632 7432 21684
rect 12808 21632 12860 21684
rect 15568 21632 15620 21684
rect 16672 21632 16724 21684
rect 19432 21632 19484 21684
rect 7932 21607 7984 21616
rect 7932 21573 7941 21607
rect 7941 21573 7975 21607
rect 7975 21573 7984 21607
rect 7932 21564 7984 21573
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 2228 21496 2280 21548
rect 3240 21496 3292 21548
rect 5540 21496 5592 21548
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 5816 21496 5868 21505
rect 6276 21496 6328 21548
rect 6920 21539 6972 21548
rect 6920 21505 6929 21539
rect 6929 21505 6963 21539
rect 6963 21505 6972 21539
rect 6920 21496 6972 21505
rect 7196 21539 7248 21548
rect 7196 21505 7205 21539
rect 7205 21505 7239 21539
rect 7239 21505 7248 21539
rect 9588 21564 9640 21616
rect 10416 21564 10468 21616
rect 12256 21564 12308 21616
rect 15292 21564 15344 21616
rect 7196 21496 7248 21505
rect 8484 21496 8536 21548
rect 9220 21496 9272 21548
rect 10692 21496 10744 21548
rect 15844 21564 15896 21616
rect 17040 21564 17092 21616
rect 18604 21564 18656 21616
rect 19892 21564 19944 21616
rect 20444 21564 20496 21616
rect 21548 21564 21600 21616
rect 22008 21607 22060 21616
rect 22008 21573 22017 21607
rect 22017 21573 22051 21607
rect 22051 21573 22060 21607
rect 22008 21564 22060 21573
rect 22468 21564 22520 21616
rect 15660 21496 15712 21548
rect 17132 21496 17184 21548
rect 11520 21428 11572 21480
rect 15108 21428 15160 21480
rect 2780 21360 2832 21412
rect 8944 21360 8996 21412
rect 11244 21360 11296 21412
rect 17500 21360 17552 21412
rect 3056 21335 3108 21344
rect 3056 21301 3065 21335
rect 3065 21301 3099 21335
rect 3099 21301 3108 21335
rect 3056 21292 3108 21301
rect 6460 21292 6512 21344
rect 7932 21292 7984 21344
rect 10048 21335 10100 21344
rect 10048 21301 10057 21335
rect 10057 21301 10091 21335
rect 10091 21301 10100 21335
rect 10048 21292 10100 21301
rect 18052 21496 18104 21548
rect 19064 21539 19116 21548
rect 19064 21505 19073 21539
rect 19073 21505 19107 21539
rect 19107 21505 19116 21539
rect 19064 21496 19116 21505
rect 18420 21428 18472 21480
rect 18880 21428 18932 21480
rect 19340 21539 19392 21548
rect 19340 21505 19349 21539
rect 19349 21505 19383 21539
rect 19383 21505 19392 21539
rect 19616 21539 19668 21548
rect 19340 21496 19392 21505
rect 19616 21505 19625 21539
rect 19625 21505 19659 21539
rect 19659 21505 19668 21539
rect 19616 21496 19668 21505
rect 20536 21496 20588 21548
rect 18696 21360 18748 21412
rect 20444 21428 20496 21480
rect 19892 21292 19944 21344
rect 20352 21292 20404 21344
rect 5915 21190 5967 21242
rect 5979 21190 6031 21242
rect 6043 21190 6095 21242
rect 6107 21190 6159 21242
rect 6171 21190 6223 21242
rect 15846 21190 15898 21242
rect 15910 21190 15962 21242
rect 15974 21190 16026 21242
rect 16038 21190 16090 21242
rect 16102 21190 16154 21242
rect 25776 21190 25828 21242
rect 25840 21190 25892 21242
rect 25904 21190 25956 21242
rect 25968 21190 26020 21242
rect 26032 21190 26084 21242
rect 2228 21131 2280 21140
rect 2228 21097 2237 21131
rect 2237 21097 2271 21131
rect 2271 21097 2280 21131
rect 2228 21088 2280 21097
rect 6184 21020 6236 21072
rect 6552 21088 6604 21140
rect 6736 21131 6788 21140
rect 6736 21097 6745 21131
rect 6745 21097 6779 21131
rect 6779 21097 6788 21131
rect 6736 21088 6788 21097
rect 8484 21088 8536 21140
rect 10416 21131 10468 21140
rect 10416 21097 10425 21131
rect 10425 21097 10459 21131
rect 10459 21097 10468 21131
rect 10416 21088 10468 21097
rect 11336 21088 11388 21140
rect 13544 21088 13596 21140
rect 7656 21020 7708 21072
rect 12624 21020 12676 21072
rect 16580 21020 16632 21072
rect 19340 21088 19392 21140
rect 19708 21131 19760 21140
rect 19708 21097 19717 21131
rect 19717 21097 19751 21131
rect 19751 21097 19760 21131
rect 19708 21088 19760 21097
rect 20536 21131 20588 21140
rect 20536 21097 20545 21131
rect 20545 21097 20579 21131
rect 20579 21097 20588 21131
rect 20536 21088 20588 21097
rect 1492 20927 1544 20936
rect 1492 20893 1501 20927
rect 1501 20893 1535 20927
rect 1535 20893 1544 20927
rect 1492 20884 1544 20893
rect 1584 20884 1636 20936
rect 1860 20927 1912 20936
rect 1860 20893 1869 20927
rect 1869 20893 1903 20927
rect 1903 20893 1912 20927
rect 1860 20884 1912 20893
rect 3056 20927 3108 20936
rect 3056 20893 3065 20927
rect 3065 20893 3099 20927
rect 3099 20893 3108 20927
rect 3056 20884 3108 20893
rect 2964 20816 3016 20868
rect 4160 20884 4212 20936
rect 6368 20995 6420 21004
rect 6368 20961 6377 20995
rect 6377 20961 6411 20995
rect 6411 20961 6420 20995
rect 6368 20952 6420 20961
rect 9312 20952 9364 21004
rect 15016 20995 15068 21004
rect 15016 20961 15025 20995
rect 15025 20961 15059 20995
rect 15059 20961 15068 20995
rect 15016 20952 15068 20961
rect 16856 20952 16908 21004
rect 19524 21020 19576 21072
rect 7012 20884 7064 20936
rect 12900 20884 12952 20936
rect 16580 20884 16632 20936
rect 1584 20748 1636 20800
rect 3148 20791 3200 20800
rect 3148 20757 3157 20791
rect 3157 20757 3191 20791
rect 3191 20757 3200 20791
rect 3148 20748 3200 20757
rect 4436 20791 4488 20800
rect 4436 20757 4445 20791
rect 4445 20757 4479 20791
rect 4479 20757 4488 20791
rect 4436 20748 4488 20757
rect 6828 20816 6880 20868
rect 7288 20816 7340 20868
rect 8484 20816 8536 20868
rect 9036 20816 9088 20868
rect 9312 20859 9364 20868
rect 9312 20825 9321 20859
rect 9321 20825 9355 20859
rect 9355 20825 9364 20859
rect 9312 20816 9364 20825
rect 10600 20816 10652 20868
rect 11336 20816 11388 20868
rect 13452 20816 13504 20868
rect 13544 20859 13596 20868
rect 13544 20825 13553 20859
rect 13553 20825 13587 20859
rect 13587 20825 13596 20859
rect 13544 20816 13596 20825
rect 17500 20816 17552 20868
rect 18880 20952 18932 21004
rect 18696 20884 18748 20936
rect 20260 20952 20312 21004
rect 20720 20952 20772 21004
rect 19800 20927 19852 20936
rect 19800 20893 19809 20927
rect 19809 20893 19843 20927
rect 19843 20893 19852 20927
rect 19800 20884 19852 20893
rect 22376 20884 22428 20936
rect 29828 20927 29880 20936
rect 29828 20893 29837 20927
rect 29837 20893 29871 20927
rect 29871 20893 29880 20927
rect 29828 20884 29880 20893
rect 19616 20816 19668 20868
rect 20536 20816 20588 20868
rect 7380 20748 7432 20800
rect 9680 20748 9732 20800
rect 12992 20748 13044 20800
rect 15568 20791 15620 20800
rect 15568 20757 15577 20791
rect 15577 20757 15611 20791
rect 15611 20757 15620 20791
rect 15568 20748 15620 20757
rect 16764 20791 16816 20800
rect 16764 20757 16773 20791
rect 16773 20757 16807 20791
rect 16807 20757 16816 20791
rect 17132 20791 17184 20800
rect 16764 20748 16816 20757
rect 17132 20757 17141 20791
rect 17141 20757 17175 20791
rect 17175 20757 17184 20791
rect 17132 20748 17184 20757
rect 18052 20748 18104 20800
rect 18880 20748 18932 20800
rect 21824 20748 21876 20800
rect 22192 20748 22244 20800
rect 30012 20791 30064 20800
rect 30012 20757 30021 20791
rect 30021 20757 30055 20791
rect 30055 20757 30064 20791
rect 30012 20748 30064 20757
rect 10880 20646 10932 20698
rect 10944 20646 10996 20698
rect 11008 20646 11060 20698
rect 11072 20646 11124 20698
rect 11136 20646 11188 20698
rect 20811 20646 20863 20698
rect 20875 20646 20927 20698
rect 20939 20646 20991 20698
rect 21003 20646 21055 20698
rect 21067 20646 21119 20698
rect 2412 20587 2464 20596
rect 2412 20553 2421 20587
rect 2421 20553 2455 20587
rect 2455 20553 2464 20587
rect 2412 20544 2464 20553
rect 5540 20544 5592 20596
rect 8484 20544 8536 20596
rect 8852 20544 8904 20596
rect 10140 20544 10192 20596
rect 14648 20544 14700 20596
rect 15384 20587 15436 20596
rect 15384 20553 15393 20587
rect 15393 20553 15427 20587
rect 15427 20553 15436 20587
rect 15384 20544 15436 20553
rect 15568 20544 15620 20596
rect 16764 20544 16816 20596
rect 19432 20544 19484 20596
rect 20628 20544 20680 20596
rect 22284 20587 22336 20596
rect 22284 20553 22293 20587
rect 22293 20553 22327 20587
rect 22327 20553 22336 20587
rect 22284 20544 22336 20553
rect 29828 20544 29880 20596
rect 1492 20408 1544 20460
rect 4436 20476 4488 20528
rect 6368 20476 6420 20528
rect 2964 20408 3016 20460
rect 3056 20451 3108 20460
rect 3056 20417 3065 20451
rect 3065 20417 3099 20451
rect 3099 20417 3108 20451
rect 3056 20408 3108 20417
rect 4528 20408 4580 20460
rect 1584 20340 1636 20392
rect 3700 20383 3752 20392
rect 1768 20272 1820 20324
rect 3700 20349 3709 20383
rect 3709 20349 3743 20383
rect 3743 20349 3752 20383
rect 3700 20340 3752 20349
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 6552 20451 6604 20460
rect 6552 20417 6562 20451
rect 6562 20417 6596 20451
rect 6596 20417 6604 20451
rect 6736 20451 6788 20460
rect 6552 20408 6604 20417
rect 6736 20417 6745 20451
rect 6745 20417 6779 20451
rect 6779 20417 6788 20451
rect 6736 20408 6788 20417
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 9588 20476 9640 20528
rect 18144 20476 18196 20528
rect 22192 20519 22244 20528
rect 6828 20408 6880 20417
rect 8484 20451 8536 20460
rect 8484 20417 8493 20451
rect 8493 20417 8527 20451
rect 8527 20417 8536 20451
rect 8484 20408 8536 20417
rect 9036 20408 9088 20460
rect 9680 20408 9732 20460
rect 10600 20451 10652 20460
rect 6644 20340 6696 20392
rect 8760 20340 8812 20392
rect 10600 20417 10609 20451
rect 10609 20417 10643 20451
rect 10643 20417 10652 20451
rect 10600 20408 10652 20417
rect 11244 20408 11296 20460
rect 10140 20340 10192 20392
rect 11060 20340 11112 20392
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 12900 20408 12952 20460
rect 13452 20451 13504 20460
rect 13452 20417 13461 20451
rect 13461 20417 13495 20451
rect 13495 20417 13504 20451
rect 13452 20408 13504 20417
rect 13544 20408 13596 20460
rect 14556 20451 14608 20460
rect 14556 20417 14565 20451
rect 14565 20417 14599 20451
rect 14599 20417 14608 20451
rect 14556 20408 14608 20417
rect 15016 20408 15068 20460
rect 16488 20408 16540 20460
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 22192 20485 22201 20519
rect 22201 20485 22235 20519
rect 22235 20485 22244 20519
rect 22192 20476 22244 20485
rect 18696 20451 18748 20460
rect 11980 20340 12032 20392
rect 15568 20383 15620 20392
rect 6828 20272 6880 20324
rect 8944 20272 8996 20324
rect 9496 20272 9548 20324
rect 15568 20349 15577 20383
rect 15577 20349 15611 20383
rect 15611 20349 15620 20383
rect 15568 20340 15620 20349
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 18604 20340 18656 20392
rect 13728 20272 13780 20324
rect 14648 20272 14700 20324
rect 19800 20408 19852 20460
rect 20352 20451 20404 20460
rect 20352 20417 20361 20451
rect 20361 20417 20395 20451
rect 20395 20417 20404 20451
rect 20352 20408 20404 20417
rect 20536 20451 20588 20460
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20536 20408 20588 20417
rect 30104 20451 30156 20460
rect 4344 20204 4396 20256
rect 5080 20247 5132 20256
rect 5080 20213 5089 20247
rect 5089 20213 5123 20247
rect 5123 20213 5132 20247
rect 5080 20204 5132 20213
rect 6368 20204 6420 20256
rect 7104 20247 7156 20256
rect 7104 20213 7113 20247
rect 7113 20213 7147 20247
rect 7147 20213 7156 20247
rect 7104 20204 7156 20213
rect 8852 20204 8904 20256
rect 10232 20204 10284 20256
rect 12256 20247 12308 20256
rect 12256 20213 12265 20247
rect 12265 20213 12299 20247
rect 12299 20213 12308 20247
rect 12256 20204 12308 20213
rect 14096 20204 14148 20256
rect 14832 20204 14884 20256
rect 15108 20204 15160 20256
rect 19340 20272 19392 20324
rect 19984 20340 20036 20392
rect 20168 20340 20220 20392
rect 20444 20272 20496 20324
rect 30104 20417 30113 20451
rect 30113 20417 30147 20451
rect 30147 20417 30156 20451
rect 30104 20408 30156 20417
rect 22376 20383 22428 20392
rect 22376 20349 22385 20383
rect 22385 20349 22419 20383
rect 22419 20349 22428 20383
rect 22376 20340 22428 20349
rect 19432 20204 19484 20256
rect 20628 20204 20680 20256
rect 21732 20204 21784 20256
rect 5915 20102 5967 20154
rect 5979 20102 6031 20154
rect 6043 20102 6095 20154
rect 6107 20102 6159 20154
rect 6171 20102 6223 20154
rect 15846 20102 15898 20154
rect 15910 20102 15962 20154
rect 15974 20102 16026 20154
rect 16038 20102 16090 20154
rect 16102 20102 16154 20154
rect 25776 20102 25828 20154
rect 25840 20102 25892 20154
rect 25904 20102 25956 20154
rect 25968 20102 26020 20154
rect 26032 20102 26084 20154
rect 4528 20043 4580 20052
rect 4528 20009 4537 20043
rect 4537 20009 4571 20043
rect 4571 20009 4580 20043
rect 4528 20000 4580 20009
rect 6460 20000 6512 20052
rect 8392 20000 8444 20052
rect 4344 19932 4396 19984
rect 6552 19932 6604 19984
rect 1860 19796 1912 19848
rect 3700 19796 3752 19848
rect 3976 19839 4028 19848
rect 2228 19728 2280 19780
rect 3516 19728 3568 19780
rect 3976 19805 3985 19839
rect 3985 19805 4019 19839
rect 4019 19805 4028 19839
rect 3976 19796 4028 19805
rect 5080 19796 5132 19848
rect 5632 19796 5684 19848
rect 10508 20000 10560 20052
rect 12900 20043 12952 20052
rect 12900 20009 12909 20043
rect 12909 20009 12943 20043
rect 12943 20009 12952 20043
rect 12900 20000 12952 20009
rect 6276 19796 6328 19848
rect 6552 19839 6604 19848
rect 4528 19728 4580 19780
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 6920 19796 6972 19848
rect 8484 19796 8536 19848
rect 10048 19864 10100 19916
rect 10784 19864 10836 19916
rect 11520 19907 11572 19916
rect 11520 19873 11529 19907
rect 11529 19873 11563 19907
rect 11563 19873 11572 19907
rect 11520 19864 11572 19873
rect 13544 20000 13596 20052
rect 13912 20000 13964 20052
rect 13820 19932 13872 19984
rect 14280 19932 14332 19984
rect 14648 19932 14700 19984
rect 15568 19932 15620 19984
rect 16580 20000 16632 20052
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 20260 20000 20312 20052
rect 1676 19660 1728 19712
rect 2780 19660 2832 19712
rect 3148 19703 3200 19712
rect 3148 19669 3157 19703
rect 3157 19669 3191 19703
rect 3191 19669 3200 19703
rect 3148 19660 3200 19669
rect 5264 19660 5316 19712
rect 7840 19728 7892 19780
rect 8852 19728 8904 19780
rect 9864 19796 9916 19848
rect 10324 19796 10376 19848
rect 12256 19796 12308 19848
rect 13728 19864 13780 19916
rect 15844 19907 15896 19916
rect 15844 19873 15853 19907
rect 15853 19873 15887 19907
rect 15887 19873 15896 19907
rect 15844 19864 15896 19873
rect 16304 19864 16356 19916
rect 18880 19932 18932 19984
rect 19340 19864 19392 19916
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 14096 19839 14148 19848
rect 14096 19805 14105 19839
rect 14105 19805 14139 19839
rect 14139 19805 14148 19839
rect 14096 19796 14148 19805
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 15752 19839 15804 19848
rect 15752 19805 15761 19839
rect 15761 19805 15795 19839
rect 15795 19805 15804 19839
rect 15752 19796 15804 19805
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 16764 19839 16816 19848
rect 16764 19805 16773 19839
rect 16773 19805 16807 19839
rect 16807 19805 16816 19839
rect 16764 19796 16816 19805
rect 17960 19796 18012 19848
rect 19892 19796 19944 19848
rect 20812 19796 20864 19848
rect 21364 19839 21416 19848
rect 21364 19805 21373 19839
rect 21373 19805 21407 19839
rect 21407 19805 21416 19839
rect 21364 19796 21416 19805
rect 21088 19728 21140 19780
rect 7012 19660 7064 19712
rect 8392 19660 8444 19712
rect 8944 19660 8996 19712
rect 14740 19703 14792 19712
rect 14740 19669 14749 19703
rect 14749 19669 14783 19703
rect 14783 19669 14792 19703
rect 14740 19660 14792 19669
rect 15384 19660 15436 19712
rect 17316 19703 17368 19712
rect 17316 19669 17325 19703
rect 17325 19669 17359 19703
rect 17359 19669 17368 19703
rect 17316 19660 17368 19669
rect 17776 19703 17828 19712
rect 17776 19669 17785 19703
rect 17785 19669 17819 19703
rect 17819 19669 17828 19703
rect 17776 19660 17828 19669
rect 20720 19660 20772 19712
rect 10880 19558 10932 19610
rect 10944 19558 10996 19610
rect 11008 19558 11060 19610
rect 11072 19558 11124 19610
rect 11136 19558 11188 19610
rect 20811 19558 20863 19610
rect 20875 19558 20927 19610
rect 20939 19558 20991 19610
rect 21003 19558 21055 19610
rect 21067 19558 21119 19610
rect 1308 19456 1360 19508
rect 1768 19388 1820 19440
rect 2228 19431 2280 19440
rect 1492 19363 1544 19372
rect 1492 19329 1501 19363
rect 1501 19329 1535 19363
rect 1535 19329 1544 19363
rect 1492 19320 1544 19329
rect 1676 19363 1728 19372
rect 1676 19329 1685 19363
rect 1685 19329 1719 19363
rect 1719 19329 1728 19363
rect 1676 19320 1728 19329
rect 2228 19397 2237 19431
rect 2237 19397 2271 19431
rect 2271 19397 2280 19431
rect 2228 19388 2280 19397
rect 6736 19456 6788 19508
rect 8208 19499 8260 19508
rect 8208 19465 8217 19499
rect 8217 19465 8251 19499
rect 8251 19465 8260 19499
rect 8208 19456 8260 19465
rect 9864 19456 9916 19508
rect 10416 19456 10468 19508
rect 12440 19456 12492 19508
rect 13176 19499 13228 19508
rect 13176 19465 13185 19499
rect 13185 19465 13219 19499
rect 13219 19465 13228 19499
rect 13176 19456 13228 19465
rect 13544 19456 13596 19508
rect 16672 19499 16724 19508
rect 16672 19465 16681 19499
rect 16681 19465 16715 19499
rect 16715 19465 16724 19499
rect 16672 19456 16724 19465
rect 16764 19456 16816 19508
rect 17500 19456 17552 19508
rect 17776 19456 17828 19508
rect 18328 19456 18380 19508
rect 18972 19456 19024 19508
rect 20720 19499 20772 19508
rect 20720 19465 20729 19499
rect 20729 19465 20763 19499
rect 20763 19465 20772 19499
rect 20720 19456 20772 19465
rect 30012 19499 30064 19508
rect 30012 19465 30021 19499
rect 30021 19465 30055 19499
rect 30055 19465 30064 19499
rect 30012 19456 30064 19465
rect 14740 19388 14792 19440
rect 3516 19363 3568 19372
rect 1584 19252 1636 19304
rect 2044 19184 2096 19236
rect 3148 19184 3200 19236
rect 1492 19116 1544 19168
rect 3516 19329 3525 19363
rect 3525 19329 3559 19363
rect 3559 19329 3568 19363
rect 3516 19320 3568 19329
rect 3700 19320 3752 19372
rect 4804 19320 4856 19372
rect 6920 19320 6972 19372
rect 7104 19363 7156 19372
rect 7104 19329 7138 19363
rect 7138 19329 7156 19363
rect 7104 19320 7156 19329
rect 7932 19320 7984 19372
rect 9220 19363 9272 19372
rect 3792 19295 3844 19304
rect 3792 19261 3801 19295
rect 3801 19261 3835 19295
rect 3835 19261 3844 19295
rect 3792 19252 3844 19261
rect 9220 19329 9229 19363
rect 9229 19329 9263 19363
rect 9263 19329 9272 19363
rect 9220 19320 9272 19329
rect 9312 19252 9364 19304
rect 10324 19320 10376 19372
rect 10416 19363 10468 19372
rect 10416 19329 10425 19363
rect 10425 19329 10459 19363
rect 10459 19329 10468 19363
rect 19340 19388 19392 19440
rect 20628 19431 20680 19440
rect 15476 19363 15528 19372
rect 10416 19320 10468 19329
rect 15476 19329 15485 19363
rect 15485 19329 15519 19363
rect 15519 19329 15528 19363
rect 15476 19320 15528 19329
rect 16764 19320 16816 19372
rect 16212 19252 16264 19304
rect 17960 19363 18012 19372
rect 17960 19329 17969 19363
rect 17969 19329 18003 19363
rect 18003 19329 18012 19363
rect 17960 19320 18012 19329
rect 19248 19363 19300 19372
rect 19248 19329 19257 19363
rect 19257 19329 19291 19363
rect 19291 19329 19300 19363
rect 19248 19320 19300 19329
rect 6552 19184 6604 19236
rect 6828 19184 6880 19236
rect 15936 19184 15988 19236
rect 16488 19184 16540 19236
rect 18604 19252 18656 19304
rect 19340 19295 19392 19304
rect 19340 19261 19349 19295
rect 19349 19261 19383 19295
rect 19383 19261 19392 19295
rect 19340 19252 19392 19261
rect 20628 19397 20637 19431
rect 20637 19397 20671 19431
rect 20671 19397 20680 19431
rect 20628 19388 20680 19397
rect 29920 19320 29972 19372
rect 19616 19184 19668 19236
rect 5632 19159 5684 19168
rect 5632 19125 5641 19159
rect 5641 19125 5675 19159
rect 5675 19125 5684 19159
rect 5632 19116 5684 19125
rect 6460 19116 6512 19168
rect 8852 19116 8904 19168
rect 14832 19116 14884 19168
rect 20536 19184 20588 19236
rect 20260 19159 20312 19168
rect 20260 19125 20269 19159
rect 20269 19125 20303 19159
rect 20303 19125 20312 19159
rect 20260 19116 20312 19125
rect 5915 19014 5967 19066
rect 5979 19014 6031 19066
rect 6043 19014 6095 19066
rect 6107 19014 6159 19066
rect 6171 19014 6223 19066
rect 15846 19014 15898 19066
rect 15910 19014 15962 19066
rect 15974 19014 16026 19066
rect 16038 19014 16090 19066
rect 16102 19014 16154 19066
rect 25776 19014 25828 19066
rect 25840 19014 25892 19066
rect 25904 19014 25956 19066
rect 25968 19014 26020 19066
rect 26032 19014 26084 19066
rect 4804 18955 4856 18964
rect 4804 18921 4813 18955
rect 4813 18921 4847 18955
rect 4847 18921 4856 18955
rect 4804 18912 4856 18921
rect 5816 18912 5868 18964
rect 4344 18844 4396 18896
rect 1860 18819 1912 18828
rect 1860 18785 1869 18819
rect 1869 18785 1903 18819
rect 1903 18785 1912 18819
rect 1860 18776 1912 18785
rect 4528 18844 4580 18896
rect 10048 18912 10100 18964
rect 17960 18912 18012 18964
rect 18696 18912 18748 18964
rect 21364 18912 21416 18964
rect 4252 18751 4304 18760
rect 2504 18640 2556 18692
rect 4252 18717 4261 18751
rect 4261 18717 4295 18751
rect 4295 18717 4304 18751
rect 4252 18708 4304 18717
rect 5632 18776 5684 18828
rect 9404 18776 9456 18828
rect 5264 18751 5316 18760
rect 5264 18717 5273 18751
rect 5273 18717 5307 18751
rect 5307 18717 5316 18751
rect 5264 18708 5316 18717
rect 8208 18708 8260 18760
rect 8944 18751 8996 18760
rect 8944 18717 8953 18751
rect 8953 18717 8987 18751
rect 8987 18717 8996 18751
rect 8944 18708 8996 18717
rect 9312 18751 9364 18760
rect 4988 18640 5040 18692
rect 6920 18640 6972 18692
rect 7012 18683 7064 18692
rect 7012 18649 7030 18683
rect 7030 18649 7064 18683
rect 7012 18640 7064 18649
rect 8116 18640 8168 18692
rect 8760 18640 8812 18692
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 11428 18776 11480 18828
rect 16488 18776 16540 18828
rect 16672 18819 16724 18828
rect 16672 18785 16681 18819
rect 16681 18785 16715 18819
rect 16715 18785 16724 18819
rect 16672 18776 16724 18785
rect 19340 18776 19392 18828
rect 10600 18708 10652 18760
rect 12532 18751 12584 18760
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 14004 18708 14056 18760
rect 15660 18708 15712 18760
rect 16212 18751 16264 18760
rect 16212 18717 16221 18751
rect 16221 18717 16255 18751
rect 16255 18717 16264 18751
rect 16212 18708 16264 18717
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 19708 18708 19760 18760
rect 20444 18751 20496 18760
rect 20444 18717 20453 18751
rect 20453 18717 20487 18751
rect 20487 18717 20496 18751
rect 20444 18708 20496 18717
rect 16948 18640 17000 18692
rect 2320 18572 2372 18624
rect 4160 18572 4212 18624
rect 5816 18572 5868 18624
rect 9680 18615 9732 18624
rect 9680 18581 9689 18615
rect 9689 18581 9723 18615
rect 9723 18581 9732 18615
rect 9680 18572 9732 18581
rect 10324 18572 10376 18624
rect 10508 18572 10560 18624
rect 10692 18572 10744 18624
rect 11244 18572 11296 18624
rect 12624 18615 12676 18624
rect 12624 18581 12633 18615
rect 12633 18581 12667 18615
rect 12667 18581 12676 18615
rect 12624 18572 12676 18581
rect 12900 18572 12952 18624
rect 15476 18572 15528 18624
rect 19708 18615 19760 18624
rect 19708 18581 19717 18615
rect 19717 18581 19751 18615
rect 19751 18581 19760 18615
rect 19708 18572 19760 18581
rect 22192 18708 22244 18760
rect 21916 18572 21968 18624
rect 10880 18470 10932 18522
rect 10944 18470 10996 18522
rect 11008 18470 11060 18522
rect 11072 18470 11124 18522
rect 11136 18470 11188 18522
rect 20811 18470 20863 18522
rect 20875 18470 20927 18522
rect 20939 18470 20991 18522
rect 21003 18470 21055 18522
rect 21067 18470 21119 18522
rect 2504 18411 2556 18420
rect 2504 18377 2513 18411
rect 2513 18377 2547 18411
rect 2547 18377 2556 18411
rect 2504 18368 2556 18377
rect 1492 18232 1544 18284
rect 1952 18275 2004 18284
rect 1952 18241 1961 18275
rect 1961 18241 1995 18275
rect 1995 18241 2004 18275
rect 1952 18232 2004 18241
rect 2320 18275 2372 18284
rect 2044 18207 2096 18216
rect 2044 18173 2053 18207
rect 2053 18173 2087 18207
rect 2087 18173 2096 18207
rect 2044 18164 2096 18173
rect 1952 18096 2004 18148
rect 2320 18241 2329 18275
rect 2329 18241 2363 18275
rect 2363 18241 2372 18275
rect 2320 18232 2372 18241
rect 3516 18275 3568 18284
rect 3516 18241 3525 18275
rect 3525 18241 3559 18275
rect 3559 18241 3568 18275
rect 3516 18232 3568 18241
rect 3700 18275 3752 18284
rect 3700 18241 3709 18275
rect 3709 18241 3743 18275
rect 3743 18241 3752 18275
rect 3700 18232 3752 18241
rect 5724 18368 5776 18420
rect 9956 18368 10008 18420
rect 12900 18411 12952 18420
rect 4344 18300 4396 18352
rect 5448 18300 5500 18352
rect 4896 18275 4948 18284
rect 4896 18241 4905 18275
rect 4905 18241 4939 18275
rect 4939 18241 4948 18275
rect 8668 18300 8720 18352
rect 12900 18377 12909 18411
rect 12909 18377 12943 18411
rect 12943 18377 12952 18411
rect 12900 18368 12952 18377
rect 15476 18411 15528 18420
rect 15476 18377 15485 18411
rect 15485 18377 15519 18411
rect 15519 18377 15528 18411
rect 15476 18368 15528 18377
rect 18972 18411 19024 18420
rect 18972 18377 18981 18411
rect 18981 18377 19015 18411
rect 19015 18377 19024 18411
rect 18972 18368 19024 18377
rect 19616 18368 19668 18420
rect 20444 18368 20496 18420
rect 21916 18411 21968 18420
rect 21916 18377 21925 18411
rect 21925 18377 21959 18411
rect 21959 18377 21968 18411
rect 21916 18368 21968 18377
rect 13912 18343 13964 18352
rect 4896 18232 4948 18241
rect 6460 18232 6512 18284
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 9036 18232 9088 18284
rect 9404 18232 9456 18284
rect 13912 18309 13921 18343
rect 13921 18309 13955 18343
rect 13955 18309 13964 18343
rect 13912 18300 13964 18309
rect 14556 18300 14608 18352
rect 15384 18343 15436 18352
rect 15384 18309 15393 18343
rect 15393 18309 15427 18343
rect 15427 18309 15436 18343
rect 15384 18300 15436 18309
rect 9312 18207 9364 18216
rect 9312 18173 9321 18207
rect 9321 18173 9355 18207
rect 9355 18173 9364 18207
rect 9312 18164 9364 18173
rect 14280 18232 14332 18284
rect 14832 18232 14884 18284
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 18236 18232 18288 18284
rect 19340 18232 19392 18284
rect 19708 18275 19760 18284
rect 19708 18241 19718 18275
rect 19718 18241 19752 18275
rect 19752 18241 19760 18275
rect 19708 18232 19760 18241
rect 11520 18207 11572 18216
rect 11520 18173 11529 18207
rect 11529 18173 11563 18207
rect 11563 18173 11572 18207
rect 11520 18164 11572 18173
rect 15568 18207 15620 18216
rect 15568 18173 15577 18207
rect 15577 18173 15611 18207
rect 15611 18173 15620 18207
rect 15568 18164 15620 18173
rect 17500 18207 17552 18216
rect 17500 18173 17509 18207
rect 17509 18173 17543 18207
rect 17543 18173 17552 18207
rect 17500 18164 17552 18173
rect 18052 18207 18104 18216
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 20168 18232 20220 18284
rect 20536 18275 20588 18284
rect 20536 18241 20545 18275
rect 20545 18241 20579 18275
rect 20579 18241 20588 18275
rect 20536 18232 20588 18241
rect 20720 18275 20772 18284
rect 20720 18241 20729 18275
rect 20729 18241 20763 18275
rect 20763 18241 20772 18275
rect 20720 18232 20772 18241
rect 21180 18232 21232 18284
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 29828 18275 29880 18284
rect 29828 18241 29837 18275
rect 29837 18241 29871 18275
rect 29871 18241 29880 18275
rect 29828 18232 29880 18241
rect 4436 18096 4488 18148
rect 4252 18071 4304 18080
rect 4252 18037 4261 18071
rect 4261 18037 4295 18071
rect 4295 18037 4304 18071
rect 4252 18028 4304 18037
rect 4344 18028 4396 18080
rect 6460 18071 6512 18080
rect 6460 18037 6469 18071
rect 6469 18037 6503 18071
rect 6503 18037 6512 18071
rect 6460 18028 6512 18037
rect 6736 18028 6788 18080
rect 9496 18096 9548 18148
rect 13452 18096 13504 18148
rect 13728 18139 13780 18148
rect 13728 18105 13737 18139
rect 13737 18105 13771 18139
rect 13771 18105 13780 18139
rect 13728 18096 13780 18105
rect 10508 18028 10560 18080
rect 10692 18028 10744 18080
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 15016 18071 15068 18080
rect 15016 18037 15025 18071
rect 15025 18037 15059 18071
rect 15059 18037 15068 18071
rect 15016 18028 15068 18037
rect 19984 18071 20036 18080
rect 19984 18037 19993 18071
rect 19993 18037 20027 18071
rect 20027 18037 20036 18071
rect 19984 18028 20036 18037
rect 30012 18071 30064 18080
rect 30012 18037 30021 18071
rect 30021 18037 30055 18071
rect 30055 18037 30064 18071
rect 30012 18028 30064 18037
rect 5915 17926 5967 17978
rect 5979 17926 6031 17978
rect 6043 17926 6095 17978
rect 6107 17926 6159 17978
rect 6171 17926 6223 17978
rect 15846 17926 15898 17978
rect 15910 17926 15962 17978
rect 15974 17926 16026 17978
rect 16038 17926 16090 17978
rect 16102 17926 16154 17978
rect 25776 17926 25828 17978
rect 25840 17926 25892 17978
rect 25904 17926 25956 17978
rect 25968 17926 26020 17978
rect 26032 17926 26084 17978
rect 3700 17824 3752 17876
rect 11428 17824 11480 17876
rect 12992 17867 13044 17876
rect 12992 17833 13001 17867
rect 13001 17833 13035 17867
rect 13035 17833 13044 17867
rect 12992 17824 13044 17833
rect 14004 17824 14056 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 15752 17824 15804 17876
rect 16948 17824 17000 17876
rect 17500 17824 17552 17876
rect 19340 17867 19392 17876
rect 19340 17833 19349 17867
rect 19349 17833 19383 17867
rect 19383 17833 19392 17867
rect 19340 17824 19392 17833
rect 20720 17824 20772 17876
rect 29828 17824 29880 17876
rect 6276 17756 6328 17808
rect 2044 17731 2096 17740
rect 2044 17697 2053 17731
rect 2053 17697 2087 17731
rect 2087 17697 2096 17731
rect 2044 17688 2096 17697
rect 1952 17663 2004 17672
rect 1676 17484 1728 17536
rect 1952 17629 1961 17663
rect 1961 17629 1995 17663
rect 1995 17629 2004 17663
rect 1952 17620 2004 17629
rect 2872 17688 2924 17740
rect 3792 17731 3844 17740
rect 3792 17697 3801 17731
rect 3801 17697 3835 17731
rect 3835 17697 3844 17731
rect 3792 17688 3844 17697
rect 4344 17688 4396 17740
rect 2780 17663 2832 17672
rect 2780 17629 2789 17663
rect 2789 17629 2823 17663
rect 2823 17629 2832 17663
rect 2780 17620 2832 17629
rect 2872 17552 2924 17604
rect 3516 17552 3568 17604
rect 4160 17620 4212 17672
rect 6276 17620 6328 17672
rect 8944 17756 8996 17808
rect 13452 17756 13504 17808
rect 15200 17756 15252 17808
rect 8116 17688 8168 17740
rect 8300 17688 8352 17740
rect 13820 17688 13872 17740
rect 17224 17756 17276 17808
rect 16672 17688 16724 17740
rect 19248 17756 19300 17808
rect 18052 17688 18104 17740
rect 19984 17756 20036 17808
rect 19616 17688 19668 17740
rect 2412 17484 2464 17536
rect 5632 17484 5684 17536
rect 9220 17620 9272 17672
rect 9680 17620 9732 17672
rect 11520 17620 11572 17672
rect 13912 17620 13964 17672
rect 14556 17663 14608 17672
rect 14556 17629 14565 17663
rect 14565 17629 14599 17663
rect 14599 17629 14608 17663
rect 14556 17620 14608 17629
rect 16212 17663 16264 17672
rect 16212 17629 16221 17663
rect 16221 17629 16255 17663
rect 16255 17629 16264 17663
rect 16212 17620 16264 17629
rect 16856 17620 16908 17672
rect 17684 17620 17736 17672
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 19524 17620 19576 17672
rect 20168 17620 20220 17672
rect 30104 17663 30156 17672
rect 30104 17629 30113 17663
rect 30113 17629 30147 17663
rect 30147 17629 30156 17663
rect 30104 17620 30156 17629
rect 9496 17552 9548 17604
rect 9864 17552 9916 17604
rect 11980 17552 12032 17604
rect 19708 17552 19760 17604
rect 8208 17484 8260 17536
rect 8392 17527 8444 17536
rect 8392 17493 8401 17527
rect 8401 17493 8435 17527
rect 8435 17493 8444 17527
rect 8392 17484 8444 17493
rect 13636 17484 13688 17536
rect 16028 17484 16080 17536
rect 10880 17382 10932 17434
rect 10944 17382 10996 17434
rect 11008 17382 11060 17434
rect 11072 17382 11124 17434
rect 11136 17382 11188 17434
rect 20811 17382 20863 17434
rect 20875 17382 20927 17434
rect 20939 17382 20991 17434
rect 21003 17382 21055 17434
rect 21067 17382 21119 17434
rect 9220 17280 9272 17332
rect 9864 17323 9916 17332
rect 9864 17289 9873 17323
rect 9873 17289 9907 17323
rect 9907 17289 9916 17323
rect 9864 17280 9916 17289
rect 15200 17280 15252 17332
rect 16304 17280 16356 17332
rect 16856 17280 16908 17332
rect 18052 17280 18104 17332
rect 2320 17212 2372 17264
rect 7196 17212 7248 17264
rect 8392 17212 8444 17264
rect 12624 17212 12676 17264
rect 1676 17187 1728 17196
rect 1676 17153 1710 17187
rect 1710 17153 1728 17187
rect 1676 17144 1728 17153
rect 3240 17187 3292 17196
rect 3240 17153 3249 17187
rect 3249 17153 3283 17187
rect 3283 17153 3292 17187
rect 3240 17144 3292 17153
rect 4068 17187 4120 17196
rect 4068 17153 4077 17187
rect 4077 17153 4111 17187
rect 4111 17153 4120 17187
rect 4068 17144 4120 17153
rect 4344 17187 4396 17196
rect 4344 17153 4378 17187
rect 4378 17153 4396 17187
rect 4344 17144 4396 17153
rect 6276 17144 6328 17196
rect 7932 17144 7984 17196
rect 8944 17144 8996 17196
rect 9220 17144 9272 17196
rect 9772 17144 9824 17196
rect 13820 17187 13872 17196
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 7196 17076 7248 17128
rect 9404 17119 9456 17128
rect 9404 17085 9413 17119
rect 9413 17085 9447 17119
rect 9447 17085 9456 17119
rect 9404 17076 9456 17085
rect 9496 17119 9548 17128
rect 9496 17085 9505 17119
rect 9505 17085 9539 17119
rect 9539 17085 9548 17119
rect 11980 17119 12032 17128
rect 9496 17076 9548 17085
rect 11980 17085 11989 17119
rect 11989 17085 12023 17119
rect 12023 17085 12032 17119
rect 11980 17076 12032 17085
rect 2412 17008 2464 17060
rect 2320 16940 2372 16992
rect 3976 16940 4028 16992
rect 4712 16940 4764 16992
rect 4804 16940 4856 16992
rect 5448 16983 5500 16992
rect 5448 16949 5457 16983
rect 5457 16949 5491 16983
rect 5491 16949 5500 16983
rect 5448 16940 5500 16949
rect 6644 16940 6696 16992
rect 8392 16940 8444 16992
rect 10048 16940 10100 16992
rect 10324 16940 10376 16992
rect 13820 16940 13872 16992
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 14924 17119 14976 17128
rect 14924 17085 14933 17119
rect 14933 17085 14967 17119
rect 14967 17085 14976 17119
rect 15752 17212 15804 17264
rect 16028 17144 16080 17196
rect 17224 17212 17276 17264
rect 17592 17212 17644 17264
rect 17684 17144 17736 17196
rect 19248 17144 19300 17196
rect 21272 17280 21324 17332
rect 19800 17212 19852 17264
rect 19616 17144 19668 17196
rect 20260 17144 20312 17196
rect 14924 17076 14976 17085
rect 17868 17076 17920 17128
rect 19892 17119 19944 17128
rect 19892 17085 19901 17119
rect 19901 17085 19935 17119
rect 19935 17085 19944 17119
rect 19892 17076 19944 17085
rect 14740 17008 14792 17060
rect 16764 17008 16816 17060
rect 19708 17008 19760 17060
rect 13912 16940 13964 16949
rect 15108 16940 15160 16992
rect 18972 16983 19024 16992
rect 18972 16949 18981 16983
rect 18981 16949 19015 16983
rect 19015 16949 19024 16983
rect 18972 16940 19024 16949
rect 19340 16940 19392 16992
rect 19984 16940 20036 16992
rect 20720 16940 20772 16992
rect 5915 16838 5967 16890
rect 5979 16838 6031 16890
rect 6043 16838 6095 16890
rect 6107 16838 6159 16890
rect 6171 16838 6223 16890
rect 15846 16838 15898 16890
rect 15910 16838 15962 16890
rect 15974 16838 16026 16890
rect 16038 16838 16090 16890
rect 16102 16838 16154 16890
rect 25776 16838 25828 16890
rect 25840 16838 25892 16890
rect 25904 16838 25956 16890
rect 25968 16838 26020 16890
rect 26032 16838 26084 16890
rect 6276 16779 6328 16788
rect 6276 16745 6285 16779
rect 6285 16745 6319 16779
rect 6319 16745 6328 16779
rect 6276 16736 6328 16745
rect 4160 16668 4212 16720
rect 4068 16600 4120 16652
rect 7196 16736 7248 16788
rect 10048 16736 10100 16788
rect 18236 16736 18288 16788
rect 19340 16736 19392 16788
rect 13268 16711 13320 16720
rect 13268 16677 13277 16711
rect 13277 16677 13311 16711
rect 13311 16677 13320 16711
rect 13268 16668 13320 16677
rect 8116 16600 8168 16652
rect 9404 16600 9456 16652
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 2044 16532 2096 16584
rect 4252 16532 4304 16584
rect 6644 16532 6696 16584
rect 9128 16532 9180 16584
rect 10232 16532 10284 16584
rect 13084 16532 13136 16584
rect 13820 16600 13872 16652
rect 14464 16600 14516 16652
rect 19340 16600 19392 16652
rect 19800 16668 19852 16720
rect 20168 16600 20220 16652
rect 13636 16532 13688 16584
rect 15108 16575 15160 16584
rect 15108 16541 15117 16575
rect 15117 16541 15151 16575
rect 15151 16541 15160 16575
rect 15108 16532 15160 16541
rect 16764 16532 16816 16584
rect 17224 16575 17276 16584
rect 17224 16541 17233 16575
rect 17233 16541 17267 16575
rect 17267 16541 17276 16575
rect 17224 16532 17276 16541
rect 19432 16575 19484 16584
rect 19432 16541 19441 16575
rect 19441 16541 19475 16575
rect 19475 16541 19484 16575
rect 19432 16532 19484 16541
rect 19699 16575 19751 16584
rect 19699 16541 19714 16575
rect 19714 16541 19748 16575
rect 19748 16541 19751 16575
rect 19699 16532 19751 16541
rect 19892 16532 19944 16584
rect 20260 16532 20312 16584
rect 20628 16575 20680 16584
rect 20628 16541 20637 16575
rect 20637 16541 20671 16575
rect 20671 16541 20680 16575
rect 20628 16532 20680 16541
rect 20720 16532 20772 16584
rect 29920 16532 29972 16584
rect 7196 16464 7248 16516
rect 2228 16396 2280 16448
rect 5724 16439 5776 16448
rect 5724 16405 5733 16439
rect 5733 16405 5767 16439
rect 5767 16405 5776 16439
rect 5724 16396 5776 16405
rect 6828 16396 6880 16448
rect 6920 16396 6972 16448
rect 13728 16464 13780 16516
rect 8576 16396 8628 16448
rect 12532 16396 12584 16448
rect 18052 16396 18104 16448
rect 19616 16396 19668 16448
rect 22008 16439 22060 16448
rect 22008 16405 22017 16439
rect 22017 16405 22051 16439
rect 22051 16405 22060 16439
rect 22008 16396 22060 16405
rect 30012 16439 30064 16448
rect 30012 16405 30021 16439
rect 30021 16405 30055 16439
rect 30055 16405 30064 16439
rect 30012 16396 30064 16405
rect 10880 16294 10932 16346
rect 10944 16294 10996 16346
rect 11008 16294 11060 16346
rect 11072 16294 11124 16346
rect 11136 16294 11188 16346
rect 20811 16294 20863 16346
rect 20875 16294 20927 16346
rect 20939 16294 20991 16346
rect 21003 16294 21055 16346
rect 21067 16294 21119 16346
rect 7196 16235 7248 16244
rect 7196 16201 7205 16235
rect 7205 16201 7239 16235
rect 7239 16201 7248 16235
rect 7196 16192 7248 16201
rect 7288 16192 7340 16244
rect 7748 16192 7800 16244
rect 7932 16192 7984 16244
rect 13452 16235 13504 16244
rect 2780 16124 2832 16176
rect 3792 16124 3844 16176
rect 8576 16124 8628 16176
rect 1216 16056 1268 16108
rect 2872 16056 2924 16108
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 4712 16056 4764 16108
rect 6276 16056 6328 16108
rect 6920 16056 6972 16108
rect 7748 16099 7800 16108
rect 7748 16065 7757 16099
rect 7757 16065 7791 16099
rect 7791 16065 7800 16099
rect 7932 16099 7984 16108
rect 7748 16056 7800 16065
rect 7932 16065 7941 16099
rect 7941 16065 7975 16099
rect 7975 16065 7984 16099
rect 7932 16056 7984 16065
rect 2320 16031 2372 16040
rect 2320 15997 2329 16031
rect 2329 15997 2363 16031
rect 2363 15997 2372 16031
rect 2320 15988 2372 15997
rect 4160 16031 4212 16040
rect 4160 15997 4169 16031
rect 4169 15997 4203 16031
rect 4203 15997 4212 16031
rect 4160 15988 4212 15997
rect 4528 15988 4580 16040
rect 6644 15988 6696 16040
rect 7104 15988 7156 16040
rect 8116 15988 8168 16040
rect 9496 16056 9548 16108
rect 13452 16201 13461 16235
rect 13461 16201 13495 16235
rect 13495 16201 13504 16235
rect 13452 16192 13504 16201
rect 13544 16192 13596 16244
rect 9956 16124 10008 16176
rect 10784 16124 10836 16176
rect 15200 16192 15252 16244
rect 17224 16192 17276 16244
rect 3700 15963 3752 15972
rect 3700 15929 3709 15963
rect 3709 15929 3743 15963
rect 3743 15929 3752 15963
rect 3700 15920 3752 15929
rect 7472 15920 7524 15972
rect 7932 15920 7984 15972
rect 9128 15988 9180 16040
rect 9404 15920 9456 15972
rect 2964 15852 3016 15904
rect 5724 15852 5776 15904
rect 6644 15895 6696 15904
rect 6644 15861 6653 15895
rect 6653 15861 6687 15895
rect 6687 15861 6696 15895
rect 6644 15852 6696 15861
rect 10416 15852 10468 15904
rect 12532 16099 12584 16108
rect 12532 16065 12541 16099
rect 12541 16065 12575 16099
rect 12575 16065 12584 16099
rect 12532 16056 12584 16065
rect 13636 16099 13688 16108
rect 13636 16065 13645 16099
rect 13645 16065 13679 16099
rect 13679 16065 13688 16099
rect 13636 16056 13688 16065
rect 13820 16099 13872 16108
rect 13820 16065 13829 16099
rect 13829 16065 13863 16099
rect 13863 16065 13872 16099
rect 13820 16056 13872 16065
rect 14924 16124 14976 16176
rect 18604 16192 18656 16244
rect 18696 16192 18748 16244
rect 20260 16192 20312 16244
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 14832 16099 14884 16108
rect 14832 16065 14841 16099
rect 14841 16065 14875 16099
rect 14875 16065 14884 16099
rect 14832 16056 14884 16065
rect 16672 16099 16724 16108
rect 16672 16065 16681 16099
rect 16681 16065 16715 16099
rect 16715 16065 16724 16099
rect 16672 16056 16724 16065
rect 16856 16099 16908 16108
rect 16856 16065 16865 16099
rect 16865 16065 16899 16099
rect 16899 16065 16908 16099
rect 16856 16056 16908 16065
rect 19984 16124 20036 16176
rect 14556 15988 14608 16040
rect 16948 16031 17000 16040
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 17316 16056 17368 16108
rect 18052 16056 18104 16108
rect 17868 15988 17920 16040
rect 13268 15920 13320 15972
rect 13728 15963 13780 15972
rect 13728 15929 13737 15963
rect 13737 15929 13771 15963
rect 13771 15929 13780 15963
rect 13728 15920 13780 15929
rect 14740 15920 14792 15972
rect 18604 16099 18656 16108
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 18972 16056 19024 16108
rect 19248 15988 19300 16040
rect 19340 15988 19392 16040
rect 20628 16056 20680 16108
rect 19064 15920 19116 15972
rect 19708 15920 19760 15972
rect 10692 15852 10744 15904
rect 12256 15852 12308 15904
rect 19524 15852 19576 15904
rect 19892 15852 19944 15904
rect 5915 15750 5967 15802
rect 5979 15750 6031 15802
rect 6043 15750 6095 15802
rect 6107 15750 6159 15802
rect 6171 15750 6223 15802
rect 15846 15750 15898 15802
rect 15910 15750 15962 15802
rect 15974 15750 16026 15802
rect 16038 15750 16090 15802
rect 16102 15750 16154 15802
rect 25776 15750 25828 15802
rect 25840 15750 25892 15802
rect 25904 15750 25956 15802
rect 25968 15750 26020 15802
rect 26032 15750 26084 15802
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 2780 15648 2832 15700
rect 4344 15648 4396 15700
rect 3148 15580 3200 15632
rect 2872 15555 2924 15564
rect 2872 15521 2881 15555
rect 2881 15521 2915 15555
rect 2915 15521 2924 15555
rect 2872 15512 2924 15521
rect 3056 15512 3108 15564
rect 4068 15555 4120 15564
rect 4068 15521 4077 15555
rect 4077 15521 4111 15555
rect 4111 15521 4120 15555
rect 4068 15512 4120 15521
rect 4436 15512 4488 15564
rect 2228 15444 2280 15496
rect 1952 15376 2004 15428
rect 3700 15444 3752 15496
rect 3792 15487 3844 15496
rect 3792 15453 3801 15487
rect 3801 15453 3835 15487
rect 3835 15453 3844 15487
rect 3976 15487 4028 15496
rect 3792 15444 3844 15453
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 4804 15444 4856 15496
rect 5356 15444 5408 15496
rect 5908 15580 5960 15632
rect 6644 15648 6696 15700
rect 6736 15580 6788 15632
rect 6828 15580 6880 15632
rect 7104 15648 7156 15700
rect 7932 15648 7984 15700
rect 9312 15648 9364 15700
rect 13636 15648 13688 15700
rect 9772 15580 9824 15632
rect 6092 15444 6144 15496
rect 6460 15444 6512 15496
rect 7472 15487 7524 15496
rect 5264 15376 5316 15428
rect 7472 15453 7481 15487
rect 7481 15453 7515 15487
rect 7515 15453 7524 15487
rect 7472 15444 7524 15453
rect 7932 15376 7984 15428
rect 8392 15444 8444 15496
rect 9128 15487 9180 15496
rect 9128 15453 9135 15487
rect 9135 15453 9180 15487
rect 9128 15444 9180 15453
rect 9312 15512 9364 15564
rect 15752 15648 15804 15700
rect 16212 15648 16264 15700
rect 17040 15648 17092 15700
rect 17684 15691 17736 15700
rect 17684 15657 17693 15691
rect 17693 15657 17727 15691
rect 17727 15657 17736 15691
rect 17684 15648 17736 15657
rect 17776 15648 17828 15700
rect 20720 15648 20772 15700
rect 29920 15691 29972 15700
rect 29920 15657 29929 15691
rect 29929 15657 29963 15691
rect 29963 15657 29972 15691
rect 29920 15648 29972 15657
rect 30104 15648 30156 15700
rect 18604 15580 18656 15632
rect 19708 15580 19760 15632
rect 9404 15487 9456 15496
rect 9404 15453 9418 15487
rect 9418 15453 9452 15487
rect 9452 15453 9456 15487
rect 10048 15487 10100 15496
rect 9404 15444 9456 15453
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 12256 15487 12308 15496
rect 12256 15453 12290 15487
rect 12290 15453 12308 15487
rect 12256 15444 12308 15453
rect 13084 15444 13136 15496
rect 14556 15444 14608 15496
rect 14924 15512 14976 15564
rect 16856 15512 16908 15564
rect 17500 15512 17552 15564
rect 18236 15512 18288 15564
rect 14740 15487 14792 15496
rect 14740 15453 14749 15487
rect 14749 15453 14783 15487
rect 14783 15453 14792 15487
rect 15016 15487 15068 15496
rect 14740 15444 14792 15453
rect 15016 15453 15025 15487
rect 15025 15453 15059 15487
rect 15059 15453 15068 15487
rect 15016 15444 15068 15453
rect 15752 15444 15804 15496
rect 17592 15444 17644 15496
rect 19432 15444 19484 15496
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 19892 15444 19944 15496
rect 8300 15376 8352 15428
rect 4068 15308 4120 15360
rect 6276 15308 6328 15360
rect 6828 15308 6880 15360
rect 7104 15308 7156 15360
rect 7564 15351 7616 15360
rect 7564 15317 7573 15351
rect 7573 15317 7607 15351
rect 7607 15317 7616 15351
rect 7564 15308 7616 15317
rect 7656 15308 7708 15360
rect 10784 15376 10836 15428
rect 16580 15376 16632 15428
rect 17776 15376 17828 15428
rect 15200 15351 15252 15360
rect 15200 15317 15209 15351
rect 15209 15317 15243 15351
rect 15243 15317 15252 15351
rect 15200 15308 15252 15317
rect 18236 15376 18288 15428
rect 19248 15376 19300 15428
rect 21548 15444 21600 15496
rect 29920 15487 29972 15496
rect 29920 15453 29929 15487
rect 29929 15453 29963 15487
rect 29963 15453 29972 15487
rect 29920 15444 29972 15453
rect 30288 15444 30340 15496
rect 22744 15376 22796 15428
rect 18144 15308 18196 15360
rect 21824 15351 21876 15360
rect 21824 15317 21833 15351
rect 21833 15317 21867 15351
rect 21867 15317 21876 15351
rect 21824 15308 21876 15317
rect 10880 15206 10932 15258
rect 10944 15206 10996 15258
rect 11008 15206 11060 15258
rect 11072 15206 11124 15258
rect 11136 15206 11188 15258
rect 20811 15206 20863 15258
rect 20875 15206 20927 15258
rect 20939 15206 20991 15258
rect 21003 15206 21055 15258
rect 21067 15206 21119 15258
rect 5264 15147 5316 15156
rect 2780 15036 2832 15088
rect 2964 15036 3016 15088
rect 5264 15113 5273 15147
rect 5273 15113 5307 15147
rect 5307 15113 5316 15147
rect 5264 15104 5316 15113
rect 6092 15104 6144 15156
rect 6736 15104 6788 15156
rect 8852 15147 8904 15156
rect 8852 15113 8861 15147
rect 8861 15113 8895 15147
rect 8895 15113 8904 15147
rect 8852 15104 8904 15113
rect 9404 15104 9456 15156
rect 9496 15104 9548 15156
rect 4252 15036 4304 15088
rect 5540 15036 5592 15088
rect 14648 15104 14700 15156
rect 15568 15104 15620 15156
rect 16764 15104 16816 15156
rect 17868 15104 17920 15156
rect 19800 15104 19852 15156
rect 29184 15104 29236 15156
rect 1216 14900 1268 14952
rect 2780 14900 2832 14952
rect 2964 14943 3016 14952
rect 2964 14909 2973 14943
rect 2973 14909 3007 14943
rect 3007 14909 3016 14943
rect 2964 14900 3016 14909
rect 5264 14968 5316 15020
rect 6460 14968 6512 15020
rect 6736 15011 6788 15020
rect 6736 14977 6745 15011
rect 6745 14977 6779 15011
rect 6779 14977 6788 15011
rect 6736 14968 6788 14977
rect 7564 14968 7616 15020
rect 9128 14968 9180 15020
rect 10692 15011 10744 15020
rect 10692 14977 10710 15011
rect 10710 14977 10744 15011
rect 10692 14968 10744 14977
rect 11980 14968 12032 15020
rect 12440 14968 12492 15020
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12716 15011 12768 15020
rect 12532 14968 12584 14977
rect 12716 14977 12725 15011
rect 12725 14977 12759 15011
rect 12759 14977 12768 15011
rect 12716 14968 12768 14977
rect 13636 14968 13688 15020
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 15200 15036 15252 15088
rect 15752 15036 15804 15088
rect 16948 15036 17000 15088
rect 17592 15036 17644 15088
rect 17960 15036 18012 15088
rect 18144 15036 18196 15088
rect 18236 15079 18288 15088
rect 18236 15045 18245 15079
rect 18245 15045 18279 15079
rect 18279 15045 18288 15079
rect 18972 15079 19024 15088
rect 18236 15036 18288 15045
rect 18972 15045 18981 15079
rect 18981 15045 19015 15079
rect 19015 15045 19024 15079
rect 18972 15036 19024 15045
rect 22744 15036 22796 15088
rect 16580 14968 16632 15020
rect 16764 14968 16816 15020
rect 20444 14968 20496 15020
rect 20628 15011 20680 15020
rect 20628 14977 20637 15011
rect 20637 14977 20671 15011
rect 20671 14977 20680 15011
rect 20628 14968 20680 14977
rect 21456 14968 21508 15020
rect 21916 14968 21968 15020
rect 29184 15011 29236 15020
rect 29184 14977 29193 15011
rect 29193 14977 29227 15011
rect 29227 14977 29236 15011
rect 29184 14968 29236 14977
rect 29828 15011 29880 15020
rect 1492 14832 1544 14884
rect 2320 14832 2372 14884
rect 1860 14764 1912 14816
rect 1952 14764 2004 14816
rect 5908 14832 5960 14884
rect 6368 14832 6420 14884
rect 6828 14832 6880 14884
rect 9680 14900 9732 14952
rect 12808 14943 12860 14952
rect 12808 14909 12817 14943
rect 12817 14909 12851 14943
rect 12851 14909 12860 14943
rect 12808 14900 12860 14909
rect 14464 14943 14516 14952
rect 14464 14909 14473 14943
rect 14473 14909 14507 14943
rect 14507 14909 14516 14943
rect 14464 14900 14516 14909
rect 15476 14900 15528 14952
rect 17408 14900 17460 14952
rect 20260 14943 20312 14952
rect 20260 14909 20269 14943
rect 20269 14909 20303 14943
rect 20303 14909 20312 14943
rect 20260 14900 20312 14909
rect 29828 14977 29837 15011
rect 29837 14977 29871 15011
rect 29871 14977 29880 15011
rect 29828 14968 29880 14977
rect 30288 14900 30340 14952
rect 5172 14764 5224 14816
rect 6460 14764 6512 14816
rect 9496 14764 9548 14816
rect 9956 14764 10008 14816
rect 12348 14764 12400 14816
rect 12532 14764 12584 14816
rect 13728 14764 13780 14816
rect 14648 14764 14700 14816
rect 14832 14764 14884 14816
rect 29644 14832 29696 14884
rect 15752 14764 15804 14816
rect 19156 14764 19208 14816
rect 22284 14764 22336 14816
rect 30012 14807 30064 14816
rect 30012 14773 30021 14807
rect 30021 14773 30055 14807
rect 30055 14773 30064 14807
rect 30012 14764 30064 14773
rect 5915 14662 5967 14714
rect 5979 14662 6031 14714
rect 6043 14662 6095 14714
rect 6107 14662 6159 14714
rect 6171 14662 6223 14714
rect 15846 14662 15898 14714
rect 15910 14662 15962 14714
rect 15974 14662 16026 14714
rect 16038 14662 16090 14714
rect 16102 14662 16154 14714
rect 25776 14662 25828 14714
rect 25840 14662 25892 14714
rect 25904 14662 25956 14714
rect 25968 14662 26020 14714
rect 26032 14662 26084 14714
rect 3148 14560 3200 14612
rect 6460 14603 6512 14612
rect 6460 14569 6469 14603
rect 6469 14569 6503 14603
rect 6503 14569 6512 14603
rect 6460 14560 6512 14569
rect 11888 14560 11940 14612
rect 12716 14560 12768 14612
rect 14280 14560 14332 14612
rect 6092 14492 6144 14544
rect 6736 14492 6788 14544
rect 8116 14492 8168 14544
rect 9956 14492 10008 14544
rect 10784 14492 10836 14544
rect 16028 14492 16080 14544
rect 16304 14560 16356 14612
rect 29828 14560 29880 14612
rect 16580 14492 16632 14544
rect 29920 14492 29972 14544
rect 5172 14467 5224 14476
rect 5172 14433 5181 14467
rect 5181 14433 5215 14467
rect 5215 14433 5224 14467
rect 5172 14424 5224 14433
rect 1492 14399 1544 14408
rect 1492 14365 1501 14399
rect 1501 14365 1535 14399
rect 1535 14365 1544 14399
rect 1492 14356 1544 14365
rect 2596 14356 2648 14408
rect 5540 14356 5592 14408
rect 6460 14424 6512 14476
rect 7012 14424 7064 14476
rect 8300 14424 8352 14476
rect 12532 14424 12584 14476
rect 5816 14356 5868 14408
rect 1400 14288 1452 14340
rect 2412 14288 2464 14340
rect 3792 14263 3844 14272
rect 3792 14229 3801 14263
rect 3801 14229 3835 14263
rect 3835 14229 3844 14263
rect 3792 14220 3844 14229
rect 4620 14288 4672 14340
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6276 14399 6328 14408
rect 6092 14356 6144 14365
rect 6276 14365 6285 14399
rect 6285 14365 6319 14399
rect 6319 14365 6328 14399
rect 6276 14356 6328 14365
rect 6644 14356 6696 14408
rect 7104 14399 7156 14408
rect 7104 14365 7113 14399
rect 7113 14365 7147 14399
rect 7147 14365 7156 14399
rect 7104 14356 7156 14365
rect 6184 14220 6236 14272
rect 6276 14220 6328 14272
rect 7104 14220 7156 14272
rect 8024 14356 8076 14408
rect 10048 14356 10100 14408
rect 11796 14399 11848 14408
rect 11796 14365 11805 14399
rect 11805 14365 11839 14399
rect 11839 14365 11848 14399
rect 11796 14356 11848 14365
rect 13636 14424 13688 14476
rect 16120 14467 16172 14476
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 18144 14467 18196 14476
rect 18144 14433 18153 14467
rect 18153 14433 18187 14467
rect 18187 14433 18196 14467
rect 18144 14424 18196 14433
rect 18236 14424 18288 14476
rect 8116 14288 8168 14340
rect 8668 14288 8720 14340
rect 12900 14288 12952 14340
rect 13820 14356 13872 14408
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 15936 14356 15988 14408
rect 16764 14356 16816 14408
rect 16948 14399 17000 14408
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 16948 14356 17000 14365
rect 17316 14399 17368 14408
rect 15108 14288 15160 14340
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 17500 14399 17552 14408
rect 17500 14365 17509 14399
rect 17509 14365 17543 14399
rect 17543 14365 17552 14399
rect 17500 14356 17552 14365
rect 17868 14356 17920 14408
rect 18052 14399 18104 14408
rect 18052 14365 18061 14399
rect 18061 14365 18095 14399
rect 18095 14365 18104 14399
rect 18328 14399 18380 14408
rect 18052 14356 18104 14365
rect 18328 14365 18337 14399
rect 18337 14365 18371 14399
rect 18371 14365 18380 14399
rect 18328 14356 18380 14365
rect 18604 14356 18656 14408
rect 20628 14424 20680 14476
rect 30104 14492 30156 14544
rect 20536 14356 20588 14408
rect 20720 14399 20772 14408
rect 20720 14365 20729 14399
rect 20729 14365 20763 14399
rect 20763 14365 20772 14399
rect 20720 14356 20772 14365
rect 12716 14220 12768 14272
rect 15476 14220 15528 14272
rect 15844 14263 15896 14272
rect 15844 14229 15853 14263
rect 15853 14229 15887 14263
rect 15887 14229 15896 14263
rect 15844 14220 15896 14229
rect 16212 14220 16264 14272
rect 17316 14263 17368 14272
rect 17316 14229 17325 14263
rect 17325 14229 17359 14263
rect 17359 14229 17368 14263
rect 17316 14220 17368 14229
rect 17868 14220 17920 14272
rect 20260 14288 20312 14340
rect 22376 14399 22428 14408
rect 22376 14365 22385 14399
rect 22385 14365 22419 14399
rect 22419 14365 22428 14399
rect 22376 14356 22428 14365
rect 29920 14399 29972 14408
rect 29184 14288 29236 14340
rect 29920 14365 29929 14399
rect 29929 14365 29963 14399
rect 29963 14365 29972 14399
rect 29920 14356 29972 14365
rect 30288 14356 30340 14408
rect 18604 14263 18656 14272
rect 18604 14229 18613 14263
rect 18613 14229 18647 14263
rect 18647 14229 18656 14263
rect 18604 14220 18656 14229
rect 22468 14220 22520 14272
rect 28080 14220 28132 14272
rect 10880 14118 10932 14170
rect 10944 14118 10996 14170
rect 11008 14118 11060 14170
rect 11072 14118 11124 14170
rect 11136 14118 11188 14170
rect 20811 14118 20863 14170
rect 20875 14118 20927 14170
rect 20939 14118 20991 14170
rect 21003 14118 21055 14170
rect 21067 14118 21119 14170
rect 1400 14059 1452 14068
rect 1400 14025 1409 14059
rect 1409 14025 1443 14059
rect 1443 14025 1452 14059
rect 1400 14016 1452 14025
rect 4620 14059 4672 14068
rect 4620 14025 4629 14059
rect 4629 14025 4663 14059
rect 4663 14025 4672 14059
rect 4620 14016 4672 14025
rect 7564 14059 7616 14068
rect 7564 14025 7573 14059
rect 7573 14025 7607 14059
rect 7607 14025 7616 14059
rect 7564 14016 7616 14025
rect 8024 14016 8076 14068
rect 3148 13948 3200 14000
rect 3792 13948 3844 14000
rect 1952 13923 2004 13932
rect 1952 13889 1961 13923
rect 1961 13889 1995 13923
rect 1995 13889 2004 13923
rect 1952 13880 2004 13889
rect 1676 13812 1728 13864
rect 2412 13812 2464 13864
rect 4068 13923 4120 13932
rect 3332 13812 3384 13864
rect 4068 13889 4077 13923
rect 4077 13889 4111 13923
rect 4111 13889 4120 13923
rect 4068 13880 4120 13889
rect 4252 13923 4304 13932
rect 4252 13889 4261 13923
rect 4261 13889 4295 13923
rect 4295 13889 4304 13923
rect 4252 13880 4304 13889
rect 4160 13855 4212 13864
rect 4160 13821 4169 13855
rect 4169 13821 4203 13855
rect 4203 13821 4212 13855
rect 4160 13812 4212 13821
rect 6736 13880 6788 13932
rect 7012 13923 7064 13932
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7012 13880 7064 13889
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7380 13923 7432 13932
rect 7104 13880 7156 13889
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 9128 13991 9180 14000
rect 9128 13957 9137 13991
rect 9137 13957 9171 13991
rect 9171 13957 9180 13991
rect 9128 13948 9180 13957
rect 9588 14016 9640 14068
rect 17776 14016 17828 14068
rect 18604 14016 18656 14068
rect 22468 14016 22520 14068
rect 30196 14016 30248 14068
rect 9956 13948 10008 14000
rect 2964 13744 3016 13796
rect 6368 13812 6420 13864
rect 6920 13812 6972 13864
rect 7564 13812 7616 13864
rect 7932 13812 7984 13864
rect 2596 13676 2648 13728
rect 8852 13880 8904 13932
rect 9312 13923 9364 13932
rect 9312 13889 9321 13923
rect 9321 13889 9355 13923
rect 9355 13889 9364 13923
rect 9312 13880 9364 13889
rect 9588 13880 9640 13932
rect 9680 13880 9732 13932
rect 9772 13812 9824 13864
rect 10784 13880 10836 13932
rect 13268 13880 13320 13932
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13728 13923 13780 13932
rect 13360 13880 13412 13889
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 13728 13880 13780 13889
rect 14556 13923 14608 13932
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 15384 13948 15436 14000
rect 15844 13948 15896 14000
rect 15568 13923 15620 13932
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 14648 13812 14700 13864
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 19156 13948 19208 14000
rect 19340 13948 19392 14000
rect 16028 13880 16080 13932
rect 16948 13923 17000 13932
rect 16948 13889 16957 13923
rect 16957 13889 16991 13923
rect 16991 13889 17000 13923
rect 16948 13880 17000 13889
rect 17500 13923 17552 13932
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 17500 13880 17552 13889
rect 17960 13880 18012 13932
rect 18788 13880 18840 13932
rect 19524 13923 19576 13932
rect 19524 13889 19542 13923
rect 19542 13889 19576 13923
rect 19524 13880 19576 13889
rect 20536 13880 20588 13932
rect 22376 13948 22428 14000
rect 22284 13923 22336 13932
rect 22284 13889 22293 13923
rect 22293 13889 22327 13923
rect 22327 13889 22336 13923
rect 22284 13880 22336 13889
rect 28080 13880 28132 13932
rect 30288 13880 30340 13932
rect 17684 13812 17736 13864
rect 8668 13787 8720 13796
rect 8668 13753 8677 13787
rect 8677 13753 8711 13787
rect 8711 13753 8720 13787
rect 8668 13744 8720 13753
rect 8852 13744 8904 13796
rect 19984 13812 20036 13864
rect 21548 13812 21600 13864
rect 29644 13812 29696 13864
rect 8576 13676 8628 13728
rect 9128 13676 9180 13728
rect 9312 13676 9364 13728
rect 9680 13676 9732 13728
rect 10140 13676 10192 13728
rect 10324 13676 10376 13728
rect 14556 13676 14608 13728
rect 15292 13719 15344 13728
rect 15292 13685 15301 13719
rect 15301 13685 15335 13719
rect 15335 13685 15344 13719
rect 15292 13676 15344 13685
rect 18328 13676 18380 13728
rect 21824 13676 21876 13728
rect 5915 13574 5967 13626
rect 5979 13574 6031 13626
rect 6043 13574 6095 13626
rect 6107 13574 6159 13626
rect 6171 13574 6223 13626
rect 15846 13574 15898 13626
rect 15910 13574 15962 13626
rect 15974 13574 16026 13626
rect 16038 13574 16090 13626
rect 16102 13574 16154 13626
rect 25776 13574 25828 13626
rect 25840 13574 25892 13626
rect 25904 13574 25956 13626
rect 25968 13574 26020 13626
rect 26032 13574 26084 13626
rect 4252 13515 4304 13524
rect 4252 13481 4261 13515
rect 4261 13481 4295 13515
rect 4295 13481 4304 13515
rect 4252 13472 4304 13481
rect 4712 13472 4764 13524
rect 5448 13472 5500 13524
rect 7012 13404 7064 13456
rect 8484 13404 8536 13456
rect 9128 13404 9180 13456
rect 11796 13472 11848 13524
rect 15292 13472 15344 13524
rect 18052 13472 18104 13524
rect 20352 13472 20404 13524
rect 3792 13336 3844 13388
rect 5632 13336 5684 13388
rect 2596 13268 2648 13320
rect 4712 13268 4764 13320
rect 5080 13268 5132 13320
rect 4804 13200 4856 13252
rect 5908 13200 5960 13252
rect 4528 13132 4580 13184
rect 6092 13132 6144 13184
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 19892 13404 19944 13456
rect 20536 13404 20588 13456
rect 7380 13200 7432 13252
rect 8760 13200 8812 13252
rect 9588 13200 9640 13252
rect 6276 13132 6328 13184
rect 6828 13132 6880 13184
rect 8852 13132 8904 13184
rect 8944 13132 8996 13184
rect 10048 13268 10100 13320
rect 15292 13336 15344 13388
rect 15752 13336 15804 13388
rect 17224 13336 17276 13388
rect 17684 13336 17736 13388
rect 11428 13200 11480 13252
rect 12348 13268 12400 13320
rect 12624 13268 12676 13320
rect 13360 13268 13412 13320
rect 14280 13268 14332 13320
rect 15384 13311 15436 13320
rect 15384 13277 15393 13311
rect 15393 13277 15427 13311
rect 15427 13277 15436 13311
rect 15384 13268 15436 13277
rect 15016 13243 15068 13252
rect 15016 13209 15025 13243
rect 15025 13209 15059 13243
rect 15059 13209 15068 13243
rect 15016 13200 15068 13209
rect 15568 13268 15620 13320
rect 16212 13311 16264 13320
rect 16212 13277 16221 13311
rect 16221 13277 16255 13311
rect 16255 13277 16264 13311
rect 16212 13268 16264 13277
rect 17776 13311 17828 13320
rect 17776 13277 17785 13311
rect 17785 13277 17819 13311
rect 17819 13277 17828 13311
rect 17776 13268 17828 13277
rect 18236 13336 18288 13388
rect 19616 13336 19668 13388
rect 19340 13268 19392 13320
rect 19984 13268 20036 13320
rect 20260 13311 20312 13320
rect 20260 13277 20269 13311
rect 20269 13277 20303 13311
rect 20303 13277 20312 13311
rect 20260 13268 20312 13277
rect 20536 13311 20588 13320
rect 20536 13277 20545 13311
rect 20545 13277 20579 13311
rect 20579 13277 20588 13311
rect 20536 13268 20588 13277
rect 29552 13268 29604 13320
rect 29828 13311 29880 13320
rect 29828 13277 29837 13311
rect 29837 13277 29871 13311
rect 29871 13277 29880 13311
rect 29828 13268 29880 13277
rect 29920 13200 29972 13252
rect 16948 13132 17000 13184
rect 17684 13132 17736 13184
rect 30012 13175 30064 13184
rect 30012 13141 30021 13175
rect 30021 13141 30055 13175
rect 30055 13141 30064 13175
rect 30012 13132 30064 13141
rect 10880 13030 10932 13082
rect 10944 13030 10996 13082
rect 11008 13030 11060 13082
rect 11072 13030 11124 13082
rect 11136 13030 11188 13082
rect 20811 13030 20863 13082
rect 20875 13030 20927 13082
rect 20939 13030 20991 13082
rect 21003 13030 21055 13082
rect 21067 13030 21119 13082
rect 2964 12928 3016 12980
rect 4620 12971 4672 12980
rect 4620 12937 4629 12971
rect 4629 12937 4663 12971
rect 4663 12937 4672 12971
rect 4620 12928 4672 12937
rect 5172 12928 5224 12980
rect 5540 12928 5592 12980
rect 5632 12928 5684 12980
rect 7472 12928 7524 12980
rect 4988 12860 5040 12912
rect 1584 12792 1636 12844
rect 3332 12835 3384 12844
rect 3332 12801 3341 12835
rect 3341 12801 3375 12835
rect 3375 12801 3384 12835
rect 3332 12792 3384 12801
rect 3516 12835 3568 12844
rect 3516 12801 3525 12835
rect 3525 12801 3559 12835
rect 3559 12801 3568 12835
rect 3516 12792 3568 12801
rect 4528 12792 4580 12844
rect 1492 12767 1544 12776
rect 1492 12733 1501 12767
rect 1501 12733 1535 12767
rect 1535 12733 1544 12767
rect 1492 12724 1544 12733
rect 2596 12724 2648 12776
rect 4252 12724 4304 12776
rect 6828 12860 6880 12912
rect 8852 12860 8904 12912
rect 11428 12928 11480 12980
rect 12808 12971 12860 12980
rect 12808 12937 12817 12971
rect 12817 12937 12851 12971
rect 12851 12937 12860 12971
rect 12808 12928 12860 12937
rect 13728 12928 13780 12980
rect 15568 12928 15620 12980
rect 16304 12928 16356 12980
rect 6092 12792 6144 12844
rect 6368 12792 6420 12844
rect 8024 12792 8076 12844
rect 9772 12792 9824 12844
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 5172 12724 5224 12776
rect 1676 12588 1728 12640
rect 5816 12656 5868 12708
rect 5908 12656 5960 12708
rect 7932 12656 7984 12708
rect 8300 12699 8352 12708
rect 8300 12665 8309 12699
rect 8309 12665 8343 12699
rect 8343 12665 8352 12699
rect 8300 12656 8352 12665
rect 4068 12631 4120 12640
rect 4068 12597 4077 12631
rect 4077 12597 4111 12631
rect 4111 12597 4120 12631
rect 4068 12588 4120 12597
rect 7104 12588 7156 12640
rect 7748 12588 7800 12640
rect 8944 12631 8996 12640
rect 8944 12597 8953 12631
rect 8953 12597 8987 12631
rect 8987 12597 8996 12631
rect 8944 12588 8996 12597
rect 10324 12724 10376 12776
rect 10784 12656 10836 12708
rect 13268 12860 13320 12912
rect 16396 12860 16448 12912
rect 12716 12792 12768 12844
rect 13636 12835 13688 12844
rect 13636 12801 13645 12835
rect 13645 12801 13679 12835
rect 13679 12801 13688 12835
rect 13636 12792 13688 12801
rect 15016 12792 15068 12844
rect 17592 12928 17644 12980
rect 19064 12928 19116 12980
rect 19340 12928 19392 12980
rect 19800 12928 19852 12980
rect 29828 12928 29880 12980
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 17040 12835 17092 12844
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 17040 12792 17092 12801
rect 17500 12792 17552 12844
rect 17684 12835 17736 12844
rect 17684 12801 17693 12835
rect 17693 12801 17727 12835
rect 17727 12801 17736 12835
rect 17684 12792 17736 12801
rect 18420 12792 18472 12844
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 29000 12860 29052 12912
rect 18604 12792 18656 12801
rect 20168 12792 20220 12844
rect 19892 12724 19944 12776
rect 17500 12656 17552 12708
rect 20352 12835 20404 12844
rect 20352 12801 20361 12835
rect 20361 12801 20395 12835
rect 20395 12801 20404 12835
rect 20352 12792 20404 12801
rect 30288 12792 30340 12844
rect 14464 12588 14516 12640
rect 16764 12631 16816 12640
rect 16764 12597 16773 12631
rect 16773 12597 16807 12631
rect 16807 12597 16816 12631
rect 16764 12588 16816 12597
rect 17408 12588 17460 12640
rect 19524 12631 19576 12640
rect 19524 12597 19533 12631
rect 19533 12597 19567 12631
rect 19567 12597 19576 12631
rect 19524 12588 19576 12597
rect 5915 12486 5967 12538
rect 5979 12486 6031 12538
rect 6043 12486 6095 12538
rect 6107 12486 6159 12538
rect 6171 12486 6223 12538
rect 15846 12486 15898 12538
rect 15910 12486 15962 12538
rect 15974 12486 16026 12538
rect 16038 12486 16090 12538
rect 16102 12486 16154 12538
rect 25776 12486 25828 12538
rect 25840 12486 25892 12538
rect 25904 12486 25956 12538
rect 25968 12486 26020 12538
rect 26032 12486 26084 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 6552 12384 6604 12436
rect 1860 12316 1912 12368
rect 1676 12248 1728 12300
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 2964 12316 3016 12368
rect 6184 12316 6236 12368
rect 2872 12248 2924 12300
rect 3332 12248 3384 12300
rect 5724 12248 5776 12300
rect 6276 12291 6328 12300
rect 2780 12223 2832 12232
rect 2780 12189 2789 12223
rect 2789 12189 2823 12223
rect 2823 12189 2832 12223
rect 2780 12180 2832 12189
rect 4620 12180 4672 12232
rect 6276 12257 6285 12291
rect 6285 12257 6319 12291
rect 6319 12257 6328 12291
rect 6276 12248 6328 12257
rect 8024 12316 8076 12368
rect 8116 12248 8168 12300
rect 6460 12223 6512 12232
rect 4068 12155 4120 12164
rect 4068 12121 4102 12155
rect 4102 12121 4120 12155
rect 4068 12112 4120 12121
rect 5724 12112 5776 12164
rect 6460 12189 6469 12223
rect 6469 12189 6503 12223
rect 6503 12189 6512 12223
rect 6460 12180 6512 12189
rect 7104 12223 7156 12232
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 7104 12180 7156 12189
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 7656 12223 7708 12232
rect 7656 12189 7665 12223
rect 7665 12189 7699 12223
rect 7699 12189 7708 12223
rect 7656 12180 7708 12189
rect 7748 12180 7800 12232
rect 10232 12316 10284 12368
rect 9036 12248 9088 12300
rect 8300 12180 8352 12232
rect 9680 12248 9732 12300
rect 13084 12248 13136 12300
rect 6368 12112 6420 12164
rect 7564 12112 7616 12164
rect 8760 12112 8812 12164
rect 9220 12155 9272 12164
rect 9220 12121 9229 12155
rect 9229 12121 9263 12155
rect 9263 12121 9272 12155
rect 9220 12112 9272 12121
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 12440 12180 12492 12232
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 13360 12223 13412 12232
rect 9680 12112 9732 12164
rect 3516 12044 3568 12096
rect 4528 12044 4580 12096
rect 5448 12044 5500 12096
rect 10140 12087 10192 12096
rect 10140 12053 10149 12087
rect 10149 12053 10183 12087
rect 10183 12053 10192 12087
rect 10140 12044 10192 12053
rect 11244 12155 11296 12164
rect 11244 12121 11278 12155
rect 11278 12121 11296 12155
rect 11244 12112 11296 12121
rect 11520 12112 11572 12164
rect 11612 12044 11664 12096
rect 12532 12044 12584 12096
rect 12716 12112 12768 12164
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 13820 12180 13872 12232
rect 14280 12384 14332 12436
rect 14464 12384 14516 12436
rect 17224 12384 17276 12436
rect 15200 12316 15252 12368
rect 19616 12316 19668 12368
rect 16764 12248 16816 12300
rect 21180 12248 21232 12300
rect 16212 12223 16264 12232
rect 14832 12112 14884 12164
rect 14924 12112 14976 12164
rect 16212 12189 16221 12223
rect 16221 12189 16255 12223
rect 16255 12189 16264 12223
rect 16212 12180 16264 12189
rect 18236 12180 18288 12232
rect 19616 12180 19668 12232
rect 21916 12180 21968 12232
rect 29000 12180 29052 12232
rect 14556 12044 14608 12096
rect 15476 12087 15528 12096
rect 15476 12053 15485 12087
rect 15485 12053 15519 12087
rect 15519 12053 15528 12087
rect 19064 12112 19116 12164
rect 20076 12155 20128 12164
rect 20076 12121 20085 12155
rect 20085 12121 20119 12155
rect 20119 12121 20128 12155
rect 20076 12112 20128 12121
rect 29184 12112 29236 12164
rect 30288 12180 30340 12232
rect 15476 12044 15528 12053
rect 16396 12044 16448 12096
rect 18512 12044 18564 12096
rect 19800 12044 19852 12096
rect 29828 12044 29880 12096
rect 10880 11942 10932 11994
rect 10944 11942 10996 11994
rect 11008 11942 11060 11994
rect 11072 11942 11124 11994
rect 11136 11942 11188 11994
rect 20811 11942 20863 11994
rect 20875 11942 20927 11994
rect 20939 11942 20991 11994
rect 21003 11942 21055 11994
rect 21067 11942 21119 11994
rect 4988 11883 5040 11892
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 2872 11772 2924 11824
rect 4988 11849 4997 11883
rect 4997 11849 5031 11883
rect 5031 11849 5040 11883
rect 4988 11840 5040 11849
rect 5080 11840 5132 11892
rect 4620 11772 4672 11824
rect 5448 11772 5500 11824
rect 1952 11568 2004 11620
rect 2596 11568 2648 11620
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 5816 11704 5868 11756
rect 7012 11747 7064 11756
rect 7012 11713 7021 11747
rect 7021 11713 7055 11747
rect 7055 11713 7064 11747
rect 7012 11704 7064 11713
rect 7564 11747 7616 11756
rect 7564 11713 7573 11747
rect 7573 11713 7607 11747
rect 7607 11713 7616 11747
rect 7564 11704 7616 11713
rect 10048 11772 10100 11824
rect 2136 11500 2188 11552
rect 7748 11636 7800 11688
rect 10140 11704 10192 11756
rect 9956 11636 10008 11688
rect 10324 11704 10376 11756
rect 11244 11840 11296 11892
rect 12992 11840 13044 11892
rect 14188 11840 14240 11892
rect 12808 11772 12860 11824
rect 13452 11772 13504 11824
rect 17592 11840 17644 11892
rect 17868 11883 17920 11892
rect 17868 11849 17877 11883
rect 17877 11849 17911 11883
rect 17911 11849 17920 11883
rect 17868 11840 17920 11849
rect 18144 11840 18196 11892
rect 18512 11883 18564 11892
rect 18512 11849 18521 11883
rect 18521 11849 18555 11883
rect 18555 11849 18564 11883
rect 18512 11840 18564 11849
rect 20536 11883 20588 11892
rect 20536 11849 20545 11883
rect 20545 11849 20579 11883
rect 20579 11849 20588 11883
rect 20536 11840 20588 11849
rect 21180 11883 21232 11892
rect 21180 11849 21189 11883
rect 21189 11849 21223 11883
rect 21223 11849 21232 11883
rect 21180 11840 21232 11849
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 12532 11704 12584 11756
rect 13912 11704 13964 11756
rect 14280 11747 14332 11756
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 14372 11704 14424 11756
rect 11244 11636 11296 11688
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 8208 11568 8260 11620
rect 6460 11543 6512 11552
rect 6460 11509 6469 11543
rect 6469 11509 6503 11543
rect 6503 11509 6512 11543
rect 6460 11500 6512 11509
rect 7748 11543 7800 11552
rect 7748 11509 7757 11543
rect 7757 11509 7791 11543
rect 7791 11509 7800 11543
rect 7748 11500 7800 11509
rect 8024 11500 8076 11552
rect 11520 11568 11572 11620
rect 15660 11568 15712 11620
rect 16396 11568 16448 11620
rect 9404 11500 9456 11552
rect 9680 11500 9732 11552
rect 16580 11704 16632 11756
rect 18236 11772 18288 11824
rect 17684 11747 17736 11756
rect 17684 11713 17693 11747
rect 17693 11713 17727 11747
rect 17727 11713 17736 11747
rect 17684 11704 17736 11713
rect 17776 11704 17828 11756
rect 19892 11772 19944 11824
rect 19524 11704 19576 11756
rect 19984 11747 20036 11756
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 20352 11747 20404 11756
rect 20352 11713 20361 11747
rect 20361 11713 20395 11747
rect 20395 11713 20404 11747
rect 20352 11704 20404 11713
rect 21364 11704 21416 11756
rect 29184 11747 29236 11756
rect 29184 11713 29193 11747
rect 29193 11713 29227 11747
rect 29227 11713 29236 11747
rect 29184 11704 29236 11713
rect 17408 11679 17460 11688
rect 17408 11645 17417 11679
rect 17417 11645 17451 11679
rect 17451 11645 17460 11679
rect 17408 11636 17460 11645
rect 19708 11636 19760 11688
rect 20076 11679 20128 11688
rect 20076 11645 20085 11679
rect 20085 11645 20119 11679
rect 20119 11645 20128 11679
rect 20076 11636 20128 11645
rect 18052 11568 18104 11620
rect 17132 11500 17184 11552
rect 22100 11500 22152 11552
rect 30012 11543 30064 11552
rect 30012 11509 30021 11543
rect 30021 11509 30055 11543
rect 30055 11509 30064 11543
rect 30012 11500 30064 11509
rect 5915 11398 5967 11450
rect 5979 11398 6031 11450
rect 6043 11398 6095 11450
rect 6107 11398 6159 11450
rect 6171 11398 6223 11450
rect 15846 11398 15898 11450
rect 15910 11398 15962 11450
rect 15974 11398 16026 11450
rect 16038 11398 16090 11450
rect 16102 11398 16154 11450
rect 25776 11398 25828 11450
rect 25840 11398 25892 11450
rect 25904 11398 25956 11450
rect 25968 11398 26020 11450
rect 26032 11398 26084 11450
rect 5724 11296 5776 11348
rect 6276 11296 6328 11348
rect 6920 11339 6972 11348
rect 6920 11305 6929 11339
rect 6929 11305 6963 11339
rect 6963 11305 6972 11339
rect 6920 11296 6972 11305
rect 7564 11296 7616 11348
rect 7656 11296 7708 11348
rect 9404 11339 9456 11348
rect 4896 11228 4948 11280
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 11152 11296 11204 11348
rect 13084 11296 13136 11348
rect 14372 11296 14424 11348
rect 14832 11339 14884 11348
rect 14832 11305 14841 11339
rect 14841 11305 14875 11339
rect 14875 11305 14884 11339
rect 14832 11296 14884 11305
rect 16948 11296 17000 11348
rect 17684 11296 17736 11348
rect 20444 11296 20496 11348
rect 5356 11203 5408 11212
rect 5356 11169 5365 11203
rect 5365 11169 5399 11203
rect 5399 11169 5408 11203
rect 5356 11160 5408 11169
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 2872 11024 2924 11076
rect 5540 11135 5592 11144
rect 5540 11101 5585 11135
rect 5585 11101 5592 11135
rect 5540 11092 5592 11101
rect 6828 11092 6880 11144
rect 7656 11092 7708 11144
rect 7748 11092 7800 11144
rect 8208 11092 8260 11144
rect 8576 11092 8628 11144
rect 9220 11092 9272 11144
rect 9404 11092 9456 11144
rect 10784 11160 10836 11212
rect 11612 11228 11664 11280
rect 12808 11228 12860 11280
rect 11244 11203 11296 11212
rect 11244 11169 11253 11203
rect 11253 11169 11287 11203
rect 11287 11169 11296 11203
rect 11244 11160 11296 11169
rect 11520 11160 11572 11212
rect 12716 11160 12768 11212
rect 13820 11228 13872 11280
rect 13912 11228 13964 11280
rect 17040 11228 17092 11280
rect 19984 11228 20036 11280
rect 13084 11203 13136 11212
rect 13084 11169 13093 11203
rect 13093 11169 13127 11203
rect 13127 11169 13136 11203
rect 14372 11203 14424 11212
rect 13084 11160 13136 11169
rect 14372 11169 14381 11203
rect 14381 11169 14415 11203
rect 14415 11169 14424 11203
rect 14372 11160 14424 11169
rect 5356 11067 5408 11076
rect 5356 11033 5365 11067
rect 5365 11033 5399 11067
rect 5399 11033 5408 11067
rect 5356 11024 5408 11033
rect 7012 11024 7064 11076
rect 9956 11024 10008 11076
rect 1676 10956 1728 11008
rect 7472 10956 7524 11008
rect 9128 10999 9180 11008
rect 9128 10965 9137 10999
rect 9137 10965 9171 10999
rect 9171 10965 9180 10999
rect 9128 10956 9180 10965
rect 10508 11024 10560 11076
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 12164 11067 12216 11076
rect 12164 11033 12173 11067
rect 12173 11033 12207 11067
rect 12207 11033 12216 11067
rect 12164 11024 12216 11033
rect 12716 11024 12768 11076
rect 13084 11024 13136 11076
rect 13452 11092 13504 11144
rect 13912 11092 13964 11144
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 15476 11092 15528 11144
rect 15752 11092 15804 11144
rect 15200 11024 15252 11076
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16212 11135 16264 11144
rect 16028 11092 16080 11101
rect 16212 11101 16221 11135
rect 16221 11101 16255 11135
rect 16255 11101 16264 11135
rect 16212 11092 16264 11101
rect 16396 11092 16448 11144
rect 19892 11160 19944 11212
rect 17316 11092 17368 11144
rect 17960 11135 18012 11144
rect 17960 11101 17969 11135
rect 17969 11101 18003 11135
rect 18003 11101 18012 11135
rect 17960 11092 18012 11101
rect 18880 11092 18932 11144
rect 19800 11135 19852 11144
rect 19800 11101 19809 11135
rect 19809 11101 19843 11135
rect 19843 11101 19852 11135
rect 19800 11092 19852 11101
rect 11336 10956 11388 11008
rect 11888 10956 11940 11008
rect 15844 10956 15896 11008
rect 16580 10956 16632 11008
rect 17040 11067 17092 11076
rect 17040 11033 17049 11067
rect 17049 11033 17083 11067
rect 17083 11033 17092 11067
rect 17040 11024 17092 11033
rect 17132 11067 17184 11076
rect 17132 11033 17141 11067
rect 17141 11033 17175 11067
rect 17175 11033 17184 11067
rect 20076 11135 20128 11144
rect 20076 11101 20085 11135
rect 20085 11101 20119 11135
rect 20119 11101 20128 11135
rect 20076 11092 20128 11101
rect 20260 11092 20312 11144
rect 21732 11092 21784 11144
rect 17132 11024 17184 11033
rect 20720 11024 20772 11076
rect 17224 10956 17276 11008
rect 17408 10956 17460 11008
rect 10880 10854 10932 10906
rect 10944 10854 10996 10906
rect 11008 10854 11060 10906
rect 11072 10854 11124 10906
rect 11136 10854 11188 10906
rect 20811 10854 20863 10906
rect 20875 10854 20927 10906
rect 20939 10854 20991 10906
rect 21003 10854 21055 10906
rect 21067 10854 21119 10906
rect 2872 10795 2924 10804
rect 2872 10761 2881 10795
rect 2881 10761 2915 10795
rect 2915 10761 2924 10795
rect 2872 10752 2924 10761
rect 4988 10684 5040 10736
rect 5172 10684 5224 10736
rect 7288 10752 7340 10804
rect 9956 10752 10008 10804
rect 10140 10752 10192 10804
rect 11244 10752 11296 10804
rect 12164 10752 12216 10804
rect 16212 10752 16264 10804
rect 17316 10752 17368 10804
rect 17500 10795 17552 10804
rect 17500 10761 17509 10795
rect 17509 10761 17543 10795
rect 17543 10761 17552 10795
rect 17500 10752 17552 10761
rect 18052 10795 18104 10804
rect 18052 10761 18061 10795
rect 18061 10761 18095 10795
rect 18095 10761 18104 10795
rect 18052 10752 18104 10761
rect 19892 10752 19944 10804
rect 20628 10752 20680 10804
rect 20720 10752 20772 10804
rect 5816 10684 5868 10736
rect 10784 10684 10836 10736
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 2228 10616 2280 10668
rect 4896 10616 4948 10668
rect 5448 10659 5500 10668
rect 5448 10625 5462 10659
rect 5462 10625 5496 10659
rect 5496 10625 5500 10659
rect 5448 10616 5500 10625
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 7840 10616 7892 10668
rect 8852 10616 8904 10668
rect 7748 10548 7800 10600
rect 10140 10659 10192 10668
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 10324 10659 10376 10668
rect 10140 10616 10192 10625
rect 10324 10625 10333 10659
rect 10333 10625 10367 10659
rect 10367 10625 10376 10659
rect 10324 10616 10376 10625
rect 11612 10616 11664 10668
rect 15752 10684 15804 10736
rect 13084 10616 13136 10668
rect 14004 10616 14056 10668
rect 14188 10659 14240 10668
rect 14188 10625 14197 10659
rect 14197 10625 14231 10659
rect 14231 10625 14240 10659
rect 14188 10616 14240 10625
rect 15200 10659 15252 10668
rect 15200 10625 15209 10659
rect 15209 10625 15243 10659
rect 15243 10625 15252 10659
rect 15200 10616 15252 10625
rect 15660 10659 15712 10668
rect 15660 10625 15669 10659
rect 15669 10625 15703 10659
rect 15703 10625 15712 10659
rect 15660 10616 15712 10625
rect 10232 10548 10284 10600
rect 11520 10548 11572 10600
rect 15752 10591 15804 10600
rect 15752 10557 15761 10591
rect 15761 10557 15795 10591
rect 15795 10557 15804 10591
rect 15752 10548 15804 10557
rect 5264 10480 5316 10532
rect 10140 10480 10192 10532
rect 13636 10480 13688 10532
rect 14556 10480 14608 10532
rect 9680 10412 9732 10464
rect 10876 10455 10928 10464
rect 10876 10421 10885 10455
rect 10885 10421 10919 10455
rect 10919 10421 10928 10455
rect 10876 10412 10928 10421
rect 13452 10412 13504 10464
rect 16672 10616 16724 10668
rect 16948 10659 17000 10668
rect 16948 10625 16957 10659
rect 16957 10625 16991 10659
rect 16991 10625 17000 10659
rect 16948 10616 17000 10625
rect 17224 10616 17276 10668
rect 17500 10616 17552 10668
rect 17592 10616 17644 10668
rect 18788 10659 18840 10668
rect 18788 10625 18797 10659
rect 18797 10625 18831 10659
rect 18831 10625 18840 10659
rect 18788 10616 18840 10625
rect 19892 10659 19944 10668
rect 19892 10625 19901 10659
rect 19901 10625 19935 10659
rect 19935 10625 19944 10659
rect 19892 10616 19944 10625
rect 20260 10659 20312 10668
rect 20260 10625 20269 10659
rect 20269 10625 20303 10659
rect 20303 10625 20312 10659
rect 20260 10616 20312 10625
rect 21180 10616 21232 10668
rect 16028 10480 16080 10532
rect 20076 10480 20128 10532
rect 17868 10412 17920 10464
rect 19064 10455 19116 10464
rect 19064 10421 19073 10455
rect 19073 10421 19107 10455
rect 19107 10421 19116 10455
rect 19064 10412 19116 10421
rect 5915 10310 5967 10362
rect 5979 10310 6031 10362
rect 6043 10310 6095 10362
rect 6107 10310 6159 10362
rect 6171 10310 6223 10362
rect 15846 10310 15898 10362
rect 15910 10310 15962 10362
rect 15974 10310 16026 10362
rect 16038 10310 16090 10362
rect 16102 10310 16154 10362
rect 25776 10310 25828 10362
rect 25840 10310 25892 10362
rect 25904 10310 25956 10362
rect 25968 10310 26020 10362
rect 26032 10310 26084 10362
rect 2228 10251 2280 10260
rect 2228 10217 2237 10251
rect 2237 10217 2271 10251
rect 2271 10217 2280 10251
rect 2228 10208 2280 10217
rect 9496 10208 9548 10260
rect 11612 10251 11664 10260
rect 11612 10217 11621 10251
rect 11621 10217 11655 10251
rect 11655 10217 11664 10251
rect 11612 10208 11664 10217
rect 1492 10140 1544 10192
rect 1952 10072 2004 10124
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2872 10072 2924 10124
rect 6644 10072 6696 10124
rect 10048 10072 10100 10124
rect 2780 10004 2832 10056
rect 5816 10004 5868 10056
rect 6828 10004 6880 10056
rect 3332 9936 3384 9988
rect 6000 9979 6052 9988
rect 6000 9945 6009 9979
rect 6009 9945 6043 9979
rect 6043 9945 6052 9979
rect 6000 9936 6052 9945
rect 2688 9868 2740 9920
rect 2872 9911 2924 9920
rect 2872 9877 2881 9911
rect 2881 9877 2915 9911
rect 2915 9877 2924 9911
rect 2872 9868 2924 9877
rect 3148 9868 3200 9920
rect 4988 9868 5040 9920
rect 5264 9868 5316 9920
rect 6460 9868 6512 9920
rect 7656 9979 7708 9988
rect 7656 9945 7665 9979
rect 7665 9945 7699 9979
rect 7699 9945 7708 9979
rect 7656 9936 7708 9945
rect 9680 9979 9732 9988
rect 9680 9945 9689 9979
rect 9689 9945 9723 9979
rect 9723 9945 9732 9979
rect 9680 9936 9732 9945
rect 10876 10004 10928 10056
rect 12440 10208 12492 10260
rect 12716 10208 12768 10260
rect 13452 10251 13504 10260
rect 13452 10217 13461 10251
rect 13461 10217 13495 10251
rect 13495 10217 13504 10251
rect 13452 10208 13504 10217
rect 17500 10251 17552 10260
rect 11888 10072 11940 10124
rect 12624 9936 12676 9988
rect 14004 10072 14056 10124
rect 14464 10115 14516 10124
rect 14464 10081 14473 10115
rect 14473 10081 14507 10115
rect 14507 10081 14516 10115
rect 14464 10072 14516 10081
rect 13912 10004 13964 10056
rect 10232 9868 10284 9920
rect 11612 9868 11664 9920
rect 13544 9868 13596 9920
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14648 10047 14700 10056
rect 14372 10004 14424 10013
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 15016 10004 15068 10056
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 19892 10208 19944 10260
rect 18236 10140 18288 10192
rect 16672 10115 16724 10124
rect 16672 10081 16681 10115
rect 16681 10081 16715 10115
rect 16715 10081 16724 10115
rect 16672 10072 16724 10081
rect 17316 10072 17368 10124
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 18696 10072 18748 10124
rect 28632 10208 28684 10260
rect 18788 10004 18840 10056
rect 19248 10004 19300 10056
rect 20720 10004 20772 10056
rect 21824 10004 21876 10056
rect 29828 10047 29880 10056
rect 29828 10013 29837 10047
rect 29837 10013 29871 10047
rect 29871 10013 29880 10047
rect 29828 10004 29880 10013
rect 14556 9936 14608 9988
rect 15568 9979 15620 9988
rect 15568 9945 15577 9979
rect 15577 9945 15611 9979
rect 15611 9945 15620 9979
rect 15568 9936 15620 9945
rect 16396 9979 16448 9988
rect 16396 9945 16405 9979
rect 16405 9945 16439 9979
rect 16439 9945 16448 9979
rect 16396 9936 16448 9945
rect 14832 9911 14884 9920
rect 14832 9877 14841 9911
rect 14841 9877 14875 9911
rect 14875 9877 14884 9911
rect 14832 9868 14884 9877
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 22560 9936 22612 9988
rect 21272 9868 21324 9920
rect 30012 9911 30064 9920
rect 30012 9877 30021 9911
rect 30021 9877 30055 9911
rect 30055 9877 30064 9911
rect 30012 9868 30064 9877
rect 10880 9766 10932 9818
rect 10944 9766 10996 9818
rect 11008 9766 11060 9818
rect 11072 9766 11124 9818
rect 11136 9766 11188 9818
rect 20811 9766 20863 9818
rect 20875 9766 20927 9818
rect 20939 9766 20991 9818
rect 21003 9766 21055 9818
rect 21067 9766 21119 9818
rect 3332 9707 3384 9716
rect 3332 9673 3341 9707
rect 3341 9673 3375 9707
rect 3375 9673 3384 9707
rect 3332 9664 3384 9673
rect 4436 9664 4488 9716
rect 6000 9664 6052 9716
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 1492 9528 1544 9580
rect 2320 9528 2372 9580
rect 2872 9596 2924 9648
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3516 9528 3568 9580
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 10508 9664 10560 9716
rect 12348 9664 12400 9716
rect 14464 9664 14516 9716
rect 7656 9596 7708 9648
rect 10784 9596 10836 9648
rect 13176 9596 13228 9648
rect 13268 9596 13320 9648
rect 13912 9596 13964 9648
rect 14740 9596 14792 9648
rect 4804 9528 4856 9580
rect 5356 9528 5408 9580
rect 5448 9571 5500 9580
rect 5448 9537 5457 9571
rect 5457 9537 5491 9571
rect 5491 9537 5500 9571
rect 5448 9528 5500 9537
rect 2596 9392 2648 9444
rect 2688 9392 2740 9444
rect 4252 9392 4304 9444
rect 5080 9460 5132 9512
rect 6460 9460 6512 9512
rect 6828 9528 6880 9580
rect 7472 9528 7524 9580
rect 8944 9528 8996 9580
rect 9496 9528 9548 9580
rect 10048 9528 10100 9580
rect 8300 9503 8352 9512
rect 8300 9469 8309 9503
rect 8309 9469 8343 9503
rect 8343 9469 8352 9503
rect 8300 9460 8352 9469
rect 9680 9460 9732 9512
rect 2504 9324 2556 9376
rect 2780 9324 2832 9376
rect 6736 9392 6788 9444
rect 12348 9460 12400 9512
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 14556 9460 14608 9512
rect 15292 9664 15344 9716
rect 15660 9596 15712 9648
rect 18420 9664 18472 9716
rect 19248 9707 19300 9716
rect 19248 9673 19257 9707
rect 19257 9673 19291 9707
rect 19291 9673 19300 9707
rect 19248 9664 19300 9673
rect 20260 9664 20312 9716
rect 15476 9571 15528 9580
rect 15476 9537 15485 9571
rect 15485 9537 15519 9571
rect 15519 9537 15528 9571
rect 15476 9528 15528 9537
rect 13268 9392 13320 9444
rect 4620 9324 4672 9376
rect 4988 9324 5040 9376
rect 8668 9324 8720 9376
rect 14648 9324 14700 9376
rect 14832 9324 14884 9376
rect 15660 9460 15712 9512
rect 15108 9392 15160 9444
rect 16948 9460 17000 9512
rect 17040 9460 17092 9512
rect 18144 9571 18196 9580
rect 18144 9537 18178 9571
rect 18178 9537 18196 9571
rect 18144 9528 18196 9537
rect 16212 9324 16264 9376
rect 21916 9528 21968 9580
rect 21824 9503 21876 9512
rect 21824 9469 21833 9503
rect 21833 9469 21867 9503
rect 21867 9469 21876 9503
rect 21824 9460 21876 9469
rect 22008 9324 22060 9376
rect 5915 9222 5967 9274
rect 5979 9222 6031 9274
rect 6043 9222 6095 9274
rect 6107 9222 6159 9274
rect 6171 9222 6223 9274
rect 15846 9222 15898 9274
rect 15910 9222 15962 9274
rect 15974 9222 16026 9274
rect 16038 9222 16090 9274
rect 16102 9222 16154 9274
rect 25776 9222 25828 9274
rect 25840 9222 25892 9274
rect 25904 9222 25956 9274
rect 25968 9222 26020 9274
rect 26032 9222 26084 9274
rect 2688 9027 2740 9036
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 2688 8984 2740 8993
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 5264 9120 5316 9172
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 10232 9163 10284 9172
rect 10232 9129 10241 9163
rect 10241 9129 10275 9163
rect 10275 9129 10284 9163
rect 10232 9120 10284 9129
rect 3608 8984 3660 9036
rect 2596 8916 2648 8925
rect 1492 8848 1544 8900
rect 8300 8916 8352 8968
rect 8668 8916 8720 8968
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 9680 8984 9732 9036
rect 10232 8984 10284 9036
rect 9496 8959 9548 8968
rect 3884 8848 3936 8900
rect 1676 8780 1728 8832
rect 4344 8848 4396 8900
rect 4988 8848 5040 8900
rect 5448 8848 5500 8900
rect 6368 8848 6420 8900
rect 6644 8848 6696 8900
rect 7196 8848 7248 8900
rect 9220 8848 9272 8900
rect 9496 8925 9505 8959
rect 9505 8925 9539 8959
rect 9539 8925 9548 8959
rect 9496 8916 9548 8925
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 10508 8916 10560 8968
rect 12440 8984 12492 9036
rect 11612 8959 11664 8968
rect 11612 8925 11621 8959
rect 11621 8925 11655 8959
rect 11655 8925 11664 8959
rect 11612 8916 11664 8925
rect 6736 8780 6788 8832
rect 6920 8780 6972 8832
rect 7380 8780 7432 8832
rect 10784 8780 10836 8832
rect 11520 8823 11572 8832
rect 11520 8789 11529 8823
rect 11529 8789 11563 8823
rect 11563 8789 11572 8823
rect 11520 8780 11572 8789
rect 14372 8916 14424 8968
rect 16672 9120 16724 9172
rect 20168 9120 20220 9172
rect 20352 9120 20404 9172
rect 21916 9163 21968 9172
rect 21916 9129 21925 9163
rect 21925 9129 21959 9163
rect 21959 9129 21968 9163
rect 21916 9120 21968 9129
rect 17776 9052 17828 9104
rect 17868 9052 17920 9104
rect 19248 8984 19300 9036
rect 15568 8916 15620 8968
rect 17960 8916 18012 8968
rect 14096 8848 14148 8900
rect 14648 8848 14700 8900
rect 15476 8780 15528 8832
rect 17684 8848 17736 8900
rect 17040 8823 17092 8832
rect 17040 8789 17049 8823
rect 17049 8789 17083 8823
rect 17083 8789 17092 8823
rect 17040 8780 17092 8789
rect 18328 8916 18380 8968
rect 21640 8984 21692 9036
rect 21548 8959 21600 8968
rect 19156 8848 19208 8900
rect 18144 8780 18196 8832
rect 18236 8780 18288 8832
rect 18420 8780 18472 8832
rect 18788 8780 18840 8832
rect 21548 8925 21557 8959
rect 21557 8925 21591 8959
rect 21591 8925 21600 8959
rect 21548 8916 21600 8925
rect 22008 9052 22060 9104
rect 22008 8848 22060 8900
rect 21548 8780 21600 8832
rect 10880 8678 10932 8730
rect 10944 8678 10996 8730
rect 11008 8678 11060 8730
rect 11072 8678 11124 8730
rect 11136 8678 11188 8730
rect 20811 8678 20863 8730
rect 20875 8678 20927 8730
rect 20939 8678 20991 8730
rect 21003 8678 21055 8730
rect 21067 8678 21119 8730
rect 2780 8619 2832 8628
rect 2780 8585 2789 8619
rect 2789 8585 2823 8619
rect 2823 8585 2832 8619
rect 2780 8576 2832 8585
rect 4804 8576 4856 8628
rect 6644 8576 6696 8628
rect 2688 8508 2740 8560
rect 1492 8440 1544 8492
rect 2228 8440 2280 8492
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 3884 8440 3936 8492
rect 5540 8508 5592 8560
rect 6828 8508 6880 8560
rect 4620 8483 4672 8492
rect 4620 8449 4654 8483
rect 4654 8449 4672 8483
rect 4620 8440 4672 8449
rect 6276 8440 6328 8492
rect 3700 8236 3752 8288
rect 6920 8440 6972 8492
rect 7196 8551 7248 8560
rect 7196 8517 7205 8551
rect 7205 8517 7239 8551
rect 7239 8517 7248 8551
rect 7840 8551 7892 8560
rect 7196 8508 7248 8517
rect 7840 8517 7849 8551
rect 7849 8517 7883 8551
rect 7883 8517 7892 8551
rect 7840 8508 7892 8517
rect 10324 8576 10376 8628
rect 11520 8576 11572 8628
rect 14096 8619 14148 8628
rect 8484 8440 8536 8492
rect 8944 8440 8996 8492
rect 11796 8508 11848 8560
rect 14096 8585 14105 8619
rect 14105 8585 14139 8619
rect 14139 8585 14148 8619
rect 14096 8576 14148 8585
rect 16856 8576 16908 8628
rect 18144 8576 18196 8628
rect 19616 8576 19668 8628
rect 22560 8619 22612 8628
rect 22560 8585 22569 8619
rect 22569 8585 22603 8619
rect 22603 8585 22612 8619
rect 22560 8576 22612 8585
rect 14556 8508 14608 8560
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 13268 8440 13320 8492
rect 13820 8440 13872 8492
rect 14648 8440 14700 8492
rect 14832 8483 14884 8492
rect 14832 8449 14866 8483
rect 14866 8449 14884 8483
rect 14832 8440 14884 8449
rect 17040 8508 17092 8560
rect 21272 8508 21324 8560
rect 16764 8440 16816 8492
rect 18788 8483 18840 8492
rect 18788 8449 18797 8483
rect 18797 8449 18831 8483
rect 18831 8449 18840 8483
rect 18788 8440 18840 8449
rect 21548 8440 21600 8492
rect 22284 8440 22336 8492
rect 29644 8440 29696 8492
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 10140 8372 10192 8424
rect 10324 8372 10376 8424
rect 12072 8415 12124 8424
rect 12072 8381 12081 8415
rect 12081 8381 12115 8415
rect 12115 8381 12124 8415
rect 12072 8372 12124 8381
rect 7656 8347 7708 8356
rect 7656 8313 7665 8347
rect 7665 8313 7699 8347
rect 7699 8313 7708 8347
rect 7656 8304 7708 8313
rect 11336 8304 11388 8356
rect 6828 8236 6880 8288
rect 7012 8236 7064 8288
rect 10416 8236 10468 8288
rect 10692 8236 10744 8288
rect 10968 8236 11020 8288
rect 14464 8372 14516 8424
rect 14556 8415 14608 8424
rect 14556 8381 14565 8415
rect 14565 8381 14599 8415
rect 14599 8381 14608 8415
rect 14556 8372 14608 8381
rect 17776 8372 17828 8424
rect 21456 8372 21508 8424
rect 21640 8372 21692 8424
rect 21916 8372 21968 8424
rect 16212 8304 16264 8356
rect 30012 8347 30064 8356
rect 30012 8313 30021 8347
rect 30021 8313 30055 8347
rect 30055 8313 30064 8347
rect 30012 8304 30064 8313
rect 15660 8236 15712 8288
rect 16488 8236 16540 8288
rect 19156 8236 19208 8288
rect 5915 8134 5967 8186
rect 5979 8134 6031 8186
rect 6043 8134 6095 8186
rect 6107 8134 6159 8186
rect 6171 8134 6223 8186
rect 15846 8134 15898 8186
rect 15910 8134 15962 8186
rect 15974 8134 16026 8186
rect 16038 8134 16090 8186
rect 16102 8134 16154 8186
rect 25776 8134 25828 8186
rect 25840 8134 25892 8186
rect 25904 8134 25956 8186
rect 25968 8134 26020 8186
rect 26032 8134 26084 8186
rect 1584 8032 1636 8084
rect 2320 8032 2372 8084
rect 8852 8032 8904 8084
rect 13360 8032 13412 8084
rect 16764 8032 16816 8084
rect 21180 8032 21232 8084
rect 21456 8032 21508 8084
rect 9220 7964 9272 8016
rect 9588 7964 9640 8016
rect 2412 7939 2464 7948
rect 2412 7905 2421 7939
rect 2421 7905 2455 7939
rect 2455 7905 2464 7939
rect 2412 7896 2464 7905
rect 10508 7896 10560 7948
rect 10784 7896 10836 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 3792 7828 3844 7880
rect 1860 7692 1912 7744
rect 4160 7760 4212 7812
rect 4344 7828 4396 7880
rect 6276 7828 6328 7880
rect 4436 7760 4488 7812
rect 5448 7760 5500 7812
rect 7196 7760 7248 7812
rect 10140 7828 10192 7880
rect 6920 7692 6972 7744
rect 7656 7692 7708 7744
rect 10692 7760 10744 7812
rect 17960 7964 18012 8016
rect 12072 7896 12124 7948
rect 13176 7896 13228 7948
rect 15568 7896 15620 7948
rect 21916 7964 21968 8016
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 11796 7828 11848 7880
rect 11336 7760 11388 7812
rect 12348 7828 12400 7880
rect 12532 7760 12584 7812
rect 13360 7828 13412 7880
rect 15476 7828 15528 7880
rect 15752 7828 15804 7880
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 16488 7828 16540 7880
rect 16856 7828 16908 7880
rect 18052 7828 18104 7880
rect 19800 7828 19852 7880
rect 21548 7871 21600 7880
rect 21548 7837 21557 7871
rect 21557 7837 21591 7871
rect 21591 7837 21600 7871
rect 21548 7828 21600 7837
rect 17500 7760 17552 7812
rect 20076 7760 20128 7812
rect 12164 7735 12216 7744
rect 12164 7701 12173 7735
rect 12173 7701 12207 7735
rect 12207 7701 12216 7735
rect 13452 7735 13504 7744
rect 12164 7692 12216 7701
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 14924 7692 14976 7744
rect 15292 7692 15344 7744
rect 22100 7871 22152 7880
rect 22100 7837 22109 7871
rect 22109 7837 22143 7871
rect 22143 7837 22152 7871
rect 22100 7828 22152 7837
rect 22100 7692 22152 7744
rect 22284 7735 22336 7744
rect 22284 7701 22293 7735
rect 22293 7701 22327 7735
rect 22327 7701 22336 7735
rect 22284 7692 22336 7701
rect 10880 7590 10932 7642
rect 10944 7590 10996 7642
rect 11008 7590 11060 7642
rect 11072 7590 11124 7642
rect 11136 7590 11188 7642
rect 20811 7590 20863 7642
rect 20875 7590 20927 7642
rect 20939 7590 20991 7642
rect 21003 7590 21055 7642
rect 21067 7590 21119 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 6920 7488 6972 7540
rect 7012 7488 7064 7540
rect 7380 7488 7432 7540
rect 9772 7488 9824 7540
rect 11888 7488 11940 7540
rect 13452 7531 13504 7540
rect 13452 7497 13461 7531
rect 13461 7497 13495 7531
rect 13495 7497 13504 7531
rect 13452 7488 13504 7497
rect 14280 7488 14332 7540
rect 22192 7488 22244 7540
rect 1584 7420 1636 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 2596 7420 2648 7472
rect 4252 7420 4304 7472
rect 5540 7463 5592 7472
rect 2780 7352 2832 7404
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 4344 7352 4396 7404
rect 5540 7429 5549 7463
rect 5549 7429 5583 7463
rect 5583 7429 5592 7463
rect 5540 7420 5592 7429
rect 6276 7352 6328 7404
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 8484 7395 8536 7404
rect 8484 7361 8493 7395
rect 8493 7361 8527 7395
rect 8527 7361 8536 7395
rect 8484 7352 8536 7361
rect 8576 7352 8628 7404
rect 9680 7420 9732 7472
rect 10232 7352 10284 7404
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 10692 7352 10744 7404
rect 10784 7352 10836 7404
rect 11612 7352 11664 7404
rect 12348 7352 12400 7404
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 13912 7352 13964 7404
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 2688 7284 2740 7336
rect 5264 7284 5316 7336
rect 6828 7284 6880 7336
rect 7196 7284 7248 7336
rect 9220 7284 9272 7336
rect 11336 7284 11388 7336
rect 12532 7284 12584 7336
rect 13176 7327 13228 7336
rect 13176 7293 13185 7327
rect 13185 7293 13219 7327
rect 13219 7293 13228 7327
rect 13176 7284 13228 7293
rect 13360 7327 13412 7336
rect 13360 7293 13369 7327
rect 13369 7293 13403 7327
rect 13403 7293 13412 7327
rect 13360 7284 13412 7293
rect 18144 7420 18196 7472
rect 18420 7420 18472 7472
rect 22284 7420 22336 7472
rect 15384 7352 15436 7404
rect 15016 7284 15068 7336
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 16672 7352 16724 7404
rect 17960 7395 18012 7404
rect 17960 7361 17969 7395
rect 17969 7361 18003 7395
rect 18003 7361 18012 7395
rect 17960 7352 18012 7361
rect 29828 7395 29880 7404
rect 29828 7361 29837 7395
rect 29837 7361 29871 7395
rect 29871 7361 29880 7395
rect 29828 7352 29880 7361
rect 8116 7148 8168 7200
rect 9220 7191 9272 7200
rect 9220 7157 9229 7191
rect 9229 7157 9263 7191
rect 9263 7157 9272 7191
rect 9220 7148 9272 7157
rect 10508 7191 10560 7200
rect 10508 7157 10517 7191
rect 10517 7157 10551 7191
rect 10551 7157 10560 7191
rect 10508 7148 10560 7157
rect 12624 7191 12676 7200
rect 12624 7157 12633 7191
rect 12633 7157 12667 7191
rect 12667 7157 12676 7191
rect 12624 7148 12676 7157
rect 15384 7148 15436 7200
rect 16028 7284 16080 7336
rect 16948 7284 17000 7336
rect 19432 7327 19484 7336
rect 19432 7293 19441 7327
rect 19441 7293 19475 7327
rect 19475 7293 19484 7327
rect 19432 7284 19484 7293
rect 19616 7284 19668 7336
rect 20628 7284 20680 7336
rect 21640 7284 21692 7336
rect 21824 7327 21876 7336
rect 21824 7293 21833 7327
rect 21833 7293 21867 7327
rect 21867 7293 21876 7327
rect 21824 7284 21876 7293
rect 15752 7148 15804 7200
rect 18328 7148 18380 7200
rect 21272 7148 21324 7200
rect 30012 7191 30064 7200
rect 30012 7157 30021 7191
rect 30021 7157 30055 7191
rect 30055 7157 30064 7191
rect 30012 7148 30064 7157
rect 5915 7046 5967 7098
rect 5979 7046 6031 7098
rect 6043 7046 6095 7098
rect 6107 7046 6159 7098
rect 6171 7046 6223 7098
rect 15846 7046 15898 7098
rect 15910 7046 15962 7098
rect 15974 7046 16026 7098
rect 16038 7046 16090 7098
rect 16102 7046 16154 7098
rect 25776 7046 25828 7098
rect 25840 7046 25892 7098
rect 25904 7046 25956 7098
rect 25968 7046 26020 7098
rect 26032 7046 26084 7098
rect 4160 6944 4212 6996
rect 7012 6987 7064 6996
rect 7012 6953 7021 6987
rect 7021 6953 7055 6987
rect 7055 6953 7064 6987
rect 7012 6944 7064 6953
rect 7288 6944 7340 6996
rect 9312 6944 9364 6996
rect 3792 6876 3844 6928
rect 10232 6944 10284 6996
rect 18328 6944 18380 6996
rect 20076 6987 20128 6996
rect 20076 6953 20085 6987
rect 20085 6953 20119 6987
rect 20119 6953 20128 6987
rect 20076 6944 20128 6953
rect 29828 6944 29880 6996
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 5448 6808 5500 6860
rect 1584 6740 1636 6792
rect 1860 6783 1912 6792
rect 1860 6749 1869 6783
rect 1869 6749 1903 6783
rect 1903 6749 1912 6783
rect 1860 6740 1912 6749
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 3516 6740 3568 6792
rect 3884 6740 3936 6792
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 2596 6672 2648 6724
rect 2412 6647 2464 6656
rect 2412 6613 2421 6647
rect 2421 6613 2455 6647
rect 2455 6613 2464 6647
rect 2412 6604 2464 6613
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 4528 6647 4580 6656
rect 4528 6613 4537 6647
rect 4537 6613 4571 6647
rect 4571 6613 4580 6647
rect 4528 6604 4580 6613
rect 6552 6808 6604 6860
rect 15476 6876 15528 6928
rect 16212 6876 16264 6928
rect 18144 6919 18196 6928
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 6920 6672 6972 6724
rect 12072 6808 12124 6860
rect 12716 6808 12768 6860
rect 15568 6808 15620 6860
rect 8116 6783 8168 6792
rect 8116 6749 8134 6783
rect 8134 6749 8168 6783
rect 8116 6740 8168 6749
rect 8668 6740 8720 6792
rect 9220 6783 9272 6792
rect 9220 6749 9254 6783
rect 9254 6749 9272 6783
rect 9220 6740 9272 6749
rect 12624 6740 12676 6792
rect 6828 6604 6880 6656
rect 10416 6604 10468 6656
rect 14832 6672 14884 6724
rect 18144 6885 18153 6919
rect 18153 6885 18187 6919
rect 18187 6885 18196 6919
rect 18144 6876 18196 6885
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 19616 6851 19668 6860
rect 19616 6817 19625 6851
rect 19625 6817 19659 6851
rect 19659 6817 19668 6851
rect 19616 6808 19668 6817
rect 19800 6808 19852 6860
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 16764 6740 16816 6749
rect 16856 6783 16908 6792
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 16856 6740 16908 6749
rect 17408 6740 17460 6792
rect 17500 6740 17552 6792
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 19432 6672 19484 6724
rect 12072 6604 12124 6656
rect 12256 6604 12308 6656
rect 12440 6647 12492 6656
rect 12440 6613 12449 6647
rect 12449 6613 12483 6647
rect 12483 6613 12492 6647
rect 12440 6604 12492 6613
rect 12808 6604 12860 6656
rect 13544 6604 13596 6656
rect 13636 6604 13688 6656
rect 15292 6604 15344 6656
rect 15476 6604 15528 6656
rect 17316 6647 17368 6656
rect 17316 6613 17325 6647
rect 17325 6613 17359 6647
rect 17359 6613 17368 6647
rect 17316 6604 17368 6613
rect 21088 6740 21140 6792
rect 29644 6740 29696 6792
rect 30104 6783 30156 6792
rect 30104 6749 30113 6783
rect 30113 6749 30147 6783
rect 30147 6749 30156 6783
rect 30104 6740 30156 6749
rect 21180 6672 21232 6724
rect 21272 6604 21324 6656
rect 21732 6604 21784 6656
rect 10880 6502 10932 6554
rect 10944 6502 10996 6554
rect 11008 6502 11060 6554
rect 11072 6502 11124 6554
rect 11136 6502 11188 6554
rect 20811 6502 20863 6554
rect 20875 6502 20927 6554
rect 20939 6502 20991 6554
rect 21003 6502 21055 6554
rect 21067 6502 21119 6554
rect 2228 6400 2280 6452
rect 1492 6332 1544 6384
rect 2412 6264 2464 6316
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 4344 6400 4396 6452
rect 4528 6332 4580 6384
rect 6920 6400 6972 6452
rect 7748 6400 7800 6452
rect 12164 6400 12216 6452
rect 12256 6400 12308 6452
rect 7656 6332 7708 6384
rect 10968 6332 11020 6384
rect 13636 6332 13688 6384
rect 6184 6264 6236 6316
rect 6460 6307 6512 6316
rect 6460 6273 6464 6307
rect 6464 6273 6498 6307
rect 6498 6273 6512 6307
rect 6460 6264 6512 6273
rect 7012 6264 7064 6316
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 9680 6264 9732 6316
rect 10416 6264 10468 6316
rect 11796 6264 11848 6316
rect 12348 6307 12400 6316
rect 3240 6060 3292 6112
rect 7932 6128 7984 6180
rect 12348 6273 12357 6307
rect 12357 6273 12391 6307
rect 12391 6273 12400 6307
rect 12348 6264 12400 6273
rect 14372 6307 14424 6316
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 14648 6307 14700 6316
rect 14648 6273 14682 6307
rect 14682 6273 14700 6307
rect 15200 6400 15252 6452
rect 17408 6400 17460 6452
rect 18052 6400 18104 6452
rect 18880 6400 18932 6452
rect 19248 6400 19300 6452
rect 15108 6332 15160 6384
rect 14648 6264 14700 6273
rect 16304 6264 16356 6316
rect 17316 6264 17368 6316
rect 19340 6332 19392 6384
rect 19800 6332 19852 6384
rect 18236 6264 18288 6316
rect 21180 6400 21232 6452
rect 20536 6307 20588 6316
rect 20536 6273 20545 6307
rect 20545 6273 20579 6307
rect 20579 6273 20588 6307
rect 20536 6264 20588 6273
rect 20628 6307 20680 6316
rect 20628 6273 20637 6307
rect 20637 6273 20671 6307
rect 20671 6273 20680 6307
rect 20628 6264 20680 6273
rect 21732 6264 21784 6316
rect 12624 6128 12676 6180
rect 13728 6196 13780 6248
rect 13912 6239 13964 6248
rect 13912 6205 13921 6239
rect 13921 6205 13955 6239
rect 13955 6205 13964 6239
rect 13912 6196 13964 6205
rect 20444 6196 20496 6248
rect 21272 6196 21324 6248
rect 6368 6060 6420 6112
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 12440 6060 12492 6112
rect 13268 6060 13320 6112
rect 30104 6060 30156 6112
rect 5915 5958 5967 6010
rect 5979 5958 6031 6010
rect 6043 5958 6095 6010
rect 6107 5958 6159 6010
rect 6171 5958 6223 6010
rect 15846 5958 15898 6010
rect 15910 5958 15962 6010
rect 15974 5958 16026 6010
rect 16038 5958 16090 6010
rect 16102 5958 16154 6010
rect 25776 5958 25828 6010
rect 25840 5958 25892 6010
rect 25904 5958 25956 6010
rect 25968 5958 26020 6010
rect 26032 5958 26084 6010
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 5724 5856 5776 5908
rect 11336 5856 11388 5908
rect 13360 5856 13412 5908
rect 16672 5856 16724 5908
rect 18236 5899 18288 5908
rect 18236 5865 18245 5899
rect 18245 5865 18279 5899
rect 18279 5865 18288 5899
rect 18236 5856 18288 5865
rect 19708 5856 19760 5908
rect 29460 5856 29512 5908
rect 29828 5899 29880 5908
rect 29828 5865 29837 5899
rect 29837 5865 29871 5899
rect 29871 5865 29880 5899
rect 29828 5856 29880 5865
rect 1492 5720 1544 5772
rect 3976 5720 4028 5772
rect 6736 5788 6788 5840
rect 11980 5831 12032 5840
rect 11980 5797 11989 5831
rect 11989 5797 12023 5831
rect 12023 5797 12032 5831
rect 11980 5788 12032 5797
rect 12348 5788 12400 5840
rect 12256 5720 12308 5772
rect 12716 5720 12768 5772
rect 14372 5788 14424 5840
rect 15108 5720 15160 5772
rect 16948 5720 17000 5772
rect 19432 5720 19484 5772
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 2688 5584 2740 5636
rect 4712 5584 4764 5636
rect 6368 5584 6420 5636
rect 6644 5695 6696 5704
rect 6644 5661 6653 5695
rect 6653 5661 6687 5695
rect 6687 5661 6696 5695
rect 6828 5695 6880 5704
rect 6644 5652 6696 5661
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 8392 5584 8444 5636
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 13268 5652 13320 5704
rect 10232 5627 10284 5636
rect 10232 5593 10241 5627
rect 10241 5593 10275 5627
rect 10275 5593 10284 5627
rect 10232 5584 10284 5593
rect 10600 5627 10652 5636
rect 10600 5593 10609 5627
rect 10609 5593 10643 5627
rect 10643 5593 10652 5627
rect 10600 5584 10652 5593
rect 10968 5627 11020 5636
rect 10968 5593 10977 5627
rect 10977 5593 11011 5627
rect 11011 5593 11020 5627
rect 10968 5584 11020 5593
rect 11428 5584 11480 5636
rect 11796 5584 11848 5636
rect 12808 5584 12860 5636
rect 13452 5652 13504 5704
rect 13728 5652 13780 5704
rect 15752 5652 15804 5704
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 17684 5695 17736 5704
rect 17684 5661 17693 5695
rect 17693 5661 17727 5695
rect 17727 5661 17736 5695
rect 17684 5652 17736 5661
rect 18052 5695 18104 5704
rect 10784 5516 10836 5568
rect 12348 5559 12400 5568
rect 12348 5525 12357 5559
rect 12357 5525 12391 5559
rect 12391 5525 12400 5559
rect 12348 5516 12400 5525
rect 13268 5516 13320 5568
rect 16856 5584 16908 5636
rect 18052 5661 18061 5695
rect 18061 5661 18095 5695
rect 18095 5661 18104 5695
rect 18052 5652 18104 5661
rect 20720 5695 20772 5704
rect 18236 5584 18288 5636
rect 20720 5661 20729 5695
rect 20729 5661 20763 5695
rect 20763 5661 20772 5695
rect 20720 5652 20772 5661
rect 29736 5652 29788 5704
rect 19708 5584 19760 5636
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 10880 5414 10932 5466
rect 10944 5414 10996 5466
rect 11008 5414 11060 5466
rect 11072 5414 11124 5466
rect 11136 5414 11188 5466
rect 20811 5414 20863 5466
rect 20875 5414 20927 5466
rect 20939 5414 20991 5466
rect 21003 5414 21055 5466
rect 21067 5414 21119 5466
rect 2688 5355 2740 5364
rect 2688 5321 2697 5355
rect 2697 5321 2731 5355
rect 2731 5321 2740 5355
rect 2688 5312 2740 5321
rect 3240 5312 3292 5364
rect 4160 5312 4212 5364
rect 4712 5355 4764 5364
rect 4712 5321 4721 5355
rect 4721 5321 4755 5355
rect 4755 5321 4764 5355
rect 4712 5312 4764 5321
rect 6828 5312 6880 5364
rect 12348 5312 12400 5364
rect 12992 5355 13044 5364
rect 12992 5321 13001 5355
rect 13001 5321 13035 5355
rect 13035 5321 13044 5355
rect 12992 5312 13044 5321
rect 14556 5312 14608 5364
rect 14648 5312 14700 5364
rect 20628 5312 20680 5364
rect 30012 5355 30064 5364
rect 30012 5321 30021 5355
rect 30021 5321 30055 5355
rect 30055 5321 30064 5355
rect 30012 5312 30064 5321
rect 3056 5244 3108 5296
rect 3516 5176 3568 5228
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 4160 5219 4212 5228
rect 4160 5185 4169 5219
rect 4169 5185 4203 5219
rect 4203 5185 4212 5219
rect 4160 5176 4212 5185
rect 4252 5219 4304 5228
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 7012 5244 7064 5296
rect 4252 5176 4304 5185
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 3792 5108 3844 5160
rect 6460 5176 6512 5228
rect 9404 5244 9456 5296
rect 21180 5244 21232 5296
rect 8392 5176 8444 5228
rect 11336 5176 11388 5228
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11796 5176 11848 5185
rect 12716 5176 12768 5228
rect 13084 5176 13136 5228
rect 14372 5219 14424 5228
rect 5724 5108 5776 5160
rect 4068 4972 4120 5024
rect 4160 4972 4212 5024
rect 8024 4972 8076 5024
rect 12256 5108 12308 5160
rect 12440 5108 12492 5160
rect 13452 5151 13504 5160
rect 13452 5117 13461 5151
rect 13461 5117 13495 5151
rect 13495 5117 13504 5151
rect 13452 5108 13504 5117
rect 14372 5185 14381 5219
rect 14381 5185 14415 5219
rect 14415 5185 14424 5219
rect 14372 5176 14424 5185
rect 15200 5176 15252 5228
rect 15384 5176 15436 5228
rect 15568 5151 15620 5160
rect 15568 5117 15577 5151
rect 15577 5117 15611 5151
rect 15611 5117 15620 5151
rect 15568 5108 15620 5117
rect 16212 5176 16264 5228
rect 17316 5219 17368 5228
rect 17316 5185 17325 5219
rect 17325 5185 17359 5219
rect 17359 5185 17368 5219
rect 17316 5176 17368 5185
rect 19248 5176 19300 5228
rect 19616 5176 19668 5228
rect 21824 5176 21876 5228
rect 29828 5219 29880 5228
rect 29828 5185 29837 5219
rect 29837 5185 29871 5219
rect 29871 5185 29880 5219
rect 29828 5176 29880 5185
rect 16672 5108 16724 5160
rect 17960 5108 18012 5160
rect 18788 5108 18840 5160
rect 13912 5040 13964 5092
rect 18604 5040 18656 5092
rect 8668 4972 8720 5024
rect 9404 4972 9456 5024
rect 9864 5015 9916 5024
rect 9864 4981 9873 5015
rect 9873 4981 9907 5015
rect 9907 4981 9916 5015
rect 9864 4972 9916 4981
rect 10600 4972 10652 5024
rect 17132 5015 17184 5024
rect 17132 4981 17141 5015
rect 17141 4981 17175 5015
rect 17175 4981 17184 5015
rect 17132 4972 17184 4981
rect 18512 5015 18564 5024
rect 18512 4981 18521 5015
rect 18521 4981 18555 5015
rect 18555 4981 18564 5015
rect 18512 4972 18564 4981
rect 5915 4870 5967 4922
rect 5979 4870 6031 4922
rect 6043 4870 6095 4922
rect 6107 4870 6159 4922
rect 6171 4870 6223 4922
rect 15846 4870 15898 4922
rect 15910 4870 15962 4922
rect 15974 4870 16026 4922
rect 16038 4870 16090 4922
rect 16102 4870 16154 4922
rect 25776 4870 25828 4922
rect 25840 4870 25892 4922
rect 25904 4870 25956 4922
rect 25968 4870 26020 4922
rect 26032 4870 26084 4922
rect 3884 4768 3936 4820
rect 4068 4768 4120 4820
rect 4988 4768 5040 4820
rect 1216 4632 1268 4684
rect 4160 4632 4212 4684
rect 2780 4564 2832 4616
rect 5816 4768 5868 4820
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 10692 4768 10744 4820
rect 15016 4768 15068 4820
rect 5632 4700 5684 4752
rect 6644 4700 6696 4752
rect 4528 4496 4580 4548
rect 6276 4564 6328 4616
rect 6184 4496 6236 4548
rect 6460 4496 6512 4548
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 7104 4632 7156 4684
rect 8484 4700 8536 4752
rect 14464 4700 14516 4752
rect 17960 4768 18012 4820
rect 7932 4675 7984 4684
rect 7564 4564 7616 4616
rect 7932 4641 7941 4675
rect 7941 4641 7975 4675
rect 7975 4641 7984 4675
rect 7932 4632 7984 4641
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 8116 4564 8168 4616
rect 9864 4632 9916 4684
rect 8484 4564 8536 4616
rect 8852 4564 8904 4616
rect 5172 4471 5224 4480
rect 5172 4437 5181 4471
rect 5181 4437 5215 4471
rect 5215 4437 5224 4471
rect 5172 4428 5224 4437
rect 5724 4428 5776 4480
rect 8668 4496 8720 4548
rect 9312 4607 9364 4616
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 10784 4632 10836 4684
rect 12256 4632 12308 4684
rect 15108 4632 15160 4684
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 13176 4564 13228 4616
rect 16856 4632 16908 4684
rect 7104 4471 7156 4480
rect 7104 4437 7113 4471
rect 7113 4437 7147 4471
rect 7147 4437 7156 4471
rect 7104 4428 7156 4437
rect 7932 4428 7984 4480
rect 9588 4496 9640 4548
rect 11520 4539 11572 4548
rect 11520 4505 11529 4539
rect 11529 4505 11563 4539
rect 11563 4505 11572 4539
rect 11520 4496 11572 4505
rect 11704 4539 11756 4548
rect 11704 4505 11713 4539
rect 11713 4505 11747 4539
rect 11747 4505 11756 4539
rect 11704 4496 11756 4505
rect 16580 4496 16632 4548
rect 17040 4564 17092 4616
rect 16948 4496 17000 4548
rect 9772 4428 9824 4480
rect 11244 4428 11296 4480
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 16304 4471 16356 4480
rect 16304 4437 16313 4471
rect 16313 4437 16347 4471
rect 16347 4437 16356 4471
rect 16304 4428 16356 4437
rect 16396 4428 16448 4480
rect 17500 4564 17552 4616
rect 18236 4675 18288 4684
rect 18236 4641 18245 4675
rect 18245 4641 18279 4675
rect 18279 4641 18288 4675
rect 18236 4632 18288 4641
rect 19432 4632 19484 4684
rect 18144 4607 18196 4616
rect 18144 4573 18157 4607
rect 18157 4573 18191 4607
rect 18191 4573 18196 4607
rect 18144 4564 18196 4573
rect 19800 4768 19852 4820
rect 21364 4768 21416 4820
rect 19616 4675 19668 4684
rect 19616 4641 19625 4675
rect 19625 4641 19659 4675
rect 19659 4641 19668 4675
rect 19616 4632 19668 4641
rect 30104 4607 30156 4616
rect 30104 4573 30113 4607
rect 30113 4573 30147 4607
rect 30147 4573 30156 4607
rect 30104 4564 30156 4573
rect 18696 4471 18748 4480
rect 18696 4437 18705 4471
rect 18705 4437 18739 4471
rect 18739 4437 18748 4471
rect 18696 4428 18748 4437
rect 20168 4496 20220 4548
rect 20444 4428 20496 4480
rect 20720 4428 20772 4480
rect 29920 4471 29972 4480
rect 29920 4437 29929 4471
rect 29929 4437 29963 4471
rect 29963 4437 29972 4471
rect 29920 4428 29972 4437
rect 10880 4326 10932 4378
rect 10944 4326 10996 4378
rect 11008 4326 11060 4378
rect 11072 4326 11124 4378
rect 11136 4326 11188 4378
rect 20811 4326 20863 4378
rect 20875 4326 20927 4378
rect 20939 4326 20991 4378
rect 21003 4326 21055 4378
rect 21067 4326 21119 4378
rect 4252 4224 4304 4276
rect 4528 4224 4580 4276
rect 7564 4224 7616 4276
rect 12900 4224 12952 4276
rect 13176 4267 13228 4276
rect 13176 4233 13185 4267
rect 13185 4233 13219 4267
rect 13219 4233 13228 4267
rect 13176 4224 13228 4233
rect 14924 4224 14976 4276
rect 16672 4267 16724 4276
rect 16672 4233 16681 4267
rect 16681 4233 16715 4267
rect 16715 4233 16724 4267
rect 16672 4224 16724 4233
rect 19800 4267 19852 4276
rect 19800 4233 19809 4267
rect 19809 4233 19843 4267
rect 19843 4233 19852 4267
rect 19800 4224 19852 4233
rect 20444 4224 20496 4276
rect 21180 4224 21232 4276
rect 1860 4199 1912 4208
rect 1860 4165 1869 4199
rect 1869 4165 1903 4199
rect 1903 4165 1912 4199
rect 1860 4156 1912 4165
rect 3700 4156 3752 4208
rect 2780 4088 2832 4140
rect 2596 4020 2648 4072
rect 3976 4088 4028 4140
rect 7472 4156 7524 4208
rect 4896 4088 4948 4140
rect 5540 4088 5592 4140
rect 7104 4088 7156 4140
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 9036 4131 9088 4140
rect 9036 4097 9045 4131
rect 9045 4097 9079 4131
rect 9079 4097 9088 4131
rect 9036 4088 9088 4097
rect 9680 4156 9732 4208
rect 11888 4156 11940 4208
rect 15384 4199 15436 4208
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 5632 4020 5684 4072
rect 8300 4020 8352 4072
rect 9312 4088 9364 4140
rect 9496 4088 9548 4140
rect 9588 4088 9640 4140
rect 10232 4088 10284 4140
rect 11060 4088 11112 4140
rect 11980 4088 12032 4140
rect 15384 4165 15393 4199
rect 15393 4165 15427 4199
rect 15427 4165 15436 4199
rect 15384 4156 15436 4165
rect 18420 4156 18472 4208
rect 18696 4199 18748 4208
rect 18696 4165 18730 4199
rect 18730 4165 18748 4199
rect 18696 4156 18748 4165
rect 12256 4088 12308 4140
rect 11612 4020 11664 4072
rect 13360 4088 13412 4140
rect 14372 4088 14424 4140
rect 15200 4088 15252 4140
rect 15476 4131 15528 4140
rect 15476 4097 15485 4131
rect 15485 4097 15519 4131
rect 15519 4097 15528 4131
rect 15476 4088 15528 4097
rect 18328 4088 18380 4140
rect 19432 4088 19484 4140
rect 20444 4131 20496 4140
rect 20444 4097 20453 4131
rect 20453 4097 20487 4131
rect 20487 4097 20496 4131
rect 20444 4088 20496 4097
rect 20628 4156 20680 4208
rect 14464 4020 14516 4072
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 5080 3884 5132 3936
rect 6276 3884 6328 3936
rect 10692 3952 10744 4004
rect 15752 4020 15804 4072
rect 17408 4020 17460 4072
rect 16948 3952 17000 4004
rect 9680 3884 9732 3936
rect 11060 3884 11112 3936
rect 11244 3884 11296 3936
rect 12348 3884 12400 3936
rect 14096 3884 14148 3936
rect 16396 3884 16448 3936
rect 19708 4020 19760 4072
rect 19524 3952 19576 4004
rect 23572 3952 23624 4004
rect 29736 4088 29788 4140
rect 30840 4020 30892 4072
rect 31576 3952 31628 4004
rect 19340 3884 19392 3936
rect 20536 3884 20588 3936
rect 22928 3884 22980 3936
rect 28724 3927 28776 3936
rect 28724 3893 28733 3927
rect 28733 3893 28767 3927
rect 28767 3893 28776 3927
rect 28724 3884 28776 3893
rect 29552 3884 29604 3936
rect 30012 3927 30064 3936
rect 30012 3893 30021 3927
rect 30021 3893 30055 3927
rect 30055 3893 30064 3927
rect 30012 3884 30064 3893
rect 5915 3782 5967 3834
rect 5979 3782 6031 3834
rect 6043 3782 6095 3834
rect 6107 3782 6159 3834
rect 6171 3782 6223 3834
rect 15846 3782 15898 3834
rect 15910 3782 15962 3834
rect 15974 3782 16026 3834
rect 16038 3782 16090 3834
rect 16102 3782 16154 3834
rect 25776 3782 25828 3834
rect 25840 3782 25892 3834
rect 25904 3782 25956 3834
rect 25968 3782 26020 3834
rect 26032 3782 26084 3834
rect 10232 3680 10284 3732
rect 10784 3680 10836 3732
rect 11244 3680 11296 3732
rect 15660 3723 15712 3732
rect 15660 3689 15669 3723
rect 15669 3689 15703 3723
rect 15703 3689 15712 3723
rect 15660 3680 15712 3689
rect 16764 3680 16816 3732
rect 16948 3680 17000 3732
rect 18420 3680 18472 3732
rect 20168 3723 20220 3732
rect 20168 3689 20177 3723
rect 20177 3689 20211 3723
rect 20211 3689 20220 3723
rect 20168 3680 20220 3689
rect 20720 3680 20772 3732
rect 5080 3612 5132 3664
rect 13084 3655 13136 3664
rect 13084 3621 13093 3655
rect 13093 3621 13127 3655
rect 13127 3621 13136 3655
rect 13084 3612 13136 3621
rect 2964 3476 3016 3528
rect 2780 3451 2832 3460
rect 2780 3417 2789 3451
rect 2789 3417 2823 3451
rect 2823 3417 2832 3451
rect 2780 3408 2832 3417
rect 11612 3544 11664 3596
rect 3424 3476 3476 3528
rect 9404 3476 9456 3528
rect 9772 3519 9824 3528
rect 9772 3485 9806 3519
rect 9806 3485 9824 3519
rect 9772 3476 9824 3485
rect 11520 3476 11572 3528
rect 11980 3476 12032 3528
rect 13176 3544 13228 3596
rect 17040 3612 17092 3664
rect 15752 3544 15804 3596
rect 17316 3587 17368 3596
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 17408 3587 17460 3596
rect 17408 3553 17417 3587
rect 17417 3553 17451 3587
rect 17451 3553 17460 3587
rect 17408 3544 17460 3553
rect 17960 3544 18012 3596
rect 20444 3612 20496 3664
rect 22928 3723 22980 3732
rect 22928 3689 22937 3723
rect 22937 3689 22971 3723
rect 22971 3689 22980 3723
rect 22928 3680 22980 3689
rect 20996 3612 21048 3664
rect 21824 3612 21876 3664
rect 19708 3587 19760 3596
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 20352 3544 20404 3596
rect 12348 3476 12400 3528
rect 5172 3408 5224 3460
rect 5540 3408 5592 3460
rect 11336 3408 11388 3460
rect 12440 3408 12492 3460
rect 13176 3408 13228 3460
rect 5724 3340 5776 3392
rect 5816 3340 5868 3392
rect 9588 3340 9640 3392
rect 15016 3476 15068 3528
rect 16304 3476 16356 3528
rect 17132 3476 17184 3528
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 19892 3476 19944 3528
rect 20812 3476 20864 3528
rect 16672 3408 16724 3460
rect 16856 3408 16908 3460
rect 20996 3519 21048 3528
rect 20996 3485 21005 3519
rect 21005 3485 21039 3519
rect 21039 3485 21048 3519
rect 20996 3476 21048 3485
rect 21180 3476 21232 3528
rect 22560 3476 22612 3528
rect 27804 3476 27856 3528
rect 28540 3476 28592 3528
rect 29276 3476 29328 3528
rect 17132 3340 17184 3392
rect 21364 3408 21416 3460
rect 21824 3451 21876 3460
rect 21824 3417 21833 3451
rect 21833 3417 21867 3451
rect 21867 3417 21876 3451
rect 21824 3408 21876 3417
rect 22744 3408 22796 3460
rect 22468 3340 22520 3392
rect 25688 3340 25740 3392
rect 27712 3340 27764 3392
rect 27988 3340 28040 3392
rect 29920 3340 29972 3392
rect 10880 3238 10932 3290
rect 10944 3238 10996 3290
rect 11008 3238 11060 3290
rect 11072 3238 11124 3290
rect 11136 3238 11188 3290
rect 20811 3238 20863 3290
rect 20875 3238 20927 3290
rect 20939 3238 20991 3290
rect 21003 3238 21055 3290
rect 21067 3238 21119 3290
rect 2872 3068 2924 3120
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 4804 3136 4856 3188
rect 4896 3136 4948 3188
rect 9036 3136 9088 3188
rect 9496 3136 9548 3188
rect 11428 3136 11480 3188
rect 11704 3136 11756 3188
rect 13820 3179 13872 3188
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 5540 3068 5592 3120
rect 8300 3068 8352 3120
rect 4988 3000 5040 3052
rect 6460 3000 6512 3052
rect 7196 3000 7248 3052
rect 7472 3000 7524 3052
rect 8760 3000 8812 3052
rect 9128 3000 9180 3052
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 9680 3043 9732 3052
rect 9680 3009 9714 3043
rect 9714 3009 9732 3043
rect 9680 3000 9732 3009
rect 4988 2864 5040 2916
rect 7380 2864 7432 2916
rect 11888 3068 11940 3120
rect 11796 3000 11848 3052
rect 12992 3000 13044 3052
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 13360 3000 13412 3052
rect 17132 3136 17184 3188
rect 17684 3136 17736 3188
rect 17960 3136 18012 3188
rect 18512 3136 18564 3188
rect 19248 3179 19300 3188
rect 19248 3145 19257 3179
rect 19257 3145 19291 3179
rect 19291 3145 19300 3179
rect 19248 3136 19300 3145
rect 15108 3068 15160 3120
rect 15568 3068 15620 3120
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 15200 3043 15252 3052
rect 15200 3009 15209 3043
rect 15209 3009 15243 3043
rect 15243 3009 15252 3043
rect 15200 3000 15252 3009
rect 13084 2932 13136 2984
rect 15752 3000 15804 3052
rect 16488 3068 16540 3120
rect 16580 3068 16632 3120
rect 6368 2796 6420 2848
rect 8668 2796 8720 2848
rect 9312 2796 9364 2848
rect 11796 2796 11848 2848
rect 15108 2864 15160 2916
rect 14924 2796 14976 2848
rect 15568 2932 15620 2984
rect 17040 3000 17092 3052
rect 17960 3043 18012 3052
rect 17960 3009 17969 3043
rect 17969 3009 18003 3043
rect 18003 3009 18012 3043
rect 17960 3000 18012 3009
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 16764 2864 16816 2916
rect 16948 2864 17000 2916
rect 17224 2864 17276 2916
rect 20536 3068 20588 3120
rect 21364 3136 21416 3188
rect 21824 3179 21876 3188
rect 21824 3145 21833 3179
rect 21833 3145 21867 3179
rect 21867 3145 21876 3179
rect 21824 3136 21876 3145
rect 22928 3179 22980 3188
rect 22928 3145 22937 3179
rect 22937 3145 22971 3179
rect 22971 3145 22980 3179
rect 22928 3136 22980 3145
rect 23572 3179 23624 3188
rect 23572 3145 23581 3179
rect 23581 3145 23615 3179
rect 23615 3145 23624 3179
rect 23572 3136 23624 3145
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 20444 3043 20496 3052
rect 20444 3009 20453 3043
rect 20453 3009 20487 3043
rect 20487 3009 20496 3043
rect 21640 3068 21692 3120
rect 21732 3068 21784 3120
rect 20444 3000 20496 3009
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22468 3043 22520 3052
rect 22100 3000 22152 3009
rect 22468 3009 22477 3043
rect 22477 3009 22511 3043
rect 22511 3009 22520 3043
rect 22468 3000 22520 3009
rect 27988 3068 28040 3120
rect 23940 3000 23992 3052
rect 27436 3043 27488 3052
rect 27436 3009 27445 3043
rect 27445 3009 27479 3043
rect 27479 3009 27488 3043
rect 27436 3000 27488 3009
rect 28724 3000 28776 3052
rect 29920 3043 29972 3052
rect 29920 3009 29929 3043
rect 29929 3009 29963 3043
rect 29963 3009 29972 3043
rect 29920 3000 29972 3009
rect 30012 3043 30064 3052
rect 30012 3009 30021 3043
rect 30021 3009 30055 3043
rect 30055 3009 30064 3043
rect 30012 3000 30064 3009
rect 27620 2975 27672 2984
rect 20168 2864 20220 2916
rect 27620 2941 27629 2975
rect 27629 2941 27663 2975
rect 27663 2941 27672 2975
rect 27620 2932 27672 2941
rect 22100 2864 22152 2916
rect 22744 2864 22796 2916
rect 16672 2796 16724 2848
rect 18144 2796 18196 2848
rect 19524 2796 19576 2848
rect 20260 2839 20312 2848
rect 20260 2805 20269 2839
rect 20269 2805 20303 2839
rect 20303 2805 20312 2839
rect 20260 2796 20312 2805
rect 22376 2839 22428 2848
rect 22376 2805 22385 2839
rect 22385 2805 22419 2839
rect 22419 2805 22428 2839
rect 22376 2796 22428 2805
rect 27712 2839 27764 2848
rect 27712 2805 27721 2839
rect 27721 2805 27755 2839
rect 27755 2805 27764 2839
rect 27712 2796 27764 2805
rect 29552 2839 29604 2848
rect 29552 2805 29561 2839
rect 29561 2805 29595 2839
rect 29595 2805 29604 2839
rect 29552 2796 29604 2805
rect 5915 2694 5967 2746
rect 5979 2694 6031 2746
rect 6043 2694 6095 2746
rect 6107 2694 6159 2746
rect 6171 2694 6223 2746
rect 15846 2694 15898 2746
rect 15910 2694 15962 2746
rect 15974 2694 16026 2746
rect 16038 2694 16090 2746
rect 16102 2694 16154 2746
rect 25776 2694 25828 2746
rect 25840 2694 25892 2746
rect 25904 2694 25956 2746
rect 25968 2694 26020 2746
rect 26032 2694 26084 2746
rect 4436 2635 4488 2644
rect 4436 2601 4445 2635
rect 4445 2601 4479 2635
rect 4479 2601 4488 2635
rect 4436 2592 4488 2601
rect 7840 2592 7892 2644
rect 8300 2592 8352 2644
rect 11704 2592 11756 2644
rect 14188 2592 14240 2644
rect 14464 2635 14516 2644
rect 14464 2601 14473 2635
rect 14473 2601 14507 2635
rect 14507 2601 14516 2635
rect 14464 2592 14516 2601
rect 15384 2592 15436 2644
rect 15568 2592 15620 2644
rect 16672 2635 16724 2644
rect 16672 2601 16681 2635
rect 16681 2601 16715 2635
rect 16715 2601 16724 2635
rect 16672 2592 16724 2601
rect 7472 2524 7524 2576
rect 12900 2524 12952 2576
rect 12992 2524 13044 2576
rect 17960 2592 18012 2644
rect 20260 2635 20312 2644
rect 20260 2601 20269 2635
rect 20269 2601 20303 2635
rect 20303 2601 20312 2635
rect 20260 2592 20312 2601
rect 20720 2635 20772 2644
rect 20720 2601 20729 2635
rect 20729 2601 20763 2635
rect 20763 2601 20772 2635
rect 20720 2592 20772 2601
rect 21640 2592 21692 2644
rect 22100 2635 22152 2644
rect 22100 2601 22109 2635
rect 22109 2601 22143 2635
rect 22143 2601 22152 2635
rect 22100 2592 22152 2601
rect 22284 2592 22336 2644
rect 25688 2635 25740 2644
rect 25688 2601 25697 2635
rect 25697 2601 25731 2635
rect 25731 2601 25740 2635
rect 25688 2592 25740 2601
rect 27436 2592 27488 2644
rect 27620 2635 27672 2644
rect 27620 2601 27629 2635
rect 27629 2601 27663 2635
rect 27663 2601 27672 2635
rect 27620 2592 27672 2601
rect 18328 2524 18380 2576
rect 18604 2524 18656 2576
rect 1860 2388 1912 2440
rect 388 2320 440 2372
rect 4160 2363 4212 2372
rect 4160 2329 4169 2363
rect 4169 2329 4203 2363
rect 4203 2329 4212 2363
rect 4160 2320 4212 2329
rect 4896 2388 4948 2440
rect 5724 2388 5776 2440
rect 9312 2456 9364 2508
rect 10324 2456 10376 2508
rect 10508 2456 10560 2508
rect 15016 2499 15068 2508
rect 15016 2465 15025 2499
rect 15025 2465 15059 2499
rect 15059 2465 15068 2499
rect 15016 2456 15068 2465
rect 16764 2456 16816 2508
rect 7932 2388 7984 2440
rect 8760 2388 8812 2440
rect 9496 2388 9548 2440
rect 10232 2388 10284 2440
rect 8392 2320 8444 2372
rect 11336 2320 11388 2372
rect 14924 2388 14976 2440
rect 15292 2431 15344 2440
rect 15292 2397 15301 2431
rect 15301 2397 15335 2431
rect 15335 2397 15344 2431
rect 15292 2388 15344 2397
rect 15568 2388 15620 2440
rect 16396 2388 16448 2440
rect 17132 2456 17184 2508
rect 20444 2499 20496 2508
rect 17408 2388 17460 2440
rect 8944 2252 8996 2304
rect 12624 2252 12676 2304
rect 18052 2388 18104 2440
rect 18512 2388 18564 2440
rect 18788 2388 18840 2440
rect 20444 2465 20453 2499
rect 20453 2465 20487 2499
rect 20487 2465 20496 2499
rect 20444 2456 20496 2465
rect 20536 2431 20588 2440
rect 20076 2320 20128 2372
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 22652 2456 22704 2508
rect 21824 2388 21876 2440
rect 22744 2388 22796 2440
rect 23204 2456 23256 2508
rect 24768 2388 24820 2440
rect 25504 2388 25556 2440
rect 26240 2388 26292 2440
rect 27068 2388 27120 2440
rect 28724 2431 28776 2440
rect 28724 2397 28733 2431
rect 28733 2397 28767 2431
rect 28767 2397 28776 2431
rect 28724 2388 28776 2397
rect 29460 2388 29512 2440
rect 19248 2252 19300 2304
rect 19432 2252 19484 2304
rect 22652 2295 22704 2304
rect 22652 2261 22661 2295
rect 22661 2261 22695 2295
rect 22695 2261 22704 2295
rect 22652 2252 22704 2261
rect 23296 2295 23348 2304
rect 23296 2261 23305 2295
rect 23305 2261 23339 2295
rect 23339 2261 23348 2295
rect 23296 2252 23348 2261
rect 25044 2295 25096 2304
rect 25044 2261 25053 2295
rect 25053 2261 25087 2295
rect 25087 2261 25096 2295
rect 25044 2252 25096 2261
rect 28908 2295 28960 2304
rect 28908 2261 28917 2295
rect 28917 2261 28951 2295
rect 28951 2261 28960 2295
rect 28908 2252 28960 2261
rect 30012 2295 30064 2304
rect 30012 2261 30021 2295
rect 30021 2261 30055 2295
rect 30055 2261 30064 2295
rect 30012 2252 30064 2261
rect 10880 2150 10932 2202
rect 10944 2150 10996 2202
rect 11008 2150 11060 2202
rect 11072 2150 11124 2202
rect 11136 2150 11188 2202
rect 20811 2150 20863 2202
rect 20875 2150 20927 2202
rect 20939 2150 20991 2202
rect 21003 2150 21055 2202
rect 21067 2150 21119 2202
rect 22008 2048 22060 2100
rect 25044 2048 25096 2100
rect 19248 1980 19300 2032
rect 23296 1980 23348 2032
<< metal2 >>
rect 2778 47560 2834 47569
rect 2778 47495 2834 47504
rect 1400 45484 1452 45490
rect 1400 45426 1452 45432
rect 1412 36922 1440 45426
rect 2226 45384 2282 45393
rect 2226 45319 2228 45328
rect 2280 45319 2282 45328
rect 2228 45290 2280 45296
rect 2792 45286 2820 47495
rect 30194 47152 30250 47161
rect 30194 47087 30250 47096
rect 2870 46880 2926 46889
rect 2870 46815 2926 46824
rect 2884 45490 2912 46815
rect 2962 46064 3018 46073
rect 2962 45999 3018 46008
rect 2872 45484 2924 45490
rect 2872 45426 2924 45432
rect 2976 45354 3004 45999
rect 10880 45724 11188 45744
rect 10880 45722 10886 45724
rect 10942 45722 10966 45724
rect 11022 45722 11046 45724
rect 11102 45722 11126 45724
rect 11182 45722 11188 45724
rect 10942 45670 10944 45722
rect 11124 45670 11126 45722
rect 10880 45668 10886 45670
rect 10942 45668 10966 45670
rect 11022 45668 11046 45670
rect 11102 45668 11126 45670
rect 11182 45668 11188 45670
rect 10880 45648 11188 45668
rect 20811 45724 21119 45744
rect 20811 45722 20817 45724
rect 20873 45722 20897 45724
rect 20953 45722 20977 45724
rect 21033 45722 21057 45724
rect 21113 45722 21119 45724
rect 20873 45670 20875 45722
rect 21055 45670 21057 45722
rect 20811 45668 20817 45670
rect 20873 45668 20897 45670
rect 20953 45668 20977 45670
rect 21033 45668 21057 45670
rect 21113 45668 21119 45670
rect 20811 45648 21119 45668
rect 30102 45656 30158 45665
rect 30102 45591 30158 45600
rect 30116 45490 30144 45591
rect 3056 45484 3108 45490
rect 3056 45426 3108 45432
rect 3148 45484 3200 45490
rect 3148 45426 3200 45432
rect 4804 45484 4856 45490
rect 4804 45426 4856 45432
rect 30104 45484 30156 45490
rect 30104 45426 30156 45432
rect 2964 45348 3016 45354
rect 2964 45290 3016 45296
rect 2780 45280 2832 45286
rect 2780 45222 2832 45228
rect 2872 45280 2924 45286
rect 2872 45222 2924 45228
rect 2884 44878 2912 45222
rect 3068 45082 3096 45426
rect 3160 45082 3188 45426
rect 3056 45076 3108 45082
rect 3056 45018 3108 45024
rect 3148 45076 3200 45082
rect 3148 45018 3200 45024
rect 2872 44872 2924 44878
rect 2872 44814 2924 44820
rect 4528 44872 4580 44878
rect 4528 44814 4580 44820
rect 1492 44736 1544 44742
rect 1492 44678 1544 44684
rect 2872 44736 2924 44742
rect 2872 44678 2924 44684
rect 1504 44577 1532 44678
rect 1490 44568 1546 44577
rect 1490 44503 1546 44512
rect 2884 44470 2912 44678
rect 2872 44464 2924 44470
rect 2872 44406 2924 44412
rect 2320 44396 2372 44402
rect 2320 44338 2372 44344
rect 4252 44396 4304 44402
rect 4252 44338 4304 44344
rect 1492 44192 1544 44198
rect 1492 44134 1544 44140
rect 1952 44192 2004 44198
rect 1952 44134 2004 44140
rect 1504 43897 1532 44134
rect 1490 43888 1546 43897
rect 1490 43823 1546 43832
rect 1860 43784 1912 43790
rect 1860 43726 1912 43732
rect 1584 43648 1636 43654
rect 1584 43590 1636 43596
rect 1492 43104 1544 43110
rect 1490 43072 1492 43081
rect 1544 43072 1546 43081
rect 1490 43007 1546 43016
rect 1492 42560 1544 42566
rect 1492 42502 1544 42508
rect 1504 42401 1532 42502
rect 1490 42392 1546 42401
rect 1490 42327 1546 42336
rect 1492 42016 1544 42022
rect 1492 41958 1544 41964
rect 1504 41721 1532 41958
rect 1490 41712 1546 41721
rect 1490 41647 1546 41656
rect 1492 40928 1544 40934
rect 1490 40896 1492 40905
rect 1544 40896 1546 40905
rect 1490 40831 1546 40840
rect 1492 40384 1544 40390
rect 1492 40326 1544 40332
rect 1504 40225 1532 40326
rect 1490 40216 1546 40225
rect 1490 40151 1546 40160
rect 1596 39438 1624 43590
rect 1768 41608 1820 41614
rect 1768 41550 1820 41556
rect 1676 41472 1728 41478
rect 1676 41414 1728 41420
rect 1584 39432 1636 39438
rect 1584 39374 1636 39380
rect 1492 39296 1544 39302
rect 1492 39238 1544 39244
rect 1504 37913 1532 39238
rect 1490 37904 1546 37913
rect 1490 37839 1546 37848
rect 1400 36916 1452 36922
rect 1400 36858 1452 36864
rect 1400 36576 1452 36582
rect 1400 36518 1452 36524
rect 1412 35737 1440 36518
rect 1688 36174 1716 41414
rect 1676 36168 1728 36174
rect 1676 36110 1728 36116
rect 1492 36032 1544 36038
rect 1492 35974 1544 35980
rect 1398 35728 1454 35737
rect 1398 35663 1454 35672
rect 1504 35057 1532 35974
rect 1490 35048 1546 35057
rect 1490 34983 1546 34992
rect 1780 34746 1808 41550
rect 1872 38010 1900 43726
rect 1964 40526 1992 44134
rect 2136 42696 2188 42702
rect 2136 42638 2188 42644
rect 2044 42016 2096 42022
rect 2044 41958 2096 41964
rect 1952 40520 2004 40526
rect 1952 40462 2004 40468
rect 1952 38752 2004 38758
rect 1952 38694 2004 38700
rect 1964 38554 1992 38694
rect 1952 38548 2004 38554
rect 1952 38490 2004 38496
rect 1860 38004 1912 38010
rect 1860 37946 1912 37952
rect 1964 37670 1992 38490
rect 1952 37664 2004 37670
rect 1952 37606 2004 37612
rect 1964 37466 1992 37606
rect 1952 37460 2004 37466
rect 1952 37402 2004 37408
rect 2056 36786 2084 41958
rect 2148 38554 2176 42638
rect 2332 41274 2360 44338
rect 3976 44328 4028 44334
rect 3976 44270 4028 44276
rect 2964 44192 3016 44198
rect 2964 44134 3016 44140
rect 3424 44192 3476 44198
rect 3424 44134 3476 44140
rect 2504 43784 2556 43790
rect 2504 43726 2556 43732
rect 2412 42220 2464 42226
rect 2412 42162 2464 42168
rect 2320 41268 2372 41274
rect 2320 41210 2372 41216
rect 2228 40656 2280 40662
rect 2228 40598 2280 40604
rect 2240 39846 2268 40598
rect 2228 39840 2280 39846
rect 2280 39800 2360 39828
rect 2228 39782 2280 39788
rect 2226 39400 2282 39409
rect 2226 39335 2282 39344
rect 2240 39302 2268 39335
rect 2228 39296 2280 39302
rect 2228 39238 2280 39244
rect 2332 38758 2360 39800
rect 2320 38752 2372 38758
rect 2320 38694 2372 38700
rect 2136 38548 2188 38554
rect 2136 38490 2188 38496
rect 2320 37256 2372 37262
rect 2320 37198 2372 37204
rect 2044 36780 2096 36786
rect 2044 36722 2096 36728
rect 2332 36666 2360 37198
rect 2424 37126 2452 42162
rect 2516 39098 2544 43726
rect 2872 43308 2924 43314
rect 2872 43250 2924 43256
rect 2780 43104 2832 43110
rect 2780 43046 2832 43052
rect 2596 42560 2648 42566
rect 2596 42502 2648 42508
rect 2504 39092 2556 39098
rect 2504 39034 2556 39040
rect 2504 38208 2556 38214
rect 2504 38150 2556 38156
rect 2516 37942 2544 38150
rect 2504 37936 2556 37942
rect 2504 37878 2556 37884
rect 2608 37262 2636 42502
rect 2792 42226 2820 43046
rect 2780 42220 2832 42226
rect 2780 42162 2832 42168
rect 2884 41818 2912 43250
rect 2976 42770 3004 44134
rect 3148 43920 3200 43926
rect 3148 43862 3200 43868
rect 3056 43104 3108 43110
rect 3056 43046 3108 43052
rect 2964 42764 3016 42770
rect 2964 42706 3016 42712
rect 3068 42702 3096 43046
rect 3056 42696 3108 42702
rect 3056 42638 3108 42644
rect 2872 41812 2924 41818
rect 2872 41754 2924 41760
rect 2780 41608 2832 41614
rect 2780 41550 2832 41556
rect 2792 40526 2820 41550
rect 2964 41472 3016 41478
rect 2964 41414 3016 41420
rect 2976 41002 3004 41414
rect 2964 40996 3016 41002
rect 2964 40938 3016 40944
rect 2780 40520 2832 40526
rect 2780 40462 2832 40468
rect 2688 38344 2740 38350
rect 2688 38286 2740 38292
rect 2700 38010 2728 38286
rect 2688 38004 2740 38010
rect 2688 37946 2740 37952
rect 2596 37256 2648 37262
rect 2596 37198 2648 37204
rect 2792 37244 2820 40462
rect 2976 40050 3004 40938
rect 3056 40384 3108 40390
rect 3056 40326 3108 40332
rect 2964 40044 3016 40050
rect 2964 39986 3016 39992
rect 2872 39976 2924 39982
rect 2872 39918 2924 39924
rect 2884 39642 2912 39918
rect 2872 39636 2924 39642
rect 2872 39578 2924 39584
rect 2976 38894 3004 39986
rect 3068 39438 3096 40326
rect 3056 39432 3108 39438
rect 3056 39374 3108 39380
rect 3160 38962 3188 43862
rect 3240 43648 3292 43654
rect 3240 43590 3292 43596
rect 3252 41070 3280 43590
rect 3436 43382 3464 44134
rect 3424 43376 3476 43382
rect 3424 43318 3476 43324
rect 3884 43308 3936 43314
rect 3884 43250 3936 43256
rect 3424 42220 3476 42226
rect 3424 42162 3476 42168
rect 3516 42220 3568 42226
rect 3516 42162 3568 42168
rect 3436 41274 3464 42162
rect 3424 41268 3476 41274
rect 3424 41210 3476 41216
rect 3240 41064 3292 41070
rect 3240 41006 3292 41012
rect 3528 39846 3556 42162
rect 3700 42016 3752 42022
rect 3700 41958 3752 41964
rect 3712 41138 3740 41958
rect 3896 41614 3924 43250
rect 3884 41608 3936 41614
rect 3884 41550 3936 41556
rect 3988 41274 4016 44270
rect 4264 42362 4292 44338
rect 4540 43994 4568 44814
rect 4816 44538 4844 45426
rect 5264 45416 5316 45422
rect 5264 45358 5316 45364
rect 5172 45076 5224 45082
rect 5172 45018 5224 45024
rect 4804 44532 4856 44538
rect 4804 44474 4856 44480
rect 5184 44198 5212 45018
rect 5276 44538 5304 45358
rect 29920 45280 29972 45286
rect 29920 45222 29972 45228
rect 5915 45180 6223 45200
rect 5915 45178 5921 45180
rect 5977 45178 6001 45180
rect 6057 45178 6081 45180
rect 6137 45178 6161 45180
rect 6217 45178 6223 45180
rect 5977 45126 5979 45178
rect 6159 45126 6161 45178
rect 5915 45124 5921 45126
rect 5977 45124 6001 45126
rect 6057 45124 6081 45126
rect 6137 45124 6161 45126
rect 6217 45124 6223 45126
rect 5915 45104 6223 45124
rect 15846 45180 16154 45200
rect 15846 45178 15852 45180
rect 15908 45178 15932 45180
rect 15988 45178 16012 45180
rect 16068 45178 16092 45180
rect 16148 45178 16154 45180
rect 15908 45126 15910 45178
rect 16090 45126 16092 45178
rect 15846 45124 15852 45126
rect 15908 45124 15932 45126
rect 15988 45124 16012 45126
rect 16068 45124 16092 45126
rect 16148 45124 16154 45126
rect 15846 45104 16154 45124
rect 25776 45180 26084 45200
rect 25776 45178 25782 45180
rect 25838 45178 25862 45180
rect 25918 45178 25942 45180
rect 25998 45178 26022 45180
rect 26078 45178 26084 45180
rect 25838 45126 25840 45178
rect 26020 45126 26022 45178
rect 25776 45124 25782 45126
rect 25838 45124 25862 45126
rect 25918 45124 25942 45126
rect 25998 45124 26022 45126
rect 26078 45124 26084 45126
rect 25776 45104 26084 45124
rect 5724 44940 5776 44946
rect 5724 44882 5776 44888
rect 5540 44872 5592 44878
rect 5540 44814 5592 44820
rect 5264 44532 5316 44538
rect 5264 44474 5316 44480
rect 5552 44266 5580 44814
rect 5540 44260 5592 44266
rect 5540 44202 5592 44208
rect 5172 44192 5224 44198
rect 5172 44134 5224 44140
rect 4528 43988 4580 43994
rect 4528 43930 4580 43936
rect 5184 43926 5212 44134
rect 5172 43920 5224 43926
rect 5172 43862 5224 43868
rect 5080 43784 5132 43790
rect 5080 43726 5132 43732
rect 5092 43314 5120 43726
rect 4528 43308 4580 43314
rect 4528 43250 4580 43256
rect 5080 43308 5132 43314
rect 5080 43250 5132 43256
rect 4344 43104 4396 43110
rect 4344 43046 4396 43052
rect 4252 42356 4304 42362
rect 4252 42298 4304 42304
rect 4356 42294 4384 43046
rect 4436 42628 4488 42634
rect 4436 42570 4488 42576
rect 4344 42288 4396 42294
rect 4344 42230 4396 42236
rect 4068 42084 4120 42090
rect 4068 42026 4120 42032
rect 3976 41268 4028 41274
rect 3976 41210 4028 41216
rect 3700 41132 3752 41138
rect 3700 41074 3752 41080
rect 3976 41132 4028 41138
rect 3976 41074 4028 41080
rect 3988 40730 4016 41074
rect 3976 40724 4028 40730
rect 3976 40666 4028 40672
rect 3988 40610 4016 40666
rect 3896 40582 4016 40610
rect 3792 40384 3844 40390
rect 3792 40326 3844 40332
rect 3804 40118 3832 40326
rect 3792 40112 3844 40118
rect 3792 40054 3844 40060
rect 3516 39840 3568 39846
rect 3516 39782 3568 39788
rect 3792 39432 3844 39438
rect 3792 39374 3844 39380
rect 3148 38956 3200 38962
rect 3148 38898 3200 38904
rect 2964 38888 3016 38894
rect 2964 38830 3016 38836
rect 2872 38820 2924 38826
rect 2872 38762 2924 38768
rect 2884 38418 2912 38762
rect 2976 38486 3004 38830
rect 3056 38752 3108 38758
rect 3054 38720 3056 38729
rect 3108 38720 3110 38729
rect 3054 38655 3110 38664
rect 2964 38480 3016 38486
rect 2964 38422 3016 38428
rect 2872 38412 2924 38418
rect 2872 38354 2924 38360
rect 2976 37806 3004 38422
rect 3148 38344 3200 38350
rect 3148 38286 3200 38292
rect 3160 38010 3188 38286
rect 3148 38004 3200 38010
rect 3148 37946 3200 37952
rect 3700 38004 3752 38010
rect 3700 37946 3752 37952
rect 2964 37800 3016 37806
rect 2964 37742 3016 37748
rect 2964 37256 3016 37262
rect 2792 37216 2964 37244
rect 2412 37120 2464 37126
rect 2412 37062 2464 37068
rect 2596 36916 2648 36922
rect 2596 36858 2648 36864
rect 2332 36650 2452 36666
rect 2332 36644 2464 36650
rect 2332 36638 2412 36644
rect 2412 36586 2464 36592
rect 2320 36576 2372 36582
rect 2318 36544 2320 36553
rect 2372 36544 2374 36553
rect 2318 36479 2374 36488
rect 2228 36032 2280 36038
rect 2228 35974 2280 35980
rect 1860 35692 1912 35698
rect 1860 35634 1912 35640
rect 1872 35222 1900 35634
rect 2240 35494 2268 35974
rect 2424 35698 2452 36586
rect 2412 35692 2464 35698
rect 2412 35634 2464 35640
rect 2228 35488 2280 35494
rect 2228 35430 2280 35436
rect 2240 35290 2268 35430
rect 2228 35284 2280 35290
rect 2228 35226 2280 35232
rect 1860 35216 1912 35222
rect 1860 35158 1912 35164
rect 1768 34740 1820 34746
rect 1768 34682 1820 34688
rect 2240 34406 2268 35226
rect 2424 34610 2452 35634
rect 2412 34604 2464 34610
rect 2412 34546 2464 34552
rect 2228 34400 2280 34406
rect 2228 34342 2280 34348
rect 2240 34202 2268 34342
rect 2228 34196 2280 34202
rect 2228 34138 2280 34144
rect 2044 33516 2096 33522
rect 2044 33458 2096 33464
rect 1492 33312 1544 33318
rect 1492 33254 1544 33260
rect 1504 32745 1532 33254
rect 1490 32736 1546 32745
rect 1490 32671 1546 32680
rect 1492 32224 1544 32230
rect 1492 32166 1544 32172
rect 1504 31385 1532 32166
rect 1490 31376 1546 31385
rect 1490 31311 1546 31320
rect 1490 29880 1546 29889
rect 1490 29815 1492 29824
rect 1544 29815 1546 29824
rect 1492 29786 1544 29792
rect 1676 29164 1728 29170
rect 1676 29106 1728 29112
rect 1490 29064 1546 29073
rect 1490 28999 1492 29008
rect 1544 28999 1546 29008
rect 1492 28970 1544 28976
rect 1688 28762 1716 29106
rect 1676 28756 1728 28762
rect 1676 28698 1728 28704
rect 1492 28416 1544 28422
rect 1490 28384 1492 28393
rect 1544 28384 1546 28393
rect 1490 28319 1546 28328
rect 2056 28218 2084 33458
rect 2136 33312 2188 33318
rect 2136 33254 2188 33260
rect 2148 33046 2176 33254
rect 2240 33114 2268 34138
rect 2424 34134 2452 34546
rect 2412 34128 2464 34134
rect 2412 34070 2464 34076
rect 2228 33108 2280 33114
rect 2228 33050 2280 33056
rect 2136 33040 2188 33046
rect 2136 32982 2188 32988
rect 2148 31958 2176 32982
rect 2412 32768 2464 32774
rect 2412 32710 2464 32716
rect 2228 32224 2280 32230
rect 2228 32166 2280 32172
rect 2240 32065 2268 32166
rect 2226 32056 2282 32065
rect 2226 31991 2282 32000
rect 2320 32020 2372 32026
rect 2320 31962 2372 31968
rect 2136 31952 2188 31958
rect 2136 31894 2188 31900
rect 2148 31346 2176 31894
rect 2136 31340 2188 31346
rect 2136 31282 2188 31288
rect 2148 30870 2176 31282
rect 2332 31142 2360 31962
rect 2320 31136 2372 31142
rect 2320 31078 2372 31084
rect 2332 30938 2360 31078
rect 2320 30932 2372 30938
rect 2320 30874 2372 30880
rect 2136 30864 2188 30870
rect 2136 30806 2188 30812
rect 2148 30258 2176 30806
rect 2136 30252 2188 30258
rect 2136 30194 2188 30200
rect 2320 30048 2372 30054
rect 2320 29990 2372 29996
rect 2332 29646 2360 29990
rect 2320 29640 2372 29646
rect 2320 29582 2372 29588
rect 2044 28212 2096 28218
rect 2044 28154 2096 28160
rect 2424 28082 2452 32710
rect 2504 30592 2556 30598
rect 2504 30534 2556 30540
rect 2516 29170 2544 30534
rect 2504 29164 2556 29170
rect 2504 29106 2556 29112
rect 2412 28076 2464 28082
rect 2412 28018 2464 28024
rect 1492 27872 1544 27878
rect 1492 27814 1544 27820
rect 1504 27577 1532 27814
rect 1490 27568 1546 27577
rect 1490 27503 1546 27512
rect 1676 27328 1728 27334
rect 1676 27270 1728 27276
rect 1688 26994 1716 27270
rect 1676 26988 1728 26994
rect 1676 26930 1728 26936
rect 1490 26888 1546 26897
rect 1490 26823 1492 26832
rect 1544 26823 1546 26832
rect 1492 26794 1544 26800
rect 1492 26240 1544 26246
rect 1490 26208 1492 26217
rect 1544 26208 1546 26217
rect 1490 26143 1546 26152
rect 1492 25696 1544 25702
rect 1492 25638 1544 25644
rect 1504 25401 1532 25638
rect 1490 25392 1546 25401
rect 1490 25327 1546 25336
rect 1490 24712 1546 24721
rect 1490 24647 1492 24656
rect 1544 24647 1546 24656
rect 1492 24618 1544 24624
rect 1492 24064 1544 24070
rect 1492 24006 1544 24012
rect 1504 23905 1532 24006
rect 1490 23896 1546 23905
rect 1490 23831 1546 23840
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 2136 23656 2188 23662
rect 2136 23598 2188 23604
rect 1412 23225 1440 23598
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 21049 1440 23054
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1398 21040 1454 21049
rect 1398 20975 1454 20984
rect 1596 20942 1624 22918
rect 2044 22636 2096 22642
rect 2044 22578 2096 22584
rect 1952 22432 2004 22438
rect 1952 22374 2004 22380
rect 1676 22024 1728 22030
rect 1676 21966 1728 21972
rect 1688 21554 1716 21966
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1492 20936 1544 20942
rect 1492 20878 1544 20884
rect 1584 20936 1636 20942
rect 1860 20936 1912 20942
rect 1584 20878 1636 20884
rect 1780 20896 1860 20924
rect 1504 20466 1532 20878
rect 1584 20800 1636 20806
rect 1584 20742 1636 20748
rect 1492 20460 1544 20466
rect 1492 20402 1544 20408
rect 1308 19508 1360 19514
rect 1308 19450 1360 19456
rect 1216 16108 1268 16114
rect 1216 16050 1268 16056
rect 1228 15065 1256 16050
rect 1214 15056 1270 15065
rect 1214 14991 1270 15000
rect 1216 14952 1268 14958
rect 1216 14894 1268 14900
rect 1228 12889 1256 14894
rect 1214 12880 1270 12889
rect 1214 12815 1270 12824
rect 1214 5536 1270 5545
rect 1214 5471 1270 5480
rect 1228 4690 1256 5471
rect 1216 4684 1268 4690
rect 1216 4626 1268 4632
rect 1320 2774 1348 19450
rect 1504 19378 1532 20402
rect 1596 20398 1624 20742
rect 1584 20392 1636 20398
rect 1584 20334 1636 20340
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1504 19174 1532 19314
rect 1596 19310 1624 20334
rect 1780 20330 1808 20896
rect 1860 20878 1912 20884
rect 1768 20324 1820 20330
rect 1768 20266 1820 20272
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 19378 1716 19654
rect 1780 19446 1808 20266
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 1768 19440 1820 19446
rect 1768 19382 1820 19388
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 18290 1532 19110
rect 1872 18834 1900 19790
rect 1860 18828 1912 18834
rect 1860 18770 1912 18776
rect 1964 18290 1992 22374
rect 2056 21729 2084 22578
rect 2042 21720 2098 21729
rect 2042 21655 2098 21664
rect 2044 19236 2096 19242
rect 2044 19178 2096 19184
rect 1492 18284 1544 18290
rect 1492 18226 1544 18232
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 2056 18222 2084 19178
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 1952 18148 2004 18154
rect 1952 18090 2004 18096
rect 1964 17678 1992 18090
rect 2056 17746 2084 18158
rect 2044 17740 2096 17746
rect 2044 17682 2096 17688
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1688 17202 1716 17478
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1412 15881 1440 16526
rect 1398 15872 1454 15881
rect 1398 15807 1454 15816
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 14521 1440 15438
rect 1964 15434 1992 17614
rect 2056 16590 2084 17682
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 1952 15428 2004 15434
rect 1952 15370 2004 15376
rect 1492 14884 1544 14890
rect 1492 14826 1544 14832
rect 1398 14512 1454 14521
rect 1398 14447 1454 14456
rect 1504 14414 1532 14826
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1492 14408 1544 14414
rect 1492 14350 1544 14356
rect 1400 14340 1452 14346
rect 1400 14282 1452 14288
rect 1412 14074 1440 14282
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1504 12782 1532 14350
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1412 11393 1440 11698
rect 1398 11384 1454 11393
rect 1398 11319 1454 11328
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10713 1440 11086
rect 1398 10704 1454 10713
rect 1504 10674 1532 12718
rect 1596 12442 1624 12786
rect 1688 12646 1716 13806
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1688 12306 1716 12582
rect 1872 12374 1900 14758
rect 1964 13938 1992 14758
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1860 12368 1912 12374
rect 1860 12310 1912 12316
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 2044 12232 2096 12238
rect 1964 12192 2044 12220
rect 1964 11626 1992 12192
rect 2044 12174 2096 12180
rect 1952 11620 2004 11626
rect 1952 11562 2004 11568
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1398 10639 1454 10648
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1504 10198 1532 10610
rect 1492 10192 1544 10198
rect 1492 10134 1544 10140
rect 1688 10062 1716 10950
rect 1964 10130 1992 11562
rect 2148 11558 2176 23598
rect 2412 21956 2464 21962
rect 2412 21898 2464 21904
rect 2228 21548 2280 21554
rect 2228 21490 2280 21496
rect 2240 21146 2268 21490
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 2424 20602 2452 21898
rect 2412 20596 2464 20602
rect 2412 20538 2464 20544
rect 2228 19780 2280 19786
rect 2228 19722 2280 19728
rect 2240 19446 2268 19722
rect 2228 19440 2280 19446
rect 2228 19382 2280 19388
rect 2504 18692 2556 18698
rect 2504 18634 2556 18640
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 2332 18290 2360 18566
rect 2516 18426 2544 18634
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2320 17264 2372 17270
rect 2320 17206 2372 17212
rect 2332 16998 2360 17206
rect 2424 17066 2452 17478
rect 2412 17060 2464 17066
rect 2412 17002 2464 17008
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2240 15502 2268 16390
rect 2332 16046 2360 16934
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2332 14890 2360 15982
rect 2320 14884 2372 14890
rect 2320 14826 2372 14832
rect 2608 14414 2636 36858
rect 2792 36786 2820 37216
rect 2964 37198 3016 37204
rect 3054 37224 3110 37233
rect 3054 37159 3110 37168
rect 3068 37126 3096 37159
rect 2872 37120 2924 37126
rect 2872 37062 2924 37068
rect 3056 37120 3108 37126
rect 3056 37062 3108 37068
rect 2780 36780 2832 36786
rect 2780 36722 2832 36728
rect 2884 34762 2912 37062
rect 3516 36100 3568 36106
rect 3516 36042 3568 36048
rect 2964 36032 3016 36038
rect 2964 35974 3016 35980
rect 2976 35698 3004 35974
rect 2964 35692 3016 35698
rect 2964 35634 3016 35640
rect 3424 35692 3476 35698
rect 3424 35634 3476 35640
rect 2964 34944 3016 34950
rect 2964 34886 3016 34892
rect 2792 34734 2912 34762
rect 2792 33862 2820 34734
rect 2872 34604 2924 34610
rect 2872 34546 2924 34552
rect 2780 33856 2832 33862
rect 2780 33798 2832 33804
rect 2884 33658 2912 34546
rect 2976 34241 3004 34886
rect 3436 34746 3464 35634
rect 3424 34740 3476 34746
rect 3424 34682 3476 34688
rect 3056 34400 3108 34406
rect 3056 34342 3108 34348
rect 2962 34232 3018 34241
rect 2962 34167 3018 34176
rect 3068 34066 3096 34342
rect 3056 34060 3108 34066
rect 3056 34002 3108 34008
rect 2964 33856 3016 33862
rect 2964 33798 3016 33804
rect 2872 33652 2924 33658
rect 2872 33594 2924 33600
rect 2976 33561 3004 33798
rect 2962 33552 3018 33561
rect 2962 33487 3018 33496
rect 3148 33516 3200 33522
rect 3148 33458 3200 33464
rect 3160 33386 3188 33458
rect 3148 33380 3200 33386
rect 3148 33322 3200 33328
rect 3160 32910 3188 33322
rect 3148 32904 3200 32910
rect 3148 32846 3200 32852
rect 3332 32904 3384 32910
rect 3332 32846 3384 32852
rect 3148 32768 3200 32774
rect 3148 32710 3200 32716
rect 3160 32434 3188 32710
rect 3344 32570 3372 32846
rect 3332 32564 3384 32570
rect 3332 32506 3384 32512
rect 2780 32428 2832 32434
rect 2780 32370 2832 32376
rect 3148 32428 3200 32434
rect 3148 32370 3200 32376
rect 2688 30932 2740 30938
rect 2688 30874 2740 30880
rect 2700 30122 2728 30874
rect 2688 30116 2740 30122
rect 2688 30058 2740 30064
rect 2700 29186 2728 30058
rect 2792 29306 2820 32370
rect 2964 32360 3016 32366
rect 2964 32302 3016 32308
rect 2976 32026 3004 32302
rect 2964 32020 3016 32026
rect 2964 31962 3016 31968
rect 2964 31884 3016 31890
rect 2964 31826 3016 31832
rect 2872 30184 2924 30190
rect 2872 30126 2924 30132
rect 2884 29850 2912 30126
rect 2872 29844 2924 29850
rect 2872 29786 2924 29792
rect 2780 29300 2832 29306
rect 2780 29242 2832 29248
rect 2700 29158 2820 29186
rect 2976 29170 3004 31826
rect 3148 31816 3200 31822
rect 3148 31758 3200 31764
rect 3160 31482 3188 31758
rect 3528 31754 3556 36042
rect 3608 33924 3660 33930
rect 3608 33866 3660 33872
rect 3620 33658 3648 33866
rect 3608 33652 3660 33658
rect 3608 33594 3660 33600
rect 3344 31726 3556 31754
rect 3148 31476 3200 31482
rect 3148 31418 3200 31424
rect 3056 30728 3108 30734
rect 3056 30670 3108 30676
rect 2792 27878 2820 29158
rect 2964 29164 3016 29170
rect 2964 29106 3016 29112
rect 3068 29034 3096 30670
rect 3148 30592 3200 30598
rect 3146 30560 3148 30569
rect 3200 30560 3202 30569
rect 3146 30495 3202 30504
rect 3056 29028 3108 29034
rect 3056 28970 3108 28976
rect 3148 28484 3200 28490
rect 3148 28426 3200 28432
rect 3160 28014 3188 28426
rect 3344 28082 3372 31726
rect 3712 31414 3740 37946
rect 3804 37126 3832 39374
rect 3896 38196 3924 40582
rect 3976 40520 4028 40526
rect 3976 40462 4028 40468
rect 3988 40186 4016 40462
rect 3976 40180 4028 40186
rect 3976 40122 4028 40128
rect 4080 39506 4108 42026
rect 4448 41818 4476 42570
rect 4436 41812 4488 41818
rect 4436 41754 4488 41760
rect 4344 41676 4396 41682
rect 4344 41618 4396 41624
rect 4356 41414 4384 41618
rect 4436 41608 4488 41614
rect 4436 41550 4488 41556
rect 4264 41386 4384 41414
rect 4264 41070 4292 41386
rect 4448 41256 4476 41550
rect 4356 41228 4476 41256
rect 4252 41064 4304 41070
rect 4252 41006 4304 41012
rect 4160 40996 4212 41002
rect 4160 40938 4212 40944
rect 4172 40526 4200 40938
rect 4264 40594 4292 41006
rect 4252 40588 4304 40594
rect 4252 40530 4304 40536
rect 4160 40520 4212 40526
rect 4160 40462 4212 40468
rect 4172 39522 4200 40462
rect 4264 39658 4292 40530
rect 4356 39846 4384 41228
rect 4436 41132 4488 41138
rect 4436 41074 4488 41080
rect 4448 40526 4476 41074
rect 4436 40520 4488 40526
rect 4436 40462 4488 40468
rect 4540 39914 4568 43250
rect 4712 41608 4764 41614
rect 4632 41556 4712 41562
rect 4632 41550 4764 41556
rect 4632 41534 4752 41550
rect 4632 41414 4660 41534
rect 4632 41386 4752 41414
rect 4724 41070 4752 41386
rect 4712 41064 4764 41070
rect 4712 41006 4764 41012
rect 4804 40928 4856 40934
rect 4804 40870 4856 40876
rect 4620 40520 4672 40526
rect 4620 40462 4672 40468
rect 4528 39908 4580 39914
rect 4528 39850 4580 39856
rect 4344 39840 4396 39846
rect 4344 39782 4396 39788
rect 4264 39630 4384 39658
rect 4068 39500 4120 39506
rect 4172 39494 4292 39522
rect 4068 39442 4120 39448
rect 3976 39296 4028 39302
rect 3976 39238 4028 39244
rect 3988 38418 4016 39238
rect 4160 38956 4212 38962
rect 4160 38898 4212 38904
rect 4172 38554 4200 38898
rect 4264 38894 4292 39494
rect 4356 38894 4384 39630
rect 4528 39568 4580 39574
rect 4528 39510 4580 39516
rect 4436 38956 4488 38962
rect 4540 38944 4568 39510
rect 4632 38962 4660 40462
rect 4816 40186 4844 40870
rect 5092 40526 5120 43250
rect 5184 43110 5212 43862
rect 5552 43790 5580 44202
rect 5540 43784 5592 43790
rect 5540 43726 5592 43732
rect 5356 43648 5408 43654
rect 5356 43590 5408 43596
rect 5172 43104 5224 43110
rect 5172 43046 5224 43052
rect 5184 42906 5212 43046
rect 5172 42900 5224 42906
rect 5172 42842 5224 42848
rect 5264 42152 5316 42158
rect 5264 42094 5316 42100
rect 5276 41682 5304 42094
rect 5368 42022 5396 43590
rect 5356 42016 5408 42022
rect 5356 41958 5408 41964
rect 5368 41750 5396 41958
rect 5356 41744 5408 41750
rect 5356 41686 5408 41692
rect 5264 41676 5316 41682
rect 5264 41618 5316 41624
rect 5172 41608 5224 41614
rect 5172 41550 5224 41556
rect 5184 41206 5212 41550
rect 5172 41200 5224 41206
rect 5172 41142 5224 41148
rect 5080 40520 5132 40526
rect 5080 40462 5132 40468
rect 4804 40180 4856 40186
rect 4804 40122 4856 40128
rect 4896 39840 4948 39846
rect 4896 39782 4948 39788
rect 4712 39296 4764 39302
rect 4712 39238 4764 39244
rect 4724 39030 4752 39238
rect 4712 39024 4764 39030
rect 4712 38966 4764 38972
rect 4488 38916 4568 38944
rect 4436 38898 4488 38904
rect 4252 38888 4304 38894
rect 4252 38830 4304 38836
rect 4344 38888 4396 38894
rect 4344 38830 4396 38836
rect 4252 38752 4304 38758
rect 4252 38694 4304 38700
rect 4160 38548 4212 38554
rect 4160 38490 4212 38496
rect 3976 38412 4028 38418
rect 3976 38354 4028 38360
rect 4264 38350 4292 38694
rect 4068 38344 4120 38350
rect 4252 38344 4304 38350
rect 4120 38304 4200 38332
rect 4068 38286 4120 38292
rect 3896 38168 4108 38196
rect 3976 37256 4028 37262
rect 3976 37198 4028 37204
rect 3792 37120 3844 37126
rect 3792 37062 3844 37068
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 3792 35488 3844 35494
rect 3792 35430 3844 35436
rect 3804 35018 3832 35430
rect 3792 35012 3844 35018
rect 3792 34954 3844 34960
rect 3804 34610 3832 34954
rect 3792 34604 3844 34610
rect 3792 34546 3844 34552
rect 3896 33998 3924 37062
rect 3988 36650 4016 37198
rect 3976 36644 4028 36650
rect 3976 36586 4028 36592
rect 4080 34610 4108 38168
rect 4172 37670 4200 38304
rect 4252 38286 4304 38292
rect 4356 38214 4384 38830
rect 4344 38208 4396 38214
rect 4344 38150 4396 38156
rect 4356 37874 4384 38150
rect 4344 37868 4396 37874
rect 4344 37810 4396 37816
rect 4436 37800 4488 37806
rect 4436 37742 4488 37748
rect 4160 37664 4212 37670
rect 4160 37606 4212 37612
rect 4448 36922 4476 37742
rect 4436 36916 4488 36922
rect 4436 36858 4488 36864
rect 4160 36780 4212 36786
rect 4160 36722 4212 36728
rect 4068 34604 4120 34610
rect 4068 34546 4120 34552
rect 4068 34468 4120 34474
rect 4068 34410 4120 34416
rect 3976 34400 4028 34406
rect 3976 34342 4028 34348
rect 3884 33992 3936 33998
rect 3884 33934 3936 33940
rect 3792 33856 3844 33862
rect 3792 33798 3844 33804
rect 3804 33522 3832 33798
rect 3792 33516 3844 33522
rect 3792 33458 3844 33464
rect 3988 33454 4016 34342
rect 4080 33522 4108 34410
rect 4068 33516 4120 33522
rect 4068 33458 4120 33464
rect 3976 33448 4028 33454
rect 3976 33390 4028 33396
rect 3884 32836 3936 32842
rect 3884 32778 3936 32784
rect 3896 32570 3924 32778
rect 3884 32564 3936 32570
rect 3884 32506 3936 32512
rect 3988 32348 4016 33390
rect 4080 32892 4108 33458
rect 4172 33318 4200 36722
rect 4252 36168 4304 36174
rect 4252 36110 4304 36116
rect 4264 35086 4292 36110
rect 4436 35692 4488 35698
rect 4436 35634 4488 35640
rect 4448 35290 4476 35634
rect 4436 35284 4488 35290
rect 4436 35226 4488 35232
rect 4252 35080 4304 35086
rect 4252 35022 4304 35028
rect 4264 33386 4292 35022
rect 4344 34604 4396 34610
rect 4344 34546 4396 34552
rect 4356 33522 4384 34546
rect 4344 33516 4396 33522
rect 4396 33476 4476 33504
rect 4344 33458 4396 33464
rect 4252 33380 4304 33386
rect 4252 33322 4304 33328
rect 4160 33312 4212 33318
rect 4160 33254 4212 33260
rect 4080 32864 4292 32892
rect 4264 32434 4292 32864
rect 4448 32434 4476 33476
rect 4252 32428 4304 32434
rect 4252 32370 4304 32376
rect 4436 32428 4488 32434
rect 4436 32370 4488 32376
rect 4068 32360 4120 32366
rect 3988 32320 4068 32348
rect 4068 32302 4120 32308
rect 4080 31958 4108 32302
rect 3792 31952 3844 31958
rect 3792 31894 3844 31900
rect 4068 31952 4120 31958
rect 4068 31894 4120 31900
rect 3700 31408 3752 31414
rect 3700 31350 3752 31356
rect 3804 31346 3832 31894
rect 4160 31680 4212 31686
rect 4160 31622 4212 31628
rect 3792 31340 3844 31346
rect 3792 31282 3844 31288
rect 3516 31204 3568 31210
rect 3516 31146 3568 31152
rect 3424 31136 3476 31142
rect 3424 31078 3476 31084
rect 3436 30326 3464 31078
rect 3528 30802 3556 31146
rect 4172 31124 4200 31622
rect 4264 31414 4292 32370
rect 4448 31634 4476 32370
rect 4540 32298 4568 38916
rect 4620 38956 4672 38962
rect 4620 38898 4672 38904
rect 4632 37738 4660 38898
rect 4620 37732 4672 37738
rect 4620 37674 4672 37680
rect 4908 36718 4936 39782
rect 4988 38820 5040 38826
rect 4988 38762 5040 38768
rect 5000 38418 5028 38762
rect 4988 38412 5040 38418
rect 4988 38354 5040 38360
rect 4988 37256 5040 37262
rect 4988 37198 5040 37204
rect 5000 36922 5028 37198
rect 4988 36916 5040 36922
rect 4988 36858 5040 36864
rect 4896 36712 4948 36718
rect 4896 36654 4948 36660
rect 5092 36038 5120 40462
rect 5172 36780 5224 36786
rect 5172 36722 5224 36728
rect 5184 36378 5212 36722
rect 5172 36372 5224 36378
rect 5172 36314 5224 36320
rect 5080 36032 5132 36038
rect 5080 35974 5132 35980
rect 4896 35488 4948 35494
rect 4896 35430 4948 35436
rect 4908 35154 4936 35430
rect 4896 35148 4948 35154
rect 4896 35090 4948 35096
rect 4712 35012 4764 35018
rect 4712 34954 4764 34960
rect 4724 34746 4752 34954
rect 4896 34944 4948 34950
rect 4896 34886 4948 34892
rect 4712 34740 4764 34746
rect 4712 34682 4764 34688
rect 4908 34610 4936 34886
rect 5276 34610 5304 41618
rect 5368 41002 5396 41686
rect 5448 41064 5500 41070
rect 5448 41006 5500 41012
rect 5356 40996 5408 41002
rect 5356 40938 5408 40944
rect 5368 39846 5396 40938
rect 5460 40458 5488 41006
rect 5448 40452 5500 40458
rect 5448 40394 5500 40400
rect 5356 39840 5408 39846
rect 5356 39782 5408 39788
rect 5460 39658 5488 40394
rect 5368 39630 5488 39658
rect 4896 34604 4948 34610
rect 4896 34546 4948 34552
rect 5080 34604 5132 34610
rect 5080 34546 5132 34552
rect 5264 34604 5316 34610
rect 5264 34546 5316 34552
rect 5092 34406 5120 34546
rect 5080 34400 5132 34406
rect 5080 34342 5132 34348
rect 5368 34134 5396 39630
rect 5448 37664 5500 37670
rect 5448 37606 5500 37612
rect 5460 37330 5488 37606
rect 5448 37324 5500 37330
rect 5448 37266 5500 37272
rect 5552 36242 5580 43726
rect 5632 43716 5684 43722
rect 5632 43658 5684 43664
rect 5644 41818 5672 43658
rect 5736 42634 5764 44882
rect 6552 44872 6604 44878
rect 6552 44814 6604 44820
rect 8392 44872 8444 44878
rect 8392 44814 8444 44820
rect 6276 44736 6328 44742
rect 6276 44678 6328 44684
rect 5915 44092 6223 44112
rect 5915 44090 5921 44092
rect 5977 44090 6001 44092
rect 6057 44090 6081 44092
rect 6137 44090 6161 44092
rect 6217 44090 6223 44092
rect 5977 44038 5979 44090
rect 6159 44038 6161 44090
rect 5915 44036 5921 44038
rect 5977 44036 6001 44038
rect 6057 44036 6081 44038
rect 6137 44036 6161 44038
rect 6217 44036 6223 44038
rect 5915 44016 6223 44036
rect 6288 43926 6316 44678
rect 6564 44538 6592 44814
rect 7012 44804 7064 44810
rect 7012 44746 7064 44752
rect 7024 44538 7052 44746
rect 7196 44736 7248 44742
rect 7196 44678 7248 44684
rect 6552 44532 6604 44538
rect 6552 44474 6604 44480
rect 7012 44532 7064 44538
rect 7012 44474 7064 44480
rect 7208 44402 7236 44678
rect 7564 44532 7616 44538
rect 7564 44474 7616 44480
rect 7576 44402 7604 44474
rect 6368 44396 6420 44402
rect 6368 44338 6420 44344
rect 7196 44396 7248 44402
rect 7196 44338 7248 44344
rect 7564 44396 7616 44402
rect 7564 44338 7616 44344
rect 7748 44396 7800 44402
rect 7748 44338 7800 44344
rect 8300 44396 8352 44402
rect 8300 44338 8352 44344
rect 6380 43994 6408 44338
rect 7380 44328 7432 44334
rect 7380 44270 7432 44276
rect 6368 43988 6420 43994
rect 6368 43930 6420 43936
rect 6276 43920 6328 43926
rect 6276 43862 6328 43868
rect 7392 43858 7420 44270
rect 7380 43852 7432 43858
rect 7380 43794 7432 43800
rect 5908 43784 5960 43790
rect 5908 43726 5960 43732
rect 6644 43784 6696 43790
rect 6644 43726 6696 43732
rect 5920 43314 5948 43726
rect 5908 43308 5960 43314
rect 5908 43250 5960 43256
rect 5915 43004 6223 43024
rect 5915 43002 5921 43004
rect 5977 43002 6001 43004
rect 6057 43002 6081 43004
rect 6137 43002 6161 43004
rect 6217 43002 6223 43004
rect 5977 42950 5979 43002
rect 6159 42950 6161 43002
rect 5915 42948 5921 42950
rect 5977 42948 6001 42950
rect 6057 42948 6081 42950
rect 6137 42948 6161 42950
rect 6217 42948 6223 42950
rect 5915 42928 6223 42948
rect 5908 42696 5960 42702
rect 5908 42638 5960 42644
rect 5724 42628 5776 42634
rect 5724 42570 5776 42576
rect 5816 42560 5868 42566
rect 5816 42502 5868 42508
rect 5632 41812 5684 41818
rect 5632 41754 5684 41760
rect 5828 41546 5856 42502
rect 5920 42226 5948 42638
rect 6552 42288 6604 42294
rect 6552 42230 6604 42236
rect 5908 42220 5960 42226
rect 5908 42162 5960 42168
rect 6276 42220 6328 42226
rect 6276 42162 6328 42168
rect 5915 41916 6223 41936
rect 5915 41914 5921 41916
rect 5977 41914 6001 41916
rect 6057 41914 6081 41916
rect 6137 41914 6161 41916
rect 6217 41914 6223 41916
rect 5977 41862 5979 41914
rect 6159 41862 6161 41914
rect 5915 41860 5921 41862
rect 5977 41860 6001 41862
rect 6057 41860 6081 41862
rect 6137 41860 6161 41862
rect 6217 41860 6223 41862
rect 5915 41840 6223 41860
rect 6288 41750 6316 42162
rect 6276 41744 6328 41750
rect 6276 41686 6328 41692
rect 5816 41540 5868 41546
rect 5816 41482 5868 41488
rect 5816 41132 5868 41138
rect 5816 41074 5868 41080
rect 5724 40996 5776 41002
rect 5724 40938 5776 40944
rect 5736 40050 5764 40938
rect 5724 40044 5776 40050
rect 5724 39986 5776 39992
rect 5828 39642 5856 41074
rect 6288 41002 6316 41686
rect 6368 41540 6420 41546
rect 6368 41482 6420 41488
rect 6380 41414 6408 41482
rect 6380 41386 6500 41414
rect 6368 41200 6420 41206
rect 6368 41142 6420 41148
rect 6276 40996 6328 41002
rect 6276 40938 6328 40944
rect 5915 40828 6223 40848
rect 5915 40826 5921 40828
rect 5977 40826 6001 40828
rect 6057 40826 6081 40828
rect 6137 40826 6161 40828
rect 6217 40826 6223 40828
rect 5977 40774 5979 40826
rect 6159 40774 6161 40826
rect 5915 40772 5921 40774
rect 5977 40772 6001 40774
rect 6057 40772 6081 40774
rect 6137 40772 6161 40774
rect 6217 40772 6223 40774
rect 5915 40752 6223 40772
rect 5915 39740 6223 39760
rect 5915 39738 5921 39740
rect 5977 39738 6001 39740
rect 6057 39738 6081 39740
rect 6137 39738 6161 39740
rect 6217 39738 6223 39740
rect 5977 39686 5979 39738
rect 6159 39686 6161 39738
rect 5915 39684 5921 39686
rect 5977 39684 6001 39686
rect 6057 39684 6081 39686
rect 6137 39684 6161 39686
rect 6217 39684 6223 39686
rect 5915 39664 6223 39684
rect 5816 39636 5868 39642
rect 5816 39578 5868 39584
rect 5828 39438 5856 39578
rect 6380 39506 6408 41142
rect 6472 40662 6500 41386
rect 6564 41274 6592 42230
rect 6656 41614 6684 43726
rect 7196 43648 7248 43654
rect 7196 43590 7248 43596
rect 7288 43648 7340 43654
rect 7288 43590 7340 43596
rect 7208 43450 7236 43590
rect 7196 43444 7248 43450
rect 7196 43386 7248 43392
rect 7012 43308 7064 43314
rect 7012 43250 7064 43256
rect 6736 43240 6788 43246
rect 6736 43182 6788 43188
rect 6748 42362 6776 43182
rect 6920 43104 6972 43110
rect 6920 43046 6972 43052
rect 6736 42356 6788 42362
rect 6736 42298 6788 42304
rect 6932 42226 6960 43046
rect 7024 42906 7052 43250
rect 7012 42900 7064 42906
rect 7012 42842 7064 42848
rect 7208 42702 7236 43386
rect 7196 42696 7248 42702
rect 7196 42638 7248 42644
rect 6920 42220 6972 42226
rect 6920 42162 6972 42168
rect 7012 41744 7064 41750
rect 7012 41686 7064 41692
rect 6644 41608 6696 41614
rect 6644 41550 6696 41556
rect 6552 41268 6604 41274
rect 6552 41210 6604 41216
rect 6460 40656 6512 40662
rect 6460 40598 6512 40604
rect 6368 39500 6420 39506
rect 6368 39442 6420 39448
rect 5816 39432 5868 39438
rect 5816 39374 5868 39380
rect 6380 39098 6408 39442
rect 6472 39438 6500 40598
rect 6564 40526 6592 41210
rect 6656 41138 6684 41550
rect 6920 41200 6972 41206
rect 6920 41142 6972 41148
rect 6644 41132 6696 41138
rect 6644 41074 6696 41080
rect 6736 41132 6788 41138
rect 6736 41074 6788 41080
rect 6748 40730 6776 41074
rect 6932 41070 6960 41142
rect 6920 41064 6972 41070
rect 6920 41006 6972 41012
rect 6828 40996 6880 41002
rect 6828 40938 6880 40944
rect 6840 40730 6868 40938
rect 6736 40724 6788 40730
rect 6736 40666 6788 40672
rect 6828 40724 6880 40730
rect 6828 40666 6880 40672
rect 6552 40520 6604 40526
rect 6552 40462 6604 40468
rect 6920 40520 6972 40526
rect 6920 40462 6972 40468
rect 6736 40452 6788 40458
rect 6736 40394 6788 40400
rect 6748 40050 6776 40394
rect 6736 40044 6788 40050
rect 6736 39986 6788 39992
rect 6644 39636 6696 39642
rect 6644 39578 6696 39584
rect 6656 39438 6684 39578
rect 6748 39438 6776 39986
rect 6932 39846 6960 40462
rect 6920 39840 6972 39846
rect 6920 39782 6972 39788
rect 6932 39438 6960 39782
rect 7024 39574 7052 41686
rect 7196 40928 7248 40934
rect 7196 40870 7248 40876
rect 7208 40050 7236 40870
rect 7300 40662 7328 43590
rect 7392 42702 7420 43794
rect 7380 42696 7432 42702
rect 7380 42638 7432 42644
rect 7392 42362 7420 42638
rect 7380 42356 7432 42362
rect 7380 42298 7432 42304
rect 7472 41472 7524 41478
rect 7472 41414 7524 41420
rect 7288 40656 7340 40662
rect 7288 40598 7340 40604
rect 7288 40112 7340 40118
rect 7288 40054 7340 40060
rect 7196 40044 7248 40050
rect 7196 39986 7248 39992
rect 7012 39568 7064 39574
rect 7012 39510 7064 39516
rect 6460 39432 6512 39438
rect 6460 39374 6512 39380
rect 6644 39432 6696 39438
rect 6644 39374 6696 39380
rect 6736 39432 6788 39438
rect 6736 39374 6788 39380
rect 6920 39432 6972 39438
rect 6920 39374 6972 39380
rect 6368 39092 6420 39098
rect 6368 39034 6420 39040
rect 5816 38956 5868 38962
rect 5816 38898 5868 38904
rect 5724 38752 5776 38758
rect 5724 38694 5776 38700
rect 5736 37874 5764 38694
rect 5828 38350 5856 38898
rect 6472 38758 6500 39374
rect 6828 39296 6880 39302
rect 6828 39238 6880 39244
rect 6460 38752 6512 38758
rect 6460 38694 6512 38700
rect 5915 38652 6223 38672
rect 5915 38650 5921 38652
rect 5977 38650 6001 38652
rect 6057 38650 6081 38652
rect 6137 38650 6161 38652
rect 6217 38650 6223 38652
rect 5977 38598 5979 38650
rect 6159 38598 6161 38650
rect 5915 38596 5921 38598
rect 5977 38596 6001 38598
rect 6057 38596 6081 38598
rect 6137 38596 6161 38598
rect 6217 38596 6223 38598
rect 5915 38576 6223 38596
rect 5816 38344 5868 38350
rect 5816 38286 5868 38292
rect 6368 37936 6420 37942
rect 6368 37878 6420 37884
rect 6552 37936 6604 37942
rect 6552 37878 6604 37884
rect 5724 37868 5776 37874
rect 5724 37810 5776 37816
rect 6380 37806 6408 37878
rect 6368 37800 6420 37806
rect 6368 37742 6420 37748
rect 5915 37564 6223 37584
rect 5915 37562 5921 37564
rect 5977 37562 6001 37564
rect 6057 37562 6081 37564
rect 6137 37562 6161 37564
rect 6217 37562 6223 37564
rect 5977 37510 5979 37562
rect 6159 37510 6161 37562
rect 5915 37508 5921 37510
rect 5977 37508 6001 37510
rect 6057 37508 6081 37510
rect 6137 37508 6161 37510
rect 6217 37508 6223 37510
rect 5915 37488 6223 37508
rect 5632 36780 5684 36786
rect 5632 36722 5684 36728
rect 5540 36236 5592 36242
rect 5540 36178 5592 36184
rect 5448 36100 5500 36106
rect 5448 36042 5500 36048
rect 5460 35442 5488 36042
rect 5540 35488 5592 35494
rect 5460 35436 5540 35442
rect 5460 35430 5592 35436
rect 5460 35414 5580 35430
rect 4804 34128 4856 34134
rect 4804 34070 4856 34076
rect 5356 34128 5408 34134
rect 5356 34070 5408 34076
rect 4816 33590 4844 34070
rect 4804 33584 4856 33590
rect 4804 33526 4856 33532
rect 5172 32768 5224 32774
rect 5172 32710 5224 32716
rect 5184 32502 5212 32710
rect 5172 32496 5224 32502
rect 5172 32438 5224 32444
rect 4528 32292 4580 32298
rect 4528 32234 4580 32240
rect 4528 31816 4580 31822
rect 4528 31758 4580 31764
rect 5172 31816 5224 31822
rect 5172 31758 5224 31764
rect 4540 31634 4568 31758
rect 4804 31748 4856 31754
rect 4804 31690 4856 31696
rect 4448 31606 4568 31634
rect 4252 31408 4304 31414
rect 4252 31350 4304 31356
rect 4448 31346 4476 31606
rect 4436 31340 4488 31346
rect 4436 31282 4488 31288
rect 4252 31136 4304 31142
rect 4172 31096 4252 31124
rect 4252 31078 4304 31084
rect 3516 30796 3568 30802
rect 3516 30738 3568 30744
rect 4160 30592 4212 30598
rect 4160 30534 4212 30540
rect 3424 30320 3476 30326
rect 3424 30262 3476 30268
rect 4172 29238 4200 30534
rect 4264 30394 4292 31078
rect 4816 30734 4844 31690
rect 5080 31204 5132 31210
rect 5080 31146 5132 31152
rect 5092 30802 5120 31146
rect 5080 30796 5132 30802
rect 5080 30738 5132 30744
rect 4528 30728 4580 30734
rect 4528 30670 4580 30676
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 4804 30728 4856 30734
rect 4856 30688 4936 30716
rect 4804 30670 4856 30676
rect 4540 30394 4568 30670
rect 4252 30388 4304 30394
rect 4252 30330 4304 30336
rect 4528 30388 4580 30394
rect 4528 30330 4580 30336
rect 4620 30252 4672 30258
rect 4620 30194 4672 30200
rect 4632 29646 4660 30194
rect 4620 29640 4672 29646
rect 4620 29582 4672 29588
rect 4436 29504 4488 29510
rect 4436 29446 4488 29452
rect 4160 29232 4212 29238
rect 4160 29174 4212 29180
rect 3792 29096 3844 29102
rect 3792 29038 3844 29044
rect 3804 28762 3832 29038
rect 3792 28756 3844 28762
rect 3792 28698 3844 28704
rect 4448 28558 4476 29446
rect 4632 28558 4660 29582
rect 4724 29306 4752 30670
rect 4804 30320 4856 30326
rect 4804 30262 4856 30268
rect 4816 29850 4844 30262
rect 4908 30122 4936 30688
rect 5092 30190 5120 30738
rect 5184 30734 5212 31758
rect 5172 30728 5224 30734
rect 5172 30670 5224 30676
rect 5460 30326 5488 35414
rect 5644 33658 5672 36722
rect 5915 36476 6223 36496
rect 5915 36474 5921 36476
rect 5977 36474 6001 36476
rect 6057 36474 6081 36476
rect 6137 36474 6161 36476
rect 6217 36474 6223 36476
rect 5977 36422 5979 36474
rect 6159 36422 6161 36474
rect 5915 36420 5921 36422
rect 5977 36420 6001 36422
rect 6057 36420 6081 36422
rect 6137 36420 6161 36422
rect 6217 36420 6223 36422
rect 5915 36400 6223 36420
rect 6460 36236 6512 36242
rect 6460 36178 6512 36184
rect 6276 35692 6328 35698
rect 6276 35634 6328 35640
rect 5915 35388 6223 35408
rect 5915 35386 5921 35388
rect 5977 35386 6001 35388
rect 6057 35386 6081 35388
rect 6137 35386 6161 35388
rect 6217 35386 6223 35388
rect 5977 35334 5979 35386
rect 6159 35334 6161 35386
rect 5915 35332 5921 35334
rect 5977 35332 6001 35334
rect 6057 35332 6081 35334
rect 6137 35332 6161 35334
rect 6217 35332 6223 35334
rect 5915 35312 6223 35332
rect 5724 34604 5776 34610
rect 5724 34546 5776 34552
rect 5632 33652 5684 33658
rect 5632 33594 5684 33600
rect 5736 33114 5764 34546
rect 5915 34300 6223 34320
rect 5915 34298 5921 34300
rect 5977 34298 6001 34300
rect 6057 34298 6081 34300
rect 6137 34298 6161 34300
rect 6217 34298 6223 34300
rect 5977 34246 5979 34298
rect 6159 34246 6161 34298
rect 5915 34244 5921 34246
rect 5977 34244 6001 34246
rect 6057 34244 6081 34246
rect 6137 34244 6161 34246
rect 6217 34244 6223 34246
rect 5915 34224 6223 34244
rect 6288 34202 6316 35634
rect 6368 35080 6420 35086
rect 6368 35022 6420 35028
rect 6276 34196 6328 34202
rect 6276 34138 6328 34144
rect 6288 33522 6316 34138
rect 6276 33516 6328 33522
rect 6276 33458 6328 33464
rect 5915 33212 6223 33232
rect 5915 33210 5921 33212
rect 5977 33210 6001 33212
rect 6057 33210 6081 33212
rect 6137 33210 6161 33212
rect 6217 33210 6223 33212
rect 5977 33158 5979 33210
rect 6159 33158 6161 33210
rect 5915 33156 5921 33158
rect 5977 33156 6001 33158
rect 6057 33156 6081 33158
rect 6137 33156 6161 33158
rect 6217 33156 6223 33158
rect 5915 33136 6223 33156
rect 5724 33108 5776 33114
rect 5724 33050 5776 33056
rect 5632 32836 5684 32842
rect 5632 32778 5684 32784
rect 5644 32434 5672 32778
rect 6380 32450 6408 35022
rect 6472 34406 6500 36178
rect 6564 34898 6592 37878
rect 6840 36922 6868 39238
rect 6932 38418 6960 39374
rect 7196 39296 7248 39302
rect 7196 39238 7248 39244
rect 7208 39030 7236 39238
rect 7196 39024 7248 39030
rect 7196 38966 7248 38972
rect 7012 38752 7064 38758
rect 7012 38694 7064 38700
rect 7024 38486 7052 38694
rect 7012 38480 7064 38486
rect 7012 38422 7064 38428
rect 6920 38412 6972 38418
rect 6920 38354 6972 38360
rect 7024 38298 7052 38422
rect 7300 38350 7328 40054
rect 7380 40044 7432 40050
rect 7380 39986 7432 39992
rect 7392 38350 7420 39986
rect 6932 38270 7052 38298
rect 7288 38344 7340 38350
rect 7288 38286 7340 38292
rect 7380 38344 7432 38350
rect 7380 38286 7432 38292
rect 6828 36916 6880 36922
rect 6828 36858 6880 36864
rect 6736 36848 6788 36854
rect 6736 36790 6788 36796
rect 6644 36576 6696 36582
rect 6644 36518 6696 36524
rect 6656 36242 6684 36518
rect 6748 36242 6776 36790
rect 6644 36236 6696 36242
rect 6644 36178 6696 36184
rect 6736 36236 6788 36242
rect 6736 36178 6788 36184
rect 6736 35692 6788 35698
rect 6840 35680 6868 36858
rect 6788 35652 6868 35680
rect 6736 35634 6788 35640
rect 6564 34870 6684 34898
rect 6460 34400 6512 34406
rect 6460 34342 6512 34348
rect 6552 33856 6604 33862
rect 6552 33798 6604 33804
rect 6564 33522 6592 33798
rect 6552 33516 6604 33522
rect 6552 33458 6604 33464
rect 5632 32428 5684 32434
rect 6380 32422 6500 32450
rect 5632 32370 5684 32376
rect 5644 31890 5672 32370
rect 6368 32360 6420 32366
rect 6368 32302 6420 32308
rect 5915 32124 6223 32144
rect 5915 32122 5921 32124
rect 5977 32122 6001 32124
rect 6057 32122 6081 32124
rect 6137 32122 6161 32124
rect 6217 32122 6223 32124
rect 5977 32070 5979 32122
rect 6159 32070 6161 32122
rect 5915 32068 5921 32070
rect 5977 32068 6001 32070
rect 6057 32068 6081 32070
rect 6137 32068 6161 32070
rect 6217 32068 6223 32070
rect 5915 32048 6223 32068
rect 6380 32026 6408 32302
rect 6368 32020 6420 32026
rect 6368 31962 6420 31968
rect 5632 31884 5684 31890
rect 5632 31826 5684 31832
rect 6472 31822 6500 32422
rect 6656 32298 6684 34870
rect 6932 34678 6960 38270
rect 7104 38208 7156 38214
rect 7104 38150 7156 38156
rect 7116 37262 7144 38150
rect 7300 37466 7328 38286
rect 7288 37460 7340 37466
rect 7288 37402 7340 37408
rect 7196 37392 7248 37398
rect 7196 37334 7248 37340
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 7208 36786 7236 37334
rect 7196 36780 7248 36786
rect 7196 36722 7248 36728
rect 7208 36378 7236 36722
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 7012 34944 7064 34950
rect 7012 34886 7064 34892
rect 6920 34672 6972 34678
rect 6920 34614 6972 34620
rect 7024 34610 7052 34886
rect 7012 34604 7064 34610
rect 7012 34546 7064 34552
rect 7288 34536 7340 34542
rect 7288 34478 7340 34484
rect 7104 33312 7156 33318
rect 7104 33254 7156 33260
rect 6828 32768 6880 32774
rect 6828 32710 6880 32716
rect 6644 32292 6696 32298
rect 6644 32234 6696 32240
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 6368 31136 6420 31142
rect 6368 31078 6420 31084
rect 5915 31036 6223 31056
rect 5915 31034 5921 31036
rect 5977 31034 6001 31036
rect 6057 31034 6081 31036
rect 6137 31034 6161 31036
rect 6217 31034 6223 31036
rect 5977 30982 5979 31034
rect 6159 30982 6161 31034
rect 5915 30980 5921 30982
rect 5977 30980 6001 30982
rect 6057 30980 6081 30982
rect 6137 30980 6161 30982
rect 6217 30980 6223 30982
rect 5915 30960 6223 30980
rect 6380 30734 6408 31078
rect 6368 30728 6420 30734
rect 6368 30670 6420 30676
rect 6564 30598 6592 31282
rect 6552 30592 6604 30598
rect 6552 30534 6604 30540
rect 5448 30320 5500 30326
rect 5448 30262 5500 30268
rect 5356 30252 5408 30258
rect 5356 30194 5408 30200
rect 5080 30184 5132 30190
rect 5080 30126 5132 30132
rect 5368 30122 5396 30194
rect 4896 30116 4948 30122
rect 4896 30058 4948 30064
rect 5356 30116 5408 30122
rect 5356 30058 5408 30064
rect 6368 30048 6420 30054
rect 6368 29990 6420 29996
rect 5915 29948 6223 29968
rect 5915 29946 5921 29948
rect 5977 29946 6001 29948
rect 6057 29946 6081 29948
rect 6137 29946 6161 29948
rect 6217 29946 6223 29948
rect 5977 29894 5979 29946
rect 6159 29894 6161 29946
rect 5915 29892 5921 29894
rect 5977 29892 6001 29894
rect 6057 29892 6081 29894
rect 6137 29892 6161 29894
rect 6217 29892 6223 29894
rect 5915 29872 6223 29892
rect 4804 29844 4856 29850
rect 4804 29786 4856 29792
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 5828 29306 5856 29582
rect 6380 29578 6408 29990
rect 6368 29572 6420 29578
rect 6368 29514 6420 29520
rect 6552 29572 6604 29578
rect 6552 29514 6604 29520
rect 4712 29300 4764 29306
rect 4712 29242 4764 29248
rect 5816 29300 5868 29306
rect 5816 29242 5868 29248
rect 5632 29164 5684 29170
rect 5632 29106 5684 29112
rect 5644 28762 5672 29106
rect 5915 28860 6223 28880
rect 5915 28858 5921 28860
rect 5977 28858 6001 28860
rect 6057 28858 6081 28860
rect 6137 28858 6161 28860
rect 6217 28858 6223 28860
rect 5977 28806 5979 28858
rect 6159 28806 6161 28858
rect 5915 28804 5921 28806
rect 5977 28804 6001 28806
rect 6057 28804 6081 28806
rect 6137 28804 6161 28806
rect 6217 28804 6223 28806
rect 5915 28784 6223 28804
rect 5632 28756 5684 28762
rect 5632 28698 5684 28704
rect 4436 28552 4488 28558
rect 4436 28494 4488 28500
rect 4620 28552 4672 28558
rect 4620 28494 4672 28500
rect 6460 28552 6512 28558
rect 6460 28494 6512 28500
rect 3332 28076 3384 28082
rect 3332 28018 3384 28024
rect 3148 28008 3200 28014
rect 3148 27950 3200 27956
rect 2780 27872 2832 27878
rect 2780 27814 2832 27820
rect 3160 27470 3188 27950
rect 3344 27674 3372 28018
rect 3608 27872 3660 27878
rect 3608 27814 3660 27820
rect 3332 27668 3384 27674
rect 3332 27610 3384 27616
rect 3148 27464 3200 27470
rect 3148 27406 3200 27412
rect 3160 26382 3188 27406
rect 2872 26376 2924 26382
rect 2872 26318 2924 26324
rect 3148 26376 3200 26382
rect 3148 26318 3200 26324
rect 2884 26042 2912 26318
rect 2964 26240 3016 26246
rect 2964 26182 3016 26188
rect 2872 26036 2924 26042
rect 2872 25978 2924 25984
rect 2976 25906 3004 26182
rect 3160 25906 3188 26318
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 3148 25900 3200 25906
rect 3148 25842 3200 25848
rect 3160 24818 3188 25842
rect 3148 24812 3200 24818
rect 3148 24754 3200 24760
rect 3160 24274 3188 24754
rect 3148 24268 3200 24274
rect 3148 24210 3200 24216
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2792 22409 2820 22578
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 2778 22400 2834 22409
rect 2778 22335 2834 22344
rect 2780 21412 2832 21418
rect 2780 21354 2832 21360
rect 2792 19718 2820 21354
rect 2884 20346 2912 22510
rect 2964 21888 3016 21894
rect 2964 21830 3016 21836
rect 2976 20874 3004 21830
rect 3240 21548 3292 21554
rect 3240 21490 3292 21496
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 3068 20942 3096 21286
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 2976 20466 3004 20810
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 2964 20460 3016 20466
rect 2964 20402 3016 20408
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 2884 20318 3004 20346
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2780 19712 2832 19718
rect 2780 19654 2832 19660
rect 2884 17746 2912 20198
rect 2976 18737 3004 20318
rect 2962 18728 3018 18737
rect 2962 18663 3018 18672
rect 3068 18057 3096 20402
rect 3160 19961 3188 20742
rect 3146 19952 3202 19961
rect 3146 19887 3202 19896
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3160 19242 3188 19654
rect 3252 19553 3280 21490
rect 3516 19780 3568 19786
rect 3516 19722 3568 19728
rect 3238 19544 3294 19553
rect 3238 19479 3294 19488
rect 3528 19378 3556 19722
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3054 18048 3110 18057
rect 3054 17983 3110 17992
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2792 17241 2820 17614
rect 3528 17610 3556 18226
rect 2872 17604 2924 17610
rect 2872 17546 2924 17552
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 2778 17232 2834 17241
rect 2778 17167 2834 17176
rect 2884 17082 2912 17546
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 2792 17054 2912 17082
rect 2792 16182 2820 17054
rect 3252 16561 3280 17138
rect 3238 16552 3294 16561
rect 3238 16487 3294 16496
rect 2780 16176 2832 16182
rect 2780 16118 2832 16124
rect 2792 15706 2820 16118
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2792 15094 2820 15642
rect 2884 15570 2912 16050
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2976 15094 3004 15846
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2964 14952 3016 14958
rect 3068 14940 3096 15506
rect 3016 14912 3096 14940
rect 2964 14894 3016 14900
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2412 14340 2464 14346
rect 2412 14282 2464 14288
rect 2424 13870 2452 14282
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2240 10266 2268 10610
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1504 9586 1532 9998
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 1412 9217 1440 9522
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 2332 8974 2360 9522
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 1412 8401 1440 8910
rect 1492 8900 1544 8906
rect 1492 8842 1544 8848
rect 1504 8498 1532 8842
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1398 8392 1454 8401
rect 1398 8327 1454 8336
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7721 1440 7822
rect 1398 7712 1454 7721
rect 1398 7647 1454 7656
rect 1504 6390 1532 8434
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1596 7478 1624 8026
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1596 6798 1624 7414
rect 1688 7410 1716 8774
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1872 6798 1900 7686
rect 2240 7546 2268 8434
rect 2332 8090 2360 8910
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2424 7954 2452 13806
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2608 13326 2636 13670
rect 2792 13569 2820 14894
rect 3160 14618 3188 15574
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3160 14006 3188 14554
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 2778 13560 2834 13569
rect 2778 13495 2834 13504
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2608 12782 2636 13262
rect 2976 12986 3004 13738
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2608 11626 2636 12718
rect 2976 12374 3004 12922
rect 3344 12850 3372 13806
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 3344 12306 3372 12786
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2792 12073 2820 12174
rect 2778 12064 2834 12073
rect 2778 11999 2834 12008
rect 2884 11830 2912 12242
rect 3528 12102 3556 12786
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2780 11688 2832 11694
rect 2700 11636 2780 11642
rect 2700 11630 2832 11636
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2700 11614 2820 11630
rect 2700 9926 2728 11614
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2884 10810 2912 11018
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2884 10130 2912 10746
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2688 9920 2740 9926
rect 2792 9897 2820 9998
rect 3332 9988 3384 9994
rect 3332 9930 3384 9936
rect 2872 9920 2924 9926
rect 2688 9862 2740 9868
rect 2778 9888 2834 9897
rect 2700 9450 2728 9862
rect 2872 9862 2924 9868
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 2778 9823 2834 9832
rect 2884 9654 2912 9862
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 3160 9586 3188 9862
rect 3344 9722 3372 9930
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2516 8974 2544 9318
rect 2608 8974 2636 9386
rect 2700 9042 2728 9386
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2608 7478 2636 8910
rect 2700 8566 2728 8978
rect 2792 8634 2820 9318
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2240 6458 2268 6734
rect 2608 6730 2636 7414
rect 2700 7342 2728 8502
rect 2792 7410 2820 8570
rect 3528 7410 3556 9522
rect 3620 9042 3648 27814
rect 5915 27772 6223 27792
rect 5915 27770 5921 27772
rect 5977 27770 6001 27772
rect 6057 27770 6081 27772
rect 6137 27770 6161 27772
rect 6217 27770 6223 27772
rect 5977 27718 5979 27770
rect 6159 27718 6161 27770
rect 5915 27716 5921 27718
rect 5977 27716 6001 27718
rect 6057 27716 6081 27718
rect 6137 27716 6161 27718
rect 6217 27716 6223 27718
rect 5915 27696 6223 27716
rect 6366 27704 6422 27713
rect 6366 27639 6422 27648
rect 5816 27600 5868 27606
rect 5816 27542 5868 27548
rect 5724 27464 5776 27470
rect 5724 27406 5776 27412
rect 4620 27396 4672 27402
rect 4620 27338 4672 27344
rect 3792 26512 3844 26518
rect 3790 26480 3792 26489
rect 3844 26480 3846 26489
rect 3790 26415 3846 26424
rect 4160 25424 4212 25430
rect 4160 25366 4212 25372
rect 4172 24818 4200 25366
rect 4160 24812 4212 24818
rect 4160 24754 4212 24760
rect 4436 24404 4488 24410
rect 4436 24346 4488 24352
rect 3792 24200 3844 24206
rect 3792 24142 3844 24148
rect 3804 23798 3832 24142
rect 4068 24132 4120 24138
rect 4068 24074 4120 24080
rect 4080 23866 4108 24074
rect 4344 24064 4396 24070
rect 4344 24006 4396 24012
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 3792 23792 3844 23798
rect 4356 23746 4384 24006
rect 3792 23734 3844 23740
rect 3804 22642 3832 23734
rect 4264 23730 4384 23746
rect 4252 23724 4384 23730
rect 4304 23718 4384 23724
rect 4252 23666 4304 23672
rect 4344 23656 4396 23662
rect 4448 23644 4476 24346
rect 4396 23616 4476 23644
rect 4344 23598 4396 23604
rect 4448 23186 4476 23616
rect 4436 23180 4488 23186
rect 4436 23122 4488 23128
rect 4160 22976 4212 22982
rect 4160 22918 4212 22924
rect 4172 22710 4200 22918
rect 4160 22704 4212 22710
rect 4160 22646 4212 22652
rect 3792 22636 3844 22642
rect 3712 22596 3792 22624
rect 3712 22030 3740 22596
rect 3792 22578 3844 22584
rect 3976 22500 4028 22506
rect 3976 22442 4028 22448
rect 3700 22024 3752 22030
rect 3700 21966 3752 21972
rect 3712 20398 3740 21966
rect 3700 20392 3752 20398
rect 3700 20334 3752 20340
rect 3712 19854 3740 20334
rect 3988 19854 4016 22442
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 4066 20224 4122 20233
rect 4172 20210 4200 20878
rect 4122 20182 4200 20210
rect 4066 20159 4122 20168
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3712 19378 3740 19790
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3712 17882 3740 18226
rect 3700 17876 3752 17882
rect 3700 17818 3752 17824
rect 3804 17746 3832 19246
rect 4264 18766 4292 22374
rect 4448 21690 4476 23122
rect 4528 22976 4580 22982
rect 4528 22918 4580 22924
rect 4540 22778 4568 22918
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 4436 21684 4488 21690
rect 4436 21626 4488 21632
rect 4436 20800 4488 20806
rect 4436 20742 4488 20748
rect 4448 20534 4476 20742
rect 4436 20528 4488 20534
rect 4436 20470 4488 20476
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 4344 20256 4396 20262
rect 4344 20198 4396 20204
rect 4356 19990 4384 20198
rect 4540 20058 4568 20402
rect 4528 20052 4580 20058
rect 4528 19994 4580 20000
rect 4344 19984 4396 19990
rect 4344 19926 4396 19932
rect 4356 18902 4384 19926
rect 4528 19780 4580 19786
rect 4528 19722 4580 19728
rect 4540 18902 4568 19722
rect 4344 18896 4396 18902
rect 4344 18838 4396 18844
rect 4528 18896 4580 18902
rect 4528 18838 4580 18844
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 3792 17740 3844 17746
rect 3792 17682 3844 17688
rect 4172 17678 4200 18566
rect 4356 18358 4384 18838
rect 4344 18352 4396 18358
rect 4344 18294 4396 18300
rect 4436 18148 4488 18154
rect 4436 18090 4488 18096
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3712 15502 3740 15914
rect 3804 15502 3832 16118
rect 3988 15502 4016 16934
rect 4080 16658 4108 17138
rect 4160 16720 4212 16726
rect 4160 16662 4212 16668
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4172 16046 4200 16662
rect 4264 16590 4292 18022
rect 4356 17746 4384 18022
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4356 15706 4384 17138
rect 4448 16114 4476 18090
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4448 15570 4476 16050
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 4068 15564 4120 15570
rect 4436 15564 4488 15570
rect 4120 15524 4200 15552
rect 4068 15506 4120 15512
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3804 14006 3832 14214
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 3804 13394 3832 13942
rect 4080 13938 4108 15302
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4172 13870 4200 15524
rect 4436 15506 4488 15512
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 4264 13938 4292 15030
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4264 13530 4292 13874
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 4264 12782 4292 13466
rect 4540 13190 4568 15982
rect 4632 14464 4660 27338
rect 5540 26988 5592 26994
rect 5540 26930 5592 26936
rect 4896 26784 4948 26790
rect 4896 26726 4948 26732
rect 4712 26240 4764 26246
rect 4712 26182 4764 26188
rect 4724 25906 4752 26182
rect 4908 25974 4936 26726
rect 5264 26376 5316 26382
rect 5264 26318 5316 26324
rect 5356 26376 5408 26382
rect 5356 26318 5408 26324
rect 5078 26072 5134 26081
rect 5078 26007 5134 26016
rect 4896 25968 4948 25974
rect 4894 25936 4896 25945
rect 4948 25936 4950 25945
rect 4712 25900 4764 25906
rect 4712 25842 4764 25848
rect 4804 25900 4856 25906
rect 5092 25906 5120 26007
rect 5276 25922 5304 26318
rect 5368 26246 5396 26318
rect 5356 26240 5408 26246
rect 5356 26182 5408 26188
rect 5552 26042 5580 26930
rect 5736 26489 5764 27406
rect 5722 26480 5778 26489
rect 5722 26415 5778 26424
rect 5540 26036 5592 26042
rect 5540 25978 5592 25984
rect 4894 25871 4950 25880
rect 5080 25900 5132 25906
rect 4804 25842 4856 25848
rect 5276 25894 5580 25922
rect 5080 25842 5132 25848
rect 4724 24410 4752 25842
rect 4816 25809 4844 25842
rect 4802 25800 4858 25809
rect 4802 25735 4858 25744
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 5092 24313 5120 25842
rect 5552 25786 5580 25894
rect 5552 25758 5672 25786
rect 5736 25770 5764 26415
rect 5828 26330 5856 27542
rect 6380 27470 6408 27639
rect 6368 27464 6420 27470
rect 6368 27406 6420 27412
rect 6000 27396 6052 27402
rect 6000 27338 6052 27344
rect 6012 26874 6040 27338
rect 6012 26846 6408 26874
rect 5915 26684 6223 26704
rect 5915 26682 5921 26684
rect 5977 26682 6001 26684
rect 6057 26682 6081 26684
rect 6137 26682 6161 26684
rect 6217 26682 6223 26684
rect 5977 26630 5979 26682
rect 6159 26630 6161 26682
rect 5915 26628 5921 26630
rect 5977 26628 6001 26630
rect 6057 26628 6081 26630
rect 6137 26628 6161 26630
rect 6217 26628 6223 26630
rect 5915 26608 6223 26628
rect 5906 26480 5962 26489
rect 5906 26415 5908 26424
rect 5960 26415 5962 26424
rect 5908 26386 5960 26392
rect 6092 26376 6144 26382
rect 5828 26302 6040 26330
rect 6092 26318 6144 26324
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 5816 26240 5868 26246
rect 5816 26182 5868 26188
rect 5828 25906 5856 26182
rect 6012 25922 6040 26302
rect 6104 26081 6132 26318
rect 6090 26072 6146 26081
rect 6288 26042 6316 26318
rect 6090 26007 6146 26016
rect 6276 26036 6328 26042
rect 6276 25978 6328 25984
rect 5816 25900 5868 25906
rect 5816 25842 5868 25848
rect 5908 25900 5960 25906
rect 6012 25894 6316 25922
rect 5908 25842 5960 25848
rect 5920 25786 5948 25842
rect 5644 25158 5672 25758
rect 5724 25764 5776 25770
rect 5724 25706 5776 25712
rect 5828 25758 5948 25786
rect 5632 25152 5684 25158
rect 5632 25094 5684 25100
rect 5540 24812 5592 24818
rect 5644 24800 5672 25094
rect 5828 24857 5856 25758
rect 6288 25702 6316 25894
rect 6276 25696 6328 25702
rect 6276 25638 6328 25644
rect 5915 25596 6223 25616
rect 5915 25594 5921 25596
rect 5977 25594 6001 25596
rect 6057 25594 6081 25596
rect 6137 25594 6161 25596
rect 6217 25594 6223 25596
rect 5977 25542 5979 25594
rect 6159 25542 6161 25594
rect 5915 25540 5921 25542
rect 5977 25540 6001 25542
rect 6057 25540 6081 25542
rect 6137 25540 6161 25542
rect 6217 25540 6223 25542
rect 5915 25520 6223 25540
rect 6288 25294 6316 25638
rect 6276 25288 6328 25294
rect 6276 25230 6328 25236
rect 5814 24848 5870 24857
rect 5724 24812 5776 24818
rect 5644 24772 5724 24800
rect 5540 24754 5592 24760
rect 5814 24783 5870 24792
rect 5724 24754 5776 24760
rect 5552 24410 5580 24754
rect 5540 24404 5592 24410
rect 5540 24346 5592 24352
rect 5078 24304 5134 24313
rect 5078 24239 5134 24248
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 4816 23186 4844 23462
rect 4804 23180 4856 23186
rect 4804 23122 4856 23128
rect 4816 22098 4844 23122
rect 4908 23118 4936 23666
rect 5092 23526 5120 24239
rect 5172 24200 5224 24206
rect 5172 24142 5224 24148
rect 5080 23520 5132 23526
rect 5080 23462 5132 23468
rect 4896 23112 4948 23118
rect 4896 23054 4948 23060
rect 4804 22092 4856 22098
rect 4804 22034 4856 22040
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 5092 19854 5120 20198
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4816 18970 4844 19314
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4724 16114 4752 16934
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4816 15502 4844 16934
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4908 15314 4936 18226
rect 4816 15286 4936 15314
rect 4632 14436 4752 14464
rect 4620 14340 4672 14346
rect 4620 14282 4672 14288
rect 4632 14074 4660 14282
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4724 13530 4752 14436
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4080 12170 4108 12582
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 4540 12102 4568 12786
rect 4632 12238 4660 12922
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4632 11830 4660 12174
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4252 9580 4304 9586
rect 4304 9540 4384 9568
rect 4252 9522 4304 9528
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3896 8498 3924 8842
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 3528 6798 3556 7346
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 1492 6384 1544 6390
rect 1492 6326 1544 6332
rect 1504 5778 1532 6326
rect 2424 6322 2452 6598
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2778 6216 2834 6225
rect 2778 6151 2834 6160
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2700 5370 2728 5578
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1412 4729 1440 5102
rect 1398 4720 1454 4729
rect 1398 4655 1454 4664
rect 2792 4622 2820 6151
rect 3068 5302 3096 6598
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3252 5914 3280 6054
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3252 5370 3280 5850
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 3528 5234 3556 6734
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 3712 4214 3740 8230
rect 3804 7886 3832 8434
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 4172 7002 4200 7754
rect 4264 7478 4292 9386
rect 4356 8906 4384 9540
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 3974 6896 4030 6905
rect 3804 5166 3832 6870
rect 3974 6831 4030 6840
rect 4068 6860 4120 6866
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3896 4826 3924 6734
rect 3988 6644 4016 6831
rect 4264 6848 4292 7414
rect 4356 7410 4384 7822
rect 4448 7818 4476 9658
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 8498 4660 9318
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4724 7562 4752 13262
rect 4816 13258 4844 15286
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4816 12434 4844 13194
rect 5000 13138 5028 18634
rect 5184 14906 5212 24142
rect 5736 23050 5764 24754
rect 5828 24614 5856 24783
rect 5816 24608 5868 24614
rect 5816 24550 5868 24556
rect 5828 24206 5856 24550
rect 5915 24508 6223 24528
rect 5915 24506 5921 24508
rect 5977 24506 6001 24508
rect 6057 24506 6081 24508
rect 6137 24506 6161 24508
rect 6217 24506 6223 24508
rect 5977 24454 5979 24506
rect 6159 24454 6161 24506
rect 5915 24452 5921 24454
rect 5977 24452 6001 24454
rect 6057 24452 6081 24454
rect 6137 24452 6161 24454
rect 6217 24452 6223 24454
rect 5915 24432 6223 24452
rect 6092 24336 6144 24342
rect 6092 24278 6144 24284
rect 6182 24304 6238 24313
rect 6104 24206 6132 24278
rect 6182 24239 6184 24248
rect 6236 24239 6238 24248
rect 6184 24210 6236 24216
rect 5816 24200 5868 24206
rect 5816 24142 5868 24148
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 6288 24070 6316 25230
rect 6276 24064 6328 24070
rect 6276 24006 6328 24012
rect 6288 23798 6316 24006
rect 6276 23792 6328 23798
rect 6276 23734 6328 23740
rect 6380 23730 6408 26846
rect 6368 23724 6420 23730
rect 6368 23666 6420 23672
rect 5915 23420 6223 23440
rect 5915 23418 5921 23420
rect 5977 23418 6001 23420
rect 6057 23418 6081 23420
rect 6137 23418 6161 23420
rect 6217 23418 6223 23420
rect 5977 23366 5979 23418
rect 6159 23366 6161 23418
rect 5915 23364 5921 23366
rect 5977 23364 6001 23366
rect 6057 23364 6081 23366
rect 6137 23364 6161 23366
rect 6217 23364 6223 23366
rect 5915 23344 6223 23364
rect 5632 23044 5684 23050
rect 5632 22986 5684 22992
rect 5724 23044 5776 23050
rect 5724 22986 5776 22992
rect 5540 22976 5592 22982
rect 5540 22918 5592 22924
rect 5552 22094 5580 22918
rect 5644 22778 5672 22986
rect 5632 22772 5684 22778
rect 5632 22714 5684 22720
rect 5736 22098 5764 22986
rect 6276 22704 6328 22710
rect 6380 22692 6408 23666
rect 6328 22664 6408 22692
rect 6276 22646 6328 22652
rect 6368 22568 6420 22574
rect 6368 22510 6420 22516
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5552 22066 5672 22094
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5552 21554 5580 21966
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5552 20602 5580 21490
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 5644 19854 5672 22066
rect 5724 22092 5776 22098
rect 5724 22034 5776 22040
rect 5828 21554 5856 22374
rect 5915 22332 6223 22352
rect 5915 22330 5921 22332
rect 5977 22330 6001 22332
rect 6057 22330 6081 22332
rect 6137 22330 6161 22332
rect 6217 22330 6223 22332
rect 5977 22278 5979 22330
rect 6159 22278 6161 22330
rect 5915 22276 5921 22278
rect 5977 22276 6001 22278
rect 6057 22276 6081 22278
rect 6137 22276 6161 22278
rect 6217 22276 6223 22278
rect 5915 22256 6223 22276
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 6276 21548 6328 21554
rect 6276 21490 6328 21496
rect 5632 19848 5684 19854
rect 5828 19825 5856 21490
rect 5915 21244 6223 21264
rect 5915 21242 5921 21244
rect 5977 21242 6001 21244
rect 6057 21242 6081 21244
rect 6137 21242 6161 21244
rect 6217 21242 6223 21244
rect 5977 21190 5979 21242
rect 6159 21190 6161 21242
rect 5915 21188 5921 21190
rect 5977 21188 6001 21190
rect 6057 21188 6081 21190
rect 6137 21188 6161 21190
rect 6217 21188 6223 21190
rect 5915 21168 6223 21188
rect 6184 21072 6236 21078
rect 6288 21060 6316 21490
rect 6236 21032 6316 21060
rect 6184 21014 6236 21020
rect 6380 21010 6408 22510
rect 6472 21350 6500 28494
rect 6564 27130 6592 29514
rect 6552 27124 6604 27130
rect 6552 27066 6604 27072
rect 6564 25226 6592 27066
rect 6552 25220 6604 25226
rect 6552 25162 6604 25168
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6564 23866 6592 24142
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 6552 23248 6604 23254
rect 6552 23190 6604 23196
rect 6564 22642 6592 23190
rect 6552 22636 6604 22642
rect 6552 22578 6604 22584
rect 6552 22500 6604 22506
rect 6552 22442 6604 22448
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6564 21146 6592 22442
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6380 20534 6408 20946
rect 6368 20528 6420 20534
rect 6368 20470 6420 20476
rect 6380 20346 6408 20470
rect 6564 20466 6592 21082
rect 6656 20584 6684 32234
rect 6736 32224 6788 32230
rect 6736 32166 6788 32172
rect 6748 31346 6776 32166
rect 6840 31822 6868 32710
rect 7116 32502 7144 33254
rect 7104 32496 7156 32502
rect 7104 32438 7156 32444
rect 6828 31816 6880 31822
rect 6828 31758 6880 31764
rect 7104 31680 7156 31686
rect 7104 31622 7156 31628
rect 7116 31346 7144 31622
rect 7300 31346 7328 34478
rect 7392 34406 7420 38286
rect 7484 38010 7512 41414
rect 7576 41206 7604 44338
rect 7760 43994 7788 44338
rect 7840 44328 7892 44334
rect 7840 44270 7892 44276
rect 7748 43988 7800 43994
rect 7748 43930 7800 43936
rect 7852 43772 7880 44270
rect 8312 44198 8340 44338
rect 8300 44192 8352 44198
rect 8300 44134 8352 44140
rect 7932 43784 7984 43790
rect 7852 43744 7932 43772
rect 7748 43716 7800 43722
rect 7748 43658 7800 43664
rect 7760 42702 7788 43658
rect 7852 42838 7880 43744
rect 7932 43726 7984 43732
rect 7840 42832 7892 42838
rect 7840 42774 7892 42780
rect 7656 42696 7708 42702
rect 7656 42638 7708 42644
rect 7748 42696 7800 42702
rect 7748 42638 7800 42644
rect 7668 41750 7696 42638
rect 7748 42356 7800 42362
rect 7748 42298 7800 42304
rect 7656 41744 7708 41750
rect 7656 41686 7708 41692
rect 7760 41614 7788 42298
rect 7748 41608 7800 41614
rect 7748 41550 7800 41556
rect 7564 41200 7616 41206
rect 7564 41142 7616 41148
rect 7760 40594 7788 41550
rect 7852 41546 7880 42774
rect 8024 42696 8076 42702
rect 8024 42638 8076 42644
rect 7932 42560 7984 42566
rect 7932 42502 7984 42508
rect 7944 42362 7972 42502
rect 7932 42356 7984 42362
rect 7932 42298 7984 42304
rect 7944 41614 7972 42298
rect 7932 41608 7984 41614
rect 7932 41550 7984 41556
rect 7840 41540 7892 41546
rect 7840 41482 7892 41488
rect 7852 41138 7880 41482
rect 7840 41132 7892 41138
rect 7840 41074 7892 41080
rect 7932 41064 7984 41070
rect 7932 41006 7984 41012
rect 7748 40588 7800 40594
rect 7748 40530 7800 40536
rect 7944 40186 7972 41006
rect 7932 40180 7984 40186
rect 7932 40122 7984 40128
rect 8036 40118 8064 42638
rect 8116 42220 8168 42226
rect 8116 42162 8168 42168
rect 8128 41818 8156 42162
rect 8312 42158 8340 44134
rect 8404 42566 8432 44814
rect 8944 44736 8996 44742
rect 8944 44678 8996 44684
rect 29000 44736 29052 44742
rect 29000 44678 29052 44684
rect 8760 44532 8812 44538
rect 8760 44474 8812 44480
rect 8772 44198 8800 44474
rect 8852 44260 8904 44266
rect 8852 44202 8904 44208
rect 8760 44192 8812 44198
rect 8760 44134 8812 44140
rect 8864 43450 8892 44202
rect 8956 43858 8984 44678
rect 10880 44636 11188 44656
rect 10880 44634 10886 44636
rect 10942 44634 10966 44636
rect 11022 44634 11046 44636
rect 11102 44634 11126 44636
rect 11182 44634 11188 44636
rect 10942 44582 10944 44634
rect 11124 44582 11126 44634
rect 10880 44580 10886 44582
rect 10942 44580 10966 44582
rect 11022 44580 11046 44582
rect 11102 44580 11126 44582
rect 11182 44580 11188 44582
rect 10880 44560 11188 44580
rect 20811 44636 21119 44656
rect 20811 44634 20817 44636
rect 20873 44634 20897 44636
rect 20953 44634 20977 44636
rect 21033 44634 21057 44636
rect 21113 44634 21119 44636
rect 20873 44582 20875 44634
rect 21055 44582 21057 44634
rect 20811 44580 20817 44582
rect 20873 44580 20897 44582
rect 20953 44580 20977 44582
rect 21033 44580 21057 44582
rect 21113 44580 21119 44582
rect 20811 44560 21119 44580
rect 10508 44532 10560 44538
rect 10508 44474 10560 44480
rect 18144 44532 18196 44538
rect 18144 44474 18196 44480
rect 9128 44396 9180 44402
rect 9128 44338 9180 44344
rect 8944 43852 8996 43858
rect 8944 43794 8996 43800
rect 8852 43444 8904 43450
rect 8852 43386 8904 43392
rect 9140 42566 9168 44338
rect 9956 44260 10008 44266
rect 9956 44202 10008 44208
rect 9968 43382 9996 44202
rect 10232 44192 10284 44198
rect 10232 44134 10284 44140
rect 9956 43376 10008 43382
rect 9956 43318 10008 43324
rect 10244 43314 10272 44134
rect 10232 43308 10284 43314
rect 10232 43250 10284 43256
rect 10324 42628 10376 42634
rect 10324 42570 10376 42576
rect 8392 42560 8444 42566
rect 8392 42502 8444 42508
rect 9128 42560 9180 42566
rect 9128 42502 9180 42508
rect 8300 42152 8352 42158
rect 8300 42094 8352 42100
rect 9312 42152 9364 42158
rect 9312 42094 9364 42100
rect 9324 41818 9352 42094
rect 8116 41812 8168 41818
rect 8116 41754 8168 41760
rect 9312 41812 9364 41818
rect 9312 41754 9364 41760
rect 10232 41744 10284 41750
rect 10232 41686 10284 41692
rect 10140 41540 10192 41546
rect 10140 41482 10192 41488
rect 8576 40520 8628 40526
rect 8576 40462 8628 40468
rect 9772 40520 9824 40526
rect 9772 40462 9824 40468
rect 8588 40186 8616 40462
rect 8944 40384 8996 40390
rect 8944 40326 8996 40332
rect 9128 40384 9180 40390
rect 9128 40326 9180 40332
rect 8576 40180 8628 40186
rect 8576 40122 8628 40128
rect 8024 40112 8076 40118
rect 8024 40054 8076 40060
rect 8036 39642 8064 40054
rect 8024 39636 8076 39642
rect 8024 39578 8076 39584
rect 7656 38344 7708 38350
rect 7656 38286 7708 38292
rect 7472 38004 7524 38010
rect 7472 37946 7524 37952
rect 7668 36650 7696 38286
rect 8036 37874 8064 39578
rect 8852 39568 8904 39574
rect 8852 39510 8904 39516
rect 8760 38412 8812 38418
rect 8760 38354 8812 38360
rect 8668 38276 8720 38282
rect 8668 38218 8720 38224
rect 8680 37874 8708 38218
rect 8024 37868 8076 37874
rect 8024 37810 8076 37816
rect 8300 37868 8352 37874
rect 8300 37810 8352 37816
rect 8668 37868 8720 37874
rect 8668 37810 8720 37816
rect 8312 36786 8340 37810
rect 8772 37806 8800 38354
rect 8864 38214 8892 39510
rect 8956 38842 8984 40326
rect 9140 38962 9168 40326
rect 9680 39840 9732 39846
rect 9680 39782 9732 39788
rect 9692 39642 9720 39782
rect 9680 39636 9732 39642
rect 9680 39578 9732 39584
rect 9680 39364 9732 39370
rect 9680 39306 9732 39312
rect 9128 38956 9180 38962
rect 9128 38898 9180 38904
rect 9496 38956 9548 38962
rect 9496 38898 9548 38904
rect 8956 38814 9444 38842
rect 8956 38332 8984 38814
rect 9220 38752 9272 38758
rect 9220 38694 9272 38700
rect 9036 38344 9088 38350
rect 8956 38304 9036 38332
rect 9036 38286 9088 38292
rect 8852 38208 8904 38214
rect 8852 38150 8904 38156
rect 8864 37874 8892 38150
rect 9232 37874 9260 38694
rect 9416 38554 9444 38814
rect 9312 38548 9364 38554
rect 9312 38490 9364 38496
rect 9404 38548 9456 38554
rect 9404 38490 9456 38496
rect 9324 38350 9352 38490
rect 9312 38344 9364 38350
rect 9312 38286 9364 38292
rect 8852 37868 8904 37874
rect 9220 37868 9272 37874
rect 8904 37828 8984 37856
rect 8852 37810 8904 37816
rect 8484 37800 8536 37806
rect 8484 37742 8536 37748
rect 8760 37800 8812 37806
rect 8760 37742 8812 37748
rect 8300 36780 8352 36786
rect 8300 36722 8352 36728
rect 8392 36780 8444 36786
rect 8392 36722 8444 36728
rect 8404 36650 8432 36722
rect 8496 36718 8524 37742
rect 8576 37120 8628 37126
rect 8576 37062 8628 37068
rect 8760 37120 8812 37126
rect 8760 37062 8812 37068
rect 8484 36712 8536 36718
rect 8484 36654 8536 36660
rect 7656 36644 7708 36650
rect 7656 36586 7708 36592
rect 8392 36644 8444 36650
rect 8392 36586 8444 36592
rect 8024 36168 8076 36174
rect 8404 36122 8432 36586
rect 8024 36110 8076 36116
rect 7472 36032 7524 36038
rect 7472 35974 7524 35980
rect 7380 34400 7432 34406
rect 7380 34342 7432 34348
rect 6736 31340 6788 31346
rect 6736 31282 6788 31288
rect 7104 31340 7156 31346
rect 7104 31282 7156 31288
rect 7288 31340 7340 31346
rect 7288 31282 7340 31288
rect 6748 30190 6776 31282
rect 6828 31272 6880 31278
rect 6828 31214 6880 31220
rect 6840 30258 6868 31214
rect 6920 31204 6972 31210
rect 6920 31146 6972 31152
rect 6828 30252 6880 30258
rect 6828 30194 6880 30200
rect 6736 30184 6788 30190
rect 6736 30126 6788 30132
rect 6932 29510 6960 31146
rect 7116 30258 7144 31282
rect 7104 30252 7156 30258
rect 7104 30194 7156 30200
rect 7288 30048 7340 30054
rect 7288 29990 7340 29996
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 6828 29028 6880 29034
rect 6828 28970 6880 28976
rect 6734 27704 6790 27713
rect 6734 27639 6790 27648
rect 6748 25945 6776 27639
rect 6840 27334 6868 28970
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6828 26920 6880 26926
rect 6932 26908 6960 29446
rect 7012 28960 7064 28966
rect 7012 28902 7064 28908
rect 7024 28422 7052 28902
rect 7012 28416 7064 28422
rect 7012 28358 7064 28364
rect 7104 28416 7156 28422
rect 7104 28358 7156 28364
rect 7116 28218 7144 28358
rect 7104 28212 7156 28218
rect 7104 28154 7156 28160
rect 7196 27872 7248 27878
rect 7196 27814 7248 27820
rect 7104 27328 7156 27334
rect 7104 27270 7156 27276
rect 7116 26994 7144 27270
rect 7012 26988 7064 26994
rect 7012 26930 7064 26936
rect 7104 26988 7156 26994
rect 7104 26930 7156 26936
rect 6880 26880 6960 26908
rect 6828 26862 6880 26868
rect 6840 26042 6868 26862
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 7024 25974 7052 26930
rect 7012 25968 7064 25974
rect 6734 25936 6790 25945
rect 7012 25910 7064 25916
rect 6734 25871 6736 25880
rect 6788 25871 6790 25880
rect 6736 25842 6788 25848
rect 6748 25811 6776 25842
rect 6736 24268 6788 24274
rect 6736 24210 6788 24216
rect 6748 23866 6776 24210
rect 6736 23860 6788 23866
rect 6736 23802 6788 23808
rect 6748 23338 6776 23802
rect 7024 23798 7052 25910
rect 7208 25106 7236 27814
rect 7300 25226 7328 29990
rect 7484 29646 7512 35974
rect 8036 35834 8064 36110
rect 8128 36094 8432 36122
rect 8024 35828 8076 35834
rect 8024 35770 8076 35776
rect 7564 35692 7616 35698
rect 7564 35634 7616 35640
rect 7576 34202 7604 35634
rect 7656 35012 7708 35018
rect 7656 34954 7708 34960
rect 7668 34746 7696 34954
rect 7656 34740 7708 34746
rect 7656 34682 7708 34688
rect 8024 34536 8076 34542
rect 8128 34524 8156 36094
rect 8392 36032 8444 36038
rect 8392 35974 8444 35980
rect 8404 35154 8432 35974
rect 8392 35148 8444 35154
rect 8392 35090 8444 35096
rect 8208 34604 8260 34610
rect 8208 34546 8260 34552
rect 8076 34496 8156 34524
rect 8024 34478 8076 34484
rect 7564 34196 7616 34202
rect 7564 34138 7616 34144
rect 7656 34196 7708 34202
rect 7656 34138 7708 34144
rect 7576 33590 7604 34138
rect 7668 33998 7696 34138
rect 7656 33992 7708 33998
rect 7656 33934 7708 33940
rect 7668 33658 7696 33934
rect 7656 33652 7708 33658
rect 7656 33594 7708 33600
rect 7840 33652 7892 33658
rect 7840 33594 7892 33600
rect 7564 33584 7616 33590
rect 7564 33526 7616 33532
rect 7576 32910 7604 33526
rect 7852 33522 7880 33594
rect 7748 33516 7800 33522
rect 7748 33458 7800 33464
rect 7840 33516 7892 33522
rect 7840 33458 7892 33464
rect 7564 32904 7616 32910
rect 7564 32846 7616 32852
rect 7576 31822 7604 32846
rect 7760 32570 7788 33458
rect 7748 32564 7800 32570
rect 7748 32506 7800 32512
rect 7564 31816 7616 31822
rect 7564 31758 7616 31764
rect 7852 31414 7880 33458
rect 7932 33108 7984 33114
rect 7932 33050 7984 33056
rect 7944 32978 7972 33050
rect 7932 32972 7984 32978
rect 7932 32914 7984 32920
rect 7840 31408 7892 31414
rect 7840 31350 7892 31356
rect 7564 31136 7616 31142
rect 7564 31078 7616 31084
rect 7472 29640 7524 29646
rect 7472 29582 7524 29588
rect 7380 29096 7432 29102
rect 7380 29038 7432 29044
rect 7392 28762 7420 29038
rect 7380 28756 7432 28762
rect 7380 28698 7432 28704
rect 7472 27600 7524 27606
rect 7472 27542 7524 27548
rect 7380 27464 7432 27470
rect 7380 27406 7432 27412
rect 7392 25906 7420 27406
rect 7484 27169 7512 27542
rect 7470 27160 7526 27169
rect 7470 27095 7526 27104
rect 7484 27062 7512 27095
rect 7472 27056 7524 27062
rect 7472 26998 7524 27004
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 7484 26450 7512 26726
rect 7472 26444 7524 26450
rect 7472 26386 7524 26392
rect 7380 25900 7432 25906
rect 7380 25842 7432 25848
rect 7472 25356 7524 25362
rect 7472 25298 7524 25304
rect 7288 25220 7340 25226
rect 7288 25162 7340 25168
rect 7380 25152 7432 25158
rect 7208 25078 7328 25106
rect 7380 25094 7432 25100
rect 7104 24812 7156 24818
rect 7104 24754 7156 24760
rect 7116 24410 7144 24754
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 7104 24404 7156 24410
rect 7104 24346 7156 24352
rect 7208 24138 7236 24686
rect 7196 24132 7248 24138
rect 7196 24074 7248 24080
rect 6920 23792 6972 23798
rect 6920 23734 6972 23740
rect 7012 23792 7064 23798
rect 7012 23734 7064 23740
rect 6748 23310 6868 23338
rect 6736 21956 6788 21962
rect 6736 21898 6788 21904
rect 6748 21146 6776 21898
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6840 20874 6868 23310
rect 6932 22624 6960 23734
rect 7104 23588 7156 23594
rect 7104 23530 7156 23536
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 7024 22982 7052 23462
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 7116 22778 7144 23530
rect 7196 23520 7248 23526
rect 7196 23462 7248 23468
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7012 22636 7064 22642
rect 6932 22596 7012 22624
rect 6932 21554 6960 22596
rect 7012 22578 7064 22584
rect 7208 22030 7236 23462
rect 7196 22024 7248 22030
rect 7196 21966 7248 21972
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 7024 20942 7052 21830
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 6828 20868 6880 20874
rect 6828 20810 6880 20816
rect 6656 20556 6960 20584
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6380 20318 6500 20346
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 5915 20156 6223 20176
rect 5915 20154 5921 20156
rect 5977 20154 6001 20156
rect 6057 20154 6081 20156
rect 6137 20154 6161 20156
rect 6217 20154 6223 20156
rect 5977 20102 5979 20154
rect 6159 20102 6161 20154
rect 5915 20100 5921 20102
rect 5977 20100 6001 20102
rect 6057 20100 6081 20102
rect 6137 20100 6161 20102
rect 6217 20100 6223 20102
rect 5915 20080 6223 20100
rect 6276 19848 6328 19854
rect 5632 19790 5684 19796
rect 5814 19816 5870 19825
rect 6276 19790 6328 19796
rect 5814 19751 5870 19760
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5276 18766 5304 19654
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5644 18834 5672 19110
rect 5828 18970 5856 19751
rect 5915 19068 6223 19088
rect 5915 19066 5921 19068
rect 5977 19066 6001 19068
rect 6057 19066 6081 19068
rect 6137 19066 6161 19068
rect 6217 19066 6223 19068
rect 5977 19014 5979 19066
rect 6159 19014 6161 19066
rect 5915 19012 5921 19014
rect 5977 19012 6001 19014
rect 6057 19012 6081 19014
rect 6137 19012 6161 19014
rect 6217 19012 6223 19014
rect 5915 18992 6223 19012
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5460 16998 5488 18294
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5264 15428 5316 15434
rect 5264 15370 5316 15376
rect 5276 15162 5304 15370
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5092 14878 5212 14906
rect 5092 13326 5120 14878
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 14482 5212 14758
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5000 13110 5120 13138
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 4816 12406 4936 12434
rect 4908 11286 4936 12406
rect 5000 11898 5028 12854
rect 5092 11898 5120 13110
rect 5184 12986 5212 14418
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 4908 10826 4936 11222
rect 5184 11150 5212 12718
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 4908 10798 5120 10826
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4816 8634 4844 9522
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4448 7534 4752 7562
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4120 6820 4292 6848
rect 4068 6802 4120 6808
rect 3988 6616 4200 6644
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3988 5778 4016 6258
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4172 5370 4200 6616
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4264 5234 4292 6820
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4356 6458 4384 6734
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 1860 4208 1912 4214
rect 1860 4150 1912 4156
rect 3700 4208 3752 4214
rect 3700 4150 3752 4156
rect 1136 2746 1348 2774
rect 388 2372 440 2378
rect 388 2314 440 2320
rect 400 800 428 2314
rect 1136 800 1164 2746
rect 1872 2553 1900 4150
rect 3988 4146 4016 5170
rect 4172 5030 4200 5170
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4080 4826 4108 4966
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4172 4690 4200 4966
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4264 4282 4292 5170
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 2596 4072 2648 4078
rect 2792 4049 2820 4082
rect 2596 4014 2648 4020
rect 2778 4040 2834 4049
rect 1858 2544 1914 2553
rect 1858 2479 1914 2488
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1872 800 1900 2382
rect 2608 800 2636 4014
rect 2778 3975 2834 3984
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 2780 3460 2832 3466
rect 2780 3402 2832 3408
rect 2792 3233 2820 3402
rect 2778 3224 2834 3233
rect 2778 3159 2834 3168
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2792 1737 2820 2994
rect 2778 1728 2834 1737
rect 2778 1663 2834 1672
rect 386 0 442 800
rect 1122 0 1178 800
rect 1858 0 1914 800
rect 2594 0 2650 800
rect 2884 377 2912 3062
rect 2976 1057 3004 3470
rect 2962 1048 3018 1057
rect 2962 983 3018 992
rect 3436 800 3464 3470
rect 4448 2650 4476 7534
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 6390 4568 6598
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4724 5370 4752 5578
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4540 4282 4568 4490
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4540 4078 4568 4218
rect 4908 4146 4936 10610
rect 5000 9926 5028 10678
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 5092 9518 5120 10798
rect 5184 10742 5212 11086
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 5276 10538 5304 14962
rect 5368 11218 5396 15438
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5552 14414 5580 15030
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5460 13138 5488 13466
rect 5644 13394 5672 17478
rect 5736 16454 5764 18362
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5460 13110 5672 13138
rect 5644 12986 5672 13110
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5460 11830 5488 12038
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5552 11234 5580 12922
rect 5736 12306 5764 15846
rect 5828 14414 5856 18566
rect 5915 17980 6223 18000
rect 5915 17978 5921 17980
rect 5977 17978 6001 17980
rect 6057 17978 6081 17980
rect 6137 17978 6161 17980
rect 6217 17978 6223 17980
rect 5977 17926 5979 17978
rect 6159 17926 6161 17978
rect 5915 17924 5921 17926
rect 5977 17924 6001 17926
rect 6057 17924 6081 17926
rect 6137 17924 6161 17926
rect 6217 17924 6223 17926
rect 5915 17904 6223 17924
rect 6288 17814 6316 19790
rect 6276 17808 6328 17814
rect 6276 17750 6328 17756
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 6288 17202 6316 17614
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 5915 16892 6223 16912
rect 5915 16890 5921 16892
rect 5977 16890 6001 16892
rect 6057 16890 6081 16892
rect 6137 16890 6161 16892
rect 6217 16890 6223 16892
rect 5977 16838 5979 16890
rect 6159 16838 6161 16890
rect 5915 16836 5921 16838
rect 5977 16836 6001 16838
rect 6057 16836 6081 16838
rect 6137 16836 6161 16838
rect 6217 16836 6223 16838
rect 5915 16816 6223 16836
rect 6288 16794 6316 17138
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 6288 16017 6316 16050
rect 6274 16008 6330 16017
rect 6274 15943 6330 15952
rect 5915 15804 6223 15824
rect 5915 15802 5921 15804
rect 5977 15802 6001 15804
rect 6057 15802 6081 15804
rect 6137 15802 6161 15804
rect 6217 15802 6223 15804
rect 5977 15750 5979 15802
rect 6159 15750 6161 15802
rect 5915 15748 5921 15750
rect 5977 15748 6001 15750
rect 6057 15748 6081 15750
rect 6137 15748 6161 15750
rect 6217 15748 6223 15750
rect 5915 15728 6223 15748
rect 5908 15632 5960 15638
rect 5908 15574 5960 15580
rect 5920 14890 5948 15574
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6104 15162 6132 15438
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 5908 14884 5960 14890
rect 5908 14826 5960 14832
rect 5915 14716 6223 14736
rect 5915 14714 5921 14716
rect 5977 14714 6001 14716
rect 6057 14714 6081 14716
rect 6137 14714 6161 14716
rect 6217 14714 6223 14716
rect 5977 14662 5979 14714
rect 6159 14662 6161 14714
rect 5915 14660 5921 14662
rect 5977 14660 6001 14662
rect 6057 14660 6081 14662
rect 6137 14660 6161 14662
rect 6217 14660 6223 14662
rect 5915 14640 6223 14660
rect 6092 14544 6144 14550
rect 6092 14486 6144 14492
rect 6104 14414 6132 14486
rect 6288 14414 6316 15302
rect 6380 15008 6408 20198
rect 6472 20058 6500 20318
rect 6460 20052 6512 20058
rect 6460 19994 6512 20000
rect 6472 19836 6500 19994
rect 6564 19990 6592 20402
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6552 19984 6604 19990
rect 6552 19926 6604 19932
rect 6552 19848 6604 19854
rect 6472 19808 6552 19836
rect 6552 19790 6604 19796
rect 6552 19236 6604 19242
rect 6552 19178 6604 19184
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6472 18290 6500 19110
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6472 15502 6500 18022
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6460 15020 6512 15026
rect 6380 14980 6460 15008
rect 6460 14962 6512 14968
rect 6368 14884 6420 14890
rect 6368 14826 6420 14832
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 6092 14408 6144 14414
rect 6276 14408 6328 14414
rect 6092 14350 6144 14356
rect 6182 14376 6238 14385
rect 6276 14350 6328 14356
rect 6182 14311 6238 14320
rect 6196 14278 6224 14311
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6276 14272 6328 14278
rect 6380 14260 6408 14826
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 14618 6500 14758
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6328 14232 6408 14260
rect 6276 14214 6328 14220
rect 5915 13628 6223 13648
rect 5915 13626 5921 13628
rect 5977 13626 6001 13628
rect 6057 13626 6081 13628
rect 6137 13626 6161 13628
rect 6217 13626 6223 13628
rect 5977 13574 5979 13626
rect 6159 13574 6161 13626
rect 5915 13572 5921 13574
rect 5977 13572 6001 13574
rect 6057 13572 6081 13574
rect 6137 13572 6161 13574
rect 6217 13572 6223 13574
rect 5915 13552 6223 13572
rect 6288 13410 6316 14214
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6104 13382 6316 13410
rect 5908 13252 5960 13258
rect 5908 13194 5960 13200
rect 5920 12714 5948 13194
rect 6104 13190 6132 13382
rect 6380 13326 6408 13806
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6104 12850 6132 13126
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 5816 12708 5868 12714
rect 5816 12650 5868 12656
rect 5908 12708 5960 12714
rect 5908 12650 5960 12656
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5736 11354 5764 12106
rect 5828 11762 5856 12650
rect 5915 12540 6223 12560
rect 5915 12538 5921 12540
rect 5977 12538 6001 12540
rect 6057 12538 6081 12540
rect 6137 12538 6161 12540
rect 6217 12538 6223 12540
rect 5977 12486 5979 12538
rect 6159 12486 6161 12538
rect 5915 12484 5921 12486
rect 5977 12484 6001 12486
rect 6057 12484 6081 12486
rect 6137 12484 6161 12486
rect 6217 12484 6223 12486
rect 5915 12464 6223 12484
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5356 11212 5408 11218
rect 5552 11206 5764 11234
rect 5356 11154 5408 11160
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 8906 5028 9318
rect 5276 9178 5304 9862
rect 5368 9586 5396 11018
rect 5448 10668 5500 10674
rect 5552 10656 5580 11086
rect 5500 10628 5580 10656
rect 5448 10610 5500 10616
rect 5736 10248 5764 11206
rect 5828 10742 5856 11698
rect 6196 11642 6224 12310
rect 6288 12306 6316 13126
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6380 12170 6408 12786
rect 6472 12322 6500 14418
rect 6564 12442 6592 19178
rect 6656 18329 6684 20334
rect 6748 19514 6776 20402
rect 6840 20330 6868 20402
rect 6828 20324 6880 20330
rect 6828 20266 6880 20272
rect 6932 19938 6960 20556
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 6840 19910 6960 19938
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6840 19242 6868 19910
rect 6920 19848 6972 19854
rect 6918 19816 6920 19825
rect 6972 19816 6974 19825
rect 6918 19751 6974 19760
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6828 19236 6880 19242
rect 6828 19178 6880 19184
rect 6932 18698 6960 19314
rect 7024 18698 7052 19654
rect 7116 19378 7144 20198
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 6642 18320 6698 18329
rect 6642 18255 6698 18264
rect 6736 18080 6788 18086
rect 6642 18048 6698 18057
rect 6736 18022 6788 18028
rect 6642 17983 6698 17992
rect 6656 16998 6684 17983
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6656 16590 6684 16934
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6656 15910 6684 15982
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6656 15706 6684 15846
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6748 15638 6776 18022
rect 7208 17270 7236 21490
rect 7300 21026 7328 25078
rect 7392 24954 7420 25094
rect 7380 24948 7432 24954
rect 7380 24890 7432 24896
rect 7484 24834 7512 25298
rect 7392 24806 7512 24834
rect 7392 24274 7420 24806
rect 7472 24608 7524 24614
rect 7472 24550 7524 24556
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 7380 24064 7432 24070
rect 7380 24006 7432 24012
rect 7392 23322 7420 24006
rect 7380 23316 7432 23322
rect 7380 23258 7432 23264
rect 7484 23254 7512 24550
rect 7576 24206 7604 31078
rect 7944 30734 7972 32914
rect 7932 30728 7984 30734
rect 7932 30670 7984 30676
rect 7932 30592 7984 30598
rect 7932 30534 7984 30540
rect 7944 30258 7972 30534
rect 8036 30326 8064 34478
rect 8220 33998 8248 34546
rect 8300 34060 8352 34066
rect 8300 34002 8352 34008
rect 8208 33992 8260 33998
rect 8208 33934 8260 33940
rect 8220 33454 8248 33934
rect 8208 33448 8260 33454
rect 8128 33408 8208 33436
rect 8128 32910 8156 33408
rect 8208 33390 8260 33396
rect 8116 32904 8168 32910
rect 8116 32846 8168 32852
rect 8116 32564 8168 32570
rect 8116 32506 8168 32512
rect 8128 30734 8156 32506
rect 8312 31346 8340 34002
rect 8392 33924 8444 33930
rect 8392 33866 8444 33872
rect 8404 31482 8432 33866
rect 8484 33856 8536 33862
rect 8484 33798 8536 33804
rect 8496 33386 8524 33798
rect 8484 33380 8536 33386
rect 8484 33322 8536 33328
rect 8496 32978 8524 33322
rect 8484 32972 8536 32978
rect 8484 32914 8536 32920
rect 8588 31754 8616 37062
rect 8772 36786 8800 37062
rect 8760 36780 8812 36786
rect 8760 36722 8812 36728
rect 8772 35630 8800 36722
rect 8956 36122 8984 37828
rect 9220 37810 9272 37816
rect 9324 37806 9352 38286
rect 9128 37800 9180 37806
rect 9128 37742 9180 37748
rect 9312 37800 9364 37806
rect 9312 37742 9364 37748
rect 9036 37188 9088 37194
rect 9036 37130 9088 37136
rect 9048 36922 9076 37130
rect 9036 36916 9088 36922
rect 9036 36858 9088 36864
rect 9140 36802 9168 37742
rect 9312 37664 9364 37670
rect 9312 37606 9364 37612
rect 9048 36774 9168 36802
rect 9048 36718 9076 36774
rect 9036 36712 9088 36718
rect 9036 36654 9088 36660
rect 8864 36094 8984 36122
rect 8760 35624 8812 35630
rect 8760 35566 8812 35572
rect 8864 35306 8892 36094
rect 9048 36038 9076 36654
rect 9220 36576 9272 36582
rect 9220 36518 9272 36524
rect 9128 36168 9180 36174
rect 9128 36110 9180 36116
rect 8944 36032 8996 36038
rect 8944 35974 8996 35980
rect 9036 36032 9088 36038
rect 9036 35974 9088 35980
rect 8668 35284 8720 35290
rect 8668 35226 8720 35232
rect 8772 35278 8892 35306
rect 8680 34610 8708 35226
rect 8668 34604 8720 34610
rect 8668 34546 8720 34552
rect 8680 33522 8708 34546
rect 8772 33658 8800 35278
rect 8852 35216 8904 35222
rect 8852 35158 8904 35164
rect 8760 33652 8812 33658
rect 8760 33594 8812 33600
rect 8668 33516 8720 33522
rect 8668 33458 8720 33464
rect 8680 32842 8708 33458
rect 8668 32836 8720 32842
rect 8668 32778 8720 32784
rect 8760 32768 8812 32774
rect 8760 32710 8812 32716
rect 8772 32434 8800 32710
rect 8760 32428 8812 32434
rect 8760 32370 8812 32376
rect 8668 32360 8720 32366
rect 8668 32302 8720 32308
rect 8680 32026 8708 32302
rect 8668 32020 8720 32026
rect 8668 31962 8720 31968
rect 8864 31822 8892 35158
rect 8956 35154 8984 35974
rect 9140 35834 9168 36110
rect 9128 35828 9180 35834
rect 9128 35770 9180 35776
rect 9232 35714 9260 36518
rect 9324 36174 9352 37606
rect 9312 36168 9364 36174
rect 9312 36110 9364 36116
rect 9048 35686 9260 35714
rect 8944 35148 8996 35154
rect 8944 35090 8996 35096
rect 8944 34536 8996 34542
rect 8944 34478 8996 34484
rect 8956 33862 8984 34478
rect 8944 33856 8996 33862
rect 8944 33798 8996 33804
rect 8852 31816 8904 31822
rect 8852 31758 8904 31764
rect 8496 31726 8616 31754
rect 8392 31476 8444 31482
rect 8392 31418 8444 31424
rect 8300 31340 8352 31346
rect 8300 31282 8352 31288
rect 8116 30728 8168 30734
rect 8116 30670 8168 30676
rect 8024 30320 8076 30326
rect 8024 30262 8076 30268
rect 7932 30252 7984 30258
rect 7932 30194 7984 30200
rect 7840 30048 7892 30054
rect 7840 29990 7892 29996
rect 7656 29504 7708 29510
rect 7656 29446 7708 29452
rect 7668 28558 7696 29446
rect 7748 29096 7800 29102
rect 7748 29038 7800 29044
rect 7760 28626 7788 29038
rect 7748 28620 7800 28626
rect 7748 28562 7800 28568
rect 7656 28552 7708 28558
rect 7656 28494 7708 28500
rect 7656 26444 7708 26450
rect 7760 26432 7788 28562
rect 7708 26404 7788 26432
rect 7656 26386 7708 26392
rect 7668 25945 7696 26386
rect 7852 26382 7880 29990
rect 8496 29170 8524 31726
rect 9048 31346 9076 35686
rect 9220 35488 9272 35494
rect 9220 35430 9272 35436
rect 9232 35086 9260 35430
rect 9220 35080 9272 35086
rect 9220 35022 9272 35028
rect 9416 33946 9444 38490
rect 9508 38010 9536 38898
rect 9588 38412 9640 38418
rect 9588 38354 9640 38360
rect 9600 38214 9628 38354
rect 9692 38350 9720 39306
rect 9680 38344 9732 38350
rect 9680 38286 9732 38292
rect 9588 38208 9640 38214
rect 9588 38150 9640 38156
rect 9496 38004 9548 38010
rect 9496 37946 9548 37952
rect 9784 37346 9812 40462
rect 9956 38208 10008 38214
rect 9956 38150 10008 38156
rect 9968 37874 9996 38150
rect 9956 37868 10008 37874
rect 9956 37810 10008 37816
rect 10048 37868 10100 37874
rect 10048 37810 10100 37816
rect 9600 37318 9812 37346
rect 9600 36582 9628 37318
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 9772 37256 9824 37262
rect 9772 37198 9824 37204
rect 9692 36854 9720 37198
rect 9680 36848 9732 36854
rect 9680 36790 9732 36796
rect 9588 36576 9640 36582
rect 9588 36518 9640 36524
rect 9784 36378 9812 37198
rect 9864 36916 9916 36922
rect 9864 36858 9916 36864
rect 9772 36372 9824 36378
rect 9772 36314 9824 36320
rect 9680 36304 9732 36310
rect 9680 36246 9732 36252
rect 9692 36145 9720 36246
rect 9678 36136 9734 36145
rect 9678 36071 9734 36080
rect 9680 35760 9732 35766
rect 9680 35702 9732 35708
rect 9692 34950 9720 35702
rect 9680 34944 9732 34950
rect 9680 34886 9732 34892
rect 9772 34672 9824 34678
rect 9772 34614 9824 34620
rect 9680 34536 9732 34542
rect 9680 34478 9732 34484
rect 9692 34134 9720 34478
rect 9680 34128 9732 34134
rect 9680 34070 9732 34076
rect 9784 34066 9812 34614
rect 9772 34060 9824 34066
rect 9772 34002 9824 34008
rect 9232 33918 9444 33946
rect 9680 33992 9732 33998
rect 9680 33934 9732 33940
rect 9232 33114 9260 33918
rect 9404 33856 9456 33862
rect 9404 33798 9456 33804
rect 9312 33312 9364 33318
rect 9312 33254 9364 33260
rect 9220 33108 9272 33114
rect 9220 33050 9272 33056
rect 9324 32978 9352 33254
rect 9312 32972 9364 32978
rect 9312 32914 9364 32920
rect 9416 32910 9444 33798
rect 9496 33584 9548 33590
rect 9496 33526 9548 33532
rect 9220 32904 9272 32910
rect 9220 32846 9272 32852
rect 9404 32904 9456 32910
rect 9404 32846 9456 32852
rect 9232 32570 9260 32846
rect 9220 32564 9272 32570
rect 9220 32506 9272 32512
rect 9128 31884 9180 31890
rect 9128 31826 9180 31832
rect 9036 31340 9088 31346
rect 9036 31282 9088 31288
rect 8852 31136 8904 31142
rect 8852 31078 8904 31084
rect 8864 30938 8892 31078
rect 8852 30932 8904 30938
rect 8852 30874 8904 30880
rect 8576 30592 8628 30598
rect 8576 30534 8628 30540
rect 8588 30258 8616 30534
rect 9048 30433 9076 31282
rect 9034 30424 9090 30433
rect 9034 30359 9090 30368
rect 9140 30258 9168 31826
rect 9232 30734 9260 32506
rect 9220 30728 9272 30734
rect 9220 30670 9272 30676
rect 9220 30592 9272 30598
rect 9220 30534 9272 30540
rect 8576 30252 8628 30258
rect 8576 30194 8628 30200
rect 9128 30252 9180 30258
rect 9128 30194 9180 30200
rect 8484 29164 8536 29170
rect 8484 29106 8536 29112
rect 8668 28416 8720 28422
rect 8668 28358 8720 28364
rect 8944 28416 8996 28422
rect 8944 28358 8996 28364
rect 8680 28082 8708 28358
rect 8956 28150 8984 28358
rect 8944 28144 8996 28150
rect 8944 28086 8996 28092
rect 8668 28076 8720 28082
rect 8668 28018 8720 28024
rect 8760 28076 8812 28082
rect 8760 28018 8812 28024
rect 7932 27872 7984 27878
rect 7932 27814 7984 27820
rect 7944 26926 7972 27814
rect 8772 27606 8800 28018
rect 9128 27668 9180 27674
rect 9128 27610 9180 27616
rect 8760 27600 8812 27606
rect 9036 27600 9088 27606
rect 8760 27542 8812 27548
rect 9034 27568 9036 27577
rect 9088 27568 9090 27577
rect 8208 27532 8260 27538
rect 9034 27503 9090 27512
rect 8208 27474 8260 27480
rect 8024 27056 8076 27062
rect 8024 26998 8076 27004
rect 7932 26920 7984 26926
rect 7932 26862 7984 26868
rect 7840 26376 7892 26382
rect 7840 26318 7892 26324
rect 7654 25936 7710 25945
rect 7654 25871 7710 25880
rect 7668 25362 7696 25871
rect 7656 25356 7708 25362
rect 7656 25298 7708 25304
rect 7748 25356 7800 25362
rect 7748 25298 7800 25304
rect 7656 24948 7708 24954
rect 7760 24936 7788 25298
rect 7840 25288 7892 25294
rect 7944 25265 7972 26862
rect 8036 25974 8064 26998
rect 8116 26308 8168 26314
rect 8116 26250 8168 26256
rect 8024 25968 8076 25974
rect 8024 25910 8076 25916
rect 7840 25230 7892 25236
rect 7930 25256 7986 25265
rect 7708 24908 7788 24936
rect 7656 24890 7708 24896
rect 7564 24200 7616 24206
rect 7564 24142 7616 24148
rect 7656 24200 7708 24206
rect 7656 24142 7708 24148
rect 7668 24052 7696 24142
rect 7576 24024 7696 24052
rect 7472 23248 7524 23254
rect 7472 23190 7524 23196
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7392 21690 7420 23054
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 7300 20998 7512 21026
rect 7288 20868 7340 20874
rect 7288 20810 7340 20816
rect 7196 17264 7248 17270
rect 7196 17206 7248 17212
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7208 16794 7236 17070
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6840 15638 6868 16390
rect 6932 16114 6960 16390
rect 7208 16250 7236 16458
rect 7300 16250 7328 20810
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7300 16130 7328 16186
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7208 16102 7328 16130
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7116 15706 7144 15982
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6748 15026 6776 15098
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6748 14550 6776 14962
rect 6840 14890 6868 15302
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6472 12294 6592 12322
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6196 11614 6408 11642
rect 5915 11452 6223 11472
rect 5915 11450 5921 11452
rect 5977 11450 6001 11452
rect 6057 11450 6081 11452
rect 6137 11450 6161 11452
rect 6217 11450 6223 11452
rect 5977 11398 5979 11450
rect 6159 11398 6161 11450
rect 5915 11396 5921 11398
rect 5977 11396 6001 11398
rect 6057 11396 6081 11398
rect 6137 11396 6161 11398
rect 6217 11396 6223 11398
rect 5915 11376 6223 11396
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5915 10364 6223 10384
rect 5915 10362 5921 10364
rect 5977 10362 6001 10364
rect 6057 10362 6081 10364
rect 6137 10362 6161 10364
rect 6217 10362 6223 10364
rect 5977 10310 5979 10362
rect 6159 10310 6161 10362
rect 5915 10308 5921 10310
rect 5977 10308 6001 10310
rect 6057 10308 6081 10310
rect 6137 10308 6161 10310
rect 6217 10308 6223 10310
rect 5915 10288 6223 10308
rect 5644 10220 5764 10248
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5262 9072 5318 9081
rect 5262 9007 5318 9016
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 5000 4826 5028 8842
rect 5276 7342 5304 9007
rect 5460 8906 5488 9522
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5460 7818 5488 8842
rect 5644 8650 5672 10220
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5644 8622 5708 8650
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5680 8514 5708 8622
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5276 6798 5304 7278
rect 5460 6866 5488 7754
rect 5552 7478 5580 8502
rect 5680 8486 5764 8514
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4908 3194 4936 4082
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4816 3074 4844 3130
rect 4816 3046 4936 3074
rect 5000 3058 5028 3878
rect 5092 3670 5120 3878
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 5184 3466 5212 4422
rect 5552 4146 5580 7414
rect 5736 5914 5764 8486
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5736 5166 5764 5850
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5828 4826 5856 9998
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 6012 9722 6040 9930
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 5915 9276 6223 9296
rect 5915 9274 5921 9276
rect 5977 9274 6001 9276
rect 6057 9274 6081 9276
rect 6137 9274 6161 9276
rect 6217 9274 6223 9276
rect 5977 9222 5979 9274
rect 6159 9222 6161 9274
rect 5915 9220 5921 9222
rect 5977 9220 6001 9222
rect 6057 9220 6081 9222
rect 6137 9220 6161 9222
rect 6217 9220 6223 9222
rect 5915 9200 6223 9220
rect 6288 8650 6316 11290
rect 6380 8906 6408 11614
rect 6472 11558 6500 12174
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 9518 6500 9862
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6288 8622 6408 8650
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 5915 8188 6223 8208
rect 5915 8186 5921 8188
rect 5977 8186 6001 8188
rect 6057 8186 6081 8188
rect 6137 8186 6161 8188
rect 6217 8186 6223 8188
rect 5977 8134 5979 8186
rect 6159 8134 6161 8186
rect 5915 8132 5921 8134
rect 5977 8132 6001 8134
rect 6057 8132 6081 8134
rect 6137 8132 6161 8134
rect 6217 8132 6223 8134
rect 5915 8112 6223 8132
rect 6288 7886 6316 8434
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6288 7410 6316 7822
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 5915 7100 6223 7120
rect 5915 7098 5921 7100
rect 5977 7098 6001 7100
rect 6057 7098 6081 7100
rect 6137 7098 6161 7100
rect 6217 7098 6223 7100
rect 5977 7046 5979 7098
rect 6159 7046 6161 7098
rect 5915 7044 5921 7046
rect 5977 7044 6001 7046
rect 6057 7044 6081 7046
rect 6137 7044 6161 7046
rect 6217 7044 6223 7046
rect 5915 7024 6223 7044
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6196 6322 6224 6734
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 5915 6012 6223 6032
rect 5915 6010 5921 6012
rect 5977 6010 6001 6012
rect 6057 6010 6081 6012
rect 6137 6010 6161 6012
rect 6217 6010 6223 6012
rect 5977 5958 5979 6010
rect 6159 5958 6161 6010
rect 5915 5956 5921 5958
rect 5977 5956 6001 5958
rect 6057 5956 6081 5958
rect 6137 5956 6161 5958
rect 6217 5956 6223 5958
rect 5915 5936 6223 5956
rect 6288 5710 6316 7346
rect 6380 6118 6408 8622
rect 6472 6798 6500 9454
rect 6564 6866 6592 12294
rect 6656 10130 6684 14350
rect 7024 14090 7052 14418
rect 7116 14414 7144 15302
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 6932 14062 7052 14090
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6748 9450 6776 13874
rect 6932 13870 6960 14062
rect 7116 13938 7144 14214
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 7024 13462 7052 13874
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6840 12918 6868 13126
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6840 11150 6868 12854
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7116 12238 7144 12582
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7208 12084 7236 16102
rect 7392 13938 7420 20742
rect 7484 16153 7512 20998
rect 7470 16144 7526 16153
rect 7470 16079 7526 16088
rect 7576 15994 7604 24024
rect 7760 23882 7788 24908
rect 7668 23854 7788 23882
rect 7668 23186 7696 23854
rect 7748 23248 7800 23254
rect 7748 23190 7800 23196
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 7668 21078 7696 23122
rect 7656 21072 7708 21078
rect 7656 21014 7708 21020
rect 7760 19768 7788 23190
rect 7852 21894 7880 25230
rect 7930 25191 7986 25200
rect 7944 24138 7972 25191
rect 8128 24954 8156 26250
rect 8116 24948 8168 24954
rect 8116 24890 8168 24896
rect 8114 24848 8170 24857
rect 8114 24783 8116 24792
rect 8168 24783 8170 24792
rect 8116 24754 8168 24760
rect 8220 24274 8248 27474
rect 8392 27464 8444 27470
rect 8390 27432 8392 27441
rect 8852 27464 8904 27470
rect 8444 27432 8446 27441
rect 8852 27406 8904 27412
rect 8390 27367 8446 27376
rect 8576 27124 8628 27130
rect 8576 27066 8628 27072
rect 8300 26988 8352 26994
rect 8300 26930 8352 26936
rect 8312 26586 8340 26930
rect 8392 26852 8444 26858
rect 8392 26794 8444 26800
rect 8300 26580 8352 26586
rect 8300 26522 8352 26528
rect 8300 26376 8352 26382
rect 8300 26318 8352 26324
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 7932 24132 7984 24138
rect 7932 24074 7984 24080
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7944 21622 7972 24074
rect 8114 23624 8170 23633
rect 8114 23559 8170 23568
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 8036 22642 8064 23462
rect 8128 22778 8156 23559
rect 8220 23254 8248 24210
rect 8208 23248 8260 23254
rect 8208 23190 8260 23196
rect 8312 22794 8340 26318
rect 8404 25362 8432 26794
rect 8588 26382 8616 27066
rect 8668 26920 8720 26926
rect 8668 26862 8720 26868
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 8574 25936 8630 25945
rect 8574 25871 8576 25880
rect 8628 25871 8630 25880
rect 8576 25842 8628 25848
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 8576 24812 8628 24818
rect 8576 24754 8628 24760
rect 8588 24410 8616 24754
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8576 24132 8628 24138
rect 8576 24074 8628 24080
rect 8484 23588 8536 23594
rect 8484 23530 8536 23536
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8404 23322 8432 23462
rect 8392 23316 8444 23322
rect 8392 23258 8444 23264
rect 8496 23118 8524 23530
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 8484 23112 8536 23118
rect 8484 23054 8536 23060
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8220 22766 8340 22794
rect 8024 22636 8076 22642
rect 8024 22578 8076 22584
rect 7932 21616 7984 21622
rect 7932 21558 7984 21564
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7840 19780 7892 19786
rect 7760 19740 7840 19768
rect 7840 19722 7892 19728
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7760 16114 7788 16186
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7472 15972 7524 15978
rect 7576 15966 7788 15994
rect 7472 15914 7524 15920
rect 7484 15502 7512 15914
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7576 15026 7604 15302
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7562 14104 7618 14113
rect 7562 14039 7564 14048
rect 7616 14039 7618 14048
rect 7564 14010 7616 14016
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7116 12056 7236 12084
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6840 10062 6868 11086
rect 6932 10674 6960 11290
rect 7024 11082 7052 11698
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6840 9178 6868 9522
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 6656 8634 6684 8842
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6748 8378 6776 8774
rect 6840 8566 6868 9114
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6932 8498 6960 8774
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6828 8424 6880 8430
rect 6656 8372 6828 8378
rect 6656 8366 6880 8372
rect 6656 8350 6868 8366
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6472 6322 6500 6734
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6656 5710 6684 8350
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6840 7342 6868 8230
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7546 6960 7686
rect 7024 7546 7052 8230
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 6828 7336 6880 7342
rect 6748 7296 6828 7324
rect 6748 5846 6776 7296
rect 6828 7278 6880 7284
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 5915 4924 6223 4944
rect 5915 4922 5921 4924
rect 5977 4922 6001 4924
rect 6057 4922 6081 4924
rect 6137 4922 6161 4924
rect 6217 4922 6223 4924
rect 5977 4870 5979 4922
rect 6159 4870 6161 4922
rect 5915 4868 5921 4870
rect 5977 4868 6001 4870
rect 6057 4868 6081 4870
rect 6137 4868 6161 4870
rect 6217 4868 6223 4870
rect 5915 4848 6223 4868
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5552 3466 5580 4082
rect 5644 4078 5672 4694
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5552 3126 5580 3402
rect 5736 3398 5764 4422
rect 5828 3398 5856 4762
rect 6288 4622 6316 5646
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 6196 4026 6224 4490
rect 6196 3998 6316 4026
rect 6288 3942 6316 3998
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 5915 3836 6223 3856
rect 5915 3834 5921 3836
rect 5977 3834 6001 3836
rect 6057 3834 6081 3836
rect 6137 3834 6161 3836
rect 6217 3834 6223 3836
rect 5977 3782 5979 3834
rect 6159 3782 6161 3834
rect 5915 3780 5921 3782
rect 5977 3780 6001 3782
rect 6057 3780 6081 3782
rect 6137 3780 6161 3782
rect 6217 3780 6223 3782
rect 5915 3760 6223 3780
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 4908 2938 4936 3046
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 4908 2922 5028 2938
rect 4908 2916 5040 2922
rect 4908 2910 4988 2916
rect 4988 2858 5040 2864
rect 6380 2854 6408 5578
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6472 4554 6500 5170
rect 6656 4758 6684 5646
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6644 4616 6696 4622
rect 6748 4570 6776 5782
rect 6840 5710 6868 6598
rect 6932 6458 6960 6666
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 7024 6322 7052 6938
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6840 5370 6868 5646
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 7024 5302 7052 5510
rect 7012 5296 7064 5302
rect 7012 5238 7064 5244
rect 7116 4690 7144 12056
rect 7300 10810 7328 12174
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7208 8566 7236 8842
rect 7392 8838 7420 13194
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7484 11014 7512 12922
rect 7576 12170 7604 13806
rect 7668 12238 7696 15302
rect 7760 12646 7788 15966
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7576 11354 7604 11698
rect 7760 11694 7788 12174
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7668 11150 7696 11290
rect 7760 11150 7788 11494
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7472 11008 7524 11014
rect 7852 10996 7880 19722
rect 7944 19378 7972 21286
rect 8022 19952 8078 19961
rect 8022 19887 8078 19896
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7944 16250 7972 17138
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7944 16114 7972 16186
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7944 15706 7972 15914
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7932 15428 7984 15434
rect 7932 15370 7984 15376
rect 7944 13870 7972 15370
rect 8036 14414 8064 19887
rect 8128 18698 8156 22714
rect 8220 22166 8248 22766
rect 8300 22704 8352 22710
rect 8300 22646 8352 22652
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 8206 21992 8262 22001
rect 8312 21962 8340 22646
rect 8206 21927 8262 21936
rect 8300 21956 8352 21962
rect 8220 19514 8248 21927
rect 8300 21898 8352 21904
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8208 18760 8260 18766
rect 8312 18748 8340 21898
rect 8404 20058 8432 23054
rect 8496 21554 8524 23054
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 8496 21146 8524 21490
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8484 20868 8536 20874
rect 8484 20810 8536 20816
rect 8496 20602 8524 20810
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8496 19854 8524 20402
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8260 18720 8340 18748
rect 8208 18702 8260 18708
rect 8116 18692 8168 18698
rect 8116 18634 8168 18640
rect 8312 17746 8340 18720
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8128 16658 8156 17682
rect 8404 17626 8432 19654
rect 8312 17598 8432 17626
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8128 16046 8156 16594
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8128 14346 8156 14486
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8036 13977 8064 14010
rect 8022 13968 8078 13977
rect 8022 13903 8078 13912
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 8128 13326 8156 14282
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7472 10950 7524 10956
rect 7760 10968 7880 10996
rect 7760 10606 7788 10968
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7668 9654 7696 9930
rect 7656 9648 7708 9654
rect 7708 9608 7788 9636
rect 7656 9590 7708 9596
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7208 7342 7236 7754
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7300 7002 7328 7346
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 6696 4564 6776 4570
rect 6644 4558 6776 4564
rect 6460 4548 6512 4554
rect 6656 4542 6776 4558
rect 6460 4490 6512 4496
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7116 4146 7144 4422
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 5915 2748 6223 2768
rect 5915 2746 5921 2748
rect 5977 2746 6001 2748
rect 6057 2746 6081 2748
rect 6137 2746 6161 2748
rect 6217 2746 6223 2748
rect 5977 2694 5979 2746
rect 6159 2694 6161 2746
rect 5915 2692 5921 2694
rect 5977 2692 6001 2694
rect 6057 2692 6081 2694
rect 6137 2692 6161 2694
rect 6217 2692 6223 2694
rect 5915 2672 6223 2692
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 4172 800 4200 2314
rect 4908 800 4936 2382
rect 5736 800 5764 2382
rect 6472 800 6500 2994
rect 7208 800 7236 2994
rect 7392 2922 7420 7482
rect 7484 4214 7512 9522
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7668 7750 7696 8298
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7668 6390 7696 7686
rect 7760 6458 7788 9608
rect 7852 8566 7880 10610
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7760 6322 7788 6394
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7576 4622 7604 6258
rect 7944 6186 7972 12650
rect 8036 12374 8064 12786
rect 8024 12368 8076 12374
rect 8024 12310 8076 12316
rect 8036 11558 8064 12310
rect 8128 12306 8156 13262
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8220 11744 8248 17478
rect 8312 15434 8340 17598
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8404 17270 8432 17478
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 15502 8432 16934
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8312 15314 8340 15370
rect 8312 15286 8432 15314
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8312 12714 8340 14418
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8312 12238 8340 12650
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8128 11716 8248 11744
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8128 7290 8156 11716
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 8220 11150 8248 11562
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8312 8974 8340 9454
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8036 7262 8156 7290
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 8036 5030 8064 7262
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 6798 8156 7142
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8404 5642 8432 15286
rect 8496 13462 8524 19790
rect 8588 16454 8616 24074
rect 8680 18358 8708 26862
rect 8760 25832 8812 25838
rect 8760 25774 8812 25780
rect 8772 25294 8800 25774
rect 8760 25288 8812 25294
rect 8760 25230 8812 25236
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 8772 23730 8800 24754
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8772 20398 8800 23666
rect 8864 20602 8892 27406
rect 8944 26988 8996 26994
rect 8944 26930 8996 26936
rect 8956 26382 8984 26930
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 8956 25752 8984 26318
rect 9048 25820 9076 27503
rect 9140 27470 9168 27610
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9232 27146 9260 30534
rect 9312 30048 9364 30054
rect 9312 29990 9364 29996
rect 9324 28558 9352 29990
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 9508 28490 9536 33526
rect 9692 33114 9720 33934
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 9772 32224 9824 32230
rect 9772 32166 9824 32172
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 9692 31142 9720 31962
rect 9784 31686 9812 32166
rect 9876 31958 9904 36858
rect 9956 36576 10008 36582
rect 10060 36564 10088 37810
rect 10008 36536 10088 36564
rect 9956 36518 10008 36524
rect 9968 35086 9996 36518
rect 10046 36272 10102 36281
rect 10046 36207 10048 36216
rect 10100 36207 10102 36216
rect 10048 36178 10100 36184
rect 10048 35692 10100 35698
rect 10048 35634 10100 35640
rect 10060 35290 10088 35634
rect 10048 35284 10100 35290
rect 10048 35226 10100 35232
rect 9956 35080 10008 35086
rect 9956 35022 10008 35028
rect 10152 34134 10180 41482
rect 10244 35630 10272 41686
rect 10336 36922 10364 42570
rect 10324 36916 10376 36922
rect 10324 36858 10376 36864
rect 10520 36786 10548 44474
rect 18052 44260 18104 44266
rect 18052 44202 18104 44208
rect 17960 44192 18012 44198
rect 17960 44134 18012 44140
rect 15846 44092 16154 44112
rect 15846 44090 15852 44092
rect 15908 44090 15932 44092
rect 15988 44090 16012 44092
rect 16068 44090 16092 44092
rect 16148 44090 16154 44092
rect 15908 44038 15910 44090
rect 16090 44038 16092 44090
rect 15846 44036 15852 44038
rect 15908 44036 15932 44038
rect 15988 44036 16012 44038
rect 16068 44036 16092 44038
rect 16148 44036 16154 44038
rect 15846 44016 16154 44036
rect 17972 43722 18000 44134
rect 10692 43716 10744 43722
rect 10692 43658 10744 43664
rect 17960 43716 18012 43722
rect 17960 43658 18012 43664
rect 10600 38344 10652 38350
rect 10600 38286 10652 38292
rect 10612 37874 10640 38286
rect 10600 37868 10652 37874
rect 10600 37810 10652 37816
rect 10704 37754 10732 43658
rect 10880 43548 11188 43568
rect 10880 43546 10886 43548
rect 10942 43546 10966 43548
rect 11022 43546 11046 43548
rect 11102 43546 11126 43548
rect 11182 43546 11188 43548
rect 10942 43494 10944 43546
rect 11124 43494 11126 43546
rect 10880 43492 10886 43494
rect 10942 43492 10966 43494
rect 11022 43492 11046 43494
rect 11102 43492 11126 43494
rect 11182 43492 11188 43494
rect 10880 43472 11188 43492
rect 18064 43450 18092 44202
rect 18156 43994 18184 44474
rect 18328 44396 18380 44402
rect 18328 44338 18380 44344
rect 18144 43988 18196 43994
rect 18144 43930 18196 43936
rect 18340 43790 18368 44338
rect 25776 44092 26084 44112
rect 25776 44090 25782 44092
rect 25838 44090 25862 44092
rect 25918 44090 25942 44092
rect 25998 44090 26022 44092
rect 26078 44090 26084 44092
rect 25838 44038 25840 44090
rect 26020 44038 26022 44090
rect 25776 44036 25782 44038
rect 25838 44036 25862 44038
rect 25918 44036 25942 44038
rect 25998 44036 26022 44038
rect 26078 44036 26084 44038
rect 25776 44016 26084 44036
rect 29012 43790 29040 44678
rect 29932 44334 29960 45222
rect 30208 44878 30236 47087
rect 30196 44872 30248 44878
rect 30196 44814 30248 44820
rect 30104 44396 30156 44402
rect 30104 44338 30156 44344
rect 29920 44328 29972 44334
rect 29920 44270 29972 44276
rect 29920 44192 29972 44198
rect 29920 44134 29972 44140
rect 18328 43784 18380 43790
rect 18328 43726 18380 43732
rect 29000 43784 29052 43790
rect 29000 43726 29052 43732
rect 18052 43444 18104 43450
rect 18052 43386 18104 43392
rect 18340 43314 18368 43726
rect 20811 43548 21119 43568
rect 20811 43546 20817 43548
rect 20873 43546 20897 43548
rect 20953 43546 20977 43548
rect 21033 43546 21057 43548
rect 21113 43546 21119 43548
rect 20873 43494 20875 43546
rect 21055 43494 21057 43546
rect 20811 43492 20817 43494
rect 20873 43492 20897 43494
rect 20953 43492 20977 43494
rect 21033 43492 21057 43494
rect 21113 43492 21119 43494
rect 20811 43472 21119 43492
rect 18328 43308 18380 43314
rect 18328 43250 18380 43256
rect 19064 43308 19116 43314
rect 19064 43250 19116 43256
rect 15846 43004 16154 43024
rect 15846 43002 15852 43004
rect 15908 43002 15932 43004
rect 15988 43002 16012 43004
rect 16068 43002 16092 43004
rect 16148 43002 16154 43004
rect 15908 42950 15910 43002
rect 16090 42950 16092 43002
rect 15846 42948 15852 42950
rect 15908 42948 15932 42950
rect 15988 42948 16012 42950
rect 16068 42948 16092 42950
rect 16148 42948 16154 42950
rect 15846 42928 16154 42948
rect 10880 42460 11188 42480
rect 10880 42458 10886 42460
rect 10942 42458 10966 42460
rect 11022 42458 11046 42460
rect 11102 42458 11126 42460
rect 11182 42458 11188 42460
rect 10942 42406 10944 42458
rect 11124 42406 11126 42458
rect 10880 42404 10886 42406
rect 10942 42404 10966 42406
rect 11022 42404 11046 42406
rect 11102 42404 11126 42406
rect 11182 42404 11188 42406
rect 10880 42384 11188 42404
rect 15846 41916 16154 41936
rect 15846 41914 15852 41916
rect 15908 41914 15932 41916
rect 15988 41914 16012 41916
rect 16068 41914 16092 41916
rect 16148 41914 16154 41916
rect 15908 41862 15910 41914
rect 16090 41862 16092 41914
rect 15846 41860 15852 41862
rect 15908 41860 15932 41862
rect 15988 41860 16012 41862
rect 16068 41860 16092 41862
rect 16148 41860 16154 41862
rect 15846 41840 16154 41860
rect 12992 41608 13044 41614
rect 12992 41550 13044 41556
rect 15752 41608 15804 41614
rect 15752 41550 15804 41556
rect 12624 41472 12676 41478
rect 12624 41414 12676 41420
rect 10880 41372 11188 41392
rect 10880 41370 10886 41372
rect 10942 41370 10966 41372
rect 11022 41370 11046 41372
rect 11102 41370 11126 41372
rect 11182 41370 11188 41372
rect 10942 41318 10944 41370
rect 11124 41318 11126 41370
rect 10880 41316 10886 41318
rect 10942 41316 10966 41318
rect 11022 41316 11046 41318
rect 11102 41316 11126 41318
rect 11182 41316 11188 41318
rect 10880 41296 11188 41316
rect 12636 41070 12664 41414
rect 12624 41064 12676 41070
rect 12624 41006 12676 41012
rect 12900 41064 12952 41070
rect 12900 41006 12952 41012
rect 10880 40284 11188 40304
rect 10880 40282 10886 40284
rect 10942 40282 10966 40284
rect 11022 40282 11046 40284
rect 11102 40282 11126 40284
rect 11182 40282 11188 40284
rect 10942 40230 10944 40282
rect 11124 40230 11126 40282
rect 10880 40228 10886 40230
rect 10942 40228 10966 40230
rect 11022 40228 11046 40230
rect 11102 40228 11126 40230
rect 11182 40228 11188 40230
rect 10880 40208 11188 40228
rect 12636 40050 12664 41006
rect 12912 40050 12940 41006
rect 13004 40730 13032 41550
rect 14464 41132 14516 41138
rect 14464 41074 14516 41080
rect 15568 41132 15620 41138
rect 15568 41074 15620 41080
rect 13544 41064 13596 41070
rect 13544 41006 13596 41012
rect 13728 41064 13780 41070
rect 14004 41064 14056 41070
rect 13780 41012 13860 41018
rect 13728 41006 13860 41012
rect 14004 41006 14056 41012
rect 12992 40724 13044 40730
rect 12992 40666 13044 40672
rect 13556 40594 13584 41006
rect 13740 40990 13860 41006
rect 13544 40588 13596 40594
rect 13544 40530 13596 40536
rect 12992 40520 13044 40526
rect 12992 40462 13044 40468
rect 12624 40044 12676 40050
rect 12624 39986 12676 39992
rect 12900 40044 12952 40050
rect 12900 39986 12952 39992
rect 12912 39438 12940 39986
rect 13004 39642 13032 40462
rect 13556 39982 13584 40530
rect 13832 40390 13860 40990
rect 13820 40384 13872 40390
rect 13820 40326 13872 40332
rect 13832 39982 13860 40326
rect 14016 39982 14044 41006
rect 13544 39976 13596 39982
rect 13544 39918 13596 39924
rect 13820 39976 13872 39982
rect 13820 39918 13872 39924
rect 14004 39976 14056 39982
rect 14004 39918 14056 39924
rect 12992 39636 13044 39642
rect 12992 39578 13044 39584
rect 12900 39432 12952 39438
rect 12900 39374 12952 39380
rect 10784 39296 10836 39302
rect 10784 39238 10836 39244
rect 10796 38486 10824 39238
rect 10880 39196 11188 39216
rect 10880 39194 10886 39196
rect 10942 39194 10966 39196
rect 11022 39194 11046 39196
rect 11102 39194 11126 39196
rect 11182 39194 11188 39196
rect 10942 39142 10944 39194
rect 11124 39142 11126 39194
rect 10880 39140 10886 39142
rect 10942 39140 10966 39142
rect 11022 39140 11046 39142
rect 11102 39140 11126 39142
rect 11182 39140 11188 39142
rect 10880 39120 11188 39140
rect 12624 38956 12676 38962
rect 12624 38898 12676 38904
rect 10784 38480 10836 38486
rect 10784 38422 10836 38428
rect 12532 38208 12584 38214
rect 12532 38150 12584 38156
rect 10880 38108 11188 38128
rect 10880 38106 10886 38108
rect 10942 38106 10966 38108
rect 11022 38106 11046 38108
rect 11102 38106 11126 38108
rect 11182 38106 11188 38108
rect 10942 38054 10944 38106
rect 11124 38054 11126 38106
rect 10880 38052 10886 38054
rect 10942 38052 10966 38054
rect 11022 38052 11046 38054
rect 11102 38052 11126 38054
rect 11182 38052 11188 38054
rect 10880 38032 11188 38052
rect 12544 37942 12572 38150
rect 12532 37936 12584 37942
rect 12532 37878 12584 37884
rect 12636 37874 12664 38898
rect 12912 38554 12940 39374
rect 13556 39098 13584 39918
rect 13544 39092 13596 39098
rect 13544 39034 13596 39040
rect 13832 39030 13860 39918
rect 14280 39500 14332 39506
rect 14280 39442 14332 39448
rect 14096 39364 14148 39370
rect 14096 39306 14148 39312
rect 13820 39024 13872 39030
rect 13820 38966 13872 38972
rect 14004 38888 14056 38894
rect 14004 38830 14056 38836
rect 12900 38548 12952 38554
rect 12900 38490 12952 38496
rect 12716 38344 12768 38350
rect 12716 38286 12768 38292
rect 13176 38344 13228 38350
rect 13176 38286 13228 38292
rect 12728 38010 12756 38286
rect 12716 38004 12768 38010
rect 12716 37946 12768 37952
rect 12624 37868 12676 37874
rect 12624 37810 12676 37816
rect 13084 37868 13136 37874
rect 13084 37810 13136 37816
rect 10612 37726 10732 37754
rect 10416 36780 10468 36786
rect 10416 36722 10468 36728
rect 10508 36780 10560 36786
rect 10508 36722 10560 36728
rect 10324 36712 10376 36718
rect 10324 36654 10376 36660
rect 10336 36174 10364 36654
rect 10428 36378 10456 36722
rect 10612 36378 10640 37726
rect 10876 37664 10928 37670
rect 10876 37606 10928 37612
rect 11520 37664 11572 37670
rect 11520 37606 11572 37612
rect 10888 37330 10916 37606
rect 10876 37324 10928 37330
rect 10876 37266 10928 37272
rect 11244 37188 11296 37194
rect 11244 37130 11296 37136
rect 10880 37020 11188 37040
rect 10880 37018 10886 37020
rect 10942 37018 10966 37020
rect 11022 37018 11046 37020
rect 11102 37018 11126 37020
rect 11182 37018 11188 37020
rect 10942 36966 10944 37018
rect 11124 36966 11126 37018
rect 10880 36964 10886 36966
rect 10942 36964 10966 36966
rect 11022 36964 11046 36966
rect 11102 36964 11126 36966
rect 11182 36964 11188 36966
rect 10880 36944 11188 36964
rect 10692 36712 10744 36718
rect 10692 36654 10744 36660
rect 10704 36378 10732 36654
rect 11256 36378 11284 37130
rect 11428 37120 11480 37126
rect 11428 37062 11480 37068
rect 10416 36372 10468 36378
rect 10416 36314 10468 36320
rect 10600 36372 10652 36378
rect 10600 36314 10652 36320
rect 10692 36372 10744 36378
rect 10692 36314 10744 36320
rect 11244 36372 11296 36378
rect 11244 36314 11296 36320
rect 11336 36372 11388 36378
rect 11336 36314 11388 36320
rect 10324 36168 10376 36174
rect 10324 36110 10376 36116
rect 10336 35630 10364 36110
rect 10428 35766 10456 36314
rect 10416 35760 10468 35766
rect 10416 35702 10468 35708
rect 10232 35624 10284 35630
rect 10232 35566 10284 35572
rect 10324 35624 10376 35630
rect 10324 35566 10376 35572
rect 10336 34746 10364 35566
rect 10324 34740 10376 34746
rect 10324 34682 10376 34688
rect 10232 34604 10284 34610
rect 10336 34592 10364 34682
rect 10428 34610 10456 35702
rect 10704 35562 10732 36314
rect 11348 36038 11376 36314
rect 11440 36174 11468 37062
rect 11532 36786 11560 37606
rect 12636 37330 12664 37810
rect 12716 37664 12768 37670
rect 12716 37606 12768 37612
rect 12624 37324 12676 37330
rect 12624 37266 12676 37272
rect 11520 36780 11572 36786
rect 11520 36722 11572 36728
rect 11888 36576 11940 36582
rect 11888 36518 11940 36524
rect 11520 36304 11572 36310
rect 11518 36272 11520 36281
rect 11572 36272 11574 36281
rect 11518 36207 11574 36216
rect 11428 36168 11480 36174
rect 11704 36168 11756 36174
rect 11428 36110 11480 36116
rect 11518 36136 11574 36145
rect 11704 36110 11756 36116
rect 11518 36071 11574 36080
rect 11336 36032 11388 36038
rect 11336 35974 11388 35980
rect 10880 35932 11188 35952
rect 10880 35930 10886 35932
rect 10942 35930 10966 35932
rect 11022 35930 11046 35932
rect 11102 35930 11126 35932
rect 11182 35930 11188 35932
rect 10942 35878 10944 35930
rect 11124 35878 11126 35930
rect 10880 35876 10886 35878
rect 10942 35876 10966 35878
rect 11022 35876 11046 35878
rect 11102 35876 11126 35878
rect 11182 35876 11188 35878
rect 10880 35856 11188 35876
rect 11532 35698 11560 36071
rect 11716 35834 11744 36110
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 10784 35692 10836 35698
rect 10784 35634 10836 35640
rect 11520 35692 11572 35698
rect 11520 35634 11572 35640
rect 10692 35556 10744 35562
rect 10692 35498 10744 35504
rect 10600 35488 10652 35494
rect 10600 35430 10652 35436
rect 10508 34944 10560 34950
rect 10508 34886 10560 34892
rect 10284 34564 10364 34592
rect 10416 34604 10468 34610
rect 10232 34546 10284 34552
rect 10416 34546 10468 34552
rect 10140 34128 10192 34134
rect 10140 34070 10192 34076
rect 10428 33930 10456 34546
rect 10416 33924 10468 33930
rect 10416 33866 10468 33872
rect 10428 33522 10456 33866
rect 10416 33516 10468 33522
rect 10416 33458 10468 33464
rect 10324 33108 10376 33114
rect 10324 33050 10376 33056
rect 9956 32496 10008 32502
rect 9956 32438 10008 32444
rect 9864 31952 9916 31958
rect 9864 31894 9916 31900
rect 9968 31770 9996 32438
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 10048 31816 10100 31822
rect 9968 31764 10048 31770
rect 9968 31758 10100 31764
rect 9968 31742 10088 31758
rect 9772 31680 9824 31686
rect 9772 31622 9824 31628
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9692 29322 9720 29990
rect 9772 29572 9824 29578
rect 9772 29514 9824 29520
rect 9600 29294 9720 29322
rect 9496 28484 9548 28490
rect 9496 28426 9548 28432
rect 9404 28416 9456 28422
rect 9404 28358 9456 28364
rect 9416 28218 9444 28358
rect 9404 28212 9456 28218
rect 9404 28154 9456 28160
rect 9508 27878 9536 28426
rect 9496 27872 9548 27878
rect 9416 27832 9496 27860
rect 9312 27600 9364 27606
rect 9310 27568 9312 27577
rect 9364 27568 9366 27577
rect 9310 27503 9366 27512
rect 9312 27442 9364 27448
rect 9312 27384 9364 27390
rect 9140 27118 9260 27146
rect 9140 25974 9168 27118
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 9232 26382 9260 26930
rect 9324 26790 9352 27384
rect 9416 27112 9444 27832
rect 9496 27814 9548 27820
rect 9494 27704 9550 27713
rect 9494 27639 9496 27648
rect 9548 27639 9550 27648
rect 9496 27610 9548 27616
rect 9600 27418 9628 29294
rect 9680 29232 9732 29238
rect 9680 29174 9732 29180
rect 9692 27606 9720 29174
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9600 27390 9720 27418
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 9600 27169 9628 27270
rect 9413 27084 9444 27112
rect 9586 27160 9642 27169
rect 9586 27095 9642 27104
rect 9413 27010 9441 27084
rect 9413 26994 9444 27010
rect 9404 26988 9456 26994
rect 9588 26988 9640 26994
rect 9404 26930 9456 26936
rect 9508 26948 9588 26976
rect 9312 26784 9364 26790
rect 9312 26726 9364 26732
rect 9508 26382 9536 26948
rect 9588 26930 9640 26936
rect 9692 26466 9720 27390
rect 9784 26586 9812 29514
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 9876 26790 9904 28018
rect 9864 26784 9916 26790
rect 9864 26726 9916 26732
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 9692 26438 9812 26466
rect 9220 26376 9272 26382
rect 9220 26318 9272 26324
rect 9496 26376 9548 26382
rect 9680 26376 9732 26382
rect 9496 26318 9548 26324
rect 9586 26344 9642 26353
rect 9128 25968 9180 25974
rect 9128 25910 9180 25916
rect 9048 25792 9168 25820
rect 8956 25724 9076 25752
rect 8944 25152 8996 25158
rect 8944 25094 8996 25100
rect 8956 24206 8984 25094
rect 9048 24818 9076 25724
rect 9036 24812 9088 24818
rect 9036 24754 9088 24760
rect 9140 24206 9168 25792
rect 9232 24818 9260 26318
rect 9404 26308 9456 26314
rect 9404 26250 9456 26256
rect 9416 25809 9444 26250
rect 9402 25800 9458 25809
rect 9402 25735 9458 25744
rect 9312 25288 9364 25294
rect 9310 25256 9312 25265
rect 9364 25256 9366 25265
rect 9310 25191 9366 25200
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 9140 24070 9168 24142
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9128 23792 9180 23798
rect 9128 23734 9180 23740
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 8944 23656 8996 23662
rect 8942 23624 8944 23633
rect 8996 23624 8998 23633
rect 8942 23559 8998 23568
rect 9048 23526 9076 23666
rect 9036 23520 9088 23526
rect 9036 23462 9088 23468
rect 8944 23316 8996 23322
rect 8944 23258 8996 23264
rect 8956 22098 8984 23258
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 9048 22710 9076 23054
rect 9140 22778 9168 23734
rect 9232 23594 9260 24754
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 9220 23588 9272 23594
rect 9220 23530 9272 23536
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 9036 22704 9088 22710
rect 9036 22646 9088 22652
rect 9128 22636 9180 22642
rect 9128 22578 9180 22584
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 8944 21412 8996 21418
rect 8944 21354 8996 21360
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8956 20482 8984 21354
rect 9036 20868 9088 20874
rect 9036 20810 9088 20816
rect 8864 20454 8984 20482
rect 9048 20466 9076 20810
rect 9036 20460 9088 20466
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8864 20262 8892 20454
rect 9036 20402 9088 20408
rect 8944 20324 8996 20330
rect 8944 20266 8996 20272
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8864 19786 8892 20198
rect 8852 19780 8904 19786
rect 8852 19722 8904 19728
rect 8864 19174 8892 19722
rect 8956 19718 8984 20266
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8668 18352 8720 18358
rect 8668 18294 8720 18300
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 8588 16182 8616 16390
rect 8576 16176 8628 16182
rect 8576 16118 8628 16124
rect 8668 14340 8720 14346
rect 8668 14282 8720 14288
rect 8680 13802 8708 14282
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 8588 12356 8616 13670
rect 8772 13258 8800 18634
rect 8864 17082 8892 19110
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 8956 18290 8984 18702
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 8956 17814 8984 18226
rect 8944 17808 8996 17814
rect 8944 17750 8996 17756
rect 8956 17202 8984 17750
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8864 17054 8984 17082
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8864 13938 8892 15098
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8864 13190 8892 13738
rect 8956 13190 8984 17054
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8588 12328 8708 12356
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8496 7410 8524 8434
rect 8588 7410 8616 11086
rect 8680 9382 8708 12328
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 8404 4826 8432 5170
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8496 4758 8524 7346
rect 8484 4752 8536 4758
rect 8484 4694 8536 4700
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7576 4282 7604 4558
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7484 2582 7512 2994
rect 7852 2650 7880 4558
rect 7944 4486 7972 4626
rect 8496 4622 8524 4694
rect 8116 4616 8168 4622
rect 8484 4616 8536 4622
rect 8168 4564 8340 4570
rect 8116 4558 8340 4564
rect 8484 4558 8536 4564
rect 8128 4542 8340 4558
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 8312 4078 8340 4542
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8312 2650 8340 3062
rect 8588 2774 8616 7346
rect 8680 6798 8708 8910
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8680 6118 8708 6734
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5030 8708 6054
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8680 2854 8708 4490
rect 8772 3058 8800 12106
rect 8864 10674 8892 12854
rect 8956 12646 8984 13126
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 9048 12434 9076 18226
rect 9140 17218 9168 22578
rect 9232 21962 9260 23530
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 9232 21554 9260 21898
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 9324 21010 9352 24006
rect 9416 22642 9444 25735
rect 9508 24818 9536 26318
rect 9680 26318 9732 26324
rect 9586 26279 9588 26288
rect 9640 26279 9642 26288
rect 9588 26250 9640 26256
rect 9692 26194 9720 26318
rect 9784 26246 9812 26438
rect 9600 26166 9720 26194
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9600 25906 9628 26166
rect 9784 26042 9812 26182
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 9588 25900 9640 25906
rect 9588 25842 9640 25848
rect 9772 25900 9824 25906
rect 9772 25842 9824 25848
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9588 24880 9640 24886
rect 9588 24822 9640 24828
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9508 23662 9536 24754
rect 9496 23656 9548 23662
rect 9600 23644 9628 24822
rect 9692 24410 9720 25230
rect 9784 24954 9812 25842
rect 9864 25492 9916 25498
rect 9864 25434 9916 25440
rect 9772 24948 9824 24954
rect 9772 24890 9824 24896
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9876 24206 9904 25434
rect 9864 24200 9916 24206
rect 9770 24168 9826 24177
rect 9864 24142 9916 24148
rect 9770 24103 9772 24112
rect 9824 24103 9826 24112
rect 9772 24074 9824 24080
rect 9600 23616 9720 23644
rect 9496 23598 9548 23604
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9404 22160 9456 22166
rect 9404 22102 9456 22108
rect 9312 21004 9364 21010
rect 9312 20946 9364 20952
rect 9312 20868 9364 20874
rect 9312 20810 9364 20816
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 9232 17678 9260 19314
rect 9324 19310 9352 20810
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9416 18986 9444 22102
rect 9508 22098 9536 23598
rect 9588 23520 9640 23526
rect 9588 23462 9640 23468
rect 9496 22092 9548 22098
rect 9496 22034 9548 22040
rect 9600 22030 9628 23462
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9600 21622 9628 21966
rect 9588 21616 9640 21622
rect 9588 21558 9640 21564
rect 9692 20890 9720 23616
rect 9864 23520 9916 23526
rect 9864 23462 9916 23468
rect 9876 23118 9904 23462
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 9968 22642 9996 31742
rect 10048 31136 10100 31142
rect 10048 31078 10100 31084
rect 10060 30734 10088 31078
rect 10048 30728 10100 30734
rect 10048 30670 10100 30676
rect 10048 28212 10100 28218
rect 10048 28154 10100 28160
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 10060 22094 10088 28154
rect 10152 26874 10180 31962
rect 10336 31346 10364 33050
rect 10416 33040 10468 33046
rect 10416 32982 10468 32988
rect 10428 32298 10456 32982
rect 10416 32292 10468 32298
rect 10416 32234 10468 32240
rect 10520 31346 10548 34886
rect 10612 34066 10640 35430
rect 10704 34610 10732 35498
rect 10796 35290 10824 35634
rect 10784 35284 10836 35290
rect 10784 35226 10836 35232
rect 10880 34844 11188 34864
rect 10880 34842 10886 34844
rect 10942 34842 10966 34844
rect 11022 34842 11046 34844
rect 11102 34842 11126 34844
rect 11182 34842 11188 34844
rect 10942 34790 10944 34842
rect 11124 34790 11126 34842
rect 10880 34788 10886 34790
rect 10942 34788 10966 34790
rect 11022 34788 11046 34790
rect 11102 34788 11126 34790
rect 11182 34788 11188 34790
rect 10880 34768 11188 34788
rect 10692 34604 10744 34610
rect 10692 34546 10744 34552
rect 11244 34604 11296 34610
rect 11244 34546 11296 34552
rect 11520 34604 11572 34610
rect 11520 34546 11572 34552
rect 10876 34400 10928 34406
rect 10876 34342 10928 34348
rect 10600 34060 10652 34066
rect 10600 34002 10652 34008
rect 10888 33998 10916 34342
rect 10692 33992 10744 33998
rect 10692 33934 10744 33940
rect 10876 33992 10928 33998
rect 10876 33934 10928 33940
rect 10704 33658 10732 33934
rect 11256 33862 11284 34546
rect 11244 33856 11296 33862
rect 11244 33798 11296 33804
rect 10880 33756 11188 33776
rect 10880 33754 10886 33756
rect 10942 33754 10966 33756
rect 11022 33754 11046 33756
rect 11102 33754 11126 33756
rect 11182 33754 11188 33756
rect 10942 33702 10944 33754
rect 11124 33702 11126 33754
rect 10880 33700 10886 33702
rect 10942 33700 10966 33702
rect 11022 33700 11046 33702
rect 11102 33700 11126 33702
rect 11182 33700 11188 33702
rect 10880 33680 11188 33700
rect 10692 33652 10744 33658
rect 10692 33594 10744 33600
rect 10704 33522 10732 33594
rect 10692 33516 10744 33522
rect 10692 33458 10744 33464
rect 10784 32972 10836 32978
rect 10784 32914 10836 32920
rect 10324 31340 10376 31346
rect 10324 31282 10376 31288
rect 10508 31340 10560 31346
rect 10508 31282 10560 31288
rect 10232 31272 10284 31278
rect 10232 31214 10284 31220
rect 10244 30054 10272 31214
rect 10692 31136 10744 31142
rect 10692 31078 10744 31084
rect 10324 30864 10376 30870
rect 10324 30806 10376 30812
rect 10232 30048 10284 30054
rect 10232 29990 10284 29996
rect 10336 28558 10364 30806
rect 10600 30796 10652 30802
rect 10600 30738 10652 30744
rect 10508 30592 10560 30598
rect 10508 30534 10560 30540
rect 10416 30252 10468 30258
rect 10416 30194 10468 30200
rect 10324 28552 10376 28558
rect 10324 28494 10376 28500
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 10244 27470 10272 28358
rect 10324 28076 10376 28082
rect 10324 28018 10376 28024
rect 10336 27538 10364 28018
rect 10324 27532 10376 27538
rect 10324 27474 10376 27480
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 10322 27432 10378 27441
rect 10322 27367 10378 27376
rect 10336 27130 10364 27367
rect 10324 27124 10376 27130
rect 10324 27066 10376 27072
rect 10230 27024 10286 27033
rect 10230 26959 10232 26968
rect 10284 26959 10286 26968
rect 10324 26988 10376 26994
rect 10232 26930 10284 26936
rect 10324 26930 10376 26936
rect 10152 26846 10272 26874
rect 10140 26308 10192 26314
rect 10140 26250 10192 26256
rect 10152 24206 10180 26250
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 9600 20862 9720 20890
rect 9968 22066 10088 22094
rect 9600 20618 9628 20862
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9508 20590 9628 20618
rect 9508 20330 9536 20590
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 9496 20324 9548 20330
rect 9496 20266 9548 20272
rect 9416 18958 9536 18986
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9324 18222 9352 18702
rect 9416 18290 9444 18770
rect 9508 18329 9536 18958
rect 9494 18320 9550 18329
rect 9404 18284 9456 18290
rect 9494 18255 9550 18264
rect 9404 18226 9456 18232
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9310 18048 9366 18057
rect 9310 17983 9366 17992
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9232 17338 9260 17614
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9140 17202 9260 17218
rect 9140 17196 9272 17202
rect 9140 17190 9220 17196
rect 9220 17138 9272 17144
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9140 16046 9168 16526
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 9140 15502 9168 15982
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9140 15026 9168 15438
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9140 14006 9168 14962
rect 9128 14000 9180 14006
rect 9126 13968 9128 13977
rect 9180 13968 9182 13977
rect 9126 13903 9182 13912
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9140 13462 9168 13670
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 8956 12406 9076 12434
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8864 8090 8892 10610
rect 8956 9586 8984 12406
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9048 9674 9076 12242
rect 9140 11014 9168 13398
rect 9232 12434 9260 17138
rect 9324 15706 9352 17983
rect 9416 17134 9444 18226
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9508 17610 9536 18090
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9508 17134 9536 17546
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9416 16658 9444 17070
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9508 16114 9536 17070
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9404 15972 9456 15978
rect 9404 15914 9456 15920
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9324 15570 9352 15642
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9416 15502 9444 15914
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9416 15162 9444 15438
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9508 14822 9536 15098
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9600 14634 9628 20470
rect 9692 20466 9720 20742
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9692 18714 9720 20402
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9876 19514 9904 19790
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9692 18686 9812 18714
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9692 17678 9720 18566
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9784 17202 9812 18686
rect 9876 18306 9904 19450
rect 9968 18426 9996 22066
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 10060 19922 10088 21286
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10152 20398 10180 20538
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 9876 18278 9996 18306
rect 9864 17604 9916 17610
rect 9864 17546 9916 17552
rect 9876 17338 9904 17546
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9968 16266 9996 18278
rect 10060 16998 10088 18906
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 9876 16238 9996 16266
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9508 14606 9628 14634
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9324 13734 9352 13874
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9232 12406 9352 12434
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 9232 11150 9260 12106
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9048 9646 9168 9674
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8956 8498 8984 8910
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8864 4146 8892 4558
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9048 3194 9076 4082
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9140 3058 9168 9646
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9232 8022 9260 8842
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 9232 7342 9260 7958
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9324 7154 9352 12406
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9416 11354 9444 11494
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9416 8786 9444 11086
rect 9508 10266 9536 14606
rect 9586 14104 9642 14113
rect 9586 14039 9588 14048
rect 9640 14039 9642 14048
rect 9588 14010 9640 14016
rect 9692 13938 9720 14894
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9600 13258 9628 13874
rect 9784 13870 9812 15574
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9508 8974 9536 9522
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9416 8758 9536 8786
rect 9232 6798 9260 7142
rect 9324 7126 9444 7154
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9324 4622 9352 6938
rect 9416 5302 9444 7126
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9324 4146 9352 4558
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9416 3534 9444 4966
rect 9508 4434 9536 8758
rect 9600 8022 9628 13194
rect 9692 12306 9720 13670
rect 9772 12844 9824 12850
rect 9876 12832 9904 16238
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9968 14822 9996 16118
rect 10060 15502 10088 16730
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9956 14544 10008 14550
rect 9956 14486 10008 14492
rect 9968 14006 9996 14486
rect 10060 14414 10088 15438
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 10060 13326 10088 14350
rect 10152 13734 10180 20334
rect 10244 20262 10272 26846
rect 10336 26586 10364 26930
rect 10324 26580 10376 26586
rect 10324 26522 10376 26528
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10336 24750 10364 25978
rect 10428 25498 10456 30194
rect 10520 29306 10548 30534
rect 10612 30190 10640 30738
rect 10704 30734 10732 31078
rect 10692 30728 10744 30734
rect 10692 30670 10744 30676
rect 10796 30308 10824 32914
rect 10880 32668 11188 32688
rect 10880 32666 10886 32668
rect 10942 32666 10966 32668
rect 11022 32666 11046 32668
rect 11102 32666 11126 32668
rect 11182 32666 11188 32668
rect 10942 32614 10944 32666
rect 11124 32614 11126 32666
rect 10880 32612 10886 32614
rect 10942 32612 10966 32614
rect 11022 32612 11046 32614
rect 11102 32612 11126 32614
rect 11182 32612 11188 32614
rect 10880 32592 11188 32612
rect 10876 32428 10928 32434
rect 10876 32370 10928 32376
rect 10888 32026 10916 32370
rect 10876 32020 10928 32026
rect 10876 31962 10928 31968
rect 11256 31958 11284 33798
rect 11532 33454 11560 34546
rect 11520 33448 11572 33454
rect 11520 33390 11572 33396
rect 11532 32502 11560 33390
rect 11900 32910 11928 36518
rect 12440 35284 12492 35290
rect 12440 35226 12492 35232
rect 12072 35012 12124 35018
rect 12072 34954 12124 34960
rect 12084 33114 12112 34954
rect 12452 34678 12480 35226
rect 12440 34672 12492 34678
rect 12440 34614 12492 34620
rect 12348 33516 12400 33522
rect 12348 33458 12400 33464
rect 12072 33108 12124 33114
rect 12072 33050 12124 33056
rect 11796 32904 11848 32910
rect 11796 32846 11848 32852
rect 11888 32904 11940 32910
rect 11888 32846 11940 32852
rect 12072 32904 12124 32910
rect 12072 32846 12124 32852
rect 11520 32496 11572 32502
rect 11520 32438 11572 32444
rect 11336 32360 11388 32366
rect 11336 32302 11388 32308
rect 11152 31952 11204 31958
rect 11152 31894 11204 31900
rect 11244 31952 11296 31958
rect 11244 31894 11296 31900
rect 11164 31754 11192 31894
rect 11348 31822 11376 32302
rect 11336 31816 11388 31822
rect 11336 31758 11388 31764
rect 11164 31726 11284 31754
rect 10880 31580 11188 31600
rect 10880 31578 10886 31580
rect 10942 31578 10966 31580
rect 11022 31578 11046 31580
rect 11102 31578 11126 31580
rect 11182 31578 11188 31580
rect 10942 31526 10944 31578
rect 11124 31526 11126 31578
rect 10880 31524 10886 31526
rect 10942 31524 10966 31526
rect 11022 31524 11046 31526
rect 11102 31524 11126 31526
rect 11182 31524 11188 31526
rect 10880 31504 11188 31524
rect 10880 30492 11188 30512
rect 10880 30490 10886 30492
rect 10942 30490 10966 30492
rect 11022 30490 11046 30492
rect 11102 30490 11126 30492
rect 11182 30490 11188 30492
rect 10942 30438 10944 30490
rect 11124 30438 11126 30490
rect 10880 30436 10886 30438
rect 10942 30436 10966 30438
rect 11022 30436 11046 30438
rect 11102 30436 11126 30438
rect 11182 30436 11188 30438
rect 10880 30416 11188 30436
rect 10876 30320 10928 30326
rect 10796 30280 10876 30308
rect 10876 30262 10928 30268
rect 10600 30184 10652 30190
rect 10600 30126 10652 30132
rect 10692 30184 10744 30190
rect 10692 30126 10744 30132
rect 10508 29300 10560 29306
rect 10508 29242 10560 29248
rect 10508 27396 10560 27402
rect 10508 27338 10560 27344
rect 10520 26994 10548 27338
rect 10508 26988 10560 26994
rect 10508 26930 10560 26936
rect 10506 26888 10562 26897
rect 10506 26823 10562 26832
rect 10520 26194 10548 26823
rect 10612 26382 10640 30126
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10520 26166 10640 26194
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 10508 25288 10560 25294
rect 10508 25230 10560 25236
rect 10520 24818 10548 25230
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 10324 24744 10376 24750
rect 10324 24686 10376 24692
rect 10428 22778 10456 24754
rect 10520 23798 10548 24754
rect 10612 23866 10640 26166
rect 10704 24682 10732 30126
rect 10880 29404 11188 29424
rect 10880 29402 10886 29404
rect 10942 29402 10966 29404
rect 11022 29402 11046 29404
rect 11102 29402 11126 29404
rect 11182 29402 11188 29404
rect 10942 29350 10944 29402
rect 11124 29350 11126 29402
rect 10880 29348 10886 29350
rect 10942 29348 10966 29350
rect 11022 29348 11046 29350
rect 11102 29348 11126 29350
rect 11182 29348 11188 29350
rect 10880 29328 11188 29348
rect 11060 29232 11112 29238
rect 11060 29174 11112 29180
rect 11072 28558 11100 29174
rect 10784 28552 10836 28558
rect 10784 28494 10836 28500
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 10796 27674 10824 28494
rect 10880 28316 11188 28336
rect 10880 28314 10886 28316
rect 10942 28314 10966 28316
rect 11022 28314 11046 28316
rect 11102 28314 11126 28316
rect 11182 28314 11188 28316
rect 10942 28262 10944 28314
rect 11124 28262 11126 28314
rect 10880 28260 10886 28262
rect 10942 28260 10966 28262
rect 11022 28260 11046 28262
rect 11102 28260 11126 28262
rect 11182 28260 11188 28262
rect 10880 28240 11188 28260
rect 10784 27668 10836 27674
rect 10784 27610 10836 27616
rect 10796 27554 10824 27610
rect 10796 27526 10916 27554
rect 10888 27470 10916 27526
rect 10784 27464 10836 27470
rect 10782 27432 10784 27441
rect 10876 27464 10928 27470
rect 10836 27432 10838 27441
rect 10876 27406 10928 27412
rect 11256 27418 11284 31726
rect 11348 29646 11376 31758
rect 11428 30728 11480 30734
rect 11428 30670 11480 30676
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 11348 28150 11376 29582
rect 11440 28762 11468 30670
rect 11520 30592 11572 30598
rect 11520 30534 11572 30540
rect 11532 30258 11560 30534
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 11428 28756 11480 28762
rect 11428 28698 11480 28704
rect 11336 28144 11388 28150
rect 11336 28086 11388 28092
rect 11348 27538 11376 28086
rect 11336 27532 11388 27538
rect 11336 27474 11388 27480
rect 11256 27390 11376 27418
rect 10782 27367 10838 27376
rect 10784 27328 10836 27334
rect 10784 27270 10836 27276
rect 10796 26994 10824 27270
rect 10880 27228 11188 27248
rect 10880 27226 10886 27228
rect 10942 27226 10966 27228
rect 11022 27226 11046 27228
rect 11102 27226 11126 27228
rect 11182 27226 11188 27228
rect 10942 27174 10944 27226
rect 11124 27174 11126 27226
rect 10880 27172 10886 27174
rect 10942 27172 10966 27174
rect 11022 27172 11046 27174
rect 11102 27172 11126 27174
rect 11182 27172 11188 27174
rect 10880 27152 11188 27172
rect 10784 26988 10836 26994
rect 10784 26930 10836 26936
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 10796 24818 10824 26318
rect 10880 26140 11188 26160
rect 10880 26138 10886 26140
rect 10942 26138 10966 26140
rect 11022 26138 11046 26140
rect 11102 26138 11126 26140
rect 11182 26138 11188 26140
rect 10942 26086 10944 26138
rect 11124 26086 11126 26138
rect 10880 26084 10886 26086
rect 10942 26084 10966 26086
rect 11022 26084 11046 26086
rect 11102 26084 11126 26086
rect 11182 26084 11188 26086
rect 10880 26064 11188 26084
rect 11244 25152 11296 25158
rect 11244 25094 11296 25100
rect 10880 25052 11188 25072
rect 10880 25050 10886 25052
rect 10942 25050 10966 25052
rect 11022 25050 11046 25052
rect 11102 25050 11126 25052
rect 11182 25050 11188 25052
rect 10942 24998 10944 25050
rect 11124 24998 11126 25050
rect 10880 24996 10886 24998
rect 10942 24996 10966 24998
rect 11022 24996 11046 24998
rect 11102 24996 11126 24998
rect 11182 24996 11188 24998
rect 10880 24976 11188 24996
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10690 24168 10746 24177
rect 10690 24103 10692 24112
rect 10744 24103 10746 24112
rect 10692 24074 10744 24080
rect 10600 23860 10652 23866
rect 10600 23802 10652 23808
rect 10508 23792 10560 23798
rect 10508 23734 10560 23740
rect 10612 23662 10640 23802
rect 10796 23712 10824 24754
rect 11256 24342 11284 25094
rect 11244 24336 11296 24342
rect 11244 24278 11296 24284
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 10880 23964 11188 23984
rect 10880 23962 10886 23964
rect 10942 23962 10966 23964
rect 11022 23962 11046 23964
rect 11102 23962 11126 23964
rect 11182 23962 11188 23964
rect 10942 23910 10944 23962
rect 11124 23910 11126 23962
rect 10880 23908 10886 23910
rect 10942 23908 10966 23910
rect 11022 23908 11046 23910
rect 11102 23908 11126 23910
rect 11182 23908 11188 23910
rect 10880 23888 11188 23908
rect 10876 23724 10928 23730
rect 10796 23684 10876 23712
rect 10876 23666 10928 23672
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10416 22772 10468 22778
rect 10468 22732 10548 22760
rect 10416 22714 10468 22720
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10336 21026 10364 21966
rect 10428 21622 10456 22578
rect 10520 22094 10548 22732
rect 10692 22636 10744 22642
rect 10796 22624 10824 23462
rect 10888 23322 10916 23666
rect 10876 23316 10928 23322
rect 10876 23258 10928 23264
rect 10880 22876 11188 22896
rect 10880 22874 10886 22876
rect 10942 22874 10966 22876
rect 11022 22874 11046 22876
rect 11102 22874 11126 22876
rect 11182 22874 11188 22876
rect 10942 22822 10944 22874
rect 11124 22822 11126 22874
rect 10880 22820 10886 22822
rect 10942 22820 10966 22822
rect 11022 22820 11046 22822
rect 11102 22820 11126 22822
rect 11182 22820 11188 22822
rect 10880 22800 11188 22820
rect 11152 22704 11204 22710
rect 11152 22646 11204 22652
rect 10876 22636 10928 22642
rect 10796 22596 10876 22624
rect 10692 22578 10744 22584
rect 10876 22578 10928 22584
rect 10704 22234 10732 22578
rect 11164 22420 11192 22646
rect 11256 22522 11284 24142
rect 11348 22710 11376 27390
rect 11428 27396 11480 27402
rect 11428 27338 11480 27344
rect 11440 27130 11468 27338
rect 11428 27124 11480 27130
rect 11428 27066 11480 27072
rect 11428 25832 11480 25838
rect 11428 25774 11480 25780
rect 11440 24206 11468 25774
rect 11532 24800 11560 30194
rect 11704 29844 11756 29850
rect 11704 29786 11756 29792
rect 11612 29640 11664 29646
rect 11612 29582 11664 29588
rect 11624 29306 11652 29582
rect 11612 29300 11664 29306
rect 11612 29242 11664 29248
rect 11716 28082 11744 29786
rect 11808 29782 11836 32846
rect 12084 32502 12112 32846
rect 12072 32496 12124 32502
rect 12072 32438 12124 32444
rect 12256 32428 12308 32434
rect 12256 32370 12308 32376
rect 12164 32224 12216 32230
rect 12164 32166 12216 32172
rect 11888 31748 11940 31754
rect 11888 31690 11940 31696
rect 11900 30938 11928 31690
rect 11888 30932 11940 30938
rect 11888 30874 11940 30880
rect 11888 30796 11940 30802
rect 11888 30738 11940 30744
rect 11900 30190 11928 30738
rect 12176 30258 12204 32166
rect 12268 30326 12296 32370
rect 12256 30320 12308 30326
rect 12256 30262 12308 30268
rect 12164 30252 12216 30258
rect 12164 30194 12216 30200
rect 11888 30184 11940 30190
rect 11888 30126 11940 30132
rect 11796 29776 11848 29782
rect 11796 29718 11848 29724
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11808 28558 11836 29106
rect 11900 28626 11928 30126
rect 12360 29850 12388 33458
rect 12452 33454 12480 34614
rect 12532 34128 12584 34134
rect 12532 34070 12584 34076
rect 12544 33998 12572 34070
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 12440 33448 12492 33454
rect 12440 33390 12492 33396
rect 12544 32842 12572 33934
rect 12532 32836 12584 32842
rect 12532 32778 12584 32784
rect 12532 32496 12584 32502
rect 12532 32438 12584 32444
rect 12544 31482 12572 32438
rect 12636 31958 12664 37266
rect 12728 37262 12756 37606
rect 13096 37398 13124 37810
rect 13188 37466 13216 38286
rect 14016 37874 14044 38830
rect 14004 37868 14056 37874
rect 14004 37810 14056 37816
rect 13176 37460 13228 37466
rect 13176 37402 13228 37408
rect 13084 37392 13136 37398
rect 13084 37334 13136 37340
rect 12716 37256 12768 37262
rect 12716 37198 12768 37204
rect 13096 37194 13124 37334
rect 13084 37188 13136 37194
rect 13084 37130 13136 37136
rect 13096 36854 13124 37130
rect 13084 36848 13136 36854
rect 13084 36790 13136 36796
rect 13096 35290 13124 36790
rect 13268 36780 13320 36786
rect 13268 36722 13320 36728
rect 13280 36038 13308 36722
rect 14016 36378 14044 37810
rect 14108 37262 14136 39306
rect 14292 38962 14320 39442
rect 14476 39370 14504 41074
rect 14924 40996 14976 41002
rect 14924 40938 14976 40944
rect 14740 40928 14792 40934
rect 14740 40870 14792 40876
rect 14752 40594 14780 40870
rect 14740 40588 14792 40594
rect 14740 40530 14792 40536
rect 14832 40384 14884 40390
rect 14832 40326 14884 40332
rect 14844 40186 14872 40326
rect 14832 40180 14884 40186
rect 14832 40122 14884 40128
rect 14832 39432 14884 39438
rect 14832 39374 14884 39380
rect 14464 39364 14516 39370
rect 14464 39306 14516 39312
rect 14280 38956 14332 38962
rect 14280 38898 14332 38904
rect 14844 38894 14872 39374
rect 14832 38888 14884 38894
rect 14832 38830 14884 38836
rect 14844 38554 14872 38830
rect 14936 38758 14964 40938
rect 15580 40118 15608 41074
rect 15568 40112 15620 40118
rect 15568 40054 15620 40060
rect 15660 40044 15712 40050
rect 15660 39986 15712 39992
rect 15672 39846 15700 39986
rect 15764 39914 15792 41550
rect 16304 41472 16356 41478
rect 16304 41414 16356 41420
rect 16316 41138 16344 41414
rect 16304 41132 16356 41138
rect 16304 41074 16356 41080
rect 17408 41132 17460 41138
rect 17408 41074 17460 41080
rect 15846 40828 16154 40848
rect 15846 40826 15852 40828
rect 15908 40826 15932 40828
rect 15988 40826 16012 40828
rect 16068 40826 16092 40828
rect 16148 40826 16154 40828
rect 15908 40774 15910 40826
rect 16090 40774 16092 40826
rect 15846 40772 15852 40774
rect 15908 40772 15932 40774
rect 15988 40772 16012 40774
rect 16068 40772 16092 40774
rect 16148 40772 16154 40774
rect 15846 40752 16154 40772
rect 16316 40526 16344 41074
rect 16488 40928 16540 40934
rect 16488 40870 16540 40876
rect 16672 40928 16724 40934
rect 16672 40870 16724 40876
rect 17040 40928 17092 40934
rect 17040 40870 17092 40876
rect 16304 40520 16356 40526
rect 16304 40462 16356 40468
rect 16500 40118 16528 40870
rect 16684 40594 16712 40870
rect 16856 40656 16908 40662
rect 16856 40598 16908 40604
rect 16672 40588 16724 40594
rect 16672 40530 16724 40536
rect 16764 40588 16816 40594
rect 16764 40530 16816 40536
rect 16580 40180 16632 40186
rect 16580 40122 16632 40128
rect 16488 40112 16540 40118
rect 16488 40054 16540 40060
rect 16212 39976 16264 39982
rect 16212 39918 16264 39924
rect 15752 39908 15804 39914
rect 15752 39850 15804 39856
rect 15660 39840 15712 39846
rect 15660 39782 15712 39788
rect 15672 39642 15700 39782
rect 15846 39740 16154 39760
rect 15846 39738 15852 39740
rect 15908 39738 15932 39740
rect 15988 39738 16012 39740
rect 16068 39738 16092 39740
rect 16148 39738 16154 39740
rect 15908 39686 15910 39738
rect 16090 39686 16092 39738
rect 15846 39684 15852 39686
rect 15908 39684 15932 39686
rect 15988 39684 16012 39686
rect 16068 39684 16092 39686
rect 16148 39684 16154 39686
rect 15846 39664 16154 39684
rect 15660 39636 15712 39642
rect 15660 39578 15712 39584
rect 15016 39500 15068 39506
rect 15016 39442 15068 39448
rect 15384 39500 15436 39506
rect 15384 39442 15436 39448
rect 15028 39302 15056 39442
rect 15396 39386 15424 39442
rect 15304 39358 15424 39386
rect 15568 39432 15620 39438
rect 15568 39374 15620 39380
rect 15016 39296 15068 39302
rect 15016 39238 15068 39244
rect 15028 38842 15056 39238
rect 15304 39098 15332 39358
rect 15580 39302 15608 39374
rect 15568 39296 15620 39302
rect 15568 39238 15620 39244
rect 15672 39114 15700 39578
rect 15844 39432 15896 39438
rect 15844 39374 15896 39380
rect 15292 39092 15344 39098
rect 15292 39034 15344 39040
rect 15580 39086 15700 39114
rect 15304 38962 15332 39034
rect 15292 38956 15344 38962
rect 15292 38898 15344 38904
rect 15200 38888 15252 38894
rect 15028 38836 15200 38842
rect 15028 38830 15252 38836
rect 15028 38814 15240 38830
rect 14924 38752 14976 38758
rect 14924 38694 14976 38700
rect 14832 38548 14884 38554
rect 14832 38490 14884 38496
rect 14936 38026 14964 38694
rect 14936 37998 15056 38026
rect 15120 38010 15148 38814
rect 14924 37868 14976 37874
rect 14924 37810 14976 37816
rect 14280 37800 14332 37806
rect 14280 37742 14332 37748
rect 14188 37664 14240 37670
rect 14188 37606 14240 37612
rect 14200 37466 14228 37606
rect 14188 37460 14240 37466
rect 14188 37402 14240 37408
rect 14096 37256 14148 37262
rect 14096 37198 14148 37204
rect 14108 36718 14136 37198
rect 14200 36786 14228 37402
rect 14188 36780 14240 36786
rect 14188 36722 14240 36728
rect 14096 36712 14148 36718
rect 14096 36654 14148 36660
rect 14004 36372 14056 36378
rect 14004 36314 14056 36320
rect 14200 36174 14228 36722
rect 14292 36666 14320 37742
rect 14936 37618 14964 37810
rect 14844 37590 14964 37618
rect 14556 37188 14608 37194
rect 14556 37130 14608 37136
rect 14568 36786 14596 37130
rect 14844 36786 14872 37590
rect 14556 36780 14608 36786
rect 14556 36722 14608 36728
rect 14832 36780 14884 36786
rect 14832 36722 14884 36728
rect 14648 36712 14700 36718
rect 14292 36650 14412 36666
rect 14648 36654 14700 36660
rect 14292 36644 14424 36650
rect 14292 36638 14372 36644
rect 14292 36174 14320 36638
rect 14372 36586 14424 36592
rect 14188 36168 14240 36174
rect 14188 36110 14240 36116
rect 14280 36168 14332 36174
rect 14280 36110 14332 36116
rect 13268 36032 13320 36038
rect 13268 35974 13320 35980
rect 14464 35624 14516 35630
rect 14464 35566 14516 35572
rect 13084 35284 13136 35290
rect 13084 35226 13136 35232
rect 13728 35148 13780 35154
rect 13728 35090 13780 35096
rect 13740 34678 13768 35090
rect 14372 35080 14424 35086
rect 14372 35022 14424 35028
rect 13728 34672 13780 34678
rect 13728 34614 13780 34620
rect 14096 34604 14148 34610
rect 14096 34546 14148 34552
rect 14108 34134 14136 34546
rect 14384 34134 14412 35022
rect 14476 34406 14504 35566
rect 14660 35086 14688 36654
rect 14648 35080 14700 35086
rect 14648 35022 14700 35028
rect 14660 34542 14688 35022
rect 14648 34536 14700 34542
rect 14648 34478 14700 34484
rect 14464 34400 14516 34406
rect 14464 34342 14516 34348
rect 14096 34128 14148 34134
rect 14096 34070 14148 34076
rect 14372 34128 14424 34134
rect 14372 34070 14424 34076
rect 13452 34060 13504 34066
rect 13452 34002 13504 34008
rect 12992 33992 13044 33998
rect 12992 33934 13044 33940
rect 12716 33924 12768 33930
rect 12716 33866 12768 33872
rect 12808 33924 12860 33930
rect 12808 33866 12860 33872
rect 12728 33658 12756 33866
rect 12716 33652 12768 33658
rect 12716 33594 12768 33600
rect 12820 33522 12848 33866
rect 12808 33516 12860 33522
rect 12808 33458 12860 33464
rect 12900 33448 12952 33454
rect 12900 33390 12952 33396
rect 12912 32434 12940 33390
rect 13004 32978 13032 33934
rect 13464 33862 13492 34002
rect 14476 33930 14504 34342
rect 14372 33924 14424 33930
rect 14372 33866 14424 33872
rect 14464 33924 14516 33930
rect 14464 33866 14516 33872
rect 13176 33856 13228 33862
rect 13176 33798 13228 33804
rect 13452 33856 13504 33862
rect 13452 33798 13504 33804
rect 13188 33522 13216 33798
rect 13464 33522 13492 33798
rect 14384 33590 14412 33866
rect 14372 33584 14424 33590
rect 14372 33526 14424 33532
rect 13176 33516 13228 33522
rect 13176 33458 13228 33464
rect 13452 33516 13504 33522
rect 13452 33458 13504 33464
rect 12992 32972 13044 32978
rect 12992 32914 13044 32920
rect 12992 32836 13044 32842
rect 12992 32778 13044 32784
rect 12900 32428 12952 32434
rect 12900 32370 12952 32376
rect 12912 31958 12940 32370
rect 12624 31952 12676 31958
rect 12624 31894 12676 31900
rect 12900 31952 12952 31958
rect 12900 31894 12952 31900
rect 12532 31476 12584 31482
rect 12532 31418 12584 31424
rect 12440 31340 12492 31346
rect 12440 31282 12492 31288
rect 12452 30326 12480 31282
rect 12636 30734 12664 31894
rect 12900 31476 12952 31482
rect 12900 31418 12952 31424
rect 12716 31408 12768 31414
rect 12716 31350 12768 31356
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 12440 30320 12492 30326
rect 12440 30262 12492 30268
rect 12348 29844 12400 29850
rect 12348 29786 12400 29792
rect 12164 29776 12216 29782
rect 12164 29718 12216 29724
rect 11888 28620 11940 28626
rect 11888 28562 11940 28568
rect 11796 28552 11848 28558
rect 11796 28494 11848 28500
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 11610 26752 11666 26761
rect 11610 26687 11666 26696
rect 11624 26364 11652 26687
rect 11716 26518 11744 28018
rect 11808 28014 11836 28494
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 11900 27554 11928 28562
rect 11980 28552 12032 28558
rect 11980 28494 12032 28500
rect 11992 27674 12020 28494
rect 12176 28490 12204 29718
rect 12728 29714 12756 31350
rect 12912 31346 12940 31418
rect 13004 31346 13032 32778
rect 13464 31482 13492 33458
rect 13912 32496 13964 32502
rect 13912 32438 13964 32444
rect 13820 31748 13872 31754
rect 13820 31690 13872 31696
rect 13832 31482 13860 31690
rect 13452 31476 13504 31482
rect 13452 31418 13504 31424
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 12992 31340 13044 31346
rect 12992 31282 13044 31288
rect 13268 31340 13320 31346
rect 13268 31282 13320 31288
rect 12808 30796 12860 30802
rect 12808 30738 12860 30744
rect 12820 30190 12848 30738
rect 12808 30184 12860 30190
rect 12808 30126 12860 30132
rect 12716 29708 12768 29714
rect 12716 29650 12768 29656
rect 12728 29238 12756 29650
rect 12820 29306 12848 30126
rect 12808 29300 12860 29306
rect 12808 29242 12860 29248
rect 12716 29232 12768 29238
rect 12716 29174 12768 29180
rect 12348 29028 12400 29034
rect 12348 28970 12400 28976
rect 12256 28756 12308 28762
rect 12256 28698 12308 28704
rect 12164 28484 12216 28490
rect 12164 28426 12216 28432
rect 12072 27940 12124 27946
rect 12072 27882 12124 27888
rect 11980 27668 12032 27674
rect 11980 27610 12032 27616
rect 11900 27526 12020 27554
rect 11796 27124 11848 27130
rect 11796 27066 11848 27072
rect 11704 26512 11756 26518
rect 11704 26454 11756 26460
rect 11704 26376 11756 26382
rect 11624 26336 11704 26364
rect 11704 26318 11756 26324
rect 11716 25906 11744 26318
rect 11808 26246 11836 27066
rect 11796 26240 11848 26246
rect 11796 26182 11848 26188
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11612 24812 11664 24818
rect 11532 24772 11612 24800
rect 11612 24754 11664 24760
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11428 23724 11480 23730
rect 11532 23712 11560 24142
rect 11480 23684 11560 23712
rect 11428 23666 11480 23672
rect 11440 22778 11468 23666
rect 11520 23112 11572 23118
rect 11520 23054 11572 23060
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11336 22704 11388 22710
rect 11336 22646 11388 22652
rect 11428 22636 11480 22642
rect 11532 22624 11560 23054
rect 11480 22596 11560 22624
rect 11428 22578 11480 22584
rect 11256 22494 11468 22522
rect 11532 22506 11560 22596
rect 11164 22392 11376 22420
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 10520 22066 10824 22094
rect 10796 22030 10824 22066
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 10416 21616 10468 21622
rect 10416 21558 10468 21564
rect 10428 21146 10456 21558
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10336 20998 10548 21026
rect 10232 20256 10284 20262
rect 10232 20198 10284 20204
rect 10244 16590 10272 20198
rect 10520 20058 10548 20998
rect 10600 20868 10652 20874
rect 10600 20810 10652 20816
rect 10612 20466 10640 20810
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10508 20052 10560 20058
rect 10508 19994 10560 20000
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10336 19378 10364 19790
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10428 19378 10456 19450
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10336 18630 10364 19314
rect 10520 19224 10548 19994
rect 10428 19196 10548 19224
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10336 13734 10364 16934
rect 10428 15910 10456 19196
rect 10612 18766 10640 20402
rect 10704 19802 10732 21490
rect 10796 19922 10824 21966
rect 10880 21788 11188 21808
rect 10880 21786 10886 21788
rect 10942 21786 10966 21788
rect 11022 21786 11046 21788
rect 11102 21786 11126 21788
rect 11182 21786 11188 21788
rect 10942 21734 10944 21786
rect 11124 21734 11126 21786
rect 10880 21732 10886 21734
rect 10942 21732 10966 21734
rect 11022 21732 11046 21734
rect 11102 21732 11126 21734
rect 11182 21732 11188 21734
rect 10880 21712 11188 21732
rect 11256 21418 11284 21966
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 10880 20700 11188 20720
rect 10880 20698 10886 20700
rect 10942 20698 10966 20700
rect 11022 20698 11046 20700
rect 11102 20698 11126 20700
rect 11182 20698 11188 20700
rect 10942 20646 10944 20698
rect 11124 20646 11126 20698
rect 10880 20644 10886 20646
rect 10942 20644 10966 20646
rect 11022 20644 11046 20646
rect 11102 20644 11126 20646
rect 11182 20644 11188 20646
rect 10880 20624 11188 20644
rect 11256 20466 11284 21354
rect 11348 21146 11376 22392
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11336 20868 11388 20874
rect 11336 20810 11388 20816
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 11072 19802 11100 20334
rect 10704 19774 11100 19802
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10508 18624 10560 18630
rect 10692 18624 10744 18630
rect 10560 18584 10640 18612
rect 10508 18566 10560 18572
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10140 13728 10192 13734
rect 10324 13728 10376 13734
rect 10140 13670 10192 13676
rect 10244 13688 10324 13716
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 9824 12804 9904 12832
rect 9772 12786 9824 12792
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 11558 9720 12106
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9692 9994 9720 10406
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9692 9178 9720 9454
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9692 7478 9720 8978
rect 9784 7546 9812 12786
rect 10060 11830 10088 13262
rect 10244 12374 10272 13688
rect 10324 13670 10376 13676
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9968 11082 9996 11630
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9968 10810 9996 11018
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10060 10130 10088 11766
rect 10152 11762 10180 12038
rect 10244 11801 10272 12310
rect 10336 12238 10364 12718
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10230 11792 10286 11801
rect 10140 11756 10192 11762
rect 10230 11727 10286 11736
rect 10324 11756 10376 11762
rect 10140 11698 10192 11704
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10152 10674 10180 10746
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10244 10606 10272 11727
rect 10324 11698 10376 11704
rect 10336 11257 10364 11698
rect 10322 11248 10378 11257
rect 10322 11183 10378 11192
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10046 9616 10102 9625
rect 10046 9551 10048 9560
rect 10100 9551 10102 9560
rect 10048 9522 10100 9528
rect 10152 8974 10180 10474
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10244 9178 10272 9862
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10244 9042 10272 9114
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10152 8430 10180 8910
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10140 7880 10192 7886
rect 10244 7868 10272 8978
rect 10336 8634 10364 10610
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10192 7840 10272 7868
rect 10140 7822 10192 7828
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9692 6322 9720 7414
rect 10336 7410 10364 8366
rect 10428 8294 10456 15846
rect 10520 14804 10548 18022
rect 10612 14906 10640 18584
rect 10692 18566 10744 18572
rect 10704 18086 10732 18566
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10796 16182 10824 19774
rect 10880 19612 11188 19632
rect 10880 19610 10886 19612
rect 10942 19610 10966 19612
rect 11022 19610 11046 19612
rect 11102 19610 11126 19612
rect 11182 19610 11188 19612
rect 10942 19558 10944 19610
rect 11124 19558 11126 19610
rect 10880 19556 10886 19558
rect 10942 19556 10966 19558
rect 11022 19556 11046 19558
rect 11102 19556 11126 19558
rect 11182 19556 11188 19558
rect 10880 19536 11188 19556
rect 11244 18624 11296 18630
rect 11348 18612 11376 20810
rect 11440 18834 11468 22494
rect 11520 22500 11572 22506
rect 11520 22442 11572 22448
rect 11532 21486 11560 22442
rect 11624 22030 11652 24754
rect 11716 24206 11744 25842
rect 11888 25764 11940 25770
rect 11888 25706 11940 25712
rect 11900 25226 11928 25706
rect 11796 25220 11848 25226
rect 11796 25162 11848 25168
rect 11888 25220 11940 25226
rect 11888 25162 11940 25168
rect 11808 24954 11836 25162
rect 11796 24948 11848 24954
rect 11796 24890 11848 24896
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11900 23798 11928 25162
rect 11992 24750 12020 27526
rect 12084 26586 12112 27882
rect 12072 26580 12124 26586
rect 12072 26522 12124 26528
rect 12084 26382 12112 26522
rect 12072 26376 12124 26382
rect 12072 26318 12124 26324
rect 11980 24744 12032 24750
rect 11980 24686 12032 24692
rect 11888 23792 11940 23798
rect 11888 23734 11940 23740
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 11808 22094 11836 23666
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11900 22098 11928 22646
rect 11716 22066 11836 22094
rect 11888 22092 11940 22098
rect 11612 22024 11664 22030
rect 11612 21966 11664 21972
rect 11520 21480 11572 21486
rect 11520 21422 11572 21428
rect 11532 19922 11560 21422
rect 11716 21298 11744 22066
rect 11888 22034 11940 22040
rect 11992 22030 12020 24686
rect 12084 24682 12112 26318
rect 12072 24676 12124 24682
rect 12072 24618 12124 24624
rect 12084 22778 12112 24618
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 12176 22574 12204 28426
rect 12268 25906 12296 28698
rect 12360 26926 12388 28970
rect 12912 28694 12940 31282
rect 13004 30734 13032 31282
rect 13084 31272 13136 31278
rect 13084 31214 13136 31220
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 13004 30394 13032 30670
rect 12992 30388 13044 30394
rect 12992 30330 13044 30336
rect 13096 30258 13124 31214
rect 13280 30870 13308 31282
rect 13268 30864 13320 30870
rect 13268 30806 13320 30812
rect 13360 30320 13412 30326
rect 13360 30262 13412 30268
rect 13084 30252 13136 30258
rect 13084 30194 13136 30200
rect 12900 28688 12952 28694
rect 12900 28630 12952 28636
rect 12532 28620 12584 28626
rect 12532 28562 12584 28568
rect 12544 28150 12572 28562
rect 13176 28416 13228 28422
rect 13176 28358 13228 28364
rect 12532 28144 12584 28150
rect 12532 28086 12584 28092
rect 13188 28082 13216 28358
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 12532 28008 12584 28014
rect 12532 27950 12584 27956
rect 12348 26920 12400 26926
rect 12348 26862 12400 26868
rect 12360 26246 12388 26862
rect 12440 26852 12492 26858
rect 12440 26794 12492 26800
rect 12348 26240 12400 26246
rect 12348 26182 12400 26188
rect 12256 25900 12308 25906
rect 12256 25842 12308 25848
rect 12268 24342 12296 25842
rect 12360 25838 12388 26182
rect 12348 25832 12400 25838
rect 12348 25774 12400 25780
rect 12256 24336 12308 24342
rect 12256 24278 12308 24284
rect 12268 23798 12296 24278
rect 12360 24206 12388 25774
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 12256 23656 12308 23662
rect 12360 23644 12388 24142
rect 12308 23616 12388 23644
rect 12256 23598 12308 23604
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11716 21270 11836 21298
rect 11808 20466 11836 21270
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11992 20398 12020 21966
rect 12268 21622 12296 22374
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 12268 19854 12296 20198
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12452 19514 12480 26794
rect 12544 23644 12572 27950
rect 12636 26994 12664 28018
rect 13372 27062 13400 30262
rect 13452 30184 13504 30190
rect 13452 30126 13504 30132
rect 13464 29170 13492 30126
rect 13636 29844 13688 29850
rect 13636 29786 13688 29792
rect 13648 29238 13676 29786
rect 13636 29232 13688 29238
rect 13636 29174 13688 29180
rect 13452 29164 13504 29170
rect 13452 29106 13504 29112
rect 13728 29164 13780 29170
rect 13728 29106 13780 29112
rect 13464 28626 13492 29106
rect 13452 28620 13504 28626
rect 13452 28562 13504 28568
rect 13544 28552 13596 28558
rect 13544 28494 13596 28500
rect 13556 28082 13584 28494
rect 13544 28076 13596 28082
rect 13544 28018 13596 28024
rect 13740 27130 13768 29106
rect 13728 27124 13780 27130
rect 13728 27066 13780 27072
rect 13360 27056 13412 27062
rect 13360 26998 13412 27004
rect 12624 26988 12676 26994
rect 12624 26930 12676 26936
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 12728 26586 12756 26930
rect 12716 26580 12768 26586
rect 12716 26522 12768 26528
rect 13372 25974 13400 26998
rect 13360 25968 13412 25974
rect 13360 25910 13412 25916
rect 12900 25900 12952 25906
rect 12900 25842 12952 25848
rect 12624 25424 12676 25430
rect 12624 25366 12676 25372
rect 12636 24818 12664 25366
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12624 24812 12676 24818
rect 12624 24754 12676 24760
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12636 23798 12664 24006
rect 12624 23792 12676 23798
rect 12624 23734 12676 23740
rect 12728 23730 12756 25230
rect 12912 24954 12940 25842
rect 12900 24948 12952 24954
rect 12900 24890 12952 24896
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 13096 24206 13124 24686
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13556 23730 13584 24142
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 12544 23616 12664 23644
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12544 23050 12572 23462
rect 12532 23044 12584 23050
rect 12532 22986 12584 22992
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 12544 22098 12572 22646
rect 12532 22092 12584 22098
rect 12532 22034 12584 22040
rect 12636 21078 12664 23616
rect 12728 22642 12756 23666
rect 13556 23322 13584 23666
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12820 21690 12848 22714
rect 13728 22432 13780 22438
rect 13728 22374 13780 22380
rect 13740 22030 13768 22374
rect 13924 22094 13952 32438
rect 14660 32230 14688 34478
rect 14648 32224 14700 32230
rect 14648 32166 14700 32172
rect 14740 32224 14792 32230
rect 14844 32212 14872 36722
rect 15028 36174 15056 37998
rect 15108 38004 15160 38010
rect 15108 37946 15160 37952
rect 15120 37466 15148 37946
rect 15108 37460 15160 37466
rect 15108 37402 15160 37408
rect 15580 37330 15608 39086
rect 15856 38894 15884 39374
rect 16120 39296 16172 39302
rect 16120 39238 16172 39244
rect 16132 39098 16160 39238
rect 16120 39092 16172 39098
rect 16120 39034 16172 39040
rect 16224 38894 16252 39918
rect 15844 38888 15896 38894
rect 15844 38830 15896 38836
rect 16212 38888 16264 38894
rect 16212 38830 16264 38836
rect 15846 38652 16154 38672
rect 15846 38650 15852 38652
rect 15908 38650 15932 38652
rect 15988 38650 16012 38652
rect 16068 38650 16092 38652
rect 16148 38650 16154 38652
rect 15908 38598 15910 38650
rect 16090 38598 16092 38650
rect 15846 38596 15852 38598
rect 15908 38596 15932 38598
rect 15988 38596 16012 38598
rect 16068 38596 16092 38598
rect 16148 38596 16154 38598
rect 15846 38576 16154 38596
rect 15846 37564 16154 37584
rect 15846 37562 15852 37564
rect 15908 37562 15932 37564
rect 15988 37562 16012 37564
rect 16068 37562 16092 37564
rect 16148 37562 16154 37564
rect 15908 37510 15910 37562
rect 16090 37510 16092 37562
rect 15846 37508 15852 37510
rect 15908 37508 15932 37510
rect 15988 37508 16012 37510
rect 16068 37508 16092 37510
rect 16148 37508 16154 37510
rect 15846 37488 16154 37508
rect 15200 37324 15252 37330
rect 15200 37266 15252 37272
rect 15568 37324 15620 37330
rect 15568 37266 15620 37272
rect 15108 37256 15160 37262
rect 15108 37198 15160 37204
rect 15120 36922 15148 37198
rect 15108 36916 15160 36922
rect 15108 36858 15160 36864
rect 15120 36242 15148 36858
rect 15212 36582 15240 37266
rect 15292 37120 15344 37126
rect 15292 37062 15344 37068
rect 15304 36718 15332 37062
rect 15292 36712 15344 36718
rect 15292 36654 15344 36660
rect 15200 36576 15252 36582
rect 15200 36518 15252 36524
rect 15212 36310 15240 36518
rect 15200 36304 15252 36310
rect 15200 36246 15252 36252
rect 15108 36236 15160 36242
rect 15108 36178 15160 36184
rect 15016 36168 15068 36174
rect 15016 36110 15068 36116
rect 15028 34474 15056 36110
rect 15212 35170 15240 36246
rect 15580 35290 15608 37266
rect 16120 37256 16172 37262
rect 16224 37210 16252 38830
rect 16304 37460 16356 37466
rect 16304 37402 16356 37408
rect 16316 37330 16344 37402
rect 16304 37324 16356 37330
rect 16304 37266 16356 37272
rect 16172 37204 16252 37210
rect 16120 37198 16252 37204
rect 16132 37182 16252 37198
rect 16224 37126 16252 37182
rect 16212 37120 16264 37126
rect 16212 37062 16264 37068
rect 15846 36476 16154 36496
rect 15846 36474 15852 36476
rect 15908 36474 15932 36476
rect 15988 36474 16012 36476
rect 16068 36474 16092 36476
rect 16148 36474 16154 36476
rect 15908 36422 15910 36474
rect 16090 36422 16092 36474
rect 15846 36420 15852 36422
rect 15908 36420 15932 36422
rect 15988 36420 16012 36422
rect 16068 36420 16092 36422
rect 16148 36420 16154 36422
rect 15846 36400 16154 36420
rect 16224 36258 16252 37062
rect 16132 36230 16252 36258
rect 16316 36242 16344 37266
rect 16304 36236 16356 36242
rect 16132 36174 16160 36230
rect 16304 36178 16356 36184
rect 16120 36168 16172 36174
rect 15764 36116 16120 36122
rect 15764 36110 16172 36116
rect 15764 36094 16160 36110
rect 15568 35284 15620 35290
rect 15568 35226 15620 35232
rect 15212 35154 15332 35170
rect 15212 35148 15344 35154
rect 15212 35142 15292 35148
rect 15212 34592 15240 35142
rect 15292 35090 15344 35096
rect 15476 35080 15528 35086
rect 15476 35022 15528 35028
rect 15488 34950 15516 35022
rect 15476 34944 15528 34950
rect 15476 34886 15528 34892
rect 15292 34604 15344 34610
rect 15212 34564 15292 34592
rect 15292 34546 15344 34552
rect 15016 34468 15068 34474
rect 15016 34410 15068 34416
rect 15028 34218 15056 34410
rect 14936 34190 15056 34218
rect 14936 33658 14964 34190
rect 15016 34128 15068 34134
rect 15016 34070 15068 34076
rect 14924 33652 14976 33658
rect 14924 33594 14976 33600
rect 15028 32978 15056 34070
rect 15580 33590 15608 35226
rect 15764 35086 15792 36094
rect 16396 35692 16448 35698
rect 16396 35634 16448 35640
rect 15846 35388 16154 35408
rect 15846 35386 15852 35388
rect 15908 35386 15932 35388
rect 15988 35386 16012 35388
rect 16068 35386 16092 35388
rect 16148 35386 16154 35388
rect 15908 35334 15910 35386
rect 16090 35334 16092 35386
rect 15846 35332 15852 35334
rect 15908 35332 15932 35334
rect 15988 35332 16012 35334
rect 16068 35332 16092 35334
rect 16148 35332 16154 35334
rect 15846 35312 16154 35332
rect 16408 35290 16436 35634
rect 16396 35284 16448 35290
rect 16396 35226 16448 35232
rect 15752 35080 15804 35086
rect 15672 35028 15752 35034
rect 15672 35022 15804 35028
rect 15672 35006 15792 35022
rect 15672 34542 15700 35006
rect 15660 34536 15712 34542
rect 15660 34478 15712 34484
rect 15846 34300 16154 34320
rect 15846 34298 15852 34300
rect 15908 34298 15932 34300
rect 15988 34298 16012 34300
rect 16068 34298 16092 34300
rect 16148 34298 16154 34300
rect 15908 34246 15910 34298
rect 16090 34246 16092 34298
rect 15846 34244 15852 34246
rect 15908 34244 15932 34246
rect 15988 34244 16012 34246
rect 16068 34244 16092 34246
rect 16148 34244 16154 34246
rect 15846 34224 16154 34244
rect 15568 33584 15620 33590
rect 15568 33526 15620 33532
rect 16396 33584 16448 33590
rect 16396 33526 16448 33532
rect 15292 33516 15344 33522
rect 15292 33458 15344 33464
rect 15476 33516 15528 33522
rect 15476 33458 15528 33464
rect 15016 32972 15068 32978
rect 15016 32914 15068 32920
rect 15304 32434 15332 33458
rect 15488 32570 15516 33458
rect 15660 33312 15712 33318
rect 15660 33254 15712 33260
rect 15672 32910 15700 33254
rect 15846 33212 16154 33232
rect 15846 33210 15852 33212
rect 15908 33210 15932 33212
rect 15988 33210 16012 33212
rect 16068 33210 16092 33212
rect 16148 33210 16154 33212
rect 15908 33158 15910 33210
rect 16090 33158 16092 33210
rect 15846 33156 15852 33158
rect 15908 33156 15932 33158
rect 15988 33156 16012 33158
rect 16068 33156 16092 33158
rect 16148 33156 16154 33158
rect 15846 33136 16154 33156
rect 16408 33046 16436 33526
rect 16396 33040 16448 33046
rect 16396 32982 16448 32988
rect 15660 32904 15712 32910
rect 15660 32846 15712 32852
rect 15476 32564 15528 32570
rect 15476 32506 15528 32512
rect 15292 32428 15344 32434
rect 15292 32370 15344 32376
rect 14792 32184 14872 32212
rect 14740 32166 14792 32172
rect 14752 31210 14780 32166
rect 15304 31482 15332 32370
rect 15846 32124 16154 32144
rect 15846 32122 15852 32124
rect 15908 32122 15932 32124
rect 15988 32122 16012 32124
rect 16068 32122 16092 32124
rect 16148 32122 16154 32124
rect 15908 32070 15910 32122
rect 16090 32070 16092 32122
rect 15846 32068 15852 32070
rect 15908 32068 15932 32070
rect 15988 32068 16012 32070
rect 16068 32068 16092 32070
rect 16148 32068 16154 32070
rect 15846 32048 16154 32068
rect 15476 31816 15528 31822
rect 15476 31758 15528 31764
rect 15384 31680 15436 31686
rect 15384 31622 15436 31628
rect 15292 31476 15344 31482
rect 15292 31418 15344 31424
rect 15396 31278 15424 31622
rect 15016 31272 15068 31278
rect 15016 31214 15068 31220
rect 15384 31272 15436 31278
rect 15384 31214 15436 31220
rect 14740 31204 14792 31210
rect 14740 31146 14792 31152
rect 14188 30728 14240 30734
rect 14188 30670 14240 30676
rect 14096 30252 14148 30258
rect 14096 30194 14148 30200
rect 14004 29572 14056 29578
rect 14004 29514 14056 29520
rect 14016 29306 14044 29514
rect 14004 29300 14056 29306
rect 14004 29242 14056 29248
rect 14108 29238 14136 30194
rect 14200 29646 14228 30670
rect 14740 30660 14792 30666
rect 14740 30602 14792 30608
rect 14752 30394 14780 30602
rect 14740 30388 14792 30394
rect 14740 30330 14792 30336
rect 14464 30252 14516 30258
rect 14292 30212 14464 30240
rect 14188 29640 14240 29646
rect 14188 29582 14240 29588
rect 14096 29232 14148 29238
rect 14096 29174 14148 29180
rect 14108 28626 14136 29174
rect 14200 29034 14228 29582
rect 14188 29028 14240 29034
rect 14188 28970 14240 28976
rect 14096 28620 14148 28626
rect 14096 28562 14148 28568
rect 14096 28484 14148 28490
rect 14096 28426 14148 28432
rect 14108 28218 14136 28426
rect 14096 28212 14148 28218
rect 14096 28154 14148 28160
rect 14108 27538 14136 28154
rect 14200 28150 14228 28970
rect 14188 28144 14240 28150
rect 14188 28086 14240 28092
rect 14292 27577 14320 30212
rect 14464 30194 14516 30200
rect 14648 30252 14700 30258
rect 14648 30194 14700 30200
rect 14660 29170 14688 30194
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14832 29096 14884 29102
rect 14832 29038 14884 29044
rect 14844 28490 14872 29038
rect 14832 28484 14884 28490
rect 14832 28426 14884 28432
rect 14844 28082 14872 28426
rect 14464 28076 14516 28082
rect 14464 28018 14516 28024
rect 14832 28076 14884 28082
rect 14832 28018 14884 28024
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14278 27568 14334 27577
rect 14096 27532 14148 27538
rect 14278 27503 14334 27512
rect 14096 27474 14148 27480
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 14016 26790 14044 26930
rect 14004 26784 14056 26790
rect 14004 26726 14056 26732
rect 14016 26450 14044 26726
rect 14004 26444 14056 26450
rect 14004 26386 14056 26392
rect 14108 26382 14136 27474
rect 14384 27470 14412 27950
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14384 26994 14412 27406
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 14004 25696 14056 25702
rect 14004 25638 14056 25644
rect 14016 24818 14044 25638
rect 14280 25424 14332 25430
rect 14280 25366 14332 25372
rect 14292 24818 14320 25366
rect 14004 24812 14056 24818
rect 14004 24754 14056 24760
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14372 24812 14424 24818
rect 14372 24754 14424 24760
rect 14384 24342 14412 24754
rect 14372 24336 14424 24342
rect 14372 24278 14424 24284
rect 14384 23866 14412 24278
rect 14372 23860 14424 23866
rect 14372 23802 14424 23808
rect 13832 22066 13952 22094
rect 14476 22094 14504 28018
rect 14740 27396 14792 27402
rect 14740 27338 14792 27344
rect 14752 26926 14780 27338
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 14740 26920 14792 26926
rect 14740 26862 14792 26868
rect 14752 26586 14780 26862
rect 14936 26586 14964 26930
rect 14740 26580 14792 26586
rect 14740 26522 14792 26528
rect 14924 26580 14976 26586
rect 14924 26522 14976 26528
rect 14924 26308 14976 26314
rect 14924 26250 14976 26256
rect 14556 26240 14608 26246
rect 14556 26182 14608 26188
rect 14568 24800 14596 26182
rect 14936 26058 14964 26250
rect 15028 26194 15056 31214
rect 15384 31136 15436 31142
rect 15384 31078 15436 31084
rect 15200 30048 15252 30054
rect 15200 29990 15252 29996
rect 15212 28558 15240 29990
rect 15292 29640 15344 29646
rect 15292 29582 15344 29588
rect 15304 28762 15332 29582
rect 15292 28756 15344 28762
rect 15292 28698 15344 28704
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 15108 26920 15160 26926
rect 15108 26862 15160 26868
rect 15120 26314 15148 26862
rect 15108 26308 15160 26314
rect 15108 26250 15160 26256
rect 15028 26166 15148 26194
rect 14936 26030 15056 26058
rect 14832 24812 14884 24818
rect 14568 24772 14832 24800
rect 14568 24206 14596 24772
rect 14832 24754 14884 24760
rect 15028 24274 15056 26030
rect 15120 24886 15148 26166
rect 15108 24880 15160 24886
rect 15108 24822 15160 24828
rect 15016 24268 15068 24274
rect 15016 24210 15068 24216
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14568 23798 14596 24142
rect 14740 24064 14792 24070
rect 14740 24006 14792 24012
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 14752 23118 14780 24006
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 14844 23118 14872 23802
rect 15028 23254 15056 24210
rect 15120 24206 15148 24822
rect 15304 24614 15332 27406
rect 15396 26874 15424 31078
rect 15488 30326 15516 31758
rect 15568 31340 15620 31346
rect 15568 31282 15620 31288
rect 15476 30320 15528 30326
rect 15476 30262 15528 30268
rect 15488 28558 15516 30262
rect 15580 29238 15608 31282
rect 15846 31036 16154 31056
rect 15846 31034 15852 31036
rect 15908 31034 15932 31036
rect 15988 31034 16012 31036
rect 16068 31034 16092 31036
rect 16148 31034 16154 31036
rect 15908 30982 15910 31034
rect 16090 30982 16092 31034
rect 15846 30980 15852 30982
rect 15908 30980 15932 30982
rect 15988 30980 16012 30982
rect 16068 30980 16092 30982
rect 16148 30980 16154 30982
rect 15846 30960 16154 30980
rect 15660 30592 15712 30598
rect 15660 30534 15712 30540
rect 15672 30122 15700 30534
rect 15660 30116 15712 30122
rect 15660 30058 15712 30064
rect 15846 29948 16154 29968
rect 15846 29946 15852 29948
rect 15908 29946 15932 29948
rect 15988 29946 16012 29948
rect 16068 29946 16092 29948
rect 16148 29946 16154 29948
rect 15908 29894 15910 29946
rect 16090 29894 16092 29946
rect 15846 29892 15852 29894
rect 15908 29892 15932 29894
rect 15988 29892 16012 29894
rect 16068 29892 16092 29894
rect 16148 29892 16154 29894
rect 15846 29872 16154 29892
rect 15568 29232 15620 29238
rect 15568 29174 15620 29180
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15580 27962 15608 29174
rect 15660 29028 15712 29034
rect 15660 28970 15712 28976
rect 15672 28762 15700 28970
rect 15846 28860 16154 28880
rect 15846 28858 15852 28860
rect 15908 28858 15932 28860
rect 15988 28858 16012 28860
rect 16068 28858 16092 28860
rect 16148 28858 16154 28860
rect 15908 28806 15910 28858
rect 16090 28806 16092 28858
rect 15846 28804 15852 28806
rect 15908 28804 15932 28806
rect 15988 28804 16012 28806
rect 16068 28804 16092 28806
rect 16148 28804 16154 28806
rect 15846 28784 16154 28804
rect 15660 28756 15712 28762
rect 15660 28698 15712 28704
rect 15580 27934 15700 27962
rect 15568 27872 15620 27878
rect 15568 27814 15620 27820
rect 15580 27062 15608 27814
rect 15568 27056 15620 27062
rect 15568 26998 15620 27004
rect 15396 26846 15608 26874
rect 15476 24744 15528 24750
rect 15476 24686 15528 24692
rect 15292 24608 15344 24614
rect 15292 24550 15344 24556
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15304 23866 15332 24142
rect 15384 24132 15436 24138
rect 15384 24074 15436 24080
rect 15292 23860 15344 23866
rect 15292 23802 15344 23808
rect 15108 23656 15160 23662
rect 15108 23598 15160 23604
rect 15016 23248 15068 23254
rect 15016 23190 15068 23196
rect 15028 23118 15056 23190
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15016 22500 15068 22506
rect 15016 22442 15068 22448
rect 14476 22066 14688 22094
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 12624 21072 12676 21078
rect 12624 21014 12676 21020
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12912 20466 12940 20878
rect 13556 20874 13584 21082
rect 13452 20868 13504 20874
rect 13452 20810 13504 20816
rect 13544 20868 13596 20874
rect 13544 20810 13596 20816
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12912 20058 12940 20402
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11296 18584 11376 18612
rect 11244 18566 11296 18572
rect 10880 18524 11188 18544
rect 10880 18522 10886 18524
rect 10942 18522 10966 18524
rect 11022 18522 11046 18524
rect 11102 18522 11126 18524
rect 11182 18522 11188 18524
rect 10942 18470 10944 18522
rect 11124 18470 11126 18522
rect 10880 18468 10886 18470
rect 10942 18468 10966 18470
rect 11022 18468 11046 18470
rect 11102 18468 11126 18470
rect 11182 18468 11188 18470
rect 10880 18448 11188 18468
rect 10880 17436 11188 17456
rect 10880 17434 10886 17436
rect 10942 17434 10966 17436
rect 11022 17434 11046 17436
rect 11102 17434 11126 17436
rect 11182 17434 11188 17436
rect 10942 17382 10944 17434
rect 11124 17382 11126 17434
rect 10880 17380 10886 17382
rect 10942 17380 10966 17382
rect 11022 17380 11046 17382
rect 11102 17380 11126 17382
rect 11182 17380 11188 17382
rect 10880 17360 11188 17380
rect 10880 16348 11188 16368
rect 10880 16346 10886 16348
rect 10942 16346 10966 16348
rect 11022 16346 11046 16348
rect 11102 16346 11126 16348
rect 11182 16346 11188 16348
rect 10942 16294 10944 16346
rect 11124 16294 11126 16346
rect 10880 16292 10886 16294
rect 10942 16292 10966 16294
rect 11022 16292 11046 16294
rect 11102 16292 11126 16294
rect 11182 16292 11188 16294
rect 10880 16272 11188 16292
rect 10784 16176 10836 16182
rect 10690 16144 10746 16153
rect 10784 16118 10836 16124
rect 10690 16079 10746 16088
rect 10704 16028 10732 16079
rect 10704 16000 10824 16028
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 15026 10732 15846
rect 10796 15434 10824 16000
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10612 14878 10732 14906
rect 10520 14776 10640 14804
rect 10506 11792 10562 11801
rect 10506 11727 10562 11736
rect 10520 11694 10548 11727
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10508 11076 10560 11082
rect 10612 11064 10640 14776
rect 10560 11036 10640 11064
rect 10508 11018 10560 11024
rect 10520 9722 10548 11018
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10520 8537 10548 8910
rect 10506 8528 10562 8537
rect 10506 8463 10562 8472
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10520 7954 10548 8463
rect 10704 8294 10732 14878
rect 10796 14550 10824 15370
rect 10880 15260 11188 15280
rect 10880 15258 10886 15260
rect 10942 15258 10966 15260
rect 11022 15258 11046 15260
rect 11102 15258 11126 15260
rect 11182 15258 11188 15260
rect 10942 15206 10944 15258
rect 11124 15206 11126 15258
rect 10880 15204 10886 15206
rect 10942 15204 10966 15206
rect 11022 15204 11046 15206
rect 11102 15204 11126 15206
rect 11182 15204 11188 15206
rect 10880 15184 11188 15204
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 11256 14385 11284 18566
rect 11440 17882 11468 18770
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11532 17678 11560 18158
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11992 17134 12020 17546
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11992 15502 12020 17070
rect 12544 16454 12572 18702
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12636 17270 12664 18566
rect 12912 18426 12940 18566
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 13004 17882 13032 20742
rect 13464 20466 13492 20810
rect 13556 20584 13584 20810
rect 13556 20556 13676 20584
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 16114 12572 16390
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12268 15502 12296 15846
rect 13096 15502 13124 16526
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 11992 15026 12020 15438
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11796 14408 11848 14414
rect 11242 14376 11298 14385
rect 11900 14385 11928 14554
rect 12360 14521 12388 14758
rect 12346 14512 12402 14521
rect 12346 14447 12402 14456
rect 11796 14350 11848 14356
rect 11886 14376 11942 14385
rect 11242 14311 11298 14320
rect 10880 14172 11188 14192
rect 10880 14170 10886 14172
rect 10942 14170 10966 14172
rect 11022 14170 11046 14172
rect 11102 14170 11126 14172
rect 11182 14170 11188 14172
rect 10942 14118 10944 14170
rect 11124 14118 11126 14170
rect 10880 14116 10886 14118
rect 10942 14116 10966 14118
rect 11022 14116 11046 14118
rect 11102 14116 11126 14118
rect 11182 14116 11188 14118
rect 10880 14096 11188 14116
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10796 12850 10824 13874
rect 11808 13530 11836 14350
rect 11886 14311 11942 14320
rect 12452 13870 12480 14962
rect 12544 14822 12572 14962
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12544 14482 12572 14758
rect 12728 14618 12756 14962
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 10880 13084 11188 13104
rect 10880 13082 10886 13084
rect 10942 13082 10966 13084
rect 11022 13082 11046 13084
rect 11102 13082 11126 13084
rect 11182 13082 11188 13084
rect 10942 13030 10944 13082
rect 11124 13030 11126 13082
rect 10880 13028 10886 13030
rect 10942 13028 10966 13030
rect 11022 13028 11046 13030
rect 11102 13028 11126 13030
rect 11182 13028 11188 13030
rect 10880 13008 11188 13028
rect 11440 12986 11468 13194
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10796 11218 10824 12650
rect 12360 12434 12388 13262
rect 12268 12406 12388 12434
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11520 12164 11572 12170
rect 11520 12106 11572 12112
rect 10880 11996 11188 12016
rect 10880 11994 10886 11996
rect 10942 11994 10966 11996
rect 11022 11994 11046 11996
rect 11102 11994 11126 11996
rect 11182 11994 11188 11996
rect 10942 11942 10944 11994
rect 11124 11942 11126 11994
rect 10880 11940 10886 11942
rect 10942 11940 10966 11942
rect 11022 11940 11046 11942
rect 11102 11940 11126 11942
rect 11182 11940 11188 11942
rect 10880 11920 11188 11940
rect 11256 11898 11284 12106
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 11164 11098 11192 11290
rect 11256 11218 11284 11630
rect 11532 11626 11560 12106
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11624 11286 11652 12038
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11978 11248 12034 11257
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11520 11212 11572 11218
rect 11978 11183 12034 11192
rect 11520 11154 11572 11160
rect 11164 11070 11284 11098
rect 10880 10908 11188 10928
rect 10880 10906 10886 10908
rect 10942 10906 10966 10908
rect 11022 10906 11046 10908
rect 11102 10906 11126 10908
rect 11182 10906 11188 10908
rect 10942 10854 10944 10906
rect 11124 10854 11126 10906
rect 10880 10852 10886 10854
rect 10942 10852 10966 10854
rect 11022 10852 11046 10854
rect 11102 10852 11126 10854
rect 11182 10852 11188 10854
rect 10880 10832 11188 10852
rect 11256 10810 11284 11070
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 10784 10736 10836 10742
rect 10784 10678 10836 10684
rect 10796 9654 10824 10678
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10888 10062 10916 10406
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10880 9820 11188 9840
rect 10880 9818 10886 9820
rect 10942 9818 10966 9820
rect 11022 9818 11046 9820
rect 11102 9818 11126 9820
rect 11182 9818 11188 9820
rect 10942 9766 10944 9818
rect 11124 9766 11126 9818
rect 10880 9764 10886 9766
rect 10942 9764 10966 9766
rect 11022 9764 11046 9766
rect 11102 9764 11126 9766
rect 11182 9764 11188 9766
rect 10880 9744 11188 9764
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10796 7954 10824 8774
rect 10880 8732 11188 8752
rect 10880 8730 10886 8732
rect 10942 8730 10966 8732
rect 11022 8730 11046 8732
rect 11102 8730 11126 8732
rect 11182 8730 11188 8732
rect 10942 8678 10944 8730
rect 11124 8678 11126 8730
rect 10880 8676 10886 8678
rect 10942 8676 10966 8678
rect 11022 8676 11046 8678
rect 11102 8676 11126 8678
rect 11182 8676 11188 8678
rect 10880 8656 11188 8676
rect 11348 8362 11376 10950
rect 11532 10606 11560 11154
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11624 10266 11652 10610
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11624 9926 11652 10202
rect 11900 10130 11928 10950
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11532 8634 11560 8774
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10244 7002 10272 7346
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9692 4570 9720 6258
rect 10244 5642 10272 6938
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9876 4690 9904 4966
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9600 4554 9720 4570
rect 9588 4548 9720 4554
rect 9640 4542 9720 4548
rect 9588 4490 9640 4496
rect 9508 4406 9628 4434
rect 9600 4146 9628 4406
rect 9692 4214 9720 4542
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9416 3058 9444 3470
rect 9508 3194 9536 4082
rect 9600 3398 9628 4082
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9692 3058 9720 3878
rect 9784 3534 9812 4422
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10244 3738 10272 4082
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8404 2746 8616 2774
rect 8772 2774 8800 2994
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 8772 2746 8984 2774
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7944 800 7972 2382
rect 8404 2378 8432 2746
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8772 800 8800 2382
rect 8956 2310 8984 2746
rect 9324 2514 9352 2790
rect 10336 2514 10364 7346
rect 10520 7206 10548 7890
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10704 7410 10732 7754
rect 10796 7410 10824 7890
rect 10980 7886 11008 8230
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 10880 7644 11188 7664
rect 10880 7642 10886 7644
rect 10942 7642 10966 7644
rect 11022 7642 11046 7644
rect 11102 7642 11126 7644
rect 11182 7642 11188 7644
rect 10942 7590 10944 7642
rect 11124 7590 11126 7642
rect 10880 7588 10886 7590
rect 10942 7588 10966 7590
rect 11022 7588 11046 7590
rect 11102 7588 11126 7590
rect 11182 7588 11188 7590
rect 10880 7568 11188 7588
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 6322 10456 6598
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10520 2514 10548 7142
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10612 5030 10640 5578
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10704 4826 10732 7346
rect 11348 7342 11376 7754
rect 11624 7410 11652 8910
rect 11796 8560 11848 8566
rect 11794 8528 11796 8537
rect 11848 8528 11850 8537
rect 11794 8463 11850 8472
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 10880 6556 11188 6576
rect 10880 6554 10886 6556
rect 10942 6554 10966 6556
rect 11022 6554 11046 6556
rect 11102 6554 11126 6556
rect 11182 6554 11188 6556
rect 10942 6502 10944 6554
rect 11124 6502 11126 6554
rect 10880 6500 10886 6502
rect 10942 6500 10966 6502
rect 11022 6500 11046 6502
rect 11102 6500 11126 6502
rect 11182 6500 11188 6502
rect 10880 6480 11188 6500
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10980 5642 11008 6326
rect 11348 5914 11376 7278
rect 11808 6322 11836 7822
rect 11900 7546 11928 8434
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11992 5846 12020 11183
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12176 10810 12204 11018
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12084 7954 12112 8366
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12084 6866 12112 7890
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10796 4690 10824 5510
rect 10880 5468 11188 5488
rect 10880 5466 10886 5468
rect 10942 5466 10966 5468
rect 11022 5466 11046 5468
rect 11102 5466 11126 5468
rect 11182 5466 11188 5468
rect 10942 5414 10944 5466
rect 11124 5414 11126 5466
rect 10880 5412 10886 5414
rect 10942 5412 10966 5414
rect 11022 5412 11046 5414
rect 11102 5412 11126 5414
rect 11182 5412 11188 5414
rect 10880 5392 11188 5412
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10704 4010 10732 4558
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10796 3738 10824 4626
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 10880 4380 11188 4400
rect 10880 4378 10886 4380
rect 10942 4378 10966 4380
rect 11022 4378 11046 4380
rect 11102 4378 11126 4380
rect 11182 4378 11188 4380
rect 10942 4326 10944 4378
rect 11124 4326 11126 4378
rect 10880 4324 10886 4326
rect 10942 4324 10966 4326
rect 11022 4324 11046 4326
rect 11102 4324 11126 4326
rect 11182 4324 11188 4326
rect 10880 4304 11188 4324
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11072 3942 11100 4082
rect 11256 3942 11284 4422
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11256 3738 11284 3878
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11348 3466 11376 5170
rect 11336 3460 11388 3466
rect 11336 3402 11388 3408
rect 10880 3292 11188 3312
rect 10880 3290 10886 3292
rect 10942 3290 10966 3292
rect 11022 3290 11046 3292
rect 11102 3290 11126 3292
rect 11182 3290 11188 3292
rect 10942 3238 10944 3290
rect 11124 3238 11126 3290
rect 10880 3236 10886 3238
rect 10942 3236 10966 3238
rect 11022 3236 11046 3238
rect 11102 3236 11126 3238
rect 11182 3236 11188 3238
rect 10880 3216 11188 3236
rect 11440 3194 11468 5578
rect 11808 5234 11836 5578
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11704 4548 11756 4554
rect 11704 4490 11756 4496
rect 11532 3534 11560 4490
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11624 3602 11652 4014
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11716 3194 11744 4490
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11808 3074 11836 5170
rect 11888 4208 11940 4214
rect 12084 4162 12112 6598
rect 12176 6458 12204 7686
rect 12268 6662 12296 12406
rect 12452 12238 12480 13806
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12452 11694 12480 12174
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 11762 12572 12038
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12452 10266 12480 11630
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12636 9994 12664 13262
rect 12728 12850 12756 14214
rect 12820 12986 12848 14894
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12728 11218 12756 12106
rect 12820 11830 12848 12174
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12806 11384 12862 11393
rect 12806 11319 12862 11328
rect 12820 11286 12848 11319
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12728 10266 12756 11018
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12360 9518 12388 9658
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12452 9042 12480 9454
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12360 7410 12388 7822
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12268 5778 12296 6394
rect 12360 6322 12388 7346
rect 12452 6662 12480 7346
rect 12544 7342 12572 7754
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12544 6440 12572 7278
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12636 6798 12664 7142
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12452 6412 12572 6440
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12360 5846 12388 6258
rect 12452 6118 12480 6412
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12360 5658 12388 5782
rect 12268 5630 12388 5658
rect 12268 5166 12296 5630
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12360 5370 12388 5510
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12452 5166 12480 6054
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12268 4690 12296 5102
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 11888 4150 11940 4156
rect 11900 4049 11928 4150
rect 11992 4146 12296 4162
rect 11980 4140 12308 4146
rect 12032 4134 12256 4140
rect 11980 4082 12032 4088
rect 12256 4082 12308 4088
rect 11886 4040 11942 4049
rect 11886 3975 11942 3984
rect 11900 3126 11928 3975
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12360 3534 12388 3878
rect 11980 3528 12032 3534
rect 11978 3496 11980 3505
rect 12348 3528 12400 3534
rect 12032 3496 12034 3505
rect 12348 3470 12400 3476
rect 11978 3431 12034 3440
rect 12440 3460 12492 3466
rect 12492 3420 12572 3448
rect 12440 3402 12492 3408
rect 11716 3058 11836 3074
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11716 3052 11848 3058
rect 11716 3046 11796 3052
rect 11716 2650 11744 3046
rect 11796 2994 11848 3000
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 10508 2508 10560 2514
rect 10508 2450 10560 2456
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 9508 800 9536 2382
rect 10244 800 10272 2382
rect 11336 2372 11388 2378
rect 11336 2314 11388 2320
rect 10880 2204 11188 2224
rect 10880 2202 10886 2204
rect 10942 2202 10966 2204
rect 11022 2202 11046 2204
rect 11102 2202 11126 2204
rect 11182 2202 11188 2204
rect 10942 2150 10944 2202
rect 11124 2150 11126 2202
rect 10880 2148 10886 2150
rect 10942 2148 10966 2150
rect 11022 2148 11046 2150
rect 11102 2148 11126 2150
rect 11182 2148 11188 2150
rect 10880 2128 11188 2148
rect 11072 870 11192 898
rect 11072 800 11100 870
rect 2870 368 2926 377
rect 2870 303 2926 312
rect 3422 0 3478 800
rect 4158 0 4214 800
rect 4894 0 4950 800
rect 5722 0 5778 800
rect 6458 0 6514 800
rect 7194 0 7250 800
rect 7930 0 7986 800
rect 8758 0 8814 800
rect 9494 0 9550 800
rect 10230 0 10286 800
rect 11058 0 11114 800
rect 11164 762 11192 870
rect 11348 762 11376 2314
rect 11808 800 11836 2790
rect 12544 800 12572 3420
rect 12636 2310 12664 6122
rect 12728 5778 12756 6802
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12728 5234 12756 5714
rect 12820 5642 12848 6598
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12820 2774 12848 5578
rect 12912 4282 12940 14282
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13004 11898 13032 12174
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 13096 11354 13124 12242
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13096 11218 13124 11290
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13004 5370 13032 11086
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13096 10674 13124 11018
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 13188 9654 13216 19450
rect 13464 19122 13492 20402
rect 13556 20058 13584 20402
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13556 19514 13584 19790
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13464 19094 13584 19122
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 13464 17814 13492 18090
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 13268 16720 13320 16726
rect 13268 16662 13320 16668
rect 13280 15978 13308 16662
rect 13464 16250 13492 17750
rect 13556 16250 13584 19094
rect 13648 17542 13676 20556
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13740 19922 13768 20266
rect 13832 19990 13860 22066
rect 14660 20602 14688 22066
rect 15028 21010 15056 22442
rect 15120 22438 15148 23598
rect 15396 23322 15424 24074
rect 15384 23316 15436 23322
rect 15384 23258 15436 23264
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 15120 21486 15148 22374
rect 15384 22160 15436 22166
rect 15384 22102 15436 22108
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 15028 20466 15056 20946
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13740 18154 13768 19858
rect 13924 18358 13952 19994
rect 14108 19854 14136 20198
rect 14280 19984 14332 19990
rect 14280 19926 14332 19932
rect 14292 19854 14320 19926
rect 14568 19854 14596 20402
rect 14648 20324 14700 20330
rect 14648 20266 14700 20272
rect 14660 19990 14688 20266
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 14648 19984 14700 19990
rect 14648 19926 14700 19932
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14752 19446 14780 19654
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14844 19174 14872 20198
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 13728 18148 13780 18154
rect 13728 18090 13780 18096
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13832 17746 13860 18022
rect 14016 17882 14044 18702
rect 14556 18352 14608 18358
rect 14556 18294 14608 18300
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13648 16674 13676 17478
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13832 16998 13860 17138
rect 13924 16998 13952 17614
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13648 16646 13768 16674
rect 13832 16658 13860 16934
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13648 16114 13676 16526
rect 13740 16522 13768 16646
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13832 16114 13860 16594
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13648 15706 13676 16050
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13648 15026 13676 15642
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13648 14482 13676 14962
rect 13740 14822 13768 15914
rect 13820 15020 13872 15026
rect 13924 15008 13952 16934
rect 13872 14980 13952 15008
rect 13820 14962 13872 14968
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13832 14414 13860 14962
rect 14292 14618 14320 18226
rect 14568 17678 14596 18294
rect 14844 18290 14872 19110
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14476 14958 14504 16594
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14568 15502 14596 15982
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14660 15162 14688 16050
rect 14752 15978 14780 17002
rect 14936 16182 14964 17070
rect 14924 16176 14976 16182
rect 14924 16118 14976 16124
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14752 15502 14780 15914
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13726 13968 13782 13977
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13360 13932 13412 13938
rect 13726 13903 13728 13912
rect 13360 13874 13412 13880
rect 13780 13903 13782 13912
rect 13728 13874 13780 13880
rect 13280 12918 13308 13874
rect 13372 13326 13400 13874
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13740 12986 13768 13874
rect 14292 13326 14320 14554
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13280 9450 13308 9590
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13280 8498 13308 9386
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13372 8090 13400 12174
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13464 11150 13492 11766
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13648 10538 13676 12786
rect 14476 12646 14504 14894
rect 14844 14822 14872 16050
rect 14936 15570 14964 16118
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 15028 15502 15056 18022
rect 15120 17202 15148 20198
rect 15212 17814 15240 21966
rect 15292 21616 15344 21622
rect 15292 21558 15344 21564
rect 15304 17882 15332 21558
rect 15396 20602 15424 22102
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15396 18358 15424 19654
rect 15488 19378 15516 24686
rect 15580 22574 15608 26846
rect 15672 24052 15700 27934
rect 15846 27772 16154 27792
rect 15846 27770 15852 27772
rect 15908 27770 15932 27772
rect 15988 27770 16012 27772
rect 16068 27770 16092 27772
rect 16148 27770 16154 27772
rect 15908 27718 15910 27770
rect 16090 27718 16092 27770
rect 15846 27716 15852 27718
rect 15908 27716 15932 27718
rect 15988 27716 16012 27718
rect 16068 27716 16092 27718
rect 16148 27716 16154 27718
rect 15846 27696 16154 27716
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16304 26784 16356 26790
rect 16304 26726 16356 26732
rect 15846 26684 16154 26704
rect 15846 26682 15852 26684
rect 15908 26682 15932 26684
rect 15988 26682 16012 26684
rect 16068 26682 16092 26684
rect 16148 26682 16154 26684
rect 15908 26630 15910 26682
rect 16090 26630 16092 26682
rect 15846 26628 15852 26630
rect 15908 26628 15932 26630
rect 15988 26628 16012 26630
rect 16068 26628 16092 26630
rect 16148 26628 16154 26630
rect 15846 26608 16154 26628
rect 16316 26382 16344 26726
rect 16500 26586 16528 27270
rect 16488 26580 16540 26586
rect 16488 26522 16540 26528
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 15752 26240 15804 26246
rect 15752 26182 15804 26188
rect 15764 26042 15792 26182
rect 15752 26036 15804 26042
rect 15752 25978 15804 25984
rect 16488 25900 16540 25906
rect 16488 25842 16540 25848
rect 16212 25696 16264 25702
rect 16212 25638 16264 25644
rect 15846 25596 16154 25616
rect 15846 25594 15852 25596
rect 15908 25594 15932 25596
rect 15988 25594 16012 25596
rect 16068 25594 16092 25596
rect 16148 25594 16154 25596
rect 15908 25542 15910 25594
rect 16090 25542 16092 25594
rect 15846 25540 15852 25542
rect 15908 25540 15932 25542
rect 15988 25540 16012 25542
rect 16068 25540 16092 25542
rect 16148 25540 16154 25542
rect 15846 25520 16154 25540
rect 16224 25294 16252 25638
rect 16212 25288 16264 25294
rect 16212 25230 16264 25236
rect 16500 25226 16528 25842
rect 16592 25294 16620 40122
rect 16776 39982 16804 40530
rect 16764 39976 16816 39982
rect 16764 39918 16816 39924
rect 16868 39506 16896 40598
rect 17052 40594 17080 40870
rect 17316 40724 17368 40730
rect 17316 40666 17368 40672
rect 17040 40588 17092 40594
rect 17040 40530 17092 40536
rect 17328 40526 17356 40666
rect 17420 40610 17448 41074
rect 17420 40594 17540 40610
rect 17420 40588 17552 40594
rect 17420 40582 17500 40588
rect 17316 40520 17368 40526
rect 17316 40462 17368 40468
rect 17420 40186 17448 40582
rect 17500 40530 17552 40536
rect 18604 40520 18656 40526
rect 18604 40462 18656 40468
rect 17960 40384 18012 40390
rect 17960 40326 18012 40332
rect 18420 40384 18472 40390
rect 18420 40326 18472 40332
rect 17408 40180 17460 40186
rect 17408 40122 17460 40128
rect 17972 40118 18000 40326
rect 18432 40186 18460 40326
rect 18420 40180 18472 40186
rect 18420 40122 18472 40128
rect 17960 40112 18012 40118
rect 17960 40054 18012 40060
rect 18052 40112 18104 40118
rect 18052 40054 18104 40060
rect 16856 39500 16908 39506
rect 16856 39442 16908 39448
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 16776 36922 16804 37062
rect 16764 36916 16816 36922
rect 16764 36858 16816 36864
rect 16868 36802 16896 39442
rect 17972 39438 18000 40054
rect 17960 39432 18012 39438
rect 17960 39374 18012 39380
rect 18064 39370 18092 40054
rect 18616 39642 18644 40462
rect 18696 40044 18748 40050
rect 18696 39986 18748 39992
rect 18604 39636 18656 39642
rect 18604 39578 18656 39584
rect 18052 39364 18104 39370
rect 18052 39306 18104 39312
rect 17408 38548 17460 38554
rect 17408 38490 17460 38496
rect 17316 38208 17368 38214
rect 17316 38150 17368 38156
rect 17328 38010 17356 38150
rect 17316 38004 17368 38010
rect 17316 37946 17368 37952
rect 17420 37942 17448 38490
rect 17592 38344 17644 38350
rect 17592 38286 17644 38292
rect 17408 37936 17460 37942
rect 17408 37878 17460 37884
rect 17604 37738 17632 38286
rect 18064 37942 18092 39306
rect 18708 39302 18736 39986
rect 18880 39976 18932 39982
rect 18880 39918 18932 39924
rect 18892 39370 18920 39918
rect 18880 39364 18932 39370
rect 18880 39306 18932 39312
rect 18696 39296 18748 39302
rect 18696 39238 18748 39244
rect 18708 39030 18736 39238
rect 18696 39024 18748 39030
rect 18696 38966 18748 38972
rect 18892 38894 18920 39306
rect 18880 38888 18932 38894
rect 18880 38830 18932 38836
rect 18420 38344 18472 38350
rect 18420 38286 18472 38292
rect 18432 37942 18460 38286
rect 18972 38208 19024 38214
rect 18972 38150 19024 38156
rect 18052 37936 18104 37942
rect 18052 37878 18104 37884
rect 18420 37936 18472 37942
rect 18420 37878 18472 37884
rect 17868 37868 17920 37874
rect 17868 37810 17920 37816
rect 17592 37732 17644 37738
rect 17592 37674 17644 37680
rect 17880 37330 17908 37810
rect 17960 37664 18012 37670
rect 17960 37606 18012 37612
rect 17868 37324 17920 37330
rect 17868 37266 17920 37272
rect 17880 36922 17908 37266
rect 17972 37262 18000 37606
rect 17960 37256 18012 37262
rect 17960 37198 18012 37204
rect 18064 37074 18092 37878
rect 18984 37874 19012 38150
rect 18972 37868 19024 37874
rect 18972 37810 19024 37816
rect 17972 37046 18092 37074
rect 18144 37120 18196 37126
rect 18144 37062 18196 37068
rect 18420 37120 18472 37126
rect 18420 37062 18472 37068
rect 17868 36916 17920 36922
rect 17868 36858 17920 36864
rect 16776 36774 16896 36802
rect 16776 36718 16804 36774
rect 16764 36712 16816 36718
rect 16764 36654 16816 36660
rect 17040 36712 17092 36718
rect 17040 36654 17092 36660
rect 16776 35630 16804 36654
rect 17052 36378 17080 36654
rect 17040 36372 17092 36378
rect 17040 36314 17092 36320
rect 17224 36032 17276 36038
rect 17224 35974 17276 35980
rect 16764 35624 16816 35630
rect 16764 35566 16816 35572
rect 16856 35624 16908 35630
rect 16856 35566 16908 35572
rect 16868 34746 16896 35566
rect 17132 35556 17184 35562
rect 17132 35498 17184 35504
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 17040 34740 17092 34746
rect 17040 34682 17092 34688
rect 16948 33856 17000 33862
rect 16948 33798 17000 33804
rect 16960 32978 16988 33798
rect 16948 32972 17000 32978
rect 16948 32914 17000 32920
rect 17052 31482 17080 34682
rect 17144 32434 17172 35498
rect 17236 34746 17264 35974
rect 17972 35698 18000 37046
rect 18052 36100 18104 36106
rect 18052 36042 18104 36048
rect 17960 35692 18012 35698
rect 17960 35634 18012 35640
rect 17316 35488 17368 35494
rect 17316 35430 17368 35436
rect 17408 35488 17460 35494
rect 17408 35430 17460 35436
rect 17328 35154 17356 35430
rect 17316 35148 17368 35154
rect 17316 35090 17368 35096
rect 17420 34746 17448 35430
rect 17224 34740 17276 34746
rect 17224 34682 17276 34688
rect 17408 34740 17460 34746
rect 17408 34682 17460 34688
rect 18064 34610 18092 36042
rect 18052 34604 18104 34610
rect 18052 34546 18104 34552
rect 17592 34536 17644 34542
rect 17592 34478 17644 34484
rect 17408 33992 17460 33998
rect 17408 33934 17460 33940
rect 17316 33584 17368 33590
rect 17316 33526 17368 33532
rect 17328 32434 17356 33526
rect 17132 32428 17184 32434
rect 17132 32370 17184 32376
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 17420 32366 17448 33934
rect 17408 32360 17460 32366
rect 17408 32302 17460 32308
rect 17420 31958 17448 32302
rect 17408 31952 17460 31958
rect 17408 31894 17460 31900
rect 17040 31476 17092 31482
rect 17040 31418 17092 31424
rect 17224 31340 17276 31346
rect 17224 31282 17276 31288
rect 17132 31272 17184 31278
rect 17132 31214 17184 31220
rect 17144 30802 17172 31214
rect 17132 30796 17184 30802
rect 17132 30738 17184 30744
rect 17040 30728 17092 30734
rect 17040 30670 17092 30676
rect 16856 30252 16908 30258
rect 16856 30194 16908 30200
rect 16764 29640 16816 29646
rect 16764 29582 16816 29588
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16684 27878 16712 28018
rect 16672 27872 16724 27878
rect 16672 27814 16724 27820
rect 16684 25362 16712 27814
rect 16776 26382 16804 29582
rect 16868 29186 16896 30194
rect 17052 30122 17080 30670
rect 17236 30598 17264 31282
rect 17224 30592 17276 30598
rect 17224 30534 17276 30540
rect 17132 30184 17184 30190
rect 17132 30126 17184 30132
rect 17040 30116 17092 30122
rect 17040 30058 17092 30064
rect 16948 29640 17000 29646
rect 16948 29582 17000 29588
rect 16960 29306 16988 29582
rect 17052 29306 17080 30058
rect 17144 29850 17172 30126
rect 17236 29850 17264 30534
rect 17132 29844 17184 29850
rect 17132 29786 17184 29792
rect 17224 29844 17276 29850
rect 17224 29786 17276 29792
rect 17132 29640 17184 29646
rect 17132 29582 17184 29588
rect 16948 29300 17000 29306
rect 16948 29242 17000 29248
rect 17040 29300 17092 29306
rect 17040 29242 17092 29248
rect 16868 29158 16988 29186
rect 16960 28558 16988 29158
rect 17040 29164 17092 29170
rect 17040 29106 17092 29112
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 16868 27674 16896 28018
rect 16856 27668 16908 27674
rect 16856 27610 16908 27616
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 16488 25220 16540 25226
rect 16488 25162 16540 25168
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15764 24206 15792 25094
rect 16212 24744 16264 24750
rect 16212 24686 16264 24692
rect 15846 24508 16154 24528
rect 15846 24506 15852 24508
rect 15908 24506 15932 24508
rect 15988 24506 16012 24508
rect 16068 24506 16092 24508
rect 16148 24506 16154 24508
rect 15908 24454 15910 24506
rect 16090 24454 16092 24506
rect 15846 24452 15852 24454
rect 15908 24452 15932 24454
rect 15988 24452 16012 24454
rect 16068 24452 16092 24454
rect 16148 24452 16154 24454
rect 15846 24432 16154 24452
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 15672 24024 15792 24052
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 15672 22778 15700 23598
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15764 22137 15792 24024
rect 16132 23866 16160 24142
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 15846 23420 16154 23440
rect 15846 23418 15852 23420
rect 15908 23418 15932 23420
rect 15988 23418 16012 23420
rect 16068 23418 16092 23420
rect 16148 23418 16154 23420
rect 15908 23366 15910 23418
rect 16090 23366 16092 23418
rect 15846 23364 15852 23366
rect 15908 23364 15932 23366
rect 15988 23364 16012 23366
rect 16068 23364 16092 23366
rect 16148 23364 16154 23366
rect 15846 23344 16154 23364
rect 16224 22506 16252 24686
rect 16396 24676 16448 24682
rect 16396 24618 16448 24624
rect 16304 23520 16356 23526
rect 16304 23462 16356 23468
rect 16212 22500 16264 22506
rect 16212 22442 16264 22448
rect 15846 22332 16154 22352
rect 15846 22330 15852 22332
rect 15908 22330 15932 22332
rect 15988 22330 16012 22332
rect 16068 22330 16092 22332
rect 16148 22330 16154 22332
rect 15908 22278 15910 22330
rect 16090 22278 16092 22330
rect 15846 22276 15852 22278
rect 15908 22276 15932 22278
rect 15988 22276 16012 22278
rect 16068 22276 16092 22278
rect 16148 22276 16154 22278
rect 15846 22256 16154 22276
rect 15750 22128 15806 22137
rect 15660 22092 15712 22098
rect 15750 22063 15806 22072
rect 15660 22034 15712 22040
rect 15568 21956 15620 21962
rect 15568 21898 15620 21904
rect 15580 21690 15608 21898
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15672 21554 15700 22034
rect 15752 22024 15804 22030
rect 15752 21966 15804 21972
rect 16210 21992 16266 22001
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15580 20602 15608 20742
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15580 19990 15608 20334
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 15764 19938 15792 21966
rect 15844 21956 15896 21962
rect 16210 21927 16266 21936
rect 15844 21898 15896 21904
rect 15856 21622 15884 21898
rect 15844 21616 15896 21622
rect 15844 21558 15896 21564
rect 15846 21244 16154 21264
rect 15846 21242 15852 21244
rect 15908 21242 15932 21244
rect 15988 21242 16012 21244
rect 16068 21242 16092 21244
rect 16148 21242 16154 21244
rect 15908 21190 15910 21242
rect 16090 21190 16092 21242
rect 15846 21188 15852 21190
rect 15908 21188 15932 21190
rect 15988 21188 16012 21190
rect 16068 21188 16092 21190
rect 16148 21188 16154 21190
rect 15846 21168 16154 21188
rect 15846 20156 16154 20176
rect 15846 20154 15852 20156
rect 15908 20154 15932 20156
rect 15988 20154 16012 20156
rect 16068 20154 16092 20156
rect 16148 20154 16154 20156
rect 15908 20102 15910 20154
rect 16090 20102 16092 20154
rect 15846 20100 15852 20102
rect 15908 20100 15932 20102
rect 15988 20100 16012 20102
rect 16068 20100 16092 20102
rect 16148 20100 16154 20102
rect 15846 20080 16154 20100
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15488 18426 15516 18566
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15580 18222 15608 19926
rect 15764 19922 15884 19938
rect 15764 19916 15896 19922
rect 15764 19910 15844 19916
rect 15844 19858 15896 19864
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16224 19802 16252 21927
rect 16316 19922 16344 23462
rect 16408 23118 16436 24618
rect 16500 23798 16528 25162
rect 16776 24818 16804 26318
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 16868 25362 16896 25774
rect 16856 25356 16908 25362
rect 16856 25298 16908 25304
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16580 24608 16632 24614
rect 16580 24550 16632 24556
rect 16592 24342 16620 24550
rect 16580 24336 16632 24342
rect 16580 24278 16632 24284
rect 16776 24274 16804 24754
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16580 24200 16632 24206
rect 16868 24154 16896 25298
rect 16580 24142 16632 24148
rect 16488 23792 16540 23798
rect 16488 23734 16540 23740
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16408 22710 16436 23054
rect 16396 22704 16448 22710
rect 16396 22646 16448 22652
rect 16500 22642 16528 23734
rect 16592 22778 16620 24142
rect 16776 24126 16896 24154
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16684 23730 16712 24006
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16776 23610 16804 24126
rect 16684 23582 16804 23610
rect 16856 23588 16908 23594
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 16578 22672 16634 22681
rect 16488 22636 16540 22642
rect 16578 22607 16634 22616
rect 16488 22578 16540 22584
rect 16396 22568 16448 22574
rect 16396 22510 16448 22516
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15120 16590 15148 16934
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15212 16250 15240 17274
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15212 15094 15240 15302
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14660 14414 14688 14758
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14568 13734 14596 13874
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14476 12442 14504 12582
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14464 12436 14516 12442
rect 14660 12434 14688 13806
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 15028 12850 15056 13194
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 14464 12378 14516 12384
rect 14568 12406 14872 12434
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13832 11286 13860 12174
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13924 11286 13952 11698
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13832 11132 13860 11222
rect 13912 11144 13964 11150
rect 13832 11104 13912 11132
rect 13912 11086 13964 11092
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13464 10266 13492 10406
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13924 10062 13952 11086
rect 14200 10674 14228 11834
rect 14292 11762 14320 12378
rect 14568 12102 14596 12406
rect 14844 12288 14872 12406
rect 14844 12260 14964 12288
rect 14936 12170 14964 12260
rect 14832 12164 14884 12170
rect 14832 12106 14884 12112
rect 14924 12164 14976 12170
rect 14924 12106 14976 12112
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14384 11354 14412 11698
rect 14844 11354 14872 12106
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14016 10130 14044 10610
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13188 7342 13216 7890
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13372 7342 13400 7822
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7546 13492 7686
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 13280 5710 13308 6054
rect 13372 5914 13400 7278
rect 13556 6662 13584 9862
rect 13924 9654 13952 9998
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 14096 8900 14148 8906
rect 14096 8842 14148 8848
rect 14108 8634 14136 8842
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13648 6390 13676 6598
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13740 5710 13768 6190
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 13096 3670 13124 5170
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13188 4282 13216 4558
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12820 2746 12940 2774
rect 12912 2582 12940 2746
rect 13004 2582 13032 2994
rect 13096 2990 13124 3606
rect 13188 3602 13216 4218
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13176 3460 13228 3466
rect 13176 3402 13228 3408
rect 13188 3058 13216 3402
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 12900 2576 12952 2582
rect 12900 2518 12952 2524
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 13280 800 13308 5510
rect 13464 5166 13492 5646
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13372 3058 13400 4082
rect 13832 3194 13860 8434
rect 14292 7546 14320 11086
rect 14384 10062 14412 11154
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14476 10130 14504 11086
rect 15120 11064 15148 14282
rect 15304 13734 15332 17818
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14278 15516 14894
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 13530 15332 13670
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15304 12434 15332 13330
rect 15396 13326 15424 13942
rect 15580 13938 15608 15098
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15580 13326 15608 13874
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15580 12986 15608 13262
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15304 12406 15424 12434
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15212 11393 15240 12310
rect 15198 11384 15254 11393
rect 15198 11319 15254 11328
rect 15200 11076 15252 11082
rect 15120 11036 15200 11064
rect 15200 11018 15252 11024
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 14556 10532 14608 10538
rect 14556 10474 14608 10480
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14476 9722 14504 10066
rect 14568 9994 14596 10474
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13924 6254 13952 7346
rect 14384 6322 14412 8910
rect 14476 8430 14504 9658
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14568 8566 14596 9454
rect 14660 9382 14688 9998
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14844 9674 14872 9862
rect 15028 9738 15056 9998
rect 15028 9710 15148 9738
rect 14752 9654 14872 9674
rect 14740 9648 14872 9654
rect 14792 9646 14872 9648
rect 14740 9590 14792 9596
rect 15120 9450 15148 9710
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14556 8560 14608 8566
rect 14556 8502 14608 8508
rect 14568 8430 14596 8502
rect 14660 8498 14688 8842
rect 14844 8498 14872 9318
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13924 5098 13952 6190
rect 14384 5846 14412 6258
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 14384 4146 14412 5170
rect 14476 4758 14504 7346
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14568 5370 14596 5510
rect 14660 5370 14688 6258
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14464 4752 14516 4758
rect 14464 4694 14516 4700
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 14108 800 14136 3878
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14200 2650 14228 2994
rect 14476 2650 14504 4014
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14844 800 14872 6666
rect 14936 4282 14964 7686
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15028 4826 15056 7278
rect 15212 6458 15240 10610
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15304 7750 15332 9658
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15396 7528 15424 12406
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15488 11150 15516 12038
rect 15672 11626 15700 18702
rect 15764 17882 15792 19790
rect 15948 19242 15976 19790
rect 16224 19774 16344 19802
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 15936 19236 15988 19242
rect 15936 19178 15988 19184
rect 15846 19068 16154 19088
rect 15846 19066 15852 19068
rect 15908 19066 15932 19068
rect 15988 19066 16012 19068
rect 16068 19066 16092 19068
rect 16148 19066 16154 19068
rect 15908 19014 15910 19066
rect 16090 19014 16092 19066
rect 15846 19012 15852 19014
rect 15908 19012 15932 19014
rect 15988 19012 16012 19014
rect 16068 19012 16092 19014
rect 16148 19012 16154 19014
rect 15846 18992 16154 19012
rect 16224 18766 16252 19246
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 15846 17980 16154 18000
rect 15846 17978 15852 17980
rect 15908 17978 15932 17980
rect 15988 17978 16012 17980
rect 16068 17978 16092 17980
rect 16148 17978 16154 17980
rect 15908 17926 15910 17978
rect 16090 17926 16092 17978
rect 15846 17924 15852 17926
rect 15908 17924 15932 17926
rect 15988 17924 16012 17926
rect 16068 17924 16092 17926
rect 16148 17924 16154 17926
rect 15846 17904 16154 17924
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15764 17270 15792 17818
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 16040 17202 16068 17478
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 15846 16892 16154 16912
rect 15846 16890 15852 16892
rect 15908 16890 15932 16892
rect 15988 16890 16012 16892
rect 16068 16890 16092 16892
rect 16148 16890 16154 16892
rect 15908 16838 15910 16890
rect 16090 16838 16092 16890
rect 15846 16836 15852 16838
rect 15908 16836 15932 16838
rect 15988 16836 16012 16838
rect 16068 16836 16092 16838
rect 16148 16836 16154 16838
rect 15846 16816 16154 16836
rect 15846 15804 16154 15824
rect 15846 15802 15852 15804
rect 15908 15802 15932 15804
rect 15988 15802 16012 15804
rect 16068 15802 16092 15804
rect 16148 15802 16154 15804
rect 15908 15750 15910 15802
rect 16090 15750 16092 15802
rect 15846 15748 15852 15750
rect 15908 15748 15932 15750
rect 15988 15748 16012 15750
rect 16068 15748 16092 15750
rect 16148 15748 16154 15750
rect 15846 15728 16154 15748
rect 16224 15706 16252 17614
rect 16316 17338 16344 19774
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 15764 15502 15792 15642
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15764 15094 15792 15438
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15764 14822 15792 15030
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15764 13394 15792 14758
rect 15846 14716 16154 14736
rect 15846 14714 15852 14716
rect 15908 14714 15932 14716
rect 15988 14714 16012 14716
rect 16068 14714 16092 14716
rect 16148 14714 16154 14716
rect 15908 14662 15910 14714
rect 16090 14662 16092 14714
rect 15846 14660 15852 14662
rect 15908 14660 15932 14662
rect 15988 14660 16012 14662
rect 16068 14660 16092 14662
rect 16148 14660 16154 14662
rect 15846 14640 16154 14660
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 15936 14408 15988 14414
rect 16040 14396 16068 14486
rect 16120 14476 16172 14482
rect 16224 14464 16252 15642
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16316 14521 16344 14554
rect 16172 14436 16252 14464
rect 16302 14512 16358 14521
rect 16302 14447 16358 14456
rect 16120 14418 16172 14424
rect 15988 14368 16068 14396
rect 15936 14350 15988 14356
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15856 14006 15884 14214
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 16040 13938 16068 14368
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 15846 13628 16154 13648
rect 15846 13626 15852 13628
rect 15908 13626 15932 13628
rect 15988 13626 16012 13628
rect 16068 13626 16092 13628
rect 16148 13626 16154 13628
rect 15908 13574 15910 13626
rect 16090 13574 16092 13626
rect 15846 13572 15852 13574
rect 15908 13572 15932 13574
rect 15988 13572 16012 13574
rect 16068 13572 16092 13574
rect 16148 13572 16154 13574
rect 15846 13552 16154 13572
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 16224 13326 16252 14214
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 15846 12540 16154 12560
rect 15846 12538 15852 12540
rect 15908 12538 15932 12540
rect 15988 12538 16012 12540
rect 16068 12538 16092 12540
rect 16148 12538 16154 12540
rect 15908 12486 15910 12538
rect 16090 12486 16092 12538
rect 15846 12484 15852 12486
rect 15908 12484 15932 12486
rect 15988 12484 16012 12486
rect 16068 12484 16092 12486
rect 16148 12484 16154 12486
rect 15846 12464 16154 12484
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15672 10674 15700 11562
rect 15846 11452 16154 11472
rect 15846 11450 15852 11452
rect 15908 11450 15932 11452
rect 15988 11450 16012 11452
rect 16068 11450 16092 11452
rect 16148 11450 16154 11452
rect 15908 11398 15910 11450
rect 16090 11398 16092 11450
rect 15846 11396 15852 11398
rect 15908 11396 15932 11398
rect 15988 11396 16012 11398
rect 16068 11396 16092 11398
rect 16148 11396 16154 11398
rect 15846 11376 16154 11396
rect 16224 11336 16252 12174
rect 16040 11308 16252 11336
rect 16040 11150 16068 11308
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 15764 10742 15792 11086
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15752 10600 15804 10606
rect 15856 10554 15884 10950
rect 15804 10548 15884 10554
rect 15752 10542 15884 10548
rect 15764 10526 15884 10542
rect 16040 10538 16068 11086
rect 16224 10810 16252 11086
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 15846 10364 16154 10384
rect 15846 10362 15852 10364
rect 15908 10362 15932 10364
rect 15988 10362 16012 10364
rect 16068 10362 16092 10364
rect 16148 10362 16154 10364
rect 15908 10310 15910 10362
rect 16090 10310 16092 10362
rect 15846 10308 15852 10310
rect 15908 10308 15932 10310
rect 15988 10308 16012 10310
rect 16068 10308 16092 10310
rect 16148 10308 16154 10310
rect 15846 10288 16154 10308
rect 15568 9988 15620 9994
rect 15568 9930 15620 9936
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15488 8838 15516 9522
rect 15580 8974 15608 9930
rect 15660 9648 15712 9654
rect 15658 9616 15660 9625
rect 15712 9616 15714 9625
rect 15658 9551 15714 9560
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15488 7886 15516 8774
rect 15672 8294 15700 9454
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 15846 9276 16154 9296
rect 15846 9274 15852 9276
rect 15908 9274 15932 9276
rect 15988 9274 16012 9276
rect 16068 9274 16092 9276
rect 16148 9274 16154 9276
rect 15908 9222 15910 9274
rect 16090 9222 16092 9274
rect 15846 9220 15852 9222
rect 15908 9220 15932 9222
rect 15988 9220 16012 9222
rect 16068 9220 16092 9222
rect 16148 9220 16154 9222
rect 15846 9200 16154 9220
rect 16224 8362 16252 9318
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15568 7948 15620 7954
rect 15672 7936 15700 8230
rect 15846 8188 16154 8208
rect 15846 8186 15852 8188
rect 15908 8186 15932 8188
rect 15988 8186 16012 8188
rect 16068 8186 16092 8188
rect 16148 8186 16154 8188
rect 15908 8134 15910 8186
rect 16090 8134 16092 8186
rect 15846 8132 15852 8134
rect 15908 8132 15932 8134
rect 15988 8132 16012 8134
rect 16068 8132 16092 8134
rect 16148 8132 16154 8134
rect 15846 8112 16154 8132
rect 15620 7908 15700 7936
rect 15568 7890 15620 7896
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15304 7500 15424 7528
rect 15304 6662 15332 7500
rect 15384 7404 15436 7410
rect 15488 7392 15516 7822
rect 15580 7410 15608 7890
rect 15752 7880 15804 7886
rect 15672 7840 15752 7868
rect 15436 7364 15516 7392
rect 15384 7346 15436 7352
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 15120 5778 15148 6326
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15212 5234 15240 6394
rect 15396 5234 15424 7142
rect 15488 6934 15516 7364
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15580 6866 15608 7346
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14936 2446 14964 2790
rect 15028 2774 15056 3470
rect 15120 3126 15148 4626
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 15120 2922 15148 3062
rect 15212 3058 15240 4082
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 15212 2774 15240 2994
rect 15028 2746 15148 2774
rect 15212 2746 15332 2774
rect 15016 2508 15068 2514
rect 15120 2496 15148 2746
rect 15068 2468 15148 2496
rect 15016 2450 15068 2456
rect 15304 2446 15332 2746
rect 15396 2650 15424 4150
rect 15488 4146 15516 6598
rect 15580 5166 15608 6802
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15580 3126 15608 4422
rect 15672 3738 15700 7840
rect 15752 7822 15804 7828
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16040 7342 16068 7822
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15764 5710 15792 7142
rect 15846 7100 16154 7120
rect 15846 7098 15852 7100
rect 15908 7098 15932 7100
rect 15988 7098 16012 7100
rect 16068 7098 16092 7100
rect 16148 7098 16154 7100
rect 15908 7046 15910 7098
rect 16090 7046 16092 7098
rect 15846 7044 15852 7046
rect 15908 7044 15932 7046
rect 15988 7044 16012 7046
rect 16068 7044 16092 7046
rect 16148 7044 16154 7046
rect 15846 7024 16154 7044
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 15846 6012 16154 6032
rect 15846 6010 15852 6012
rect 15908 6010 15932 6012
rect 15988 6010 16012 6012
rect 16068 6010 16092 6012
rect 16148 6010 16154 6012
rect 15908 5958 15910 6010
rect 16090 5958 16092 6010
rect 15846 5956 15852 5958
rect 15908 5956 15932 5958
rect 15988 5956 16012 5958
rect 16068 5956 16092 5958
rect 16148 5956 16154 5958
rect 15846 5936 16154 5956
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 16224 5234 16252 6870
rect 16316 6322 16344 12922
rect 16408 12918 16436 22510
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16500 22030 16528 22442
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16592 21078 16620 22607
rect 16684 22438 16712 23582
rect 16856 23530 16908 23536
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 16776 22817 16804 23122
rect 16762 22808 16818 22817
rect 16762 22743 16818 22752
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16684 21690 16712 21966
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16776 20890 16804 22578
rect 16868 22506 16896 23530
rect 16960 23526 16988 28494
rect 17052 27130 17080 29106
rect 17144 28218 17172 29582
rect 17236 28762 17264 29786
rect 17420 29714 17448 31894
rect 17500 30796 17552 30802
rect 17500 30738 17552 30744
rect 17512 30190 17540 30738
rect 17500 30184 17552 30190
rect 17500 30126 17552 30132
rect 17512 29714 17540 30126
rect 17408 29708 17460 29714
rect 17408 29650 17460 29656
rect 17500 29708 17552 29714
rect 17500 29650 17552 29656
rect 17224 28756 17276 28762
rect 17224 28698 17276 28704
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 17236 27470 17264 28698
rect 17224 27464 17276 27470
rect 17224 27406 17276 27412
rect 17236 27130 17264 27406
rect 17040 27124 17092 27130
rect 17040 27066 17092 27072
rect 17224 27124 17276 27130
rect 17224 27066 17276 27072
rect 17052 25906 17080 27066
rect 17316 26920 17368 26926
rect 17316 26862 17368 26868
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 17224 25152 17276 25158
rect 17224 25094 17276 25100
rect 17132 24200 17184 24206
rect 17132 24142 17184 24148
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16948 22976 17000 22982
rect 16948 22918 17000 22924
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16868 21010 16896 21966
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16500 19242 16528 20402
rect 16592 20058 16620 20878
rect 16776 20862 16896 20890
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16776 20602 16804 20742
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16578 19816 16634 19825
rect 16578 19751 16634 19760
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 16500 18834 16528 19178
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16592 15434 16620 19751
rect 16684 19514 16712 20402
rect 16776 19854 16804 20538
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16776 19378 16804 19450
rect 16764 19372 16816 19378
rect 16764 19314 16816 19320
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 16684 17746 16712 18770
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16776 17066 16804 19314
rect 16868 17678 16896 20862
rect 16960 18698 16988 22918
rect 17052 22234 17080 23666
rect 17040 22228 17092 22234
rect 17040 22170 17092 22176
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 17052 21622 17080 21966
rect 17144 21729 17172 24142
rect 17236 23662 17264 25094
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 17224 23520 17276 23526
rect 17224 23462 17276 23468
rect 17130 21720 17186 21729
rect 17130 21655 17186 21664
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 16960 17882 16988 18634
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16868 17338 16896 17614
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16776 16590 16804 17002
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16670 16280 16726 16289
rect 16670 16215 16726 16224
rect 16684 16114 16712 16215
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16776 15162 16804 16526
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16868 15570 16896 16050
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16960 15881 16988 15982
rect 16946 15872 17002 15881
rect 16946 15807 17002 15816
rect 17052 15706 17080 21558
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 17144 20806 17172 21490
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 17236 18290 17264 23462
rect 17328 22094 17356 26862
rect 17420 23798 17448 29650
rect 17500 28552 17552 28558
rect 17500 28494 17552 28500
rect 17512 27538 17540 28494
rect 17500 27532 17552 27538
rect 17500 27474 17552 27480
rect 17512 26926 17540 27474
rect 17604 27402 17632 34478
rect 17960 33516 18012 33522
rect 17960 33458 18012 33464
rect 17868 32836 17920 32842
rect 17868 32778 17920 32784
rect 17880 32570 17908 32778
rect 17868 32564 17920 32570
rect 17868 32506 17920 32512
rect 17776 32292 17828 32298
rect 17776 32234 17828 32240
rect 17592 27396 17644 27402
rect 17592 27338 17644 27344
rect 17500 26920 17552 26926
rect 17500 26862 17552 26868
rect 17512 25770 17540 26862
rect 17788 26466 17816 32234
rect 17868 31136 17920 31142
rect 17868 31078 17920 31084
rect 17880 30734 17908 31078
rect 17972 30802 18000 33458
rect 17960 30796 18012 30802
rect 17960 30738 18012 30744
rect 17868 30728 17920 30734
rect 17868 30670 17920 30676
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 17880 28626 17908 30194
rect 17868 28620 17920 28626
rect 17868 28562 17920 28568
rect 17868 28076 17920 28082
rect 17868 28018 17920 28024
rect 17880 26586 17908 28018
rect 17972 28014 18000 30738
rect 18064 30054 18092 34546
rect 18052 30048 18104 30054
rect 18050 30016 18052 30025
rect 18104 30016 18106 30025
rect 18050 29951 18106 29960
rect 18156 29714 18184 37062
rect 18432 36786 18460 37062
rect 19076 36854 19104 43250
rect 29932 43246 29960 44134
rect 30116 44033 30144 44338
rect 30102 44024 30158 44033
rect 30102 43959 30158 43968
rect 29920 43240 29972 43246
rect 29920 43182 29972 43188
rect 25776 43004 26084 43024
rect 25776 43002 25782 43004
rect 25838 43002 25862 43004
rect 25918 43002 25942 43004
rect 25998 43002 26022 43004
rect 26078 43002 26084 43004
rect 25838 42950 25840 43002
rect 26020 42950 26022 43002
rect 25776 42948 25782 42950
rect 25838 42948 25862 42950
rect 25918 42948 25942 42950
rect 25998 42948 26022 42950
rect 26078 42948 26084 42950
rect 25776 42928 26084 42948
rect 30104 42696 30156 42702
rect 30104 42638 30156 42644
rect 29920 42560 29972 42566
rect 30116 42537 30144 42638
rect 29920 42502 29972 42508
rect 30102 42528 30158 42537
rect 20811 42460 21119 42480
rect 20811 42458 20817 42460
rect 20873 42458 20897 42460
rect 20953 42458 20977 42460
rect 21033 42458 21057 42460
rect 21113 42458 21119 42460
rect 20873 42406 20875 42458
rect 21055 42406 21057 42458
rect 20811 42404 20817 42406
rect 20873 42404 20897 42406
rect 20953 42404 20977 42406
rect 21033 42404 21057 42406
rect 21113 42404 21119 42406
rect 20811 42384 21119 42404
rect 25776 41916 26084 41936
rect 25776 41914 25782 41916
rect 25838 41914 25862 41916
rect 25918 41914 25942 41916
rect 25998 41914 26022 41916
rect 26078 41914 26084 41916
rect 25838 41862 25840 41914
rect 26020 41862 26022 41914
rect 25776 41860 25782 41862
rect 25838 41860 25862 41862
rect 25918 41860 25942 41862
rect 25998 41860 26022 41862
rect 26078 41860 26084 41862
rect 25776 41840 26084 41860
rect 29932 41614 29960 42502
rect 30102 42463 30158 42472
rect 29920 41608 29972 41614
rect 29920 41550 29972 41556
rect 22008 41540 22060 41546
rect 22008 41482 22060 41488
rect 21916 41472 21968 41478
rect 21916 41414 21968 41420
rect 20811 41372 21119 41392
rect 20811 41370 20817 41372
rect 20873 41370 20897 41372
rect 20953 41370 20977 41372
rect 21033 41370 21057 41372
rect 21113 41370 21119 41372
rect 20873 41318 20875 41370
rect 21055 41318 21057 41370
rect 20811 41316 20817 41318
rect 20873 41316 20897 41318
rect 20953 41316 20977 41318
rect 21033 41316 21057 41318
rect 21113 41316 21119 41318
rect 20811 41296 21119 41316
rect 21928 41274 21956 41414
rect 21916 41268 21968 41274
rect 21916 41210 21968 41216
rect 22020 41138 22048 41482
rect 22008 41132 22060 41138
rect 22008 41074 22060 41080
rect 30104 41132 30156 41138
rect 30104 41074 30156 41080
rect 19800 40452 19852 40458
rect 19800 40394 19852 40400
rect 19812 40118 19840 40394
rect 20811 40284 21119 40304
rect 20811 40282 20817 40284
rect 20873 40282 20897 40284
rect 20953 40282 20977 40284
rect 21033 40282 21057 40284
rect 21113 40282 21119 40284
rect 20873 40230 20875 40282
rect 21055 40230 21057 40282
rect 20811 40228 20817 40230
rect 20873 40228 20897 40230
rect 20953 40228 20977 40230
rect 21033 40228 21057 40230
rect 21113 40228 21119 40230
rect 20811 40208 21119 40228
rect 19800 40112 19852 40118
rect 19800 40054 19852 40060
rect 19432 39840 19484 39846
rect 19432 39782 19484 39788
rect 19444 39438 19472 39782
rect 19432 39432 19484 39438
rect 19432 39374 19484 39380
rect 19812 39302 19840 40054
rect 20076 39840 20128 39846
rect 20076 39782 20128 39788
rect 19156 39296 19208 39302
rect 19156 39238 19208 39244
rect 19800 39296 19852 39302
rect 19800 39238 19852 39244
rect 19168 39098 19196 39238
rect 19156 39092 19208 39098
rect 19156 39034 19208 39040
rect 20088 38962 20116 39782
rect 22020 39370 22048 41074
rect 30116 41041 30144 41074
rect 30102 41032 30158 41041
rect 30102 40967 30158 40976
rect 25776 40828 26084 40848
rect 25776 40826 25782 40828
rect 25838 40826 25862 40828
rect 25918 40826 25942 40828
rect 25998 40826 26022 40828
rect 26078 40826 26084 40828
rect 25838 40774 25840 40826
rect 26020 40774 26022 40826
rect 25776 40772 25782 40774
rect 25838 40772 25862 40774
rect 25918 40772 25942 40774
rect 25998 40772 26022 40774
rect 26078 40772 26084 40774
rect 25776 40752 26084 40772
rect 25776 39740 26084 39760
rect 25776 39738 25782 39740
rect 25838 39738 25862 39740
rect 25918 39738 25942 39740
rect 25998 39738 26022 39740
rect 26078 39738 26084 39740
rect 25838 39686 25840 39738
rect 26020 39686 26022 39738
rect 25776 39684 25782 39686
rect 25838 39684 25862 39686
rect 25918 39684 25942 39686
rect 25998 39684 26022 39686
rect 26078 39684 26084 39686
rect 25776 39664 26084 39684
rect 22284 39568 22336 39574
rect 22284 39510 22336 39516
rect 20260 39364 20312 39370
rect 20260 39306 20312 39312
rect 22008 39364 22060 39370
rect 22008 39306 22060 39312
rect 20272 39098 20300 39306
rect 21548 39296 21600 39302
rect 21548 39238 21600 39244
rect 20811 39196 21119 39216
rect 20811 39194 20817 39196
rect 20873 39194 20897 39196
rect 20953 39194 20977 39196
rect 21033 39194 21057 39196
rect 21113 39194 21119 39196
rect 20873 39142 20875 39194
rect 21055 39142 21057 39194
rect 20811 39140 20817 39142
rect 20873 39140 20897 39142
rect 20953 39140 20977 39142
rect 21033 39140 21057 39142
rect 21113 39140 21119 39142
rect 20811 39120 21119 39140
rect 20260 39092 20312 39098
rect 20260 39034 20312 39040
rect 20076 38956 20128 38962
rect 20076 38898 20128 38904
rect 20260 38752 20312 38758
rect 20260 38694 20312 38700
rect 19432 38548 19484 38554
rect 19432 38490 19484 38496
rect 19248 37868 19300 37874
rect 19248 37810 19300 37816
rect 19064 36848 19116 36854
rect 19064 36790 19116 36796
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 18604 36780 18656 36786
rect 18604 36722 18656 36728
rect 18616 36378 18644 36722
rect 18604 36372 18656 36378
rect 18604 36314 18656 36320
rect 18236 36168 18288 36174
rect 18236 36110 18288 36116
rect 18604 36168 18656 36174
rect 18604 36110 18656 36116
rect 18248 35834 18276 36110
rect 18616 35834 18644 36110
rect 18236 35828 18288 35834
rect 18236 35770 18288 35776
rect 18604 35828 18656 35834
rect 18604 35770 18656 35776
rect 19156 35828 19208 35834
rect 19156 35770 19208 35776
rect 18972 35692 19024 35698
rect 18972 35634 19024 35640
rect 18236 35012 18288 35018
rect 18236 34954 18288 34960
rect 18248 34746 18276 34954
rect 18236 34740 18288 34746
rect 18236 34682 18288 34688
rect 18512 33992 18564 33998
rect 18512 33934 18564 33940
rect 18328 33584 18380 33590
rect 18328 33526 18380 33532
rect 18340 32774 18368 33526
rect 18328 32768 18380 32774
rect 18328 32710 18380 32716
rect 18420 32768 18472 32774
rect 18420 32710 18472 32716
rect 18340 32434 18368 32710
rect 18328 32428 18380 32434
rect 18328 32370 18380 32376
rect 18432 32366 18460 32710
rect 18524 32484 18552 33934
rect 18880 33924 18932 33930
rect 18880 33866 18932 33872
rect 18696 33312 18748 33318
rect 18696 33254 18748 33260
rect 18604 32496 18656 32502
rect 18524 32456 18604 32484
rect 18420 32360 18472 32366
rect 18340 32308 18420 32314
rect 18340 32302 18472 32308
rect 18340 32286 18460 32302
rect 18340 31482 18368 32286
rect 18432 32237 18460 32286
rect 18524 32026 18552 32456
rect 18604 32438 18656 32444
rect 18708 32298 18736 33254
rect 18892 32434 18920 33866
rect 18880 32428 18932 32434
rect 18880 32370 18932 32376
rect 18696 32292 18748 32298
rect 18696 32234 18748 32240
rect 18512 32020 18564 32026
rect 18512 31962 18564 31968
rect 18420 31884 18472 31890
rect 18420 31826 18472 31832
rect 18328 31476 18380 31482
rect 18328 31418 18380 31424
rect 18432 31414 18460 31826
rect 18708 31822 18736 32234
rect 18696 31816 18748 31822
rect 18696 31758 18748 31764
rect 18984 31754 19012 35634
rect 19168 34746 19196 35770
rect 19156 34740 19208 34746
rect 19156 34682 19208 34688
rect 19168 33114 19196 34682
rect 19064 33108 19116 33114
rect 19064 33050 19116 33056
rect 19156 33108 19208 33114
rect 19156 33050 19208 33056
rect 19076 32026 19104 33050
rect 19168 32366 19196 33050
rect 19260 32570 19288 37810
rect 19340 37664 19392 37670
rect 19340 37606 19392 37612
rect 19352 37262 19380 37606
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19444 37074 19472 38490
rect 19984 37256 20036 37262
rect 19984 37198 20036 37204
rect 19352 37046 19472 37074
rect 19352 34474 19380 37046
rect 19996 36650 20024 37198
rect 20076 37188 20128 37194
rect 20076 37130 20128 37136
rect 19984 36644 20036 36650
rect 19984 36586 20036 36592
rect 19800 36576 19852 36582
rect 19800 36518 19852 36524
rect 19616 36304 19668 36310
rect 19616 36246 19668 36252
rect 19524 35624 19576 35630
rect 19524 35566 19576 35572
rect 19432 35488 19484 35494
rect 19432 35430 19484 35436
rect 19444 34542 19472 35430
rect 19536 34678 19564 35566
rect 19524 34672 19576 34678
rect 19524 34614 19576 34620
rect 19432 34536 19484 34542
rect 19432 34478 19484 34484
rect 19340 34468 19392 34474
rect 19340 34410 19392 34416
rect 19444 34134 19472 34478
rect 19432 34128 19484 34134
rect 19432 34070 19484 34076
rect 19340 33856 19392 33862
rect 19340 33798 19392 33804
rect 19352 33522 19380 33798
rect 19340 33516 19392 33522
rect 19340 33458 19392 33464
rect 19248 32564 19300 32570
rect 19248 32506 19300 32512
rect 19156 32360 19208 32366
rect 19156 32302 19208 32308
rect 19064 32020 19116 32026
rect 19064 31962 19116 31968
rect 18984 31726 19104 31754
rect 18420 31408 18472 31414
rect 18420 31350 18472 31356
rect 18236 30116 18288 30122
rect 18236 30058 18288 30064
rect 18052 29708 18104 29714
rect 18052 29650 18104 29656
rect 18144 29708 18196 29714
rect 18144 29650 18196 29656
rect 18064 28558 18092 29650
rect 18248 29306 18276 30058
rect 18512 29640 18564 29646
rect 18512 29582 18564 29588
rect 18420 29504 18472 29510
rect 18420 29446 18472 29452
rect 18236 29300 18288 29306
rect 18236 29242 18288 29248
rect 18144 29164 18196 29170
rect 18144 29106 18196 29112
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 17960 28008 18012 28014
rect 17960 27950 18012 27956
rect 17972 27554 18000 27950
rect 18064 27674 18092 28018
rect 18052 27668 18104 27674
rect 18052 27610 18104 27616
rect 17972 27526 18092 27554
rect 17868 26580 17920 26586
rect 17868 26522 17920 26528
rect 17788 26438 17908 26466
rect 17592 26308 17644 26314
rect 17592 26250 17644 26256
rect 17604 26042 17632 26250
rect 17592 26036 17644 26042
rect 17592 25978 17644 25984
rect 17500 25764 17552 25770
rect 17500 25706 17552 25712
rect 17684 25696 17736 25702
rect 17684 25638 17736 25644
rect 17696 24954 17724 25638
rect 17684 24948 17736 24954
rect 17684 24890 17736 24896
rect 17684 24676 17736 24682
rect 17684 24618 17736 24624
rect 17408 23792 17460 23798
rect 17460 23752 17540 23780
rect 17408 23734 17460 23740
rect 17408 23656 17460 23662
rect 17408 23598 17460 23604
rect 17420 23322 17448 23598
rect 17408 23316 17460 23322
rect 17408 23258 17460 23264
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17420 22778 17448 22986
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17328 22066 17448 22094
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17328 19825 17356 21966
rect 17314 19816 17370 19825
rect 17314 19751 17370 19760
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17224 17808 17276 17814
rect 17224 17750 17276 17756
rect 17236 17270 17264 17750
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17236 16250 17264 16526
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17328 16114 17356 19654
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16776 15026 16804 15098
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16592 14550 16620 14962
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16764 14408 16816 14414
rect 16868 14396 16896 15506
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 16960 14414 16988 15030
rect 17420 14958 17448 22066
rect 17512 21418 17540 23752
rect 17696 22030 17724 24618
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17788 24274 17816 24550
rect 17776 24268 17828 24274
rect 17776 24210 17828 24216
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17590 21720 17646 21729
rect 17590 21655 17646 21664
rect 17500 21412 17552 21418
rect 17500 21354 17552 21360
rect 17500 20868 17552 20874
rect 17500 20810 17552 20816
rect 17512 19514 17540 20810
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17512 17882 17540 18158
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17604 17762 17632 21655
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17788 19514 17816 19654
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 17604 17734 17816 17762
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17592 17264 17644 17270
rect 17592 17206 17644 17212
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 16816 14368 16896 14396
rect 16948 14408 17000 14414
rect 16764 14350 16816 14356
rect 16948 14350 17000 14356
rect 17316 14408 17368 14414
rect 17420 14396 17448 14894
rect 17512 14414 17540 15506
rect 17604 15502 17632 17206
rect 17696 17202 17724 17614
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17696 16017 17724 17138
rect 17682 16008 17738 16017
rect 17682 15943 17738 15952
rect 17696 15706 17724 15943
rect 17788 15706 17816 17734
rect 17880 17134 17908 26438
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 17972 19854 18000 26250
rect 18064 26246 18092 27526
rect 18156 27130 18184 29106
rect 18248 29102 18276 29242
rect 18236 29096 18288 29102
rect 18236 29038 18288 29044
rect 18328 28960 18380 28966
rect 18328 28902 18380 28908
rect 18340 28558 18368 28902
rect 18328 28552 18380 28558
rect 18328 28494 18380 28500
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 18144 27124 18196 27130
rect 18144 27066 18196 27072
rect 18248 26382 18276 28358
rect 18432 28082 18460 29446
rect 18524 28422 18552 29582
rect 18696 29300 18748 29306
rect 18696 29242 18748 29248
rect 18604 28552 18656 28558
rect 18604 28494 18656 28500
rect 18512 28416 18564 28422
rect 18512 28358 18564 28364
rect 18524 28082 18552 28358
rect 18616 28218 18644 28494
rect 18604 28212 18656 28218
rect 18604 28154 18656 28160
rect 18420 28076 18472 28082
rect 18420 28018 18472 28024
rect 18512 28076 18564 28082
rect 18512 28018 18564 28024
rect 18524 27962 18552 28018
rect 18432 27934 18552 27962
rect 18604 27940 18656 27946
rect 18432 27470 18460 27934
rect 18604 27882 18656 27888
rect 18616 27538 18644 27882
rect 18604 27532 18656 27538
rect 18604 27474 18656 27480
rect 18420 27464 18472 27470
rect 18420 27406 18472 27412
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 18052 26240 18104 26246
rect 18052 26182 18104 26188
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 18052 25832 18104 25838
rect 18052 25774 18104 25780
rect 18064 25498 18092 25774
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 18064 23254 18092 25094
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18052 23248 18104 23254
rect 18052 23190 18104 23196
rect 18052 23112 18104 23118
rect 18050 23080 18052 23089
rect 18104 23080 18106 23089
rect 18050 23015 18106 23024
rect 18052 22568 18104 22574
rect 18052 22510 18104 22516
rect 18064 22030 18092 22510
rect 18156 22098 18184 23462
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 18052 21888 18104 21894
rect 18052 21830 18104 21836
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 18064 21554 18092 21830
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 18064 20806 18092 21490
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 18156 20534 18184 21830
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17972 18970 18000 19314
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 18248 18442 18276 26182
rect 18340 19514 18368 26930
rect 18432 25906 18460 27406
rect 18604 27328 18656 27334
rect 18604 27270 18656 27276
rect 18616 26926 18644 27270
rect 18708 26926 18736 29242
rect 18788 29164 18840 29170
rect 18788 29106 18840 29112
rect 18800 28218 18828 29106
rect 18788 28212 18840 28218
rect 18788 28154 18840 28160
rect 18880 28144 18932 28150
rect 18880 28086 18932 28092
rect 18604 26920 18656 26926
rect 18604 26862 18656 26868
rect 18696 26920 18748 26926
rect 18696 26862 18748 26868
rect 18616 25974 18644 26862
rect 18604 25968 18656 25974
rect 18604 25910 18656 25916
rect 18420 25900 18472 25906
rect 18420 25842 18472 25848
rect 18420 25220 18472 25226
rect 18420 25162 18472 25168
rect 18432 23202 18460 25162
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18616 23866 18644 24550
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18512 23724 18564 23730
rect 18512 23666 18564 23672
rect 18524 23322 18552 23666
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18512 23316 18564 23322
rect 18512 23258 18564 23264
rect 18432 23174 18552 23202
rect 18420 23044 18472 23050
rect 18420 22986 18472 22992
rect 18432 21486 18460 22986
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18340 18766 18368 19450
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18156 18414 18276 18442
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18064 17746 18092 18158
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 18064 17338 18092 17682
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18064 16153 18092 16390
rect 18050 16144 18106 16153
rect 18050 16079 18052 16088
rect 18104 16079 18106 16088
rect 18052 16050 18104 16056
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17604 15094 17632 15438
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17368 14368 17448 14396
rect 17316 14350 17368 14356
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16960 13190 16988 13874
rect 17038 13696 17094 13705
rect 17038 13631 17094 13640
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16408 12102 16436 12854
rect 17052 12850 17080 13631
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16776 12306 16804 12582
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16408 11150 16436 11562
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16408 9994 16436 11086
rect 16592 11014 16620 11698
rect 16960 11354 16988 12786
rect 17236 12442 17264 13330
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 17052 11082 17080 11222
rect 17144 11082 17172 11494
rect 17328 11150 17356 14214
rect 17420 12646 17448 14368
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17512 13938 17540 14350
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17512 12850 17540 13874
rect 17696 13870 17724 15642
rect 17788 15434 17816 15642
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17880 15162 17908 15982
rect 18156 15722 18184 18414
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18248 17678 18276 18226
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18248 16794 18276 17614
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18064 15694 18184 15722
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17868 14408 17920 14414
rect 17972 14396 18000 15030
rect 18064 14414 18092 15694
rect 18248 15570 18276 16730
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18156 15094 18184 15302
rect 18248 15094 18276 15370
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 18236 15088 18288 15094
rect 18236 15030 18288 15036
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 17920 14368 18000 14396
rect 18052 14408 18104 14414
rect 17868 14350 17920 14356
rect 18052 14350 18104 14356
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17696 13274 17724 13330
rect 17788 13326 17816 14010
rect 17604 13246 17724 13274
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17604 12986 17632 13246
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17696 12850 17724 13126
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17500 12708 17552 12714
rect 17500 12650 17552 12656
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17236 10674 17264 10950
rect 17328 10810 17356 11086
rect 17420 11014 17448 11630
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17512 10810 17540 12650
rect 17880 11898 17908 14214
rect 17958 13968 18014 13977
rect 17958 13903 17960 13912
rect 18012 13903 18014 13912
rect 17960 13874 18012 13880
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 16684 10130 16712 10610
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16960 9518 16988 10610
rect 17328 10130 17356 10746
rect 17604 10674 17632 11834
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17696 11354 17724 11698
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17512 10266 17540 10610
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16488 8288 16540 8294
rect 16488 8230 16540 8236
rect 16500 7886 16528 8230
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16684 7410 16712 9114
rect 17052 8838 17080 9454
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16776 8090 16804 8434
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16868 7886 16896 8570
rect 17052 8566 17080 8774
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16684 5914 16712 7346
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16960 6866 16988 7278
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 15846 4924 16154 4944
rect 15846 4922 15852 4924
rect 15908 4922 15932 4924
rect 15988 4922 16012 4924
rect 16068 4922 16092 4924
rect 16148 4922 16154 4924
rect 15908 4870 15910 4922
rect 16090 4870 16092 4922
rect 15846 4868 15852 4870
rect 15908 4868 15932 4870
rect 15988 4868 16012 4870
rect 16068 4868 16092 4870
rect 16148 4868 16154 4870
rect 15846 4848 16154 4868
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15764 4078 15792 4626
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16396 4480 16448 4486
rect 16396 4422 16448 4428
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15764 3602 15792 4014
rect 15846 3836 16154 3856
rect 15846 3834 15852 3836
rect 15908 3834 15932 3836
rect 15988 3834 16012 3836
rect 16068 3834 16092 3836
rect 16148 3834 16154 3836
rect 15908 3782 15910 3834
rect 16090 3782 16092 3834
rect 15846 3780 15852 3782
rect 15908 3780 15932 3782
rect 15988 3780 16012 3782
rect 16068 3780 16092 3782
rect 16148 3780 16154 3782
rect 15846 3760 16154 3780
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 15580 2990 15608 3062
rect 15764 3058 15792 3538
rect 16316 3534 16344 4422
rect 16408 3942 16436 4422
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16592 3126 16620 4490
rect 16684 4282 16712 5102
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16776 3738 16804 6734
rect 16868 5642 16896 6734
rect 16960 5778 16988 6802
rect 17420 6798 17448 9998
rect 17788 9674 17816 11698
rect 17972 11150 18000 13874
rect 18064 13530 18092 14350
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18156 11898 18184 14418
rect 18248 13394 18276 14418
rect 18328 14408 18380 14414
rect 18326 14376 18328 14385
rect 18380 14376 18382 14385
rect 18326 14311 18382 14320
rect 18328 13728 18380 13734
rect 18326 13696 18328 13705
rect 18380 13696 18382 13705
rect 18326 13631 18382 13640
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18432 12850 18460 21422
rect 18524 12866 18552 23174
rect 18616 23050 18644 23598
rect 18708 23186 18736 26862
rect 18892 24936 18920 28086
rect 18972 25900 19024 25906
rect 18972 25842 19024 25848
rect 18800 24908 18920 24936
rect 18800 24206 18828 24908
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18696 22228 18748 22234
rect 18696 22170 18748 22176
rect 18602 21720 18658 21729
rect 18602 21655 18658 21664
rect 18616 21622 18644 21655
rect 18604 21616 18656 21622
rect 18604 21558 18656 21564
rect 18708 21418 18736 22170
rect 18696 21412 18748 21418
rect 18696 21354 18748 21360
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 18708 20466 18736 20878
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18616 19310 18644 20334
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 18708 18970 18736 20402
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18800 17728 18828 24006
rect 18892 22982 18920 24754
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18880 22568 18932 22574
rect 18880 22510 18932 22516
rect 18892 21486 18920 22510
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18892 21010 18920 21422
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 18880 20800 18932 20806
rect 18880 20742 18932 20748
rect 18892 19990 18920 20742
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 18984 19514 19012 25842
rect 19076 23089 19104 31726
rect 19248 30796 19300 30802
rect 19248 30738 19300 30744
rect 19156 30252 19208 30258
rect 19156 30194 19208 30200
rect 19168 29782 19196 30194
rect 19156 29776 19208 29782
rect 19156 29718 19208 29724
rect 19156 24744 19208 24750
rect 19156 24686 19208 24692
rect 19168 24206 19196 24686
rect 19156 24200 19208 24206
rect 19156 24142 19208 24148
rect 19168 23254 19196 24142
rect 19156 23248 19208 23254
rect 19156 23190 19208 23196
rect 19156 23112 19208 23118
rect 19062 23080 19118 23089
rect 19156 23054 19208 23060
rect 19062 23015 19118 23024
rect 19076 22234 19104 23015
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 19076 21554 19104 21830
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18984 18426 19012 19450
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18616 17700 18828 17728
rect 18616 16250 18644 17700
rect 19168 17626 19196 23054
rect 19260 21729 19288 30738
rect 19352 30326 19380 33458
rect 19444 32910 19472 34070
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19444 29714 19472 30534
rect 19536 30394 19564 34614
rect 19628 32994 19656 36246
rect 19812 35698 19840 36518
rect 19892 36168 19944 36174
rect 19892 36110 19944 36116
rect 19800 35692 19852 35698
rect 19800 35634 19852 35640
rect 19708 34944 19760 34950
rect 19708 34886 19760 34892
rect 19720 34610 19748 34886
rect 19708 34604 19760 34610
rect 19708 34546 19760 34552
rect 19800 34604 19852 34610
rect 19800 34546 19852 34552
rect 19812 33318 19840 34546
rect 19904 33998 19932 36110
rect 19996 36038 20024 36586
rect 20088 36174 20116 37130
rect 20076 36168 20128 36174
rect 20076 36110 20128 36116
rect 19984 36032 20036 36038
rect 19984 35974 20036 35980
rect 19996 34610 20024 35974
rect 20168 35692 20220 35698
rect 20168 35634 20220 35640
rect 20180 35222 20208 35634
rect 20168 35216 20220 35222
rect 20168 35158 20220 35164
rect 20272 35170 20300 38694
rect 21560 38282 21588 39238
rect 21548 38276 21600 38282
rect 21548 38218 21600 38224
rect 20811 38108 21119 38128
rect 20811 38106 20817 38108
rect 20873 38106 20897 38108
rect 20953 38106 20977 38108
rect 21033 38106 21057 38108
rect 21113 38106 21119 38108
rect 20873 38054 20875 38106
rect 21055 38054 21057 38106
rect 20811 38052 20817 38054
rect 20873 38052 20897 38054
rect 20953 38052 20977 38054
rect 21033 38052 21057 38054
rect 21113 38052 21119 38054
rect 20811 38032 21119 38052
rect 20720 37936 20772 37942
rect 20720 37878 20772 37884
rect 20352 37664 20404 37670
rect 20352 37606 20404 37612
rect 20364 37262 20392 37606
rect 20352 37256 20404 37262
rect 20352 37198 20404 37204
rect 20352 37120 20404 37126
rect 20352 37062 20404 37068
rect 20364 36174 20392 37062
rect 20444 36848 20496 36854
rect 20444 36790 20496 36796
rect 20352 36168 20404 36174
rect 20352 36110 20404 36116
rect 20364 35698 20392 36110
rect 20456 35834 20484 36790
rect 20536 36780 20588 36786
rect 20536 36722 20588 36728
rect 20444 35828 20496 35834
rect 20444 35770 20496 35776
rect 20352 35692 20404 35698
rect 20352 35634 20404 35640
rect 20364 35290 20392 35634
rect 20352 35284 20404 35290
rect 20352 35226 20404 35232
rect 20180 35086 20208 35158
rect 20272 35142 20392 35170
rect 20456 35154 20484 35770
rect 20548 35766 20576 36722
rect 20628 36712 20680 36718
rect 20628 36654 20680 36660
rect 20640 36378 20668 36654
rect 20628 36372 20680 36378
rect 20628 36314 20680 36320
rect 20536 35760 20588 35766
rect 20536 35702 20588 35708
rect 20628 35488 20680 35494
rect 20628 35430 20680 35436
rect 20640 35154 20668 35430
rect 20168 35080 20220 35086
rect 20168 35022 20220 35028
rect 20076 34944 20128 34950
rect 20076 34886 20128 34892
rect 19984 34604 20036 34610
rect 19984 34546 20036 34552
rect 19984 34468 20036 34474
rect 19984 34410 20036 34416
rect 19892 33992 19944 33998
rect 19892 33934 19944 33940
rect 19904 33658 19932 33934
rect 19892 33652 19944 33658
rect 19892 33594 19944 33600
rect 19800 33312 19852 33318
rect 19800 33254 19852 33260
rect 19812 33114 19840 33254
rect 19800 33108 19852 33114
rect 19800 33050 19852 33056
rect 19628 32966 19748 32994
rect 19904 32978 19932 33594
rect 19616 32904 19668 32910
rect 19616 32846 19668 32852
rect 19720 32858 19748 32966
rect 19892 32972 19944 32978
rect 19892 32914 19944 32920
rect 19628 32434 19656 32846
rect 19720 32830 19840 32858
rect 19708 32564 19760 32570
rect 19708 32506 19760 32512
rect 19616 32428 19668 32434
rect 19616 32370 19668 32376
rect 19720 31754 19748 32506
rect 19812 32502 19840 32830
rect 19800 32496 19852 32502
rect 19800 32438 19852 32444
rect 19904 32230 19932 32914
rect 19892 32224 19944 32230
rect 19892 32166 19944 32172
rect 19996 32042 20024 34410
rect 19904 32014 20024 32042
rect 19720 31726 19840 31754
rect 19708 31204 19760 31210
rect 19708 31146 19760 31152
rect 19524 30388 19576 30394
rect 19524 30330 19576 30336
rect 19432 29708 19484 29714
rect 19432 29650 19484 29656
rect 19432 29572 19484 29578
rect 19432 29514 19484 29520
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 19352 24426 19380 29446
rect 19444 29170 19472 29514
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19444 28694 19472 29106
rect 19616 28960 19668 28966
rect 19616 28902 19668 28908
rect 19432 28688 19484 28694
rect 19432 28630 19484 28636
rect 19524 28008 19576 28014
rect 19524 27950 19576 27956
rect 19432 27872 19484 27878
rect 19432 27814 19484 27820
rect 19444 27470 19472 27814
rect 19536 27606 19564 27950
rect 19628 27674 19656 28902
rect 19616 27668 19668 27674
rect 19616 27610 19668 27616
rect 19524 27600 19576 27606
rect 19524 27542 19576 27548
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19444 26790 19472 27406
rect 19628 27384 19656 27610
rect 19536 27356 19656 27384
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19444 26466 19472 26726
rect 19536 26586 19564 27356
rect 19720 27282 19748 31146
rect 19812 29170 19840 31726
rect 19800 29164 19852 29170
rect 19800 29106 19852 29112
rect 19812 27674 19840 29106
rect 19904 28994 19932 32014
rect 19984 31884 20036 31890
rect 19984 31826 20036 31832
rect 19996 31414 20024 31826
rect 19984 31408 20036 31414
rect 19984 31350 20036 31356
rect 20088 30546 20116 34886
rect 20180 33522 20208 35022
rect 20260 34536 20312 34542
rect 20260 34478 20312 34484
rect 20168 33516 20220 33522
rect 20168 33458 20220 33464
rect 20180 32910 20208 33458
rect 20168 32904 20220 32910
rect 20168 32846 20220 32852
rect 20180 31346 20208 32846
rect 20272 32570 20300 34478
rect 20260 32564 20312 32570
rect 20260 32506 20312 32512
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 20272 30802 20300 32506
rect 20260 30796 20312 30802
rect 20260 30738 20312 30744
rect 19996 30518 20116 30546
rect 19996 29730 20024 30518
rect 20076 30388 20128 30394
rect 20076 30330 20128 30336
rect 20088 29850 20116 30330
rect 20272 30190 20300 30738
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 20168 30116 20220 30122
rect 20168 30058 20220 30064
rect 20076 29844 20128 29850
rect 20076 29786 20128 29792
rect 19996 29702 20116 29730
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19996 29238 20024 29582
rect 19984 29232 20036 29238
rect 19984 29174 20036 29180
rect 19904 28966 20024 28994
rect 19996 27826 20024 28966
rect 19904 27798 20024 27826
rect 19800 27668 19852 27674
rect 19800 27610 19852 27616
rect 19800 27532 19852 27538
rect 19800 27474 19852 27480
rect 19628 27254 19748 27282
rect 19524 26580 19576 26586
rect 19524 26522 19576 26528
rect 19444 26438 19564 26466
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 19444 25226 19472 26318
rect 19536 25974 19564 26438
rect 19524 25968 19576 25974
rect 19524 25910 19576 25916
rect 19524 25832 19576 25838
rect 19524 25774 19576 25780
rect 19536 25294 19564 25774
rect 19628 25702 19656 27254
rect 19708 26376 19760 26382
rect 19708 26318 19760 26324
rect 19616 25696 19668 25702
rect 19616 25638 19668 25644
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19352 24398 19472 24426
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 19352 24070 19380 24278
rect 19444 24138 19472 24398
rect 19432 24132 19484 24138
rect 19432 24074 19484 24080
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19352 22098 19380 24006
rect 19536 23662 19564 25230
rect 19628 24954 19656 25638
rect 19720 25498 19748 26318
rect 19812 25974 19840 27474
rect 19904 26518 19932 27798
rect 19984 27668 20036 27674
rect 19984 27610 20036 27616
rect 19892 26512 19944 26518
rect 19892 26454 19944 26460
rect 19892 26376 19944 26382
rect 19892 26318 19944 26324
rect 19904 26042 19932 26318
rect 19892 26036 19944 26042
rect 19892 25978 19944 25984
rect 19800 25968 19852 25974
rect 19800 25910 19852 25916
rect 19800 25832 19852 25838
rect 19800 25774 19852 25780
rect 19708 25492 19760 25498
rect 19708 25434 19760 25440
rect 19720 25294 19748 25434
rect 19708 25288 19760 25294
rect 19708 25230 19760 25236
rect 19616 24948 19668 24954
rect 19616 24890 19668 24896
rect 19812 24410 19840 25774
rect 19904 24818 19932 25978
rect 19996 25809 20024 27610
rect 20088 27606 20116 29702
rect 20076 27600 20128 27606
rect 20076 27542 20128 27548
rect 19982 25800 20038 25809
rect 19982 25735 20038 25744
rect 19984 25696 20036 25702
rect 19984 25638 20036 25644
rect 19996 25362 20024 25638
rect 19984 25356 20036 25362
rect 19984 25298 20036 25304
rect 20088 25226 20116 27542
rect 20076 25220 20128 25226
rect 20076 25162 20128 25168
rect 19892 24812 19944 24818
rect 19892 24754 19944 24760
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19708 24404 19760 24410
rect 19708 24346 19760 24352
rect 19800 24404 19852 24410
rect 19800 24346 19852 24352
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 19628 23662 19656 24142
rect 19720 24070 19748 24346
rect 19708 24064 19760 24070
rect 19708 24006 19760 24012
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19524 23656 19576 23662
rect 19524 23598 19576 23604
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19524 23112 19576 23118
rect 19524 23054 19576 23060
rect 19536 22506 19564 23054
rect 19720 22760 19748 23802
rect 19812 23730 19840 24346
rect 19996 24274 20024 24550
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19800 23724 19852 23730
rect 19800 23666 19852 23672
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19720 22732 19840 22760
rect 19708 22636 19760 22642
rect 19708 22578 19760 22584
rect 19524 22500 19576 22506
rect 19524 22442 19576 22448
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 19444 22166 19472 22374
rect 19432 22160 19484 22166
rect 19432 22102 19484 22108
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19246 21720 19302 21729
rect 19246 21655 19302 21664
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19352 21146 19380 21490
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19444 20602 19472 21626
rect 19536 21078 19564 22442
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19628 21554 19656 22374
rect 19616 21548 19668 21554
rect 19616 21490 19668 21496
rect 19720 21146 19748 22578
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 19616 20868 19668 20874
rect 19616 20810 19668 20816
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 19352 19922 19380 20266
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19352 19446 19380 19858
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19260 17814 19288 19314
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19352 18834 19380 19246
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19352 17882 19380 18226
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19248 17808 19300 17814
rect 19248 17750 19300 17756
rect 18892 17598 19196 17626
rect 18694 16280 18750 16289
rect 18604 16244 18656 16250
rect 18694 16215 18696 16224
rect 18604 16186 18656 16192
rect 18748 16215 18750 16224
rect 18696 16186 18748 16192
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18616 16017 18644 16050
rect 18602 16008 18658 16017
rect 18602 15943 18658 15952
rect 18604 15632 18656 15638
rect 18604 15574 18656 15580
rect 18616 14414 18644 15574
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18616 14074 18644 14214
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18524 12850 18644 12866
rect 18420 12844 18472 12850
rect 18524 12844 18656 12850
rect 18524 12838 18604 12844
rect 18420 12786 18472 12792
rect 18604 12786 18656 12792
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18248 11830 18276 12174
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18052 11620 18104 11626
rect 18052 11562 18104 11568
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 18064 10810 18092 11562
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17696 9646 17816 9674
rect 17696 8906 17724 9646
rect 17880 9110 17908 10406
rect 18236 10192 18288 10198
rect 18236 10134 18288 10140
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18156 9586 18184 9862
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17684 8900 17736 8906
rect 17684 8842 17736 8848
rect 17788 8430 17816 9046
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17972 8106 18000 8910
rect 18248 8838 18276 10134
rect 18432 9722 18460 12786
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11898 18552 12038
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18708 10130 18736 16186
rect 18788 13932 18840 13938
rect 18892 13920 18920 17598
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18984 16114 19012 16934
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 18984 15094 19012 16050
rect 19260 16046 19288 17138
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16794 19380 16934
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19352 16046 19380 16594
rect 19444 16590 19472 20198
rect 19628 19242 19656 20810
rect 19616 19236 19668 19242
rect 19616 19178 19668 19184
rect 19720 18766 19748 21082
rect 19812 20942 19840 22732
rect 19904 22710 19932 23666
rect 19892 22704 19944 22710
rect 19892 22646 19944 22652
rect 19892 21616 19944 21622
rect 19892 21558 19944 21564
rect 19904 21350 19932 21558
rect 19892 21344 19944 21350
rect 19892 21286 19944 21292
rect 19800 20936 19852 20942
rect 19852 20896 19932 20924
rect 19800 20878 19852 20884
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 19708 18760 19760 18766
rect 19628 18720 19708 18748
rect 19628 18426 19656 18720
rect 19708 18702 19760 18708
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19720 18290 19748 18566
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19536 16402 19564 17614
rect 19628 17202 19656 17682
rect 19720 17610 19748 18226
rect 19708 17604 19760 17610
rect 19708 17546 19760 17552
rect 19812 17270 19840 20402
rect 19904 19854 19932 20896
rect 19996 20398 20024 24210
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19996 17814 20024 18022
rect 19984 17808 20036 17814
rect 19984 17750 20036 17756
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19628 16454 19656 17138
rect 19892 17128 19944 17134
rect 19812 17088 19892 17116
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19720 16590 19748 17002
rect 19812 16726 19840 17088
rect 19892 17070 19944 17076
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 19800 16720 19852 16726
rect 19800 16662 19852 16668
rect 19699 16584 19751 16590
rect 19699 16526 19751 16532
rect 19444 16374 19564 16402
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19064 15972 19116 15978
rect 19064 15914 19116 15920
rect 19076 15881 19104 15914
rect 19062 15872 19118 15881
rect 19062 15807 19118 15816
rect 19260 15434 19288 15982
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 18972 15088 19024 15094
rect 18972 15030 19024 15036
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19168 14006 19196 14758
rect 19352 14006 19380 15982
rect 19444 15502 19472 16374
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19536 13938 19564 15846
rect 19628 15502 19656 16390
rect 19720 15978 19748 16526
rect 19708 15972 19760 15978
rect 19708 15914 19760 15920
rect 19720 15638 19748 15914
rect 19708 15632 19760 15638
rect 19708 15574 19760 15580
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19812 15162 19840 16662
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19904 15910 19932 16526
rect 19996 16182 20024 16934
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19904 15502 19932 15846
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 18840 13892 18920 13920
rect 19524 13932 19576 13938
rect 18788 13874 18840 13880
rect 19524 13874 19576 13880
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19892 13456 19944 13462
rect 19892 13398 19944 13404
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19352 12986 19380 13262
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19076 12170 19104 12922
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19064 12164 19116 12170
rect 19064 12106 19116 12112
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18800 10062 18828 10610
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18328 8968 18380 8974
rect 18380 8916 18644 8922
rect 18328 8910 18644 8916
rect 18340 8894 18644 8910
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18156 8634 18184 8774
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 17972 8078 18092 8106
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17512 6798 17540 7754
rect 17972 7410 18000 7958
rect 18064 7886 18092 8078
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 18156 6934 18184 7414
rect 18248 7188 18276 8774
rect 18432 7478 18460 8774
rect 18616 8378 18644 8894
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18800 8498 18828 8774
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18616 8350 18828 8378
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18328 7200 18380 7206
rect 18248 7160 18328 7188
rect 18328 7142 18380 7148
rect 18340 7002 18368 7142
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18144 6928 18196 6934
rect 18144 6870 18196 6876
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17328 6322 17356 6598
rect 17420 6458 17448 6734
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 17512 5710 17540 6734
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 18064 5710 18092 6394
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18248 5914 18276 6258
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16868 3466 16896 4626
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 16948 4548 17000 4554
rect 16948 4490 17000 4496
rect 16960 4010 16988 4490
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16960 3738 16988 3946
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16488 3120 16540 3126
rect 16486 3088 16488 3097
rect 16580 3120 16632 3126
rect 16540 3088 16542 3097
rect 15752 3052 15804 3058
rect 16580 3062 16632 3068
rect 16486 3023 16542 3032
rect 15752 2994 15804 3000
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15580 2650 15608 2926
rect 16684 2854 16712 3402
rect 16960 2922 16988 3674
rect 17052 3670 17080 4558
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 17052 3058 17080 3606
rect 17144 3534 17172 4966
rect 17328 3602 17356 5170
rect 17512 4622 17540 5646
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17420 3602 17448 4014
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17222 3496 17278 3505
rect 17222 3431 17278 3440
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17144 3194 17172 3334
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17236 2922 17264 3431
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 15846 2748 16154 2768
rect 15846 2746 15852 2748
rect 15908 2746 15932 2748
rect 15988 2746 16012 2748
rect 16068 2746 16092 2748
rect 16148 2746 16154 2748
rect 15908 2694 15910 2746
rect 16090 2694 16092 2746
rect 15846 2692 15852 2694
rect 15908 2692 15932 2694
rect 15988 2692 16012 2694
rect 16068 2692 16092 2694
rect 16148 2692 16154 2694
rect 15846 2672 16154 2692
rect 16684 2650 16712 2790
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16776 2514 16804 2858
rect 17328 2774 17356 3538
rect 17696 3194 17724 5646
rect 18236 5636 18288 5642
rect 18236 5578 18288 5584
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17972 4826 18000 5102
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 18248 4690 18276 5578
rect 18800 5166 18828 8350
rect 18892 6458 18920 11086
rect 19076 10470 19104 12106
rect 19536 11762 19564 12582
rect 19628 12374 19656 13330
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19812 12434 19840 12922
rect 19904 12782 19932 13398
rect 19996 13326 20024 13806
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19892 12776 19944 12782
rect 19892 12718 19944 12724
rect 19812 12406 19932 12434
rect 19616 12368 19668 12374
rect 19616 12310 19668 12316
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19260 9722 19288 9998
rect 19248 9716 19300 9722
rect 19248 9658 19300 9664
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19156 8900 19208 8906
rect 19156 8842 19208 8848
rect 19168 8294 19196 8842
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19260 6458 19288 8978
rect 19628 8634 19656 12174
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19444 6730 19472 7278
rect 19628 6866 19656 7278
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19432 6724 19484 6730
rect 19432 6666 19484 6672
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17972 3194 18000 3538
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 17866 3088 17922 3097
rect 17866 3023 17922 3032
rect 17960 3052 18012 3058
rect 17328 2746 17448 2774
rect 16764 2508 16816 2514
rect 16764 2450 16816 2456
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 15580 800 15608 2382
rect 16408 800 16436 2382
rect 17144 800 17172 2450
rect 17420 2446 17448 2746
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17880 800 17908 3023
rect 17960 2994 18012 3000
rect 17972 2650 18000 2994
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 18064 2446 18092 2926
rect 18156 2854 18184 4558
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18340 3534 18368 4082
rect 18432 3738 18460 4150
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18340 2582 18368 3470
rect 18524 3194 18552 4966
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18616 2774 18644 5034
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18708 4214 18736 4422
rect 18696 4208 18748 4214
rect 18696 4150 18748 4156
rect 18524 2746 18644 2774
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 18524 2446 18552 2746
rect 18604 2576 18656 2582
rect 18604 2518 18656 2524
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18616 800 18644 2518
rect 18800 2446 18828 5102
rect 19260 3194 19288 5170
rect 19352 3942 19380 6326
rect 19444 5778 19472 6666
rect 19432 5772 19484 5778
rect 19432 5714 19484 5720
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19444 4146 19472 4626
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19444 3534 19472 4082
rect 19536 4010 19564 6734
rect 19720 5914 19748 11630
rect 19812 11150 19840 12038
rect 19904 11830 19932 12406
rect 20088 12170 20116 25162
rect 20180 23610 20208 30058
rect 20272 29578 20300 30126
rect 20260 29572 20312 29578
rect 20260 29514 20312 29520
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20272 26994 20300 27406
rect 20260 26988 20312 26994
rect 20260 26930 20312 26936
rect 20260 26852 20312 26858
rect 20260 26794 20312 26800
rect 20272 23730 20300 26794
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20180 23594 20300 23610
rect 20180 23588 20312 23594
rect 20180 23582 20260 23588
rect 20260 23530 20312 23536
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20180 23322 20208 23462
rect 20168 23316 20220 23322
rect 20168 23258 20220 23264
rect 20272 21010 20300 23530
rect 20364 22778 20392 35142
rect 20444 35148 20496 35154
rect 20444 35090 20496 35096
rect 20628 35148 20680 35154
rect 20628 35090 20680 35096
rect 20456 34490 20484 35090
rect 20456 34462 20576 34490
rect 20444 34400 20496 34406
rect 20444 34342 20496 34348
rect 20456 34134 20484 34342
rect 20444 34128 20496 34134
rect 20444 34070 20496 34076
rect 20548 33114 20576 34462
rect 20640 33998 20668 35090
rect 20732 34202 20760 37878
rect 22020 37874 22048 39306
rect 22008 37868 22060 37874
rect 22008 37810 22060 37816
rect 20811 37020 21119 37040
rect 20811 37018 20817 37020
rect 20873 37018 20897 37020
rect 20953 37018 20977 37020
rect 21033 37018 21057 37020
rect 21113 37018 21119 37020
rect 20873 36966 20875 37018
rect 21055 36966 21057 37018
rect 20811 36964 20817 36966
rect 20873 36964 20897 36966
rect 20953 36964 20977 36966
rect 21033 36964 21057 36966
rect 21113 36964 21119 36966
rect 20811 36944 21119 36964
rect 22020 36786 22048 37810
rect 21364 36780 21416 36786
rect 21364 36722 21416 36728
rect 22008 36780 22060 36786
rect 22008 36722 22060 36728
rect 20812 36576 20864 36582
rect 20812 36518 20864 36524
rect 20824 36242 20852 36518
rect 21376 36242 21404 36722
rect 20812 36236 20864 36242
rect 20812 36178 20864 36184
rect 21364 36236 21416 36242
rect 21364 36178 21416 36184
rect 21548 36168 21600 36174
rect 21548 36110 21600 36116
rect 20811 35932 21119 35952
rect 20811 35930 20817 35932
rect 20873 35930 20897 35932
rect 20953 35930 20977 35932
rect 21033 35930 21057 35932
rect 21113 35930 21119 35932
rect 20873 35878 20875 35930
rect 21055 35878 21057 35930
rect 20811 35876 20817 35878
rect 20873 35876 20897 35878
rect 20953 35876 20977 35878
rect 21033 35876 21057 35878
rect 21113 35876 21119 35878
rect 20811 35856 21119 35876
rect 21560 35698 21588 36110
rect 21548 35692 21600 35698
rect 21548 35634 21600 35640
rect 20811 34844 21119 34864
rect 20811 34842 20817 34844
rect 20873 34842 20897 34844
rect 20953 34842 20977 34844
rect 21033 34842 21057 34844
rect 21113 34842 21119 34844
rect 20873 34790 20875 34842
rect 21055 34790 21057 34842
rect 20811 34788 20817 34790
rect 20873 34788 20897 34790
rect 20953 34788 20977 34790
rect 21033 34788 21057 34790
rect 21113 34788 21119 34790
rect 20811 34768 21119 34788
rect 20720 34196 20772 34202
rect 20720 34138 20772 34144
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 21180 33924 21232 33930
rect 21180 33866 21232 33872
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20732 33658 20760 33798
rect 20811 33756 21119 33776
rect 20811 33754 20817 33756
rect 20873 33754 20897 33756
rect 20953 33754 20977 33756
rect 21033 33754 21057 33756
rect 21113 33754 21119 33756
rect 20873 33702 20875 33754
rect 21055 33702 21057 33754
rect 20811 33700 20817 33702
rect 20873 33700 20897 33702
rect 20953 33700 20977 33702
rect 21033 33700 21057 33702
rect 21113 33700 21119 33702
rect 20811 33680 21119 33700
rect 20720 33652 20772 33658
rect 20720 33594 20772 33600
rect 21192 33590 21220 33866
rect 21272 33856 21324 33862
rect 21272 33798 21324 33804
rect 21284 33658 21312 33798
rect 21272 33652 21324 33658
rect 21272 33594 21324 33600
rect 20812 33584 20864 33590
rect 20812 33526 20864 33532
rect 21180 33584 21232 33590
rect 21180 33526 21232 33532
rect 20444 33108 20496 33114
rect 20444 33050 20496 33056
rect 20536 33108 20588 33114
rect 20536 33050 20588 33056
rect 20456 32586 20484 33050
rect 20548 32774 20576 33050
rect 20628 32836 20680 32842
rect 20628 32778 20680 32784
rect 20536 32768 20588 32774
rect 20536 32710 20588 32716
rect 20456 32558 20576 32586
rect 20444 32428 20496 32434
rect 20444 32370 20496 32376
rect 20456 31754 20484 32370
rect 20548 32298 20576 32558
rect 20640 32502 20668 32778
rect 20720 32768 20772 32774
rect 20824 32756 20852 33526
rect 21456 33516 21508 33522
rect 21456 33458 21508 33464
rect 20772 32728 20852 32756
rect 21364 32768 21416 32774
rect 20720 32710 20772 32716
rect 21364 32710 21416 32716
rect 20628 32496 20680 32502
rect 20628 32438 20680 32444
rect 20732 32366 20760 32710
rect 20811 32668 21119 32688
rect 20811 32666 20817 32668
rect 20873 32666 20897 32668
rect 20953 32666 20977 32668
rect 21033 32666 21057 32668
rect 21113 32666 21119 32668
rect 20873 32614 20875 32666
rect 21055 32614 21057 32666
rect 20811 32612 20817 32614
rect 20873 32612 20897 32614
rect 20953 32612 20977 32614
rect 21033 32612 21057 32614
rect 21113 32612 21119 32614
rect 20811 32592 21119 32612
rect 21376 32502 21404 32710
rect 21364 32496 21416 32502
rect 21364 32438 21416 32444
rect 21272 32428 21324 32434
rect 21272 32370 21324 32376
rect 20720 32360 20772 32366
rect 20720 32302 20772 32308
rect 21180 32360 21232 32366
rect 21180 32302 21232 32308
rect 20536 32292 20588 32298
rect 20536 32234 20588 32240
rect 20732 32042 20760 32302
rect 20904 32224 20956 32230
rect 20904 32166 20956 32172
rect 20640 32014 20760 32042
rect 20640 31822 20668 32014
rect 20916 31890 20944 32166
rect 20720 31884 20772 31890
rect 20720 31826 20772 31832
rect 20904 31884 20956 31890
rect 20904 31826 20956 31832
rect 20628 31816 20680 31822
rect 20628 31758 20680 31764
rect 20444 31748 20496 31754
rect 20444 31690 20496 31696
rect 20456 31210 20484 31690
rect 20444 31204 20496 31210
rect 20444 31146 20496 31152
rect 20456 29102 20484 31146
rect 20536 31136 20588 31142
rect 20536 31078 20588 31084
rect 20548 30802 20576 31078
rect 20732 30870 20760 31826
rect 21192 31754 21220 32302
rect 21284 31890 21312 32370
rect 21272 31884 21324 31890
rect 21272 31826 21324 31832
rect 21468 31754 21496 33458
rect 21088 31748 21220 31754
rect 21140 31726 21220 31748
rect 21088 31690 21140 31696
rect 20811 31580 21119 31600
rect 20811 31578 20817 31580
rect 20873 31578 20897 31580
rect 20953 31578 20977 31580
rect 21033 31578 21057 31580
rect 21113 31578 21119 31580
rect 20873 31526 20875 31578
rect 21055 31526 21057 31578
rect 20811 31524 20817 31526
rect 20873 31524 20897 31526
rect 20953 31524 20977 31526
rect 21033 31524 21057 31526
rect 21113 31524 21119 31526
rect 20811 31504 21119 31524
rect 20720 30864 20772 30870
rect 20720 30806 20772 30812
rect 20536 30796 20588 30802
rect 20536 30738 20588 30744
rect 20548 30326 20576 30738
rect 20536 30320 20588 30326
rect 20536 30262 20588 30268
rect 20732 30258 20760 30806
rect 21192 30666 21220 31726
rect 21284 31726 21496 31754
rect 21180 30660 21232 30666
rect 21180 30602 21232 30608
rect 20811 30492 21119 30512
rect 20811 30490 20817 30492
rect 20873 30490 20897 30492
rect 20953 30490 20977 30492
rect 21033 30490 21057 30492
rect 21113 30490 21119 30492
rect 20873 30438 20875 30490
rect 21055 30438 21057 30490
rect 20811 30436 20817 30438
rect 20873 30436 20897 30438
rect 20953 30436 20977 30438
rect 21033 30436 21057 30438
rect 21113 30436 21119 30438
rect 20811 30416 21119 30436
rect 20720 30252 20772 30258
rect 20720 30194 20772 30200
rect 20811 29404 21119 29424
rect 20811 29402 20817 29404
rect 20873 29402 20897 29404
rect 20953 29402 20977 29404
rect 21033 29402 21057 29404
rect 21113 29402 21119 29404
rect 20873 29350 20875 29402
rect 21055 29350 21057 29402
rect 20811 29348 20817 29350
rect 20873 29348 20897 29350
rect 20953 29348 20977 29350
rect 21033 29348 21057 29350
rect 21113 29348 21119 29350
rect 20811 29328 21119 29348
rect 20444 29096 20496 29102
rect 20444 29038 20496 29044
rect 20456 28082 20484 29038
rect 21192 28762 21220 30602
rect 21284 30054 21312 31726
rect 21272 30048 21324 30054
rect 21272 29990 21324 29996
rect 21284 29170 21312 29990
rect 21560 29714 21588 35634
rect 21640 33992 21692 33998
rect 21640 33934 21692 33940
rect 21652 32570 21680 33934
rect 21824 33516 21876 33522
rect 21824 33458 21876 33464
rect 21836 33114 21864 33458
rect 21824 33108 21876 33114
rect 21824 33050 21876 33056
rect 21916 32836 21968 32842
rect 21916 32778 21968 32784
rect 21640 32564 21692 32570
rect 21640 32506 21692 32512
rect 21928 32230 21956 32778
rect 22192 32768 22244 32774
rect 22192 32710 22244 32716
rect 22204 32502 22232 32710
rect 22192 32496 22244 32502
rect 22192 32438 22244 32444
rect 21916 32224 21968 32230
rect 21916 32166 21968 32172
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 21928 31482 21956 31758
rect 21916 31476 21968 31482
rect 21916 31418 21968 31424
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 21652 30666 21680 31282
rect 21640 30660 21692 30666
rect 21640 30602 21692 30608
rect 21548 29708 21600 29714
rect 21548 29650 21600 29656
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 21468 29238 21496 29582
rect 21560 29306 21588 29650
rect 21652 29578 21680 30602
rect 21916 29776 21968 29782
rect 21916 29718 21968 29724
rect 21640 29572 21692 29578
rect 21640 29514 21692 29520
rect 21548 29300 21600 29306
rect 21548 29242 21600 29248
rect 21456 29232 21508 29238
rect 21456 29174 21508 29180
rect 21272 29164 21324 29170
rect 21272 29106 21324 29112
rect 21180 28756 21232 28762
rect 21180 28698 21232 28704
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20640 28218 20668 28494
rect 20720 28484 20772 28490
rect 20720 28426 20772 28432
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 20444 28076 20496 28082
rect 20444 28018 20496 28024
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 20536 27940 20588 27946
rect 20536 27882 20588 27888
rect 20548 27674 20576 27882
rect 20536 27668 20588 27674
rect 20536 27610 20588 27616
rect 20640 27010 20668 28018
rect 20548 26982 20668 27010
rect 20548 26858 20576 26982
rect 20628 26920 20680 26926
rect 20628 26862 20680 26868
rect 20536 26852 20588 26858
rect 20536 26794 20588 26800
rect 20444 26580 20496 26586
rect 20444 26522 20496 26528
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20456 22030 20484 26522
rect 20640 26382 20668 26862
rect 20732 26518 20760 28426
rect 20811 28316 21119 28336
rect 20811 28314 20817 28316
rect 20873 28314 20897 28316
rect 20953 28314 20977 28316
rect 21033 28314 21057 28316
rect 21113 28314 21119 28316
rect 20873 28262 20875 28314
rect 21055 28262 21057 28314
rect 20811 28260 20817 28262
rect 20873 28260 20897 28262
rect 20953 28260 20977 28262
rect 21033 28260 21057 28262
rect 21113 28260 21119 28262
rect 20811 28240 21119 28260
rect 21180 27940 21232 27946
rect 21180 27882 21232 27888
rect 20811 27228 21119 27248
rect 20811 27226 20817 27228
rect 20873 27226 20897 27228
rect 20953 27226 20977 27228
rect 21033 27226 21057 27228
rect 21113 27226 21119 27228
rect 20873 27174 20875 27226
rect 21055 27174 21057 27226
rect 20811 27172 20817 27174
rect 20873 27172 20897 27174
rect 20953 27172 20977 27174
rect 21033 27172 21057 27174
rect 21113 27172 21119 27174
rect 20811 27152 21119 27172
rect 21088 27056 21140 27062
rect 21088 26998 21140 27004
rect 20720 26512 20772 26518
rect 20720 26454 20772 26460
rect 20536 26376 20588 26382
rect 20536 26318 20588 26324
rect 20628 26376 20680 26382
rect 20732 26353 20760 26454
rect 21100 26382 21128 26998
rect 21192 26790 21220 27882
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 21180 26444 21232 26450
rect 21180 26386 21232 26392
rect 21088 26376 21140 26382
rect 20628 26318 20680 26324
rect 20718 26344 20774 26353
rect 20548 25906 20576 26318
rect 21088 26318 21140 26324
rect 20718 26279 20774 26288
rect 20720 26240 20772 26246
rect 20720 26182 20772 26188
rect 20536 25900 20588 25906
rect 20536 25842 20588 25848
rect 20534 25800 20590 25809
rect 20534 25735 20590 25744
rect 20732 25752 20760 26182
rect 20811 26140 21119 26160
rect 20811 26138 20817 26140
rect 20873 26138 20897 26140
rect 20953 26138 20977 26140
rect 21033 26138 21057 26140
rect 21113 26138 21119 26140
rect 20873 26086 20875 26138
rect 21055 26086 21057 26138
rect 20811 26084 20817 26086
rect 20873 26084 20897 26086
rect 20953 26084 20977 26086
rect 21033 26084 21057 26086
rect 21113 26084 21119 26086
rect 20811 26064 21119 26084
rect 20810 25936 20866 25945
rect 20810 25871 20812 25880
rect 20864 25871 20866 25880
rect 21088 25900 21140 25906
rect 20812 25842 20864 25848
rect 21088 25842 21140 25848
rect 20812 25764 20864 25770
rect 20548 25362 20576 25735
rect 20732 25724 20812 25752
rect 20812 25706 20864 25712
rect 20628 25696 20680 25702
rect 20680 25656 20760 25684
rect 20628 25638 20680 25644
rect 20628 25492 20680 25498
rect 20628 25434 20680 25440
rect 20536 25356 20588 25362
rect 20536 25298 20588 25304
rect 20548 24274 20576 25298
rect 20640 24818 20668 25434
rect 20732 25294 20760 25656
rect 21100 25378 21128 25842
rect 21192 25498 21220 26386
rect 21180 25492 21232 25498
rect 21180 25434 21232 25440
rect 21100 25350 21220 25378
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20811 25052 21119 25072
rect 20811 25050 20817 25052
rect 20873 25050 20897 25052
rect 20953 25050 20977 25052
rect 21033 25050 21057 25052
rect 21113 25050 21119 25052
rect 20873 24998 20875 25050
rect 21055 24998 21057 25050
rect 20811 24996 20817 24998
rect 20873 24996 20897 24998
rect 20953 24996 20977 24998
rect 21033 24996 21057 24998
rect 21113 24996 21119 24998
rect 20811 24976 21119 24996
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20536 24268 20588 24274
rect 20536 24210 20588 24216
rect 20640 24206 20668 24754
rect 20720 24744 20772 24750
rect 20720 24686 20772 24692
rect 20628 24200 20680 24206
rect 20628 24142 20680 24148
rect 20536 24132 20588 24138
rect 20536 24074 20588 24080
rect 20548 23730 20576 24074
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20533 23724 20585 23730
rect 20533 23666 20585 23672
rect 20640 23338 20668 24006
rect 20732 23526 20760 24686
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 21100 24274 21128 24550
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 20811 23964 21119 23984
rect 20811 23962 20817 23964
rect 20873 23962 20897 23964
rect 20953 23962 20977 23964
rect 21033 23962 21057 23964
rect 21113 23962 21119 23964
rect 20873 23910 20875 23962
rect 21055 23910 21057 23962
rect 20811 23908 20817 23910
rect 20873 23908 20897 23910
rect 20953 23908 20977 23910
rect 21033 23908 21057 23910
rect 21113 23908 21119 23910
rect 20811 23888 21119 23908
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20640 23310 20760 23338
rect 21192 23322 21220 25350
rect 21284 24206 21312 29106
rect 21468 28082 21496 29174
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 21456 28076 21508 28082
rect 21456 28018 21508 28024
rect 21364 27464 21416 27470
rect 21364 27406 21416 27412
rect 21376 27130 21404 27406
rect 21364 27124 21416 27130
rect 21364 27066 21416 27072
rect 21560 26976 21588 28698
rect 21652 27470 21680 29514
rect 21824 29504 21876 29510
rect 21824 29446 21876 29452
rect 21732 29300 21784 29306
rect 21732 29242 21784 29248
rect 21640 27464 21692 27470
rect 21640 27406 21692 27412
rect 21468 26948 21588 26976
rect 21364 26376 21416 26382
rect 21364 26318 21416 26324
rect 21376 25974 21404 26318
rect 21364 25968 21416 25974
rect 21364 25910 21416 25916
rect 21468 24750 21496 26948
rect 21548 26784 21600 26790
rect 21548 26726 21600 26732
rect 21560 25226 21588 26726
rect 21548 25220 21600 25226
rect 21548 25162 21600 25168
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20444 22024 20496 22030
rect 20444 21966 20496 21972
rect 20456 21622 20484 21966
rect 20444 21616 20496 21622
rect 20444 21558 20496 21564
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20260 21004 20312 21010
rect 20260 20946 20312 20952
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 20180 20058 20208 20334
rect 20272 20058 20300 20946
rect 20364 20466 20392 21286
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20456 20330 20484 21422
rect 20548 21146 20576 21490
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20536 20868 20588 20874
rect 20536 20810 20588 20816
rect 20548 20466 20576 20810
rect 20640 20602 20668 23054
rect 20732 21010 20760 23310
rect 21180 23316 21232 23322
rect 21180 23258 21232 23264
rect 21376 23118 21404 24006
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21364 23112 21416 23118
rect 21364 23054 21416 23060
rect 20811 22876 21119 22896
rect 20811 22874 20817 22876
rect 20873 22874 20897 22876
rect 20953 22874 20977 22876
rect 21033 22874 21057 22876
rect 21113 22874 21119 22876
rect 20873 22822 20875 22874
rect 21055 22822 21057 22874
rect 20811 22820 20817 22822
rect 20873 22820 20897 22822
rect 20953 22820 20977 22822
rect 21033 22820 21057 22822
rect 21113 22820 21119 22822
rect 20811 22800 21119 22820
rect 20996 22704 21048 22710
rect 20996 22646 21048 22652
rect 21008 22098 21036 22646
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 21192 21962 21220 22578
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 20811 21788 21119 21808
rect 20811 21786 20817 21788
rect 20873 21786 20897 21788
rect 20953 21786 20977 21788
rect 21033 21786 21057 21788
rect 21113 21786 21119 21788
rect 20873 21734 20875 21786
rect 21055 21734 21057 21786
rect 20811 21732 20817 21734
rect 20873 21732 20897 21734
rect 20953 21732 20977 21734
rect 21033 21732 21057 21734
rect 21113 21732 21119 21734
rect 20811 21712 21119 21732
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20811 20700 21119 20720
rect 20811 20698 20817 20700
rect 20873 20698 20897 20700
rect 20953 20698 20977 20700
rect 21033 20698 21057 20700
rect 21113 20698 21119 20700
rect 20873 20646 20875 20698
rect 21055 20646 21057 20698
rect 20811 20644 20817 20646
rect 20873 20644 20897 20646
rect 20953 20644 20977 20646
rect 21033 20644 21057 20646
rect 21113 20644 21119 20646
rect 20811 20624 21119 20644
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20640 20346 20668 20538
rect 20444 20324 20496 20330
rect 20640 20318 20852 20346
rect 20444 20266 20496 20272
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20640 19446 20668 20198
rect 20824 19854 20852 20318
rect 21376 19938 21404 23054
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 21284 19910 21404 19938
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 21100 19786 21220 19802
rect 21088 19780 21220 19786
rect 21140 19774 21220 19780
rect 21088 19722 21140 19728
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20732 19514 20760 19654
rect 20811 19612 21119 19632
rect 20811 19610 20817 19612
rect 20873 19610 20897 19612
rect 20953 19610 20977 19612
rect 21033 19610 21057 19612
rect 21113 19610 21119 19612
rect 20873 19558 20875 19610
rect 21055 19558 21057 19610
rect 20811 19556 20817 19558
rect 20873 19556 20897 19558
rect 20953 19556 20977 19558
rect 21033 19556 21057 19558
rect 21113 19556 21119 19558
rect 20811 19536 21119 19556
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 20536 19236 20588 19242
rect 20536 19178 20588 19184
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20180 17678 20208 18226
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 20180 16658 20208 17614
rect 20272 17202 20300 19110
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20456 18426 20484 18702
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20548 18290 20576 19178
rect 20811 18524 21119 18544
rect 20811 18522 20817 18524
rect 20873 18522 20897 18524
rect 20953 18522 20977 18524
rect 21033 18522 21057 18524
rect 21113 18522 21119 18524
rect 20873 18470 20875 18522
rect 21055 18470 21057 18522
rect 20811 18468 20817 18470
rect 20873 18468 20897 18470
rect 20953 18468 20977 18470
rect 21033 18468 21057 18470
rect 21113 18468 21119 18470
rect 20811 18448 21119 18468
rect 21192 18290 21220 19774
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 20732 17882 20760 18226
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20811 17436 21119 17456
rect 20811 17434 20817 17436
rect 20873 17434 20897 17436
rect 20953 17434 20977 17436
rect 21033 17434 21057 17436
rect 21113 17434 21119 17436
rect 20873 17382 20875 17434
rect 21055 17382 21057 17434
rect 20811 17380 20817 17382
rect 20873 17380 20897 17382
rect 20953 17380 20977 17382
rect 21033 17380 21057 17382
rect 21113 17380 21119 17382
rect 20811 17360 21119 17380
rect 21284 17338 21312 19910
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21376 18970 21404 19790
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 20732 16590 20760 16934
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20272 16250 20300 16526
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20640 16114 20668 16526
rect 20811 16348 21119 16368
rect 20811 16346 20817 16348
rect 20873 16346 20897 16348
rect 20953 16346 20977 16348
rect 21033 16346 21057 16348
rect 21113 16346 21119 16348
rect 20873 16294 20875 16346
rect 21055 16294 21057 16346
rect 20811 16292 20817 16294
rect 20873 16292 20897 16294
rect 20953 16292 20977 16294
rect 21033 16292 21057 16294
rect 21113 16292 21119 16294
rect 20811 16272 21119 16292
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20444 15020 20496 15026
rect 20628 15020 20680 15026
rect 20444 14962 20496 14968
rect 20548 14980 20628 15008
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 20272 14346 20300 14894
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 20272 13326 20300 14282
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20260 13320 20312 13326
rect 20180 13280 20260 13308
rect 20180 12850 20208 13280
rect 20260 13262 20312 13268
rect 20364 12850 20392 13466
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 19892 11824 19944 11830
rect 19892 11766 19944 11772
rect 19904 11218 19932 11766
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 19996 11286 20024 11698
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 19904 10810 19932 11154
rect 20088 11150 20116 11630
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 19904 10266 19932 10610
rect 20088 10538 20116 11086
rect 20272 10826 20300 11086
rect 20180 10798 20300 10826
rect 20076 10532 20128 10538
rect 20076 10474 20128 10480
rect 19892 10260 19944 10266
rect 19892 10202 19944 10208
rect 20180 9178 20208 10798
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20272 9722 20300 10610
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 20364 9178 20392 11698
rect 20456 11354 20484 14962
rect 20548 14414 20576 14980
rect 20628 14962 20680 14968
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20536 14408 20588 14414
rect 20536 14350 20588 14356
rect 20548 13938 20576 14350
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20548 13462 20576 13874
rect 20536 13456 20588 13462
rect 20536 13398 20588 13404
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20548 11898 20576 13262
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20640 10810 20668 14418
rect 20732 14414 20760 15642
rect 20811 15260 21119 15280
rect 20811 15258 20817 15260
rect 20873 15258 20897 15260
rect 20953 15258 20977 15260
rect 21033 15258 21057 15260
rect 21113 15258 21119 15260
rect 20873 15206 20875 15258
rect 21055 15206 21057 15258
rect 20811 15204 20817 15206
rect 20873 15204 20897 15206
rect 20953 15204 20977 15206
rect 21033 15204 21057 15206
rect 21113 15204 21119 15206
rect 20811 15184 21119 15204
rect 21468 15026 21496 22170
rect 21560 21622 21588 23462
rect 21652 22030 21680 27406
rect 21744 27010 21772 29242
rect 21836 28626 21864 29446
rect 21928 28626 21956 29718
rect 22008 29096 22060 29102
rect 22008 29038 22060 29044
rect 22020 28694 22048 29038
rect 22008 28688 22060 28694
rect 22008 28630 22060 28636
rect 21824 28620 21876 28626
rect 21824 28562 21876 28568
rect 21916 28620 21968 28626
rect 21916 28562 21968 28568
rect 21916 28484 21968 28490
rect 21916 28426 21968 28432
rect 21824 28416 21876 28422
rect 21824 28358 21876 28364
rect 21836 28082 21864 28358
rect 21928 28218 21956 28426
rect 22192 28416 22244 28422
rect 22192 28358 22244 28364
rect 22204 28218 22232 28358
rect 21916 28212 21968 28218
rect 21916 28154 21968 28160
rect 22192 28212 22244 28218
rect 22192 28154 22244 28160
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 21836 27130 21864 28018
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 21744 26982 21864 27010
rect 21732 26920 21784 26926
rect 21732 26862 21784 26868
rect 21744 26450 21772 26862
rect 21732 26444 21784 26450
rect 21732 26386 21784 26392
rect 21744 25430 21772 26386
rect 21732 25424 21784 25430
rect 21732 25366 21784 25372
rect 21836 25362 21864 26982
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 21928 26042 21956 26930
rect 22008 26784 22060 26790
rect 22008 26726 22060 26732
rect 21916 26036 21968 26042
rect 21916 25978 21968 25984
rect 22020 25906 22048 26726
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 21824 25356 21876 25362
rect 21824 25298 21876 25304
rect 22020 24886 22048 25842
rect 22112 25838 22140 26930
rect 22192 26240 22244 26246
rect 22192 26182 22244 26188
rect 22100 25832 22152 25838
rect 22100 25774 22152 25780
rect 22204 25294 22232 26182
rect 22192 25288 22244 25294
rect 22192 25230 22244 25236
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 22008 24880 22060 24886
rect 22008 24822 22060 24828
rect 21916 24744 21968 24750
rect 21916 24686 21968 24692
rect 21928 24342 21956 24686
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 22020 24138 22048 24822
rect 22112 24138 22140 25162
rect 22204 24954 22232 25230
rect 22192 24948 22244 24954
rect 22192 24890 22244 24896
rect 22008 24132 22060 24138
rect 22008 24074 22060 24080
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 22008 22092 22060 22098
rect 22008 22034 22060 22040
rect 21640 22024 21692 22030
rect 21640 21966 21692 21972
rect 21824 21888 21876 21894
rect 21824 21830 21876 21836
rect 21548 21616 21600 21622
rect 21548 21558 21600 21564
rect 21560 15502 21588 21558
rect 21836 20806 21864 21830
rect 22020 21622 22048 22034
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22204 20534 22232 20742
rect 22296 20602 22324 39510
rect 30104 39432 30156 39438
rect 30102 39400 30104 39409
rect 30156 39400 30158 39409
rect 30102 39335 30158 39344
rect 25776 38652 26084 38672
rect 25776 38650 25782 38652
rect 25838 38650 25862 38652
rect 25918 38650 25942 38652
rect 25998 38650 26022 38652
rect 26078 38650 26084 38652
rect 25838 38598 25840 38650
rect 26020 38598 26022 38650
rect 25776 38596 25782 38598
rect 25838 38596 25862 38598
rect 25918 38596 25942 38598
rect 25998 38596 26022 38598
rect 26078 38596 26084 38598
rect 25776 38576 26084 38596
rect 30104 38344 30156 38350
rect 30104 38286 30156 38292
rect 29920 38208 29972 38214
rect 29920 38150 29972 38156
rect 29932 37806 29960 38150
rect 30116 37913 30144 38286
rect 30102 37904 30158 37913
rect 30102 37839 30158 37848
rect 29920 37800 29972 37806
rect 29920 37742 29972 37748
rect 25776 37564 26084 37584
rect 25776 37562 25782 37564
rect 25838 37562 25862 37564
rect 25918 37562 25942 37564
rect 25998 37562 26022 37564
rect 26078 37562 26084 37564
rect 25838 37510 25840 37562
rect 26020 37510 26022 37562
rect 25776 37508 25782 37510
rect 25838 37508 25862 37510
rect 25918 37508 25942 37510
rect 25998 37508 26022 37510
rect 26078 37508 26084 37510
rect 25776 37488 26084 37508
rect 30104 36780 30156 36786
rect 30104 36722 30156 36728
rect 25776 36476 26084 36496
rect 25776 36474 25782 36476
rect 25838 36474 25862 36476
rect 25918 36474 25942 36476
rect 25998 36474 26022 36476
rect 26078 36474 26084 36476
rect 25838 36422 25840 36474
rect 26020 36422 26022 36474
rect 25776 36420 25782 36422
rect 25838 36420 25862 36422
rect 25918 36420 25942 36422
rect 25998 36420 26022 36422
rect 26078 36420 26084 36422
rect 25776 36400 26084 36420
rect 30116 36281 30144 36722
rect 30102 36272 30158 36281
rect 30102 36207 30158 36216
rect 25776 35388 26084 35408
rect 25776 35386 25782 35388
rect 25838 35386 25862 35388
rect 25918 35386 25942 35388
rect 25998 35386 26022 35388
rect 26078 35386 26084 35388
rect 25838 35334 25840 35386
rect 26020 35334 26022 35386
rect 25776 35332 25782 35334
rect 25838 35332 25862 35334
rect 25918 35332 25942 35334
rect 25998 35332 26022 35334
rect 26078 35332 26084 35334
rect 25776 35312 26084 35332
rect 30102 34776 30158 34785
rect 30102 34711 30158 34720
rect 30116 34610 30144 34711
rect 30104 34604 30156 34610
rect 30104 34546 30156 34552
rect 29828 34536 29880 34542
rect 29828 34478 29880 34484
rect 25776 34300 26084 34320
rect 25776 34298 25782 34300
rect 25838 34298 25862 34300
rect 25918 34298 25942 34300
rect 25998 34298 26022 34300
rect 26078 34298 26084 34300
rect 25838 34246 25840 34298
rect 26020 34246 26022 34298
rect 25776 34244 25782 34246
rect 25838 34244 25862 34246
rect 25918 34244 25942 34246
rect 25998 34244 26022 34246
rect 26078 34244 26084 34246
rect 25776 34224 26084 34244
rect 22652 33856 22704 33862
rect 22652 33798 22704 33804
rect 22664 33522 22692 33798
rect 22652 33516 22704 33522
rect 22652 33458 22704 33464
rect 29840 33386 29868 34478
rect 30104 33516 30156 33522
rect 30104 33458 30156 33464
rect 29828 33380 29880 33386
rect 29828 33322 29880 33328
rect 22376 33312 22428 33318
rect 30012 33312 30064 33318
rect 22376 33254 22428 33260
rect 30010 33280 30012 33289
rect 30064 33280 30066 33289
rect 22388 29714 22416 33254
rect 25776 33212 26084 33232
rect 30010 33215 30066 33224
rect 25776 33210 25782 33212
rect 25838 33210 25862 33212
rect 25918 33210 25942 33212
rect 25998 33210 26022 33212
rect 26078 33210 26084 33212
rect 25838 33158 25840 33210
rect 26020 33158 26022 33210
rect 25776 33156 25782 33158
rect 25838 33156 25862 33158
rect 25918 33156 25942 33158
rect 25998 33156 26022 33158
rect 26078 33156 26084 33158
rect 25776 33136 26084 33156
rect 25776 32124 26084 32144
rect 25776 32122 25782 32124
rect 25838 32122 25862 32124
rect 25918 32122 25942 32124
rect 25998 32122 26022 32124
rect 26078 32122 26084 32124
rect 25838 32070 25840 32122
rect 26020 32070 26022 32122
rect 25776 32068 25782 32070
rect 25838 32068 25862 32070
rect 25918 32068 25942 32070
rect 25998 32068 26022 32070
rect 26078 32068 26084 32070
rect 25776 32048 26084 32068
rect 29828 31816 29880 31822
rect 29828 31758 29880 31764
rect 25776 31036 26084 31056
rect 25776 31034 25782 31036
rect 25838 31034 25862 31036
rect 25918 31034 25942 31036
rect 25998 31034 26022 31036
rect 26078 31034 26084 31036
rect 25838 30982 25840 31034
rect 26020 30982 26022 31034
rect 25776 30980 25782 30982
rect 25838 30980 25862 30982
rect 25918 30980 25942 30982
rect 25998 30980 26022 30982
rect 26078 30980 26084 30982
rect 25776 30960 26084 30980
rect 29840 30938 29868 31758
rect 30012 31680 30064 31686
rect 30010 31648 30012 31657
rect 30064 31648 30066 31657
rect 30010 31583 30066 31592
rect 29828 30932 29880 30938
rect 29828 30874 29880 30880
rect 30116 30734 30144 33458
rect 29552 30728 29604 30734
rect 29552 30670 29604 30676
rect 30104 30728 30156 30734
rect 30104 30670 30156 30676
rect 22928 30252 22980 30258
rect 22928 30194 22980 30200
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22376 29708 22428 29714
rect 22376 29650 22428 29656
rect 22664 29646 22692 29990
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22940 28762 22968 30194
rect 25776 29948 26084 29968
rect 25776 29946 25782 29948
rect 25838 29946 25862 29948
rect 25918 29946 25942 29948
rect 25998 29946 26022 29948
rect 26078 29946 26084 29948
rect 25838 29894 25840 29946
rect 26020 29894 26022 29946
rect 25776 29892 25782 29894
rect 25838 29892 25862 29894
rect 25918 29892 25942 29894
rect 25998 29892 26022 29894
rect 26078 29892 26084 29894
rect 25776 29872 26084 29892
rect 29368 29164 29420 29170
rect 29368 29106 29420 29112
rect 25776 28860 26084 28880
rect 25776 28858 25782 28860
rect 25838 28858 25862 28860
rect 25918 28858 25942 28860
rect 25998 28858 26022 28860
rect 26078 28858 26084 28860
rect 25838 28806 25840 28858
rect 26020 28806 26022 28858
rect 25776 28804 25782 28806
rect 25838 28804 25862 28806
rect 25918 28804 25942 28806
rect 25998 28804 26022 28806
rect 26078 28804 26084 28806
rect 25776 28784 26084 28804
rect 22928 28756 22980 28762
rect 22928 28698 22980 28704
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22376 24064 22428 24070
rect 22376 24006 22428 24012
rect 22388 23730 22416 24006
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22376 23588 22428 23594
rect 22376 23530 22428 23536
rect 22388 22574 22416 23530
rect 22480 23118 22508 23598
rect 22572 23322 22600 28494
rect 25776 27772 26084 27792
rect 25776 27770 25782 27772
rect 25838 27770 25862 27772
rect 25918 27770 25942 27772
rect 25998 27770 26022 27772
rect 26078 27770 26084 27772
rect 25838 27718 25840 27770
rect 26020 27718 26022 27770
rect 25776 27716 25782 27718
rect 25838 27716 25862 27718
rect 25918 27716 25942 27718
rect 25998 27716 26022 27718
rect 26078 27716 26084 27718
rect 25776 27696 26084 27716
rect 25776 26684 26084 26704
rect 25776 26682 25782 26684
rect 25838 26682 25862 26684
rect 25918 26682 25942 26684
rect 25998 26682 26022 26684
rect 26078 26682 26084 26684
rect 25838 26630 25840 26682
rect 26020 26630 26022 26682
rect 25776 26628 25782 26630
rect 25838 26628 25862 26630
rect 25918 26628 25942 26630
rect 25998 26628 26022 26630
rect 26078 26628 26084 26630
rect 25776 26608 26084 26628
rect 29184 25900 29236 25906
rect 29184 25842 29236 25848
rect 25776 25596 26084 25616
rect 25776 25594 25782 25596
rect 25838 25594 25862 25596
rect 25918 25594 25942 25596
rect 25998 25594 26022 25596
rect 26078 25594 26084 25596
rect 25838 25542 25840 25594
rect 26020 25542 26022 25594
rect 25776 25540 25782 25542
rect 25838 25540 25862 25542
rect 25918 25540 25942 25542
rect 25998 25540 26022 25542
rect 26078 25540 26084 25542
rect 25776 25520 26084 25540
rect 22744 24676 22796 24682
rect 22744 24618 22796 24624
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22468 23112 22520 23118
rect 22468 23054 22520 23060
rect 22480 22778 22508 23054
rect 22756 23050 22784 24618
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23768 24206 23796 24550
rect 25776 24508 26084 24528
rect 25776 24506 25782 24508
rect 25838 24506 25862 24508
rect 25918 24506 25942 24508
rect 25998 24506 26022 24508
rect 26078 24506 26084 24508
rect 25838 24454 25840 24506
rect 26020 24454 26022 24506
rect 25776 24452 25782 24454
rect 25838 24452 25862 24454
rect 25918 24452 25942 24454
rect 25998 24452 26022 24454
rect 26078 24452 26084 24454
rect 25776 24432 26084 24452
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 22940 23526 22968 24142
rect 23112 24064 23164 24070
rect 23112 24006 23164 24012
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22940 23118 22968 23462
rect 23124 23118 23152 24006
rect 25776 23420 26084 23440
rect 25776 23418 25782 23420
rect 25838 23418 25862 23420
rect 25918 23418 25942 23420
rect 25998 23418 26022 23420
rect 26078 23418 26084 23420
rect 25838 23366 25840 23418
rect 26020 23366 26022 23418
rect 25776 23364 25782 23366
rect 25838 23364 25862 23366
rect 25918 23364 25942 23366
rect 25998 23364 26022 23366
rect 26078 23364 26084 23366
rect 25776 23344 26084 23364
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 22744 23044 22796 23050
rect 22744 22986 22796 22992
rect 22468 22772 22520 22778
rect 22468 22714 22520 22720
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 22388 22098 22416 22510
rect 22376 22092 22428 22098
rect 22376 22034 22428 22040
rect 22480 22030 22508 22714
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22480 21622 22508 21966
rect 22468 21616 22520 21622
rect 22468 21558 22520 21564
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 22192 20528 22244 20534
rect 22192 20470 22244 20476
rect 21732 20256 21784 20262
rect 21784 20216 21864 20244
rect 21732 20198 21784 20204
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20811 14172 21119 14192
rect 20811 14170 20817 14172
rect 20873 14170 20897 14172
rect 20953 14170 20977 14172
rect 21033 14170 21057 14172
rect 21113 14170 21119 14172
rect 20873 14118 20875 14170
rect 21055 14118 21057 14170
rect 20811 14116 20817 14118
rect 20873 14116 20897 14118
rect 20953 14116 20977 14118
rect 21033 14116 21057 14118
rect 21113 14116 21119 14118
rect 20811 14096 21119 14116
rect 21560 13870 21588 15438
rect 21836 15366 21864 20216
rect 22204 18766 22232 20470
rect 22388 20398 22416 20878
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21928 18426 21956 18566
rect 21916 18420 21968 18426
rect 21916 18362 21968 18368
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22020 16454 22048 18226
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 22756 15434 22784 22986
rect 23124 22658 23152 23054
rect 23032 22642 23152 22658
rect 23020 22636 23152 22642
rect 23072 22630 23152 22636
rect 23020 22578 23072 22584
rect 23032 21962 23060 22578
rect 25776 22332 26084 22352
rect 25776 22330 25782 22332
rect 25838 22330 25862 22332
rect 25918 22330 25942 22332
rect 25998 22330 26022 22332
rect 26078 22330 26084 22332
rect 25838 22278 25840 22330
rect 26020 22278 26022 22330
rect 25776 22276 25782 22278
rect 25838 22276 25862 22278
rect 25918 22276 25942 22278
rect 25998 22276 26022 22278
rect 26078 22276 26084 22278
rect 25776 22256 26084 22276
rect 23020 21956 23072 21962
rect 23020 21898 23072 21904
rect 25776 21244 26084 21264
rect 25776 21242 25782 21244
rect 25838 21242 25862 21244
rect 25918 21242 25942 21244
rect 25998 21242 26022 21244
rect 26078 21242 26084 21244
rect 25838 21190 25840 21242
rect 26020 21190 26022 21242
rect 25776 21188 25782 21190
rect 25838 21188 25862 21190
rect 25918 21188 25942 21190
rect 25998 21188 26022 21190
rect 26078 21188 26084 21190
rect 25776 21168 26084 21188
rect 25776 20156 26084 20176
rect 25776 20154 25782 20156
rect 25838 20154 25862 20156
rect 25918 20154 25942 20156
rect 25998 20154 26022 20156
rect 26078 20154 26084 20156
rect 25838 20102 25840 20154
rect 26020 20102 26022 20154
rect 25776 20100 25782 20102
rect 25838 20100 25862 20102
rect 25918 20100 25942 20102
rect 25998 20100 26022 20102
rect 26078 20100 26084 20102
rect 25776 20080 26084 20100
rect 25776 19068 26084 19088
rect 25776 19066 25782 19068
rect 25838 19066 25862 19068
rect 25918 19066 25942 19068
rect 25998 19066 26022 19068
rect 26078 19066 26084 19068
rect 25838 19014 25840 19066
rect 26020 19014 26022 19066
rect 25776 19012 25782 19014
rect 25838 19012 25862 19014
rect 25918 19012 25942 19014
rect 25998 19012 26022 19014
rect 26078 19012 26084 19014
rect 25776 18992 26084 19012
rect 25776 17980 26084 18000
rect 25776 17978 25782 17980
rect 25838 17978 25862 17980
rect 25918 17978 25942 17980
rect 25998 17978 26022 17980
rect 26078 17978 26084 17980
rect 25838 17926 25840 17978
rect 26020 17926 26022 17978
rect 25776 17924 25782 17926
rect 25838 17924 25862 17926
rect 25918 17924 25942 17926
rect 25998 17924 26022 17926
rect 26078 17924 26084 17926
rect 25776 17904 26084 17924
rect 25776 16892 26084 16912
rect 25776 16890 25782 16892
rect 25838 16890 25862 16892
rect 25918 16890 25942 16892
rect 25998 16890 26022 16892
rect 26078 16890 26084 16892
rect 25838 16838 25840 16890
rect 26020 16838 26022 16890
rect 25776 16836 25782 16838
rect 25838 16836 25862 16838
rect 25918 16836 25942 16838
rect 25998 16836 26022 16838
rect 26078 16836 26084 16838
rect 25776 16816 26084 16836
rect 25776 15804 26084 15824
rect 25776 15802 25782 15804
rect 25838 15802 25862 15804
rect 25918 15802 25942 15804
rect 25998 15802 26022 15804
rect 26078 15802 26084 15804
rect 25838 15750 25840 15802
rect 26020 15750 26022 15802
rect 25776 15748 25782 15750
rect 25838 15748 25862 15750
rect 25918 15748 25942 15750
rect 25998 15748 26022 15750
rect 26078 15748 26084 15750
rect 25776 15728 26084 15748
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 21824 15360 21876 15366
rect 21824 15302 21876 15308
rect 21548 13864 21600 13870
rect 21548 13806 21600 13812
rect 21836 13734 21864 15302
rect 22756 15094 22784 15370
rect 29196 15162 29224 25842
rect 29184 15156 29236 15162
rect 29184 15098 29236 15104
rect 22744 15088 22796 15094
rect 22744 15030 22796 15036
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 29184 15020 29236 15026
rect 29184 14962 29236 14968
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 20811 13084 21119 13104
rect 20811 13082 20817 13084
rect 20873 13082 20897 13084
rect 20953 13082 20977 13084
rect 21033 13082 21057 13084
rect 21113 13082 21119 13084
rect 20873 13030 20875 13082
rect 21055 13030 21057 13082
rect 20811 13028 20817 13030
rect 20873 13028 20897 13030
rect 20953 13028 20977 13030
rect 21033 13028 21057 13030
rect 21113 13028 21119 13030
rect 20811 13008 21119 13028
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 20811 11996 21119 12016
rect 20811 11994 20817 11996
rect 20873 11994 20897 11996
rect 20953 11994 20977 11996
rect 21033 11994 21057 11996
rect 21113 11994 21119 11996
rect 20873 11942 20875 11994
rect 21055 11942 21057 11994
rect 20811 11940 20817 11942
rect 20873 11940 20897 11942
rect 20953 11940 20977 11942
rect 21033 11940 21057 11942
rect 21113 11940 21119 11942
rect 20811 11920 21119 11940
rect 21192 11898 21220 12242
rect 21928 12238 21956 14962
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22296 13938 22324 14758
rect 25776 14716 26084 14736
rect 25776 14714 25782 14716
rect 25838 14714 25862 14716
rect 25918 14714 25942 14716
rect 25998 14714 26022 14716
rect 26078 14714 26084 14716
rect 25838 14662 25840 14714
rect 26020 14662 26022 14714
rect 25776 14660 25782 14662
rect 25838 14660 25862 14662
rect 25918 14660 25942 14662
rect 25998 14660 26022 14662
rect 26078 14660 26084 14662
rect 25776 14640 26084 14660
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 22388 14006 22416 14350
rect 29196 14346 29224 14962
rect 29184 14340 29236 14346
rect 29184 14282 29236 14288
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 28080 14272 28132 14278
rect 28080 14214 28132 14220
rect 22480 14074 22508 14214
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 28092 13938 28120 14214
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 25776 13628 26084 13648
rect 25776 13626 25782 13628
rect 25838 13626 25862 13628
rect 25918 13626 25942 13628
rect 25998 13626 26022 13628
rect 26078 13626 26084 13628
rect 25838 13574 25840 13626
rect 26020 13574 26022 13626
rect 25776 13572 25782 13574
rect 25838 13572 25862 13574
rect 25918 13572 25942 13574
rect 25998 13572 26022 13574
rect 26078 13572 26084 13574
rect 25776 13552 26084 13572
rect 29000 12912 29052 12918
rect 29000 12854 29052 12860
rect 25776 12540 26084 12560
rect 25776 12538 25782 12540
rect 25838 12538 25862 12540
rect 25918 12538 25942 12540
rect 25998 12538 26022 12540
rect 26078 12538 26084 12540
rect 25838 12486 25840 12538
rect 26020 12486 26022 12538
rect 25776 12484 25782 12486
rect 25838 12484 25862 12486
rect 25918 12484 25942 12486
rect 25998 12484 26022 12486
rect 26078 12484 26084 12486
rect 25776 12464 26084 12484
rect 29012 12238 29040 12854
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 29000 12232 29052 12238
rect 29000 12174 29052 12180
rect 29184 12164 29236 12170
rect 29184 12106 29236 12112
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 29196 11762 29224 12106
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 29184 11756 29236 11762
rect 29184 11698 29236 11704
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20732 10810 20760 11018
rect 20811 10908 21119 10928
rect 20811 10906 20817 10908
rect 20873 10906 20897 10908
rect 20953 10906 20977 10908
rect 21033 10906 21057 10908
rect 21113 10906 21119 10908
rect 20873 10854 20875 10906
rect 21055 10854 21057 10906
rect 20811 10852 20817 10854
rect 20873 10852 20897 10854
rect 20953 10852 20977 10854
rect 21033 10852 21057 10854
rect 21113 10852 21119 10854
rect 20811 10832 21119 10852
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19812 6866 19840 7822
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 20088 7002 20116 7754
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19812 6390 19840 6802
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 20640 6322 20668 7278
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 19708 5908 19760 5914
rect 19708 5850 19760 5856
rect 19708 5636 19760 5642
rect 19708 5578 19760 5584
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 19628 4690 19656 5170
rect 19616 4684 19668 4690
rect 19616 4626 19668 4632
rect 19720 4078 19748 5578
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19812 4282 19840 4762
rect 20168 4548 20220 4554
rect 20168 4490 20220 4496
rect 19800 4276 19852 4282
rect 19800 4218 19852 4224
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 19524 4004 19576 4010
rect 19524 3946 19576 3952
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 19260 2310 19288 3130
rect 19536 2854 19564 3946
rect 19720 3602 19748 4014
rect 20180 3738 20208 4490
rect 20456 4486 20484 6190
rect 20444 4480 20496 4486
rect 20444 4422 20496 4428
rect 20456 4298 20484 4422
rect 20364 4282 20484 4298
rect 20364 4276 20496 4282
rect 20364 4270 20444 4276
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20364 3602 20392 4270
rect 20444 4218 20496 4224
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20456 3670 20484 4082
rect 20548 3942 20576 6258
rect 20732 5794 20760 9998
rect 20811 9820 21119 9840
rect 20811 9818 20817 9820
rect 20873 9818 20897 9820
rect 20953 9818 20977 9820
rect 21033 9818 21057 9820
rect 21113 9818 21119 9820
rect 20873 9766 20875 9818
rect 21055 9766 21057 9818
rect 20811 9764 20817 9766
rect 20873 9764 20897 9766
rect 20953 9764 20977 9766
rect 21033 9764 21057 9766
rect 21113 9764 21119 9766
rect 20811 9744 21119 9764
rect 20811 8732 21119 8752
rect 20811 8730 20817 8732
rect 20873 8730 20897 8732
rect 20953 8730 20977 8732
rect 21033 8730 21057 8732
rect 21113 8730 21119 8732
rect 20873 8678 20875 8730
rect 21055 8678 21057 8730
rect 20811 8676 20817 8678
rect 20873 8676 20897 8678
rect 20953 8676 20977 8678
rect 21033 8676 21057 8678
rect 21113 8676 21119 8678
rect 20811 8656 21119 8676
rect 21192 8090 21220 10610
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21284 8566 21312 9862
rect 21272 8560 21324 8566
rect 21272 8502 21324 8508
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 20811 7644 21119 7664
rect 20811 7642 20817 7644
rect 20873 7642 20897 7644
rect 20953 7642 20977 7644
rect 21033 7642 21057 7644
rect 21113 7642 21119 7644
rect 20873 7590 20875 7642
rect 21055 7590 21057 7642
rect 20811 7588 20817 7590
rect 20873 7588 20897 7590
rect 20953 7588 20977 7590
rect 21033 7588 21057 7590
rect 21113 7588 21119 7590
rect 20811 7568 21119 7588
rect 21192 6882 21220 8026
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 21100 6854 21220 6882
rect 21100 6798 21128 6854
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 20811 6556 21119 6576
rect 20811 6554 20817 6556
rect 20873 6554 20897 6556
rect 20953 6554 20977 6556
rect 21033 6554 21057 6556
rect 21113 6554 21119 6556
rect 20873 6502 20875 6554
rect 21055 6502 21057 6554
rect 20811 6500 20817 6502
rect 20873 6500 20897 6502
rect 20953 6500 20977 6502
rect 21033 6500 21057 6502
rect 21113 6500 21119 6502
rect 20811 6480 21119 6500
rect 21192 6458 21220 6666
rect 21284 6662 21312 7142
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21284 6254 21312 6598
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 20640 5766 20760 5794
rect 20640 5370 20668 5766
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20640 4214 20668 5306
rect 20732 4486 20760 5646
rect 20811 5468 21119 5488
rect 20811 5466 20817 5468
rect 20873 5466 20897 5468
rect 20953 5466 20977 5468
rect 21033 5466 21057 5468
rect 21113 5466 21119 5468
rect 20873 5414 20875 5466
rect 21055 5414 21057 5466
rect 20811 5412 20817 5414
rect 20873 5412 20897 5414
rect 20953 5412 20977 5414
rect 21033 5412 21057 5414
rect 21113 5412 21119 5414
rect 20811 5392 21119 5412
rect 21180 5296 21232 5302
rect 21180 5238 21232 5244
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20628 4208 20680 4214
rect 20628 4150 20680 4156
rect 20732 4162 20760 4422
rect 20811 4380 21119 4400
rect 20811 4378 20817 4380
rect 20873 4378 20897 4380
rect 20953 4378 20977 4380
rect 21033 4378 21057 4380
rect 21113 4378 21119 4380
rect 20873 4326 20875 4378
rect 21055 4326 21057 4378
rect 20811 4324 20817 4326
rect 20873 4324 20897 4326
rect 20953 4324 20977 4326
rect 21033 4324 21057 4326
rect 21113 4324 21119 4326
rect 20811 4304 21119 4324
rect 21192 4282 21220 5238
rect 21376 4826 21404 11698
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21640 9036 21692 9042
rect 21640 8978 21692 8984
rect 21548 8968 21600 8974
rect 21468 8916 21548 8922
rect 21468 8910 21600 8916
rect 21468 8894 21588 8910
rect 21468 8430 21496 8894
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 21560 8498 21588 8774
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21468 8090 21496 8366
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21560 7886 21588 8434
rect 21652 8430 21680 8978
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21652 7342 21680 8366
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21744 6662 21772 11086
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 21836 9518 21864 9998
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21836 7342 21864 9454
rect 21928 9178 21956 9522
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 22020 9110 22048 9318
rect 22008 9104 22060 9110
rect 22008 9046 22060 9052
rect 22008 8900 22060 8906
rect 22008 8842 22060 8848
rect 21916 8424 21968 8430
rect 21916 8366 21968 8372
rect 21928 8022 21956 8366
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21744 6322 21772 6598
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 21836 5234 21864 7278
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 21180 4276 21232 4282
rect 21180 4218 21232 4224
rect 20732 4134 20852 4162
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20444 3664 20496 3670
rect 20444 3606 20496 3612
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19904 3040 19932 3470
rect 20166 3088 20222 3097
rect 20456 3058 20484 3606
rect 20548 3126 20576 3878
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20536 3120 20588 3126
rect 20536 3062 20588 3068
rect 19904 3032 20166 3040
rect 19904 3012 20168 3032
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 20088 2378 20116 3012
rect 20220 3023 20222 3032
rect 20444 3052 20496 3058
rect 20168 2994 20220 3000
rect 20444 2994 20496 3000
rect 20168 2916 20220 2922
rect 20168 2858 20220 2864
rect 20076 2372 20128 2378
rect 20076 2314 20128 2320
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19260 2038 19288 2246
rect 19248 2032 19300 2038
rect 19248 1974 19300 1980
rect 19444 800 19472 2246
rect 20180 800 20208 2858
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20272 2650 20300 2790
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 20456 2514 20484 2994
rect 20548 2774 20576 3062
rect 20548 2746 20668 2774
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 20536 2440 20588 2446
rect 20640 2428 20668 2746
rect 20732 2650 20760 3674
rect 20824 3534 20852 4134
rect 20996 3664 21048 3670
rect 20996 3606 21048 3612
rect 21824 3664 21876 3670
rect 21824 3606 21876 3612
rect 21008 3534 21036 3606
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 21180 3528 21232 3534
rect 21180 3470 21232 3476
rect 20811 3292 21119 3312
rect 20811 3290 20817 3292
rect 20873 3290 20897 3292
rect 20953 3290 20977 3292
rect 21033 3290 21057 3292
rect 21113 3290 21119 3292
rect 20873 3238 20875 3290
rect 21055 3238 21057 3290
rect 20811 3236 20817 3238
rect 20873 3236 20897 3238
rect 20953 3236 20977 3238
rect 21033 3236 21057 3238
rect 21113 3236 21119 3238
rect 20811 3216 21119 3236
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20588 2400 20668 2428
rect 20536 2382 20588 2388
rect 20811 2204 21119 2224
rect 20811 2202 20817 2204
rect 20873 2202 20897 2204
rect 20953 2202 20977 2204
rect 21033 2202 21057 2204
rect 21113 2202 21119 2204
rect 20873 2150 20875 2202
rect 21055 2150 21057 2202
rect 20811 2148 20817 2150
rect 20873 2148 20897 2150
rect 20953 2148 20977 2150
rect 21033 2148 21057 2150
rect 21113 2148 21119 2150
rect 20811 2128 21119 2148
rect 20916 870 21036 898
rect 20916 800 20944 870
rect 11164 734 11376 762
rect 11794 0 11850 800
rect 12530 0 12586 800
rect 13266 0 13322 800
rect 14094 0 14150 800
rect 14830 0 14886 800
rect 15566 0 15622 800
rect 16394 0 16450 800
rect 17130 0 17186 800
rect 17866 0 17922 800
rect 18602 0 18658 800
rect 19430 0 19486 800
rect 20166 0 20222 800
rect 20902 0 20958 800
rect 21008 762 21036 870
rect 21192 762 21220 3470
rect 21836 3466 21864 3606
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21376 3194 21404 3402
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 21640 3120 21692 3126
rect 21640 3062 21692 3068
rect 21732 3120 21784 3126
rect 21732 3062 21784 3068
rect 21652 2650 21680 3062
rect 21640 2644 21692 2650
rect 21640 2586 21692 2592
rect 21744 800 21772 3062
rect 21836 2446 21864 3130
rect 22020 3058 22048 8842
rect 22112 7886 22140 11494
rect 25776 11452 26084 11472
rect 25776 11450 25782 11452
rect 25838 11450 25862 11452
rect 25918 11450 25942 11452
rect 25998 11450 26022 11452
rect 26078 11450 26084 11452
rect 25838 11398 25840 11450
rect 26020 11398 26022 11450
rect 25776 11396 25782 11398
rect 25838 11396 25862 11398
rect 25918 11396 25942 11398
rect 25998 11396 26022 11398
rect 26078 11396 26084 11398
rect 25776 11376 26084 11396
rect 25776 10364 26084 10384
rect 25776 10362 25782 10364
rect 25838 10362 25862 10364
rect 25918 10362 25942 10364
rect 25998 10362 26022 10364
rect 26078 10362 26084 10364
rect 25838 10310 25840 10362
rect 26020 10310 26022 10362
rect 25776 10308 25782 10310
rect 25838 10308 25862 10310
rect 25918 10308 25942 10310
rect 25998 10308 26022 10310
rect 26078 10308 26084 10310
rect 25776 10288 26084 10308
rect 28632 10260 28684 10266
rect 28632 10202 28684 10208
rect 22560 9988 22612 9994
rect 22560 9930 22612 9936
rect 22572 8634 22600 9930
rect 25776 9276 26084 9296
rect 25776 9274 25782 9276
rect 25838 9274 25862 9276
rect 25918 9274 25942 9276
rect 25998 9274 26022 9276
rect 26078 9274 26084 9276
rect 25838 9222 25840 9274
rect 26020 9222 26022 9274
rect 25776 9220 25782 9222
rect 25838 9220 25862 9222
rect 25918 9220 25942 9222
rect 25998 9220 26022 9222
rect 26078 9220 26084 9222
rect 25776 9200 26084 9220
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22100 7880 22152 7886
rect 22296 7834 22324 8434
rect 25776 8188 26084 8208
rect 25776 8186 25782 8188
rect 25838 8186 25862 8188
rect 25918 8186 25942 8188
rect 25998 8186 26022 8188
rect 26078 8186 26084 8188
rect 25838 8134 25840 8186
rect 26020 8134 26022 8186
rect 25776 8132 25782 8134
rect 25838 8132 25862 8134
rect 25918 8132 25942 8134
rect 25998 8132 26022 8134
rect 26078 8132 26084 8134
rect 25776 8112 26084 8132
rect 22152 7828 22232 7834
rect 22100 7822 22232 7828
rect 22112 7806 22232 7822
rect 22296 7806 22416 7834
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22112 3058 22140 7686
rect 22204 7546 22232 7806
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22296 7478 22324 7686
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 22100 3052 22152 3058
rect 22152 3012 22324 3040
rect 22100 2994 22152 3000
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 22020 2106 22048 2994
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 22112 2650 22140 2858
rect 22296 2650 22324 3012
rect 22388 2854 22416 7806
rect 25776 7100 26084 7120
rect 25776 7098 25782 7100
rect 25838 7098 25862 7100
rect 25918 7098 25942 7100
rect 25998 7098 26022 7100
rect 26078 7098 26084 7100
rect 25838 7046 25840 7098
rect 26020 7046 26022 7098
rect 25776 7044 25782 7046
rect 25838 7044 25862 7046
rect 25918 7044 25942 7046
rect 25998 7044 26022 7046
rect 26078 7044 26084 7046
rect 25776 7024 26084 7044
rect 25776 6012 26084 6032
rect 25776 6010 25782 6012
rect 25838 6010 25862 6012
rect 25918 6010 25942 6012
rect 25998 6010 26022 6012
rect 26078 6010 26084 6012
rect 25838 5958 25840 6010
rect 26020 5958 26022 6010
rect 25776 5956 25782 5958
rect 25838 5956 25862 5958
rect 25918 5956 25942 5958
rect 25998 5956 26022 5958
rect 26078 5956 26084 5958
rect 25776 5936 26084 5956
rect 25776 4924 26084 4944
rect 25776 4922 25782 4924
rect 25838 4922 25862 4924
rect 25918 4922 25942 4924
rect 25998 4922 26022 4924
rect 26078 4922 26084 4924
rect 25838 4870 25840 4922
rect 26020 4870 26022 4922
rect 25776 4868 25782 4870
rect 25838 4868 25862 4870
rect 25918 4868 25942 4870
rect 25998 4868 26022 4870
rect 26078 4868 26084 4870
rect 25776 4848 26084 4868
rect 23572 4004 23624 4010
rect 23572 3946 23624 3952
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 22940 3738 22968 3878
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 22468 3392 22520 3398
rect 22468 3334 22520 3340
rect 22480 3058 22508 3334
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 22376 2848 22428 2854
rect 22376 2790 22428 2796
rect 22572 2774 22600 3470
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 22756 2922 22784 3402
rect 23584 3194 23612 3946
rect 25776 3836 26084 3856
rect 25776 3834 25782 3836
rect 25838 3834 25862 3836
rect 25918 3834 25942 3836
rect 25998 3834 26022 3836
rect 26078 3834 26084 3836
rect 25838 3782 25840 3834
rect 26020 3782 26022 3834
rect 25776 3780 25782 3782
rect 25838 3780 25862 3782
rect 25918 3780 25942 3782
rect 25998 3780 26022 3782
rect 26078 3780 26084 3782
rect 25776 3760 26084 3780
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 25688 3392 25740 3398
rect 25688 3334 25740 3340
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 22928 3188 22980 3194
rect 22928 3130 22980 3136
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 22940 3097 22968 3130
rect 22926 3088 22982 3097
rect 22926 3023 22982 3032
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 22480 2746 22600 2774
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 22008 2100 22060 2106
rect 22008 2042 22060 2048
rect 22480 800 22508 2746
rect 22652 2508 22704 2514
rect 22652 2450 22704 2456
rect 22664 2310 22692 2450
rect 22756 2446 22784 2858
rect 23204 2508 23256 2514
rect 23204 2450 23256 2456
rect 22744 2440 22796 2446
rect 22744 2382 22796 2388
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 23216 800 23244 2450
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 23308 2038 23336 2246
rect 23296 2032 23348 2038
rect 23296 1974 23348 1980
rect 23952 800 23980 2994
rect 25700 2650 25728 3334
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 25776 2748 26084 2768
rect 25776 2746 25782 2748
rect 25838 2746 25862 2748
rect 25918 2746 25942 2748
rect 25998 2746 26022 2748
rect 26078 2746 26084 2748
rect 25838 2694 25840 2746
rect 26020 2694 26022 2746
rect 25776 2692 25782 2694
rect 25838 2692 25862 2694
rect 25918 2692 25942 2694
rect 25998 2692 26022 2694
rect 26078 2692 26084 2694
rect 25776 2672 26084 2692
rect 27448 2650 27476 2994
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 27632 2650 27660 2926
rect 27724 2854 27752 3334
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 25688 2644 25740 2650
rect 25688 2586 25740 2592
rect 27436 2644 27488 2650
rect 27436 2586 27488 2592
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 24780 800 24808 2382
rect 25044 2304 25096 2310
rect 25044 2246 25096 2252
rect 25056 2106 25084 2246
rect 25044 2100 25096 2106
rect 25044 2042 25096 2048
rect 25516 800 25544 2382
rect 26252 800 26280 2382
rect 27080 800 27108 2382
rect 27816 800 27844 3470
rect 27988 3392 28040 3398
rect 27988 3334 28040 3340
rect 28000 3126 28028 3334
rect 27988 3120 28040 3126
rect 27988 3062 28040 3068
rect 28552 800 28580 3470
rect 28644 2774 28672 10202
rect 28724 3936 28776 3942
rect 28724 3878 28776 3884
rect 28736 3058 28764 3878
rect 29276 3528 29328 3534
rect 29276 3470 29328 3476
rect 28724 3052 28776 3058
rect 28724 2994 28776 3000
rect 28644 2746 28764 2774
rect 28736 2446 28764 2746
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 28908 2304 28960 2310
rect 28908 2246 28960 2252
rect 21008 734 21220 762
rect 21730 0 21786 800
rect 22466 0 22522 800
rect 23202 0 23258 800
rect 23938 0 23994 800
rect 24766 0 24822 800
rect 25502 0 25558 800
rect 26238 0 26294 800
rect 27066 0 27122 800
rect 27802 0 27858 800
rect 28538 0 28594 800
rect 28920 785 28948 2246
rect 29288 800 29316 3470
rect 29380 2774 29408 29106
rect 29460 28212 29512 28218
rect 29460 28154 29512 28160
rect 29472 5914 29500 28154
rect 29564 13326 29592 30670
rect 30116 30326 30144 30670
rect 30104 30320 30156 30326
rect 30104 30262 30156 30268
rect 30010 30152 30066 30161
rect 30010 30087 30012 30096
rect 30064 30087 30066 30096
rect 30012 30058 30064 30064
rect 29736 29504 29788 29510
rect 29736 29446 29788 29452
rect 29644 28076 29696 28082
rect 29644 28018 29696 28024
rect 29656 14890 29684 28018
rect 29644 14884 29696 14890
rect 29644 14826 29696 14832
rect 29644 13864 29696 13870
rect 29644 13806 29696 13812
rect 29552 13320 29604 13326
rect 29552 13262 29604 13268
rect 29656 8498 29684 13806
rect 29644 8492 29696 8498
rect 29644 8434 29696 8440
rect 29656 6798 29684 8434
rect 29644 6792 29696 6798
rect 29644 6734 29696 6740
rect 29460 5908 29512 5914
rect 29460 5850 29512 5856
rect 29748 5710 29776 29446
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 30010 28520 30066 28529
rect 29840 28218 29868 28494
rect 30010 28455 30066 28464
rect 30024 28422 30052 28455
rect 30012 28416 30064 28422
rect 30012 28358 30064 28364
rect 29828 28212 29880 28218
rect 29828 28154 29880 28160
rect 30116 28082 30144 30262
rect 30104 28076 30156 28082
rect 30104 28018 30156 28024
rect 29920 27464 29972 27470
rect 29920 27406 29972 27412
rect 29932 27130 29960 27406
rect 30012 27328 30064 27334
rect 30012 27270 30064 27276
rect 29920 27124 29972 27130
rect 29920 27066 29972 27072
rect 30024 27033 30052 27270
rect 30010 27024 30066 27033
rect 30116 26994 30144 28018
rect 30010 26959 30066 26968
rect 30104 26988 30156 26994
rect 30104 26930 30156 26936
rect 30012 25696 30064 25702
rect 30012 25638 30064 25644
rect 30024 25537 30052 25638
rect 30010 25528 30066 25537
rect 30010 25463 30066 25472
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 29932 23866 29960 24142
rect 30012 24064 30064 24070
rect 30012 24006 30064 24012
rect 30024 23905 30052 24006
rect 30010 23896 30066 23905
rect 29920 23860 29972 23866
rect 30010 23831 30066 23840
rect 29920 23802 29972 23808
rect 30116 23730 30144 26930
rect 30104 23724 30156 23730
rect 30104 23666 30156 23672
rect 30116 22574 30144 23666
rect 30196 22636 30248 22642
rect 30196 22578 30248 22584
rect 30104 22568 30156 22574
rect 30104 22510 30156 22516
rect 30012 22432 30064 22438
rect 30010 22400 30012 22409
rect 30064 22400 30066 22409
rect 30010 22335 30066 22344
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 30010 20904 30066 20913
rect 29840 20602 29868 20878
rect 30010 20839 30066 20848
rect 30024 20806 30052 20839
rect 30012 20800 30064 20806
rect 30012 20742 30064 20748
rect 29828 20596 29880 20602
rect 29828 20538 29880 20544
rect 30116 20466 30144 22510
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 30012 19508 30064 19514
rect 30012 19450 30064 19456
rect 29920 19372 29972 19378
rect 29920 19314 29972 19320
rect 29828 18284 29880 18290
rect 29828 18226 29880 18232
rect 29840 17882 29868 18226
rect 29828 17876 29880 17882
rect 29828 17818 29880 17824
rect 29932 17762 29960 19314
rect 30024 19281 30052 19450
rect 30010 19272 30066 19281
rect 30010 19207 30066 19216
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 30024 17785 30052 18022
rect 29840 17734 29960 17762
rect 30010 17776 30066 17785
rect 29840 15586 29868 17734
rect 30010 17711 30066 17720
rect 30116 17678 30144 20402
rect 30104 17672 30156 17678
rect 30104 17614 30156 17620
rect 29920 16584 29972 16590
rect 29920 16526 29972 16532
rect 29932 15706 29960 16526
rect 30012 16448 30064 16454
rect 30012 16390 30064 16396
rect 30024 16153 30052 16390
rect 30010 16144 30066 16153
rect 30010 16079 30066 16088
rect 30116 15706 30144 17614
rect 29920 15700 29972 15706
rect 29920 15642 29972 15648
rect 30104 15700 30156 15706
rect 30104 15642 30156 15648
rect 29840 15558 30144 15586
rect 29920 15496 29972 15502
rect 29920 15438 29972 15444
rect 29828 15020 29880 15026
rect 29828 14962 29880 14968
rect 29840 14618 29868 14962
rect 29828 14612 29880 14618
rect 29828 14554 29880 14560
rect 29932 14550 29960 15438
rect 30012 14816 30064 14822
rect 30012 14758 30064 14764
rect 30024 14657 30052 14758
rect 30010 14648 30066 14657
rect 30010 14583 30066 14592
rect 30116 14550 30144 15558
rect 29920 14544 29972 14550
rect 29920 14486 29972 14492
rect 30104 14544 30156 14550
rect 30104 14486 30156 14492
rect 29920 14408 29972 14414
rect 29920 14350 29972 14356
rect 29828 13320 29880 13326
rect 29828 13262 29880 13268
rect 29840 12986 29868 13262
rect 29932 13258 29960 14350
rect 30208 14074 30236 22578
rect 30288 15496 30340 15502
rect 30288 15438 30340 15444
rect 30300 14958 30328 15438
rect 30288 14952 30340 14958
rect 30288 14894 30340 14900
rect 30300 14414 30328 14894
rect 30288 14408 30340 14414
rect 30288 14350 30340 14356
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 30300 13938 30328 14350
rect 30288 13932 30340 13938
rect 30288 13874 30340 13880
rect 29920 13252 29972 13258
rect 29920 13194 29972 13200
rect 30012 13184 30064 13190
rect 30010 13152 30012 13161
rect 30064 13152 30066 13161
rect 30010 13087 30066 13096
rect 29828 12980 29880 12986
rect 29828 12922 29880 12928
rect 30300 12850 30328 13874
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 30300 12238 30328 12786
rect 30288 12232 30340 12238
rect 30288 12174 30340 12180
rect 29828 12096 29880 12102
rect 29828 12038 29880 12044
rect 29840 10062 29868 12038
rect 30012 11552 30064 11558
rect 30010 11520 30012 11529
rect 30064 11520 30066 11529
rect 30010 11455 30066 11464
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 30010 10024 30066 10033
rect 30010 9959 30066 9968
rect 30024 9926 30052 9959
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 30010 8392 30066 8401
rect 30010 8327 30012 8336
rect 30064 8327 30066 8336
rect 30012 8298 30064 8304
rect 29828 7404 29880 7410
rect 29828 7346 29880 7352
rect 29840 7002 29868 7346
rect 30012 7200 30064 7206
rect 30012 7142 30064 7148
rect 29828 6996 29880 7002
rect 29828 6938 29880 6944
rect 30024 6905 30052 7142
rect 30010 6896 30066 6905
rect 30010 6831 30066 6840
rect 30104 6792 30156 6798
rect 30104 6734 30156 6740
rect 30116 6118 30144 6734
rect 30104 6112 30156 6118
rect 30104 6054 30156 6060
rect 29828 5908 29880 5914
rect 29828 5850 29880 5856
rect 29736 5704 29788 5710
rect 29736 5646 29788 5652
rect 29748 4146 29776 5646
rect 29840 5234 29868 5850
rect 30010 5400 30066 5409
rect 30010 5335 30012 5344
rect 30064 5335 30066 5344
rect 30012 5306 30064 5312
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 30104 4616 30156 4622
rect 30104 4558 30156 4564
rect 29920 4480 29972 4486
rect 29920 4422 29972 4428
rect 29736 4140 29788 4146
rect 29736 4082 29788 4088
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29564 2854 29592 3878
rect 29932 3618 29960 4422
rect 30012 3936 30064 3942
rect 30012 3878 30064 3884
rect 30024 3777 30052 3878
rect 30010 3768 30066 3777
rect 30010 3703 30066 3712
rect 29932 3590 30052 3618
rect 29920 3392 29972 3398
rect 29920 3334 29972 3340
rect 29932 3058 29960 3334
rect 30024 3058 30052 3590
rect 29920 3052 29972 3058
rect 29920 2994 29972 3000
rect 30012 3052 30064 3058
rect 30012 2994 30064 3000
rect 29552 2848 29604 2854
rect 29552 2790 29604 2796
rect 29380 2746 29500 2774
rect 29472 2446 29500 2746
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 30012 2304 30064 2310
rect 30010 2272 30012 2281
rect 30064 2272 30066 2281
rect 30010 2207 30066 2216
rect 30116 800 30144 4558
rect 30840 4072 30892 4078
rect 30840 4014 30892 4020
rect 30852 800 30880 4014
rect 31576 4004 31628 4010
rect 31576 3946 31628 3952
rect 31588 800 31616 3946
rect 28906 776 28962 785
rect 28906 711 28962 720
rect 29274 0 29330 800
rect 30102 0 30158 800
rect 30838 0 30894 800
rect 31574 0 31630 800
<< via2 >>
rect 2778 47504 2834 47560
rect 2226 45348 2282 45384
rect 2226 45328 2228 45348
rect 2228 45328 2280 45348
rect 2280 45328 2282 45348
rect 30194 47096 30250 47152
rect 2870 46824 2926 46880
rect 2962 46008 3018 46064
rect 10886 45722 10942 45724
rect 10966 45722 11022 45724
rect 11046 45722 11102 45724
rect 11126 45722 11182 45724
rect 10886 45670 10932 45722
rect 10932 45670 10942 45722
rect 10966 45670 10996 45722
rect 10996 45670 11008 45722
rect 11008 45670 11022 45722
rect 11046 45670 11060 45722
rect 11060 45670 11072 45722
rect 11072 45670 11102 45722
rect 11126 45670 11136 45722
rect 11136 45670 11182 45722
rect 10886 45668 10942 45670
rect 10966 45668 11022 45670
rect 11046 45668 11102 45670
rect 11126 45668 11182 45670
rect 20817 45722 20873 45724
rect 20897 45722 20953 45724
rect 20977 45722 21033 45724
rect 21057 45722 21113 45724
rect 20817 45670 20863 45722
rect 20863 45670 20873 45722
rect 20897 45670 20927 45722
rect 20927 45670 20939 45722
rect 20939 45670 20953 45722
rect 20977 45670 20991 45722
rect 20991 45670 21003 45722
rect 21003 45670 21033 45722
rect 21057 45670 21067 45722
rect 21067 45670 21113 45722
rect 20817 45668 20873 45670
rect 20897 45668 20953 45670
rect 20977 45668 21033 45670
rect 21057 45668 21113 45670
rect 30102 45600 30158 45656
rect 1490 44512 1546 44568
rect 1490 43832 1546 43888
rect 1490 43052 1492 43072
rect 1492 43052 1544 43072
rect 1544 43052 1546 43072
rect 1490 43016 1546 43052
rect 1490 42336 1546 42392
rect 1490 41656 1546 41712
rect 1490 40876 1492 40896
rect 1492 40876 1544 40896
rect 1544 40876 1546 40896
rect 1490 40840 1546 40876
rect 1490 40160 1546 40216
rect 1490 37848 1546 37904
rect 1398 35672 1454 35728
rect 1490 34992 1546 35048
rect 2226 39344 2282 39400
rect 5921 45178 5977 45180
rect 6001 45178 6057 45180
rect 6081 45178 6137 45180
rect 6161 45178 6217 45180
rect 5921 45126 5967 45178
rect 5967 45126 5977 45178
rect 6001 45126 6031 45178
rect 6031 45126 6043 45178
rect 6043 45126 6057 45178
rect 6081 45126 6095 45178
rect 6095 45126 6107 45178
rect 6107 45126 6137 45178
rect 6161 45126 6171 45178
rect 6171 45126 6217 45178
rect 5921 45124 5977 45126
rect 6001 45124 6057 45126
rect 6081 45124 6137 45126
rect 6161 45124 6217 45126
rect 15852 45178 15908 45180
rect 15932 45178 15988 45180
rect 16012 45178 16068 45180
rect 16092 45178 16148 45180
rect 15852 45126 15898 45178
rect 15898 45126 15908 45178
rect 15932 45126 15962 45178
rect 15962 45126 15974 45178
rect 15974 45126 15988 45178
rect 16012 45126 16026 45178
rect 16026 45126 16038 45178
rect 16038 45126 16068 45178
rect 16092 45126 16102 45178
rect 16102 45126 16148 45178
rect 15852 45124 15908 45126
rect 15932 45124 15988 45126
rect 16012 45124 16068 45126
rect 16092 45124 16148 45126
rect 25782 45178 25838 45180
rect 25862 45178 25918 45180
rect 25942 45178 25998 45180
rect 26022 45178 26078 45180
rect 25782 45126 25828 45178
rect 25828 45126 25838 45178
rect 25862 45126 25892 45178
rect 25892 45126 25904 45178
rect 25904 45126 25918 45178
rect 25942 45126 25956 45178
rect 25956 45126 25968 45178
rect 25968 45126 25998 45178
rect 26022 45126 26032 45178
rect 26032 45126 26078 45178
rect 25782 45124 25838 45126
rect 25862 45124 25918 45126
rect 25942 45124 25998 45126
rect 26022 45124 26078 45126
rect 3054 38700 3056 38720
rect 3056 38700 3108 38720
rect 3108 38700 3110 38720
rect 3054 38664 3110 38700
rect 2318 36524 2320 36544
rect 2320 36524 2372 36544
rect 2372 36524 2374 36544
rect 2318 36488 2374 36524
rect 1490 32680 1546 32736
rect 1490 31320 1546 31376
rect 1490 29844 1546 29880
rect 1490 29824 1492 29844
rect 1492 29824 1544 29844
rect 1544 29824 1546 29844
rect 1490 29028 1546 29064
rect 1490 29008 1492 29028
rect 1492 29008 1544 29028
rect 1544 29008 1546 29028
rect 1490 28364 1492 28384
rect 1492 28364 1544 28384
rect 1544 28364 1546 28384
rect 1490 28328 1546 28364
rect 2226 32000 2282 32056
rect 1490 27512 1546 27568
rect 1490 26852 1546 26888
rect 1490 26832 1492 26852
rect 1492 26832 1544 26852
rect 1544 26832 1546 26852
rect 1490 26188 1492 26208
rect 1492 26188 1544 26208
rect 1544 26188 1546 26208
rect 1490 26152 1546 26188
rect 1490 25336 1546 25392
rect 1490 24676 1546 24712
rect 1490 24656 1492 24676
rect 1492 24656 1544 24676
rect 1544 24656 1546 24676
rect 1490 23840 1546 23896
rect 1398 23160 1454 23216
rect 1398 20984 1454 21040
rect 1214 15000 1270 15056
rect 1214 12824 1270 12880
rect 1214 5480 1270 5536
rect 2042 21664 2098 21720
rect 1398 15816 1454 15872
rect 1398 14456 1454 14512
rect 1398 11328 1454 11384
rect 1398 10648 1454 10704
rect 3054 37168 3110 37224
rect 2962 34176 3018 34232
rect 2962 33496 3018 33552
rect 3146 30540 3148 30560
rect 3148 30540 3200 30560
rect 3200 30540 3202 30560
rect 3146 30504 3202 30540
rect 5921 44090 5977 44092
rect 6001 44090 6057 44092
rect 6081 44090 6137 44092
rect 6161 44090 6217 44092
rect 5921 44038 5967 44090
rect 5967 44038 5977 44090
rect 6001 44038 6031 44090
rect 6031 44038 6043 44090
rect 6043 44038 6057 44090
rect 6081 44038 6095 44090
rect 6095 44038 6107 44090
rect 6107 44038 6137 44090
rect 6161 44038 6171 44090
rect 6171 44038 6217 44090
rect 5921 44036 5977 44038
rect 6001 44036 6057 44038
rect 6081 44036 6137 44038
rect 6161 44036 6217 44038
rect 5921 43002 5977 43004
rect 6001 43002 6057 43004
rect 6081 43002 6137 43004
rect 6161 43002 6217 43004
rect 5921 42950 5967 43002
rect 5967 42950 5977 43002
rect 6001 42950 6031 43002
rect 6031 42950 6043 43002
rect 6043 42950 6057 43002
rect 6081 42950 6095 43002
rect 6095 42950 6107 43002
rect 6107 42950 6137 43002
rect 6161 42950 6171 43002
rect 6171 42950 6217 43002
rect 5921 42948 5977 42950
rect 6001 42948 6057 42950
rect 6081 42948 6137 42950
rect 6161 42948 6217 42950
rect 5921 41914 5977 41916
rect 6001 41914 6057 41916
rect 6081 41914 6137 41916
rect 6161 41914 6217 41916
rect 5921 41862 5967 41914
rect 5967 41862 5977 41914
rect 6001 41862 6031 41914
rect 6031 41862 6043 41914
rect 6043 41862 6057 41914
rect 6081 41862 6095 41914
rect 6095 41862 6107 41914
rect 6107 41862 6137 41914
rect 6161 41862 6171 41914
rect 6171 41862 6217 41914
rect 5921 41860 5977 41862
rect 6001 41860 6057 41862
rect 6081 41860 6137 41862
rect 6161 41860 6217 41862
rect 5921 40826 5977 40828
rect 6001 40826 6057 40828
rect 6081 40826 6137 40828
rect 6161 40826 6217 40828
rect 5921 40774 5967 40826
rect 5967 40774 5977 40826
rect 6001 40774 6031 40826
rect 6031 40774 6043 40826
rect 6043 40774 6057 40826
rect 6081 40774 6095 40826
rect 6095 40774 6107 40826
rect 6107 40774 6137 40826
rect 6161 40774 6171 40826
rect 6171 40774 6217 40826
rect 5921 40772 5977 40774
rect 6001 40772 6057 40774
rect 6081 40772 6137 40774
rect 6161 40772 6217 40774
rect 5921 39738 5977 39740
rect 6001 39738 6057 39740
rect 6081 39738 6137 39740
rect 6161 39738 6217 39740
rect 5921 39686 5967 39738
rect 5967 39686 5977 39738
rect 6001 39686 6031 39738
rect 6031 39686 6043 39738
rect 6043 39686 6057 39738
rect 6081 39686 6095 39738
rect 6095 39686 6107 39738
rect 6107 39686 6137 39738
rect 6161 39686 6171 39738
rect 6171 39686 6217 39738
rect 5921 39684 5977 39686
rect 6001 39684 6057 39686
rect 6081 39684 6137 39686
rect 6161 39684 6217 39686
rect 5921 38650 5977 38652
rect 6001 38650 6057 38652
rect 6081 38650 6137 38652
rect 6161 38650 6217 38652
rect 5921 38598 5967 38650
rect 5967 38598 5977 38650
rect 6001 38598 6031 38650
rect 6031 38598 6043 38650
rect 6043 38598 6057 38650
rect 6081 38598 6095 38650
rect 6095 38598 6107 38650
rect 6107 38598 6137 38650
rect 6161 38598 6171 38650
rect 6171 38598 6217 38650
rect 5921 38596 5977 38598
rect 6001 38596 6057 38598
rect 6081 38596 6137 38598
rect 6161 38596 6217 38598
rect 5921 37562 5977 37564
rect 6001 37562 6057 37564
rect 6081 37562 6137 37564
rect 6161 37562 6217 37564
rect 5921 37510 5967 37562
rect 5967 37510 5977 37562
rect 6001 37510 6031 37562
rect 6031 37510 6043 37562
rect 6043 37510 6057 37562
rect 6081 37510 6095 37562
rect 6095 37510 6107 37562
rect 6107 37510 6137 37562
rect 6161 37510 6171 37562
rect 6171 37510 6217 37562
rect 5921 37508 5977 37510
rect 6001 37508 6057 37510
rect 6081 37508 6137 37510
rect 6161 37508 6217 37510
rect 5921 36474 5977 36476
rect 6001 36474 6057 36476
rect 6081 36474 6137 36476
rect 6161 36474 6217 36476
rect 5921 36422 5967 36474
rect 5967 36422 5977 36474
rect 6001 36422 6031 36474
rect 6031 36422 6043 36474
rect 6043 36422 6057 36474
rect 6081 36422 6095 36474
rect 6095 36422 6107 36474
rect 6107 36422 6137 36474
rect 6161 36422 6171 36474
rect 6171 36422 6217 36474
rect 5921 36420 5977 36422
rect 6001 36420 6057 36422
rect 6081 36420 6137 36422
rect 6161 36420 6217 36422
rect 5921 35386 5977 35388
rect 6001 35386 6057 35388
rect 6081 35386 6137 35388
rect 6161 35386 6217 35388
rect 5921 35334 5967 35386
rect 5967 35334 5977 35386
rect 6001 35334 6031 35386
rect 6031 35334 6043 35386
rect 6043 35334 6057 35386
rect 6081 35334 6095 35386
rect 6095 35334 6107 35386
rect 6107 35334 6137 35386
rect 6161 35334 6171 35386
rect 6171 35334 6217 35386
rect 5921 35332 5977 35334
rect 6001 35332 6057 35334
rect 6081 35332 6137 35334
rect 6161 35332 6217 35334
rect 5921 34298 5977 34300
rect 6001 34298 6057 34300
rect 6081 34298 6137 34300
rect 6161 34298 6217 34300
rect 5921 34246 5967 34298
rect 5967 34246 5977 34298
rect 6001 34246 6031 34298
rect 6031 34246 6043 34298
rect 6043 34246 6057 34298
rect 6081 34246 6095 34298
rect 6095 34246 6107 34298
rect 6107 34246 6137 34298
rect 6161 34246 6171 34298
rect 6171 34246 6217 34298
rect 5921 34244 5977 34246
rect 6001 34244 6057 34246
rect 6081 34244 6137 34246
rect 6161 34244 6217 34246
rect 5921 33210 5977 33212
rect 6001 33210 6057 33212
rect 6081 33210 6137 33212
rect 6161 33210 6217 33212
rect 5921 33158 5967 33210
rect 5967 33158 5977 33210
rect 6001 33158 6031 33210
rect 6031 33158 6043 33210
rect 6043 33158 6057 33210
rect 6081 33158 6095 33210
rect 6095 33158 6107 33210
rect 6107 33158 6137 33210
rect 6161 33158 6171 33210
rect 6171 33158 6217 33210
rect 5921 33156 5977 33158
rect 6001 33156 6057 33158
rect 6081 33156 6137 33158
rect 6161 33156 6217 33158
rect 5921 32122 5977 32124
rect 6001 32122 6057 32124
rect 6081 32122 6137 32124
rect 6161 32122 6217 32124
rect 5921 32070 5967 32122
rect 5967 32070 5977 32122
rect 6001 32070 6031 32122
rect 6031 32070 6043 32122
rect 6043 32070 6057 32122
rect 6081 32070 6095 32122
rect 6095 32070 6107 32122
rect 6107 32070 6137 32122
rect 6161 32070 6171 32122
rect 6171 32070 6217 32122
rect 5921 32068 5977 32070
rect 6001 32068 6057 32070
rect 6081 32068 6137 32070
rect 6161 32068 6217 32070
rect 5921 31034 5977 31036
rect 6001 31034 6057 31036
rect 6081 31034 6137 31036
rect 6161 31034 6217 31036
rect 5921 30982 5967 31034
rect 5967 30982 5977 31034
rect 6001 30982 6031 31034
rect 6031 30982 6043 31034
rect 6043 30982 6057 31034
rect 6081 30982 6095 31034
rect 6095 30982 6107 31034
rect 6107 30982 6137 31034
rect 6161 30982 6171 31034
rect 6171 30982 6217 31034
rect 5921 30980 5977 30982
rect 6001 30980 6057 30982
rect 6081 30980 6137 30982
rect 6161 30980 6217 30982
rect 5921 29946 5977 29948
rect 6001 29946 6057 29948
rect 6081 29946 6137 29948
rect 6161 29946 6217 29948
rect 5921 29894 5967 29946
rect 5967 29894 5977 29946
rect 6001 29894 6031 29946
rect 6031 29894 6043 29946
rect 6043 29894 6057 29946
rect 6081 29894 6095 29946
rect 6095 29894 6107 29946
rect 6107 29894 6137 29946
rect 6161 29894 6171 29946
rect 6171 29894 6217 29946
rect 5921 29892 5977 29894
rect 6001 29892 6057 29894
rect 6081 29892 6137 29894
rect 6161 29892 6217 29894
rect 5921 28858 5977 28860
rect 6001 28858 6057 28860
rect 6081 28858 6137 28860
rect 6161 28858 6217 28860
rect 5921 28806 5967 28858
rect 5967 28806 5977 28858
rect 6001 28806 6031 28858
rect 6031 28806 6043 28858
rect 6043 28806 6057 28858
rect 6081 28806 6095 28858
rect 6095 28806 6107 28858
rect 6107 28806 6137 28858
rect 6161 28806 6171 28858
rect 6171 28806 6217 28858
rect 5921 28804 5977 28806
rect 6001 28804 6057 28806
rect 6081 28804 6137 28806
rect 6161 28804 6217 28806
rect 2778 22344 2834 22400
rect 2962 18672 3018 18728
rect 3146 19896 3202 19952
rect 3238 19488 3294 19544
rect 3054 17992 3110 18048
rect 2778 17176 2834 17232
rect 3238 16496 3294 16552
rect 1398 9152 1454 9208
rect 1398 8336 1454 8392
rect 1398 7656 1454 7712
rect 2778 13504 2834 13560
rect 2778 12008 2834 12064
rect 2778 9832 2834 9888
rect 5921 27770 5977 27772
rect 6001 27770 6057 27772
rect 6081 27770 6137 27772
rect 6161 27770 6217 27772
rect 5921 27718 5967 27770
rect 5967 27718 5977 27770
rect 6001 27718 6031 27770
rect 6031 27718 6043 27770
rect 6043 27718 6057 27770
rect 6081 27718 6095 27770
rect 6095 27718 6107 27770
rect 6107 27718 6137 27770
rect 6161 27718 6171 27770
rect 6171 27718 6217 27770
rect 5921 27716 5977 27718
rect 6001 27716 6057 27718
rect 6081 27716 6137 27718
rect 6161 27716 6217 27718
rect 6366 27648 6422 27704
rect 3790 26460 3792 26480
rect 3792 26460 3844 26480
rect 3844 26460 3846 26480
rect 3790 26424 3846 26460
rect 4066 20168 4122 20224
rect 5078 26016 5134 26072
rect 4894 25916 4896 25936
rect 4896 25916 4948 25936
rect 4948 25916 4950 25936
rect 4894 25880 4950 25916
rect 5722 26424 5778 26480
rect 4802 25744 4858 25800
rect 5921 26682 5977 26684
rect 6001 26682 6057 26684
rect 6081 26682 6137 26684
rect 6161 26682 6217 26684
rect 5921 26630 5967 26682
rect 5967 26630 5977 26682
rect 6001 26630 6031 26682
rect 6031 26630 6043 26682
rect 6043 26630 6057 26682
rect 6081 26630 6095 26682
rect 6095 26630 6107 26682
rect 6107 26630 6137 26682
rect 6161 26630 6171 26682
rect 6171 26630 6217 26682
rect 5921 26628 5977 26630
rect 6001 26628 6057 26630
rect 6081 26628 6137 26630
rect 6161 26628 6217 26630
rect 5906 26444 5962 26480
rect 5906 26424 5908 26444
rect 5908 26424 5960 26444
rect 5960 26424 5962 26444
rect 6090 26016 6146 26072
rect 5921 25594 5977 25596
rect 6001 25594 6057 25596
rect 6081 25594 6137 25596
rect 6161 25594 6217 25596
rect 5921 25542 5967 25594
rect 5967 25542 5977 25594
rect 6001 25542 6031 25594
rect 6031 25542 6043 25594
rect 6043 25542 6057 25594
rect 6081 25542 6095 25594
rect 6095 25542 6107 25594
rect 6107 25542 6137 25594
rect 6161 25542 6171 25594
rect 6171 25542 6217 25594
rect 5921 25540 5977 25542
rect 6001 25540 6057 25542
rect 6081 25540 6137 25542
rect 6161 25540 6217 25542
rect 5814 24792 5870 24848
rect 5078 24248 5134 24304
rect 2778 6160 2834 6216
rect 1398 4664 1454 4720
rect 3974 6840 4030 6896
rect 5921 24506 5977 24508
rect 6001 24506 6057 24508
rect 6081 24506 6137 24508
rect 6161 24506 6217 24508
rect 5921 24454 5967 24506
rect 5967 24454 5977 24506
rect 6001 24454 6031 24506
rect 6031 24454 6043 24506
rect 6043 24454 6057 24506
rect 6081 24454 6095 24506
rect 6095 24454 6107 24506
rect 6107 24454 6137 24506
rect 6161 24454 6171 24506
rect 6171 24454 6217 24506
rect 5921 24452 5977 24454
rect 6001 24452 6057 24454
rect 6081 24452 6137 24454
rect 6161 24452 6217 24454
rect 6182 24268 6238 24304
rect 6182 24248 6184 24268
rect 6184 24248 6236 24268
rect 6236 24248 6238 24268
rect 5921 23418 5977 23420
rect 6001 23418 6057 23420
rect 6081 23418 6137 23420
rect 6161 23418 6217 23420
rect 5921 23366 5967 23418
rect 5967 23366 5977 23418
rect 6001 23366 6031 23418
rect 6031 23366 6043 23418
rect 6043 23366 6057 23418
rect 6081 23366 6095 23418
rect 6095 23366 6107 23418
rect 6107 23366 6137 23418
rect 6161 23366 6171 23418
rect 6171 23366 6217 23418
rect 5921 23364 5977 23366
rect 6001 23364 6057 23366
rect 6081 23364 6137 23366
rect 6161 23364 6217 23366
rect 5921 22330 5977 22332
rect 6001 22330 6057 22332
rect 6081 22330 6137 22332
rect 6161 22330 6217 22332
rect 5921 22278 5967 22330
rect 5967 22278 5977 22330
rect 6001 22278 6031 22330
rect 6031 22278 6043 22330
rect 6043 22278 6057 22330
rect 6081 22278 6095 22330
rect 6095 22278 6107 22330
rect 6107 22278 6137 22330
rect 6161 22278 6171 22330
rect 6171 22278 6217 22330
rect 5921 22276 5977 22278
rect 6001 22276 6057 22278
rect 6081 22276 6137 22278
rect 6161 22276 6217 22278
rect 5921 21242 5977 21244
rect 6001 21242 6057 21244
rect 6081 21242 6137 21244
rect 6161 21242 6217 21244
rect 5921 21190 5967 21242
rect 5967 21190 5977 21242
rect 6001 21190 6031 21242
rect 6031 21190 6043 21242
rect 6043 21190 6057 21242
rect 6081 21190 6095 21242
rect 6095 21190 6107 21242
rect 6107 21190 6137 21242
rect 6161 21190 6171 21242
rect 6171 21190 6217 21242
rect 5921 21188 5977 21190
rect 6001 21188 6057 21190
rect 6081 21188 6137 21190
rect 6161 21188 6217 21190
rect 10886 44634 10942 44636
rect 10966 44634 11022 44636
rect 11046 44634 11102 44636
rect 11126 44634 11182 44636
rect 10886 44582 10932 44634
rect 10932 44582 10942 44634
rect 10966 44582 10996 44634
rect 10996 44582 11008 44634
rect 11008 44582 11022 44634
rect 11046 44582 11060 44634
rect 11060 44582 11072 44634
rect 11072 44582 11102 44634
rect 11126 44582 11136 44634
rect 11136 44582 11182 44634
rect 10886 44580 10942 44582
rect 10966 44580 11022 44582
rect 11046 44580 11102 44582
rect 11126 44580 11182 44582
rect 20817 44634 20873 44636
rect 20897 44634 20953 44636
rect 20977 44634 21033 44636
rect 21057 44634 21113 44636
rect 20817 44582 20863 44634
rect 20863 44582 20873 44634
rect 20897 44582 20927 44634
rect 20927 44582 20939 44634
rect 20939 44582 20953 44634
rect 20977 44582 20991 44634
rect 20991 44582 21003 44634
rect 21003 44582 21033 44634
rect 21057 44582 21067 44634
rect 21067 44582 21113 44634
rect 20817 44580 20873 44582
rect 20897 44580 20953 44582
rect 20977 44580 21033 44582
rect 21057 44580 21113 44582
rect 6734 27648 6790 27704
rect 6734 25900 6790 25936
rect 6734 25880 6736 25900
rect 6736 25880 6788 25900
rect 6788 25880 6790 25900
rect 7470 27104 7526 27160
rect 5921 20154 5977 20156
rect 6001 20154 6057 20156
rect 6081 20154 6137 20156
rect 6161 20154 6217 20156
rect 5921 20102 5967 20154
rect 5967 20102 5977 20154
rect 6001 20102 6031 20154
rect 6031 20102 6043 20154
rect 6043 20102 6057 20154
rect 6081 20102 6095 20154
rect 6095 20102 6107 20154
rect 6107 20102 6137 20154
rect 6161 20102 6171 20154
rect 6171 20102 6217 20154
rect 5921 20100 5977 20102
rect 6001 20100 6057 20102
rect 6081 20100 6137 20102
rect 6161 20100 6217 20102
rect 5814 19760 5870 19816
rect 5921 19066 5977 19068
rect 6001 19066 6057 19068
rect 6081 19066 6137 19068
rect 6161 19066 6217 19068
rect 5921 19014 5967 19066
rect 5967 19014 5977 19066
rect 6001 19014 6031 19066
rect 6031 19014 6043 19066
rect 6043 19014 6057 19066
rect 6081 19014 6095 19066
rect 6095 19014 6107 19066
rect 6107 19014 6137 19066
rect 6161 19014 6171 19066
rect 6171 19014 6217 19066
rect 5921 19012 5977 19014
rect 6001 19012 6057 19014
rect 6081 19012 6137 19014
rect 6161 19012 6217 19014
rect 1858 2488 1914 2544
rect 2778 3984 2834 4040
rect 2778 3168 2834 3224
rect 2778 1672 2834 1728
rect 2962 992 3018 1048
rect 5921 17978 5977 17980
rect 6001 17978 6057 17980
rect 6081 17978 6137 17980
rect 6161 17978 6217 17980
rect 5921 17926 5967 17978
rect 5967 17926 5977 17978
rect 6001 17926 6031 17978
rect 6031 17926 6043 17978
rect 6043 17926 6057 17978
rect 6081 17926 6095 17978
rect 6095 17926 6107 17978
rect 6107 17926 6137 17978
rect 6161 17926 6171 17978
rect 6171 17926 6217 17978
rect 5921 17924 5977 17926
rect 6001 17924 6057 17926
rect 6081 17924 6137 17926
rect 6161 17924 6217 17926
rect 5921 16890 5977 16892
rect 6001 16890 6057 16892
rect 6081 16890 6137 16892
rect 6161 16890 6217 16892
rect 5921 16838 5967 16890
rect 5967 16838 5977 16890
rect 6001 16838 6031 16890
rect 6031 16838 6043 16890
rect 6043 16838 6057 16890
rect 6081 16838 6095 16890
rect 6095 16838 6107 16890
rect 6107 16838 6137 16890
rect 6161 16838 6171 16890
rect 6171 16838 6217 16890
rect 5921 16836 5977 16838
rect 6001 16836 6057 16838
rect 6081 16836 6137 16838
rect 6161 16836 6217 16838
rect 6274 15952 6330 16008
rect 5921 15802 5977 15804
rect 6001 15802 6057 15804
rect 6081 15802 6137 15804
rect 6161 15802 6217 15804
rect 5921 15750 5967 15802
rect 5967 15750 5977 15802
rect 6001 15750 6031 15802
rect 6031 15750 6043 15802
rect 6043 15750 6057 15802
rect 6081 15750 6095 15802
rect 6095 15750 6107 15802
rect 6107 15750 6137 15802
rect 6161 15750 6171 15802
rect 6171 15750 6217 15802
rect 5921 15748 5977 15750
rect 6001 15748 6057 15750
rect 6081 15748 6137 15750
rect 6161 15748 6217 15750
rect 5921 14714 5977 14716
rect 6001 14714 6057 14716
rect 6081 14714 6137 14716
rect 6161 14714 6217 14716
rect 5921 14662 5967 14714
rect 5967 14662 5977 14714
rect 6001 14662 6031 14714
rect 6031 14662 6043 14714
rect 6043 14662 6057 14714
rect 6081 14662 6095 14714
rect 6095 14662 6107 14714
rect 6107 14662 6137 14714
rect 6161 14662 6171 14714
rect 6171 14662 6217 14714
rect 5921 14660 5977 14662
rect 6001 14660 6057 14662
rect 6081 14660 6137 14662
rect 6161 14660 6217 14662
rect 6182 14320 6238 14376
rect 5921 13626 5977 13628
rect 6001 13626 6057 13628
rect 6081 13626 6137 13628
rect 6161 13626 6217 13628
rect 5921 13574 5967 13626
rect 5967 13574 5977 13626
rect 6001 13574 6031 13626
rect 6031 13574 6043 13626
rect 6043 13574 6057 13626
rect 6081 13574 6095 13626
rect 6095 13574 6107 13626
rect 6107 13574 6137 13626
rect 6161 13574 6171 13626
rect 6171 13574 6217 13626
rect 5921 13572 5977 13574
rect 6001 13572 6057 13574
rect 6081 13572 6137 13574
rect 6161 13572 6217 13574
rect 5921 12538 5977 12540
rect 6001 12538 6057 12540
rect 6081 12538 6137 12540
rect 6161 12538 6217 12540
rect 5921 12486 5967 12538
rect 5967 12486 5977 12538
rect 6001 12486 6031 12538
rect 6031 12486 6043 12538
rect 6043 12486 6057 12538
rect 6081 12486 6095 12538
rect 6095 12486 6107 12538
rect 6107 12486 6137 12538
rect 6161 12486 6171 12538
rect 6171 12486 6217 12538
rect 5921 12484 5977 12486
rect 6001 12484 6057 12486
rect 6081 12484 6137 12486
rect 6161 12484 6217 12486
rect 6918 19796 6920 19816
rect 6920 19796 6972 19816
rect 6972 19796 6974 19816
rect 6918 19760 6974 19796
rect 6642 18264 6698 18320
rect 6642 17992 6698 18048
rect 9678 36080 9734 36136
rect 9034 30368 9090 30424
rect 9034 27548 9036 27568
rect 9036 27548 9088 27568
rect 9088 27548 9090 27568
rect 9034 27512 9090 27548
rect 7654 25880 7710 25936
rect 5921 11450 5977 11452
rect 6001 11450 6057 11452
rect 6081 11450 6137 11452
rect 6161 11450 6217 11452
rect 5921 11398 5967 11450
rect 5967 11398 5977 11450
rect 6001 11398 6031 11450
rect 6031 11398 6043 11450
rect 6043 11398 6057 11450
rect 6081 11398 6095 11450
rect 6095 11398 6107 11450
rect 6107 11398 6137 11450
rect 6161 11398 6171 11450
rect 6171 11398 6217 11450
rect 5921 11396 5977 11398
rect 6001 11396 6057 11398
rect 6081 11396 6137 11398
rect 6161 11396 6217 11398
rect 5921 10362 5977 10364
rect 6001 10362 6057 10364
rect 6081 10362 6137 10364
rect 6161 10362 6217 10364
rect 5921 10310 5967 10362
rect 5967 10310 5977 10362
rect 6001 10310 6031 10362
rect 6031 10310 6043 10362
rect 6043 10310 6057 10362
rect 6081 10310 6095 10362
rect 6095 10310 6107 10362
rect 6107 10310 6137 10362
rect 6161 10310 6171 10362
rect 6171 10310 6217 10362
rect 5921 10308 5977 10310
rect 6001 10308 6057 10310
rect 6081 10308 6137 10310
rect 6161 10308 6217 10310
rect 5262 9016 5318 9072
rect 5921 9274 5977 9276
rect 6001 9274 6057 9276
rect 6081 9274 6137 9276
rect 6161 9274 6217 9276
rect 5921 9222 5967 9274
rect 5967 9222 5977 9274
rect 6001 9222 6031 9274
rect 6031 9222 6043 9274
rect 6043 9222 6057 9274
rect 6081 9222 6095 9274
rect 6095 9222 6107 9274
rect 6107 9222 6137 9274
rect 6161 9222 6171 9274
rect 6171 9222 6217 9274
rect 5921 9220 5977 9222
rect 6001 9220 6057 9222
rect 6081 9220 6137 9222
rect 6161 9220 6217 9222
rect 5921 8186 5977 8188
rect 6001 8186 6057 8188
rect 6081 8186 6137 8188
rect 6161 8186 6217 8188
rect 5921 8134 5967 8186
rect 5967 8134 5977 8186
rect 6001 8134 6031 8186
rect 6031 8134 6043 8186
rect 6043 8134 6057 8186
rect 6081 8134 6095 8186
rect 6095 8134 6107 8186
rect 6107 8134 6137 8186
rect 6161 8134 6171 8186
rect 6171 8134 6217 8186
rect 5921 8132 5977 8134
rect 6001 8132 6057 8134
rect 6081 8132 6137 8134
rect 6161 8132 6217 8134
rect 5921 7098 5977 7100
rect 6001 7098 6057 7100
rect 6081 7098 6137 7100
rect 6161 7098 6217 7100
rect 5921 7046 5967 7098
rect 5967 7046 5977 7098
rect 6001 7046 6031 7098
rect 6031 7046 6043 7098
rect 6043 7046 6057 7098
rect 6081 7046 6095 7098
rect 6095 7046 6107 7098
rect 6107 7046 6137 7098
rect 6161 7046 6171 7098
rect 6171 7046 6217 7098
rect 5921 7044 5977 7046
rect 6001 7044 6057 7046
rect 6081 7044 6137 7046
rect 6161 7044 6217 7046
rect 5921 6010 5977 6012
rect 6001 6010 6057 6012
rect 6081 6010 6137 6012
rect 6161 6010 6217 6012
rect 5921 5958 5967 6010
rect 5967 5958 5977 6010
rect 6001 5958 6031 6010
rect 6031 5958 6043 6010
rect 6043 5958 6057 6010
rect 6081 5958 6095 6010
rect 6095 5958 6107 6010
rect 6107 5958 6137 6010
rect 6161 5958 6171 6010
rect 6171 5958 6217 6010
rect 5921 5956 5977 5958
rect 6001 5956 6057 5958
rect 6081 5956 6137 5958
rect 6161 5956 6217 5958
rect 7470 16088 7526 16144
rect 7930 25200 7986 25256
rect 8114 24812 8170 24848
rect 8114 24792 8116 24812
rect 8116 24792 8168 24812
rect 8168 24792 8170 24812
rect 8390 27412 8392 27432
rect 8392 27412 8444 27432
rect 8444 27412 8446 27432
rect 8390 27376 8446 27412
rect 8114 23568 8170 23624
rect 8574 25900 8630 25936
rect 8574 25880 8576 25900
rect 8576 25880 8628 25900
rect 8628 25880 8630 25900
rect 7562 14068 7618 14104
rect 7562 14048 7564 14068
rect 7564 14048 7616 14068
rect 7616 14048 7618 14068
rect 5921 4922 5977 4924
rect 6001 4922 6057 4924
rect 6081 4922 6137 4924
rect 6161 4922 6217 4924
rect 5921 4870 5967 4922
rect 5967 4870 5977 4922
rect 6001 4870 6031 4922
rect 6031 4870 6043 4922
rect 6043 4870 6057 4922
rect 6081 4870 6095 4922
rect 6095 4870 6107 4922
rect 6107 4870 6137 4922
rect 6161 4870 6171 4922
rect 6171 4870 6217 4922
rect 5921 4868 5977 4870
rect 6001 4868 6057 4870
rect 6081 4868 6137 4870
rect 6161 4868 6217 4870
rect 5921 3834 5977 3836
rect 6001 3834 6057 3836
rect 6081 3834 6137 3836
rect 6161 3834 6217 3836
rect 5921 3782 5967 3834
rect 5967 3782 5977 3834
rect 6001 3782 6031 3834
rect 6031 3782 6043 3834
rect 6043 3782 6057 3834
rect 6081 3782 6095 3834
rect 6095 3782 6107 3834
rect 6107 3782 6137 3834
rect 6161 3782 6171 3834
rect 6171 3782 6217 3834
rect 5921 3780 5977 3782
rect 6001 3780 6057 3782
rect 6081 3780 6137 3782
rect 6161 3780 6217 3782
rect 8022 19896 8078 19952
rect 8206 21936 8262 21992
rect 8022 13912 8078 13968
rect 5921 2746 5977 2748
rect 6001 2746 6057 2748
rect 6081 2746 6137 2748
rect 6161 2746 6217 2748
rect 5921 2694 5967 2746
rect 5967 2694 5977 2746
rect 6001 2694 6031 2746
rect 6031 2694 6043 2746
rect 6043 2694 6057 2746
rect 6081 2694 6095 2746
rect 6095 2694 6107 2746
rect 6107 2694 6137 2746
rect 6161 2694 6171 2746
rect 6171 2694 6217 2746
rect 5921 2692 5977 2694
rect 6001 2692 6057 2694
rect 6081 2692 6137 2694
rect 6161 2692 6217 2694
rect 10046 36236 10102 36272
rect 10046 36216 10048 36236
rect 10048 36216 10100 36236
rect 10100 36216 10102 36236
rect 15852 44090 15908 44092
rect 15932 44090 15988 44092
rect 16012 44090 16068 44092
rect 16092 44090 16148 44092
rect 15852 44038 15898 44090
rect 15898 44038 15908 44090
rect 15932 44038 15962 44090
rect 15962 44038 15974 44090
rect 15974 44038 15988 44090
rect 16012 44038 16026 44090
rect 16026 44038 16038 44090
rect 16038 44038 16068 44090
rect 16092 44038 16102 44090
rect 16102 44038 16148 44090
rect 15852 44036 15908 44038
rect 15932 44036 15988 44038
rect 16012 44036 16068 44038
rect 16092 44036 16148 44038
rect 10886 43546 10942 43548
rect 10966 43546 11022 43548
rect 11046 43546 11102 43548
rect 11126 43546 11182 43548
rect 10886 43494 10932 43546
rect 10932 43494 10942 43546
rect 10966 43494 10996 43546
rect 10996 43494 11008 43546
rect 11008 43494 11022 43546
rect 11046 43494 11060 43546
rect 11060 43494 11072 43546
rect 11072 43494 11102 43546
rect 11126 43494 11136 43546
rect 11136 43494 11182 43546
rect 10886 43492 10942 43494
rect 10966 43492 11022 43494
rect 11046 43492 11102 43494
rect 11126 43492 11182 43494
rect 25782 44090 25838 44092
rect 25862 44090 25918 44092
rect 25942 44090 25998 44092
rect 26022 44090 26078 44092
rect 25782 44038 25828 44090
rect 25828 44038 25838 44090
rect 25862 44038 25892 44090
rect 25892 44038 25904 44090
rect 25904 44038 25918 44090
rect 25942 44038 25956 44090
rect 25956 44038 25968 44090
rect 25968 44038 25998 44090
rect 26022 44038 26032 44090
rect 26032 44038 26078 44090
rect 25782 44036 25838 44038
rect 25862 44036 25918 44038
rect 25942 44036 25998 44038
rect 26022 44036 26078 44038
rect 20817 43546 20873 43548
rect 20897 43546 20953 43548
rect 20977 43546 21033 43548
rect 21057 43546 21113 43548
rect 20817 43494 20863 43546
rect 20863 43494 20873 43546
rect 20897 43494 20927 43546
rect 20927 43494 20939 43546
rect 20939 43494 20953 43546
rect 20977 43494 20991 43546
rect 20991 43494 21003 43546
rect 21003 43494 21033 43546
rect 21057 43494 21067 43546
rect 21067 43494 21113 43546
rect 20817 43492 20873 43494
rect 20897 43492 20953 43494
rect 20977 43492 21033 43494
rect 21057 43492 21113 43494
rect 15852 43002 15908 43004
rect 15932 43002 15988 43004
rect 16012 43002 16068 43004
rect 16092 43002 16148 43004
rect 15852 42950 15898 43002
rect 15898 42950 15908 43002
rect 15932 42950 15962 43002
rect 15962 42950 15974 43002
rect 15974 42950 15988 43002
rect 16012 42950 16026 43002
rect 16026 42950 16038 43002
rect 16038 42950 16068 43002
rect 16092 42950 16102 43002
rect 16102 42950 16148 43002
rect 15852 42948 15908 42950
rect 15932 42948 15988 42950
rect 16012 42948 16068 42950
rect 16092 42948 16148 42950
rect 10886 42458 10942 42460
rect 10966 42458 11022 42460
rect 11046 42458 11102 42460
rect 11126 42458 11182 42460
rect 10886 42406 10932 42458
rect 10932 42406 10942 42458
rect 10966 42406 10996 42458
rect 10996 42406 11008 42458
rect 11008 42406 11022 42458
rect 11046 42406 11060 42458
rect 11060 42406 11072 42458
rect 11072 42406 11102 42458
rect 11126 42406 11136 42458
rect 11136 42406 11182 42458
rect 10886 42404 10942 42406
rect 10966 42404 11022 42406
rect 11046 42404 11102 42406
rect 11126 42404 11182 42406
rect 15852 41914 15908 41916
rect 15932 41914 15988 41916
rect 16012 41914 16068 41916
rect 16092 41914 16148 41916
rect 15852 41862 15898 41914
rect 15898 41862 15908 41914
rect 15932 41862 15962 41914
rect 15962 41862 15974 41914
rect 15974 41862 15988 41914
rect 16012 41862 16026 41914
rect 16026 41862 16038 41914
rect 16038 41862 16068 41914
rect 16092 41862 16102 41914
rect 16102 41862 16148 41914
rect 15852 41860 15908 41862
rect 15932 41860 15988 41862
rect 16012 41860 16068 41862
rect 16092 41860 16148 41862
rect 10886 41370 10942 41372
rect 10966 41370 11022 41372
rect 11046 41370 11102 41372
rect 11126 41370 11182 41372
rect 10886 41318 10932 41370
rect 10932 41318 10942 41370
rect 10966 41318 10996 41370
rect 10996 41318 11008 41370
rect 11008 41318 11022 41370
rect 11046 41318 11060 41370
rect 11060 41318 11072 41370
rect 11072 41318 11102 41370
rect 11126 41318 11136 41370
rect 11136 41318 11182 41370
rect 10886 41316 10942 41318
rect 10966 41316 11022 41318
rect 11046 41316 11102 41318
rect 11126 41316 11182 41318
rect 10886 40282 10942 40284
rect 10966 40282 11022 40284
rect 11046 40282 11102 40284
rect 11126 40282 11182 40284
rect 10886 40230 10932 40282
rect 10932 40230 10942 40282
rect 10966 40230 10996 40282
rect 10996 40230 11008 40282
rect 11008 40230 11022 40282
rect 11046 40230 11060 40282
rect 11060 40230 11072 40282
rect 11072 40230 11102 40282
rect 11126 40230 11136 40282
rect 11136 40230 11182 40282
rect 10886 40228 10942 40230
rect 10966 40228 11022 40230
rect 11046 40228 11102 40230
rect 11126 40228 11182 40230
rect 10886 39194 10942 39196
rect 10966 39194 11022 39196
rect 11046 39194 11102 39196
rect 11126 39194 11182 39196
rect 10886 39142 10932 39194
rect 10932 39142 10942 39194
rect 10966 39142 10996 39194
rect 10996 39142 11008 39194
rect 11008 39142 11022 39194
rect 11046 39142 11060 39194
rect 11060 39142 11072 39194
rect 11072 39142 11102 39194
rect 11126 39142 11136 39194
rect 11136 39142 11182 39194
rect 10886 39140 10942 39142
rect 10966 39140 11022 39142
rect 11046 39140 11102 39142
rect 11126 39140 11182 39142
rect 10886 38106 10942 38108
rect 10966 38106 11022 38108
rect 11046 38106 11102 38108
rect 11126 38106 11182 38108
rect 10886 38054 10932 38106
rect 10932 38054 10942 38106
rect 10966 38054 10996 38106
rect 10996 38054 11008 38106
rect 11008 38054 11022 38106
rect 11046 38054 11060 38106
rect 11060 38054 11072 38106
rect 11072 38054 11102 38106
rect 11126 38054 11136 38106
rect 11136 38054 11182 38106
rect 10886 38052 10942 38054
rect 10966 38052 11022 38054
rect 11046 38052 11102 38054
rect 11126 38052 11182 38054
rect 10886 37018 10942 37020
rect 10966 37018 11022 37020
rect 11046 37018 11102 37020
rect 11126 37018 11182 37020
rect 10886 36966 10932 37018
rect 10932 36966 10942 37018
rect 10966 36966 10996 37018
rect 10996 36966 11008 37018
rect 11008 36966 11022 37018
rect 11046 36966 11060 37018
rect 11060 36966 11072 37018
rect 11072 36966 11102 37018
rect 11126 36966 11136 37018
rect 11136 36966 11182 37018
rect 10886 36964 10942 36966
rect 10966 36964 11022 36966
rect 11046 36964 11102 36966
rect 11126 36964 11182 36966
rect 11518 36252 11520 36272
rect 11520 36252 11572 36272
rect 11572 36252 11574 36272
rect 11518 36216 11574 36252
rect 11518 36080 11574 36136
rect 10886 35930 10942 35932
rect 10966 35930 11022 35932
rect 11046 35930 11102 35932
rect 11126 35930 11182 35932
rect 10886 35878 10932 35930
rect 10932 35878 10942 35930
rect 10966 35878 10996 35930
rect 10996 35878 11008 35930
rect 11008 35878 11022 35930
rect 11046 35878 11060 35930
rect 11060 35878 11072 35930
rect 11072 35878 11102 35930
rect 11126 35878 11136 35930
rect 11136 35878 11182 35930
rect 10886 35876 10942 35878
rect 10966 35876 11022 35878
rect 11046 35876 11102 35878
rect 11126 35876 11182 35878
rect 9310 27548 9312 27568
rect 9312 27548 9364 27568
rect 9364 27548 9366 27568
rect 9310 27512 9366 27548
rect 9494 27668 9550 27704
rect 9494 27648 9496 27668
rect 9496 27648 9548 27668
rect 9548 27648 9550 27668
rect 9586 27104 9642 27160
rect 9402 25744 9458 25800
rect 9310 25236 9312 25256
rect 9312 25236 9364 25256
rect 9364 25236 9366 25256
rect 9310 25200 9366 25236
rect 8942 23604 8944 23624
rect 8944 23604 8996 23624
rect 8996 23604 8998 23624
rect 8942 23568 8998 23604
rect 9586 26308 9642 26344
rect 9586 26288 9588 26308
rect 9588 26288 9640 26308
rect 9640 26288 9642 26308
rect 9770 24132 9826 24168
rect 9770 24112 9772 24132
rect 9772 24112 9824 24132
rect 9824 24112 9826 24132
rect 10886 34842 10942 34844
rect 10966 34842 11022 34844
rect 11046 34842 11102 34844
rect 11126 34842 11182 34844
rect 10886 34790 10932 34842
rect 10932 34790 10942 34842
rect 10966 34790 10996 34842
rect 10996 34790 11008 34842
rect 11008 34790 11022 34842
rect 11046 34790 11060 34842
rect 11060 34790 11072 34842
rect 11072 34790 11102 34842
rect 11126 34790 11136 34842
rect 11136 34790 11182 34842
rect 10886 34788 10942 34790
rect 10966 34788 11022 34790
rect 11046 34788 11102 34790
rect 11126 34788 11182 34790
rect 10886 33754 10942 33756
rect 10966 33754 11022 33756
rect 11046 33754 11102 33756
rect 11126 33754 11182 33756
rect 10886 33702 10932 33754
rect 10932 33702 10942 33754
rect 10966 33702 10996 33754
rect 10996 33702 11008 33754
rect 11008 33702 11022 33754
rect 11046 33702 11060 33754
rect 11060 33702 11072 33754
rect 11072 33702 11102 33754
rect 11126 33702 11136 33754
rect 11136 33702 11182 33754
rect 10886 33700 10942 33702
rect 10966 33700 11022 33702
rect 11046 33700 11102 33702
rect 11126 33700 11182 33702
rect 10322 27376 10378 27432
rect 10230 26988 10286 27024
rect 10230 26968 10232 26988
rect 10232 26968 10284 26988
rect 10284 26968 10286 26988
rect 9494 18264 9550 18320
rect 9310 17992 9366 18048
rect 9126 13948 9128 13968
rect 9128 13948 9180 13968
rect 9180 13948 9182 13968
rect 9126 13912 9182 13948
rect 9586 14068 9642 14104
rect 9586 14048 9588 14068
rect 9588 14048 9640 14068
rect 9640 14048 9642 14068
rect 10886 32666 10942 32668
rect 10966 32666 11022 32668
rect 11046 32666 11102 32668
rect 11126 32666 11182 32668
rect 10886 32614 10932 32666
rect 10932 32614 10942 32666
rect 10966 32614 10996 32666
rect 10996 32614 11008 32666
rect 11008 32614 11022 32666
rect 11046 32614 11060 32666
rect 11060 32614 11072 32666
rect 11072 32614 11102 32666
rect 11126 32614 11136 32666
rect 11136 32614 11182 32666
rect 10886 32612 10942 32614
rect 10966 32612 11022 32614
rect 11046 32612 11102 32614
rect 11126 32612 11182 32614
rect 10886 31578 10942 31580
rect 10966 31578 11022 31580
rect 11046 31578 11102 31580
rect 11126 31578 11182 31580
rect 10886 31526 10932 31578
rect 10932 31526 10942 31578
rect 10966 31526 10996 31578
rect 10996 31526 11008 31578
rect 11008 31526 11022 31578
rect 11046 31526 11060 31578
rect 11060 31526 11072 31578
rect 11072 31526 11102 31578
rect 11126 31526 11136 31578
rect 11136 31526 11182 31578
rect 10886 31524 10942 31526
rect 10966 31524 11022 31526
rect 11046 31524 11102 31526
rect 11126 31524 11182 31526
rect 10886 30490 10942 30492
rect 10966 30490 11022 30492
rect 11046 30490 11102 30492
rect 11126 30490 11182 30492
rect 10886 30438 10932 30490
rect 10932 30438 10942 30490
rect 10966 30438 10996 30490
rect 10996 30438 11008 30490
rect 11008 30438 11022 30490
rect 11046 30438 11060 30490
rect 11060 30438 11072 30490
rect 11072 30438 11102 30490
rect 11126 30438 11136 30490
rect 11136 30438 11182 30490
rect 10886 30436 10942 30438
rect 10966 30436 11022 30438
rect 11046 30436 11102 30438
rect 11126 30436 11182 30438
rect 10506 26832 10562 26888
rect 10886 29402 10942 29404
rect 10966 29402 11022 29404
rect 11046 29402 11102 29404
rect 11126 29402 11182 29404
rect 10886 29350 10932 29402
rect 10932 29350 10942 29402
rect 10966 29350 10996 29402
rect 10996 29350 11008 29402
rect 11008 29350 11022 29402
rect 11046 29350 11060 29402
rect 11060 29350 11072 29402
rect 11072 29350 11102 29402
rect 11126 29350 11136 29402
rect 11136 29350 11182 29402
rect 10886 29348 10942 29350
rect 10966 29348 11022 29350
rect 11046 29348 11102 29350
rect 11126 29348 11182 29350
rect 10886 28314 10942 28316
rect 10966 28314 11022 28316
rect 11046 28314 11102 28316
rect 11126 28314 11182 28316
rect 10886 28262 10932 28314
rect 10932 28262 10942 28314
rect 10966 28262 10996 28314
rect 10996 28262 11008 28314
rect 11008 28262 11022 28314
rect 11046 28262 11060 28314
rect 11060 28262 11072 28314
rect 11072 28262 11102 28314
rect 11126 28262 11136 28314
rect 11136 28262 11182 28314
rect 10886 28260 10942 28262
rect 10966 28260 11022 28262
rect 11046 28260 11102 28262
rect 11126 28260 11182 28262
rect 10782 27412 10784 27432
rect 10784 27412 10836 27432
rect 10836 27412 10838 27432
rect 10782 27376 10838 27412
rect 10886 27226 10942 27228
rect 10966 27226 11022 27228
rect 11046 27226 11102 27228
rect 11126 27226 11182 27228
rect 10886 27174 10932 27226
rect 10932 27174 10942 27226
rect 10966 27174 10996 27226
rect 10996 27174 11008 27226
rect 11008 27174 11022 27226
rect 11046 27174 11060 27226
rect 11060 27174 11072 27226
rect 11072 27174 11102 27226
rect 11126 27174 11136 27226
rect 11136 27174 11182 27226
rect 10886 27172 10942 27174
rect 10966 27172 11022 27174
rect 11046 27172 11102 27174
rect 11126 27172 11182 27174
rect 10886 26138 10942 26140
rect 10966 26138 11022 26140
rect 11046 26138 11102 26140
rect 11126 26138 11182 26140
rect 10886 26086 10932 26138
rect 10932 26086 10942 26138
rect 10966 26086 10996 26138
rect 10996 26086 11008 26138
rect 11008 26086 11022 26138
rect 11046 26086 11060 26138
rect 11060 26086 11072 26138
rect 11072 26086 11102 26138
rect 11126 26086 11136 26138
rect 11136 26086 11182 26138
rect 10886 26084 10942 26086
rect 10966 26084 11022 26086
rect 11046 26084 11102 26086
rect 11126 26084 11182 26086
rect 10886 25050 10942 25052
rect 10966 25050 11022 25052
rect 11046 25050 11102 25052
rect 11126 25050 11182 25052
rect 10886 24998 10932 25050
rect 10932 24998 10942 25050
rect 10966 24998 10996 25050
rect 10996 24998 11008 25050
rect 11008 24998 11022 25050
rect 11046 24998 11060 25050
rect 11060 24998 11072 25050
rect 11072 24998 11102 25050
rect 11126 24998 11136 25050
rect 11136 24998 11182 25050
rect 10886 24996 10942 24998
rect 10966 24996 11022 24998
rect 11046 24996 11102 24998
rect 11126 24996 11182 24998
rect 10690 24132 10746 24168
rect 10690 24112 10692 24132
rect 10692 24112 10744 24132
rect 10744 24112 10746 24132
rect 10886 23962 10942 23964
rect 10966 23962 11022 23964
rect 11046 23962 11102 23964
rect 11126 23962 11182 23964
rect 10886 23910 10932 23962
rect 10932 23910 10942 23962
rect 10966 23910 10996 23962
rect 10996 23910 11008 23962
rect 11008 23910 11022 23962
rect 11046 23910 11060 23962
rect 11060 23910 11072 23962
rect 11072 23910 11102 23962
rect 11126 23910 11136 23962
rect 11136 23910 11182 23962
rect 10886 23908 10942 23910
rect 10966 23908 11022 23910
rect 11046 23908 11102 23910
rect 11126 23908 11182 23910
rect 10886 22874 10942 22876
rect 10966 22874 11022 22876
rect 11046 22874 11102 22876
rect 11126 22874 11182 22876
rect 10886 22822 10932 22874
rect 10932 22822 10942 22874
rect 10966 22822 10996 22874
rect 10996 22822 11008 22874
rect 11008 22822 11022 22874
rect 11046 22822 11060 22874
rect 11060 22822 11072 22874
rect 11072 22822 11102 22874
rect 11126 22822 11136 22874
rect 11136 22822 11182 22874
rect 10886 22820 10942 22822
rect 10966 22820 11022 22822
rect 11046 22820 11102 22822
rect 11126 22820 11182 22822
rect 15852 40826 15908 40828
rect 15932 40826 15988 40828
rect 16012 40826 16068 40828
rect 16092 40826 16148 40828
rect 15852 40774 15898 40826
rect 15898 40774 15908 40826
rect 15932 40774 15962 40826
rect 15962 40774 15974 40826
rect 15974 40774 15988 40826
rect 16012 40774 16026 40826
rect 16026 40774 16038 40826
rect 16038 40774 16068 40826
rect 16092 40774 16102 40826
rect 16102 40774 16148 40826
rect 15852 40772 15908 40774
rect 15932 40772 15988 40774
rect 16012 40772 16068 40774
rect 16092 40772 16148 40774
rect 15852 39738 15908 39740
rect 15932 39738 15988 39740
rect 16012 39738 16068 39740
rect 16092 39738 16148 39740
rect 15852 39686 15898 39738
rect 15898 39686 15908 39738
rect 15932 39686 15962 39738
rect 15962 39686 15974 39738
rect 15974 39686 15988 39738
rect 16012 39686 16026 39738
rect 16026 39686 16038 39738
rect 16038 39686 16068 39738
rect 16092 39686 16102 39738
rect 16102 39686 16148 39738
rect 15852 39684 15908 39686
rect 15932 39684 15988 39686
rect 16012 39684 16068 39686
rect 16092 39684 16148 39686
rect 11610 26696 11666 26752
rect 10886 21786 10942 21788
rect 10966 21786 11022 21788
rect 11046 21786 11102 21788
rect 11126 21786 11182 21788
rect 10886 21734 10932 21786
rect 10932 21734 10942 21786
rect 10966 21734 10996 21786
rect 10996 21734 11008 21786
rect 11008 21734 11022 21786
rect 11046 21734 11060 21786
rect 11060 21734 11072 21786
rect 11072 21734 11102 21786
rect 11126 21734 11136 21786
rect 11136 21734 11182 21786
rect 10886 21732 10942 21734
rect 10966 21732 11022 21734
rect 11046 21732 11102 21734
rect 11126 21732 11182 21734
rect 10886 20698 10942 20700
rect 10966 20698 11022 20700
rect 11046 20698 11102 20700
rect 11126 20698 11182 20700
rect 10886 20646 10932 20698
rect 10932 20646 10942 20698
rect 10966 20646 10996 20698
rect 10996 20646 11008 20698
rect 11008 20646 11022 20698
rect 11046 20646 11060 20698
rect 11060 20646 11072 20698
rect 11072 20646 11102 20698
rect 11126 20646 11136 20698
rect 11136 20646 11182 20698
rect 10886 20644 10942 20646
rect 10966 20644 11022 20646
rect 11046 20644 11102 20646
rect 11126 20644 11182 20646
rect 10230 11736 10286 11792
rect 10322 11192 10378 11248
rect 10046 9580 10102 9616
rect 10046 9560 10048 9580
rect 10048 9560 10100 9580
rect 10100 9560 10102 9580
rect 10886 19610 10942 19612
rect 10966 19610 11022 19612
rect 11046 19610 11102 19612
rect 11126 19610 11182 19612
rect 10886 19558 10932 19610
rect 10932 19558 10942 19610
rect 10966 19558 10996 19610
rect 10996 19558 11008 19610
rect 11008 19558 11022 19610
rect 11046 19558 11060 19610
rect 11060 19558 11072 19610
rect 11072 19558 11102 19610
rect 11126 19558 11136 19610
rect 11136 19558 11182 19610
rect 10886 19556 10942 19558
rect 10966 19556 11022 19558
rect 11046 19556 11102 19558
rect 11126 19556 11182 19558
rect 15852 38650 15908 38652
rect 15932 38650 15988 38652
rect 16012 38650 16068 38652
rect 16092 38650 16148 38652
rect 15852 38598 15898 38650
rect 15898 38598 15908 38650
rect 15932 38598 15962 38650
rect 15962 38598 15974 38650
rect 15974 38598 15988 38650
rect 16012 38598 16026 38650
rect 16026 38598 16038 38650
rect 16038 38598 16068 38650
rect 16092 38598 16102 38650
rect 16102 38598 16148 38650
rect 15852 38596 15908 38598
rect 15932 38596 15988 38598
rect 16012 38596 16068 38598
rect 16092 38596 16148 38598
rect 15852 37562 15908 37564
rect 15932 37562 15988 37564
rect 16012 37562 16068 37564
rect 16092 37562 16148 37564
rect 15852 37510 15898 37562
rect 15898 37510 15908 37562
rect 15932 37510 15962 37562
rect 15962 37510 15974 37562
rect 15974 37510 15988 37562
rect 16012 37510 16026 37562
rect 16026 37510 16038 37562
rect 16038 37510 16068 37562
rect 16092 37510 16102 37562
rect 16102 37510 16148 37562
rect 15852 37508 15908 37510
rect 15932 37508 15988 37510
rect 16012 37508 16068 37510
rect 16092 37508 16148 37510
rect 15852 36474 15908 36476
rect 15932 36474 15988 36476
rect 16012 36474 16068 36476
rect 16092 36474 16148 36476
rect 15852 36422 15898 36474
rect 15898 36422 15908 36474
rect 15932 36422 15962 36474
rect 15962 36422 15974 36474
rect 15974 36422 15988 36474
rect 16012 36422 16026 36474
rect 16026 36422 16038 36474
rect 16038 36422 16068 36474
rect 16092 36422 16102 36474
rect 16102 36422 16148 36474
rect 15852 36420 15908 36422
rect 15932 36420 15988 36422
rect 16012 36420 16068 36422
rect 16092 36420 16148 36422
rect 15852 35386 15908 35388
rect 15932 35386 15988 35388
rect 16012 35386 16068 35388
rect 16092 35386 16148 35388
rect 15852 35334 15898 35386
rect 15898 35334 15908 35386
rect 15932 35334 15962 35386
rect 15962 35334 15974 35386
rect 15974 35334 15988 35386
rect 16012 35334 16026 35386
rect 16026 35334 16038 35386
rect 16038 35334 16068 35386
rect 16092 35334 16102 35386
rect 16102 35334 16148 35386
rect 15852 35332 15908 35334
rect 15932 35332 15988 35334
rect 16012 35332 16068 35334
rect 16092 35332 16148 35334
rect 15852 34298 15908 34300
rect 15932 34298 15988 34300
rect 16012 34298 16068 34300
rect 16092 34298 16148 34300
rect 15852 34246 15898 34298
rect 15898 34246 15908 34298
rect 15932 34246 15962 34298
rect 15962 34246 15974 34298
rect 15974 34246 15988 34298
rect 16012 34246 16026 34298
rect 16026 34246 16038 34298
rect 16038 34246 16068 34298
rect 16092 34246 16102 34298
rect 16102 34246 16148 34298
rect 15852 34244 15908 34246
rect 15932 34244 15988 34246
rect 16012 34244 16068 34246
rect 16092 34244 16148 34246
rect 15852 33210 15908 33212
rect 15932 33210 15988 33212
rect 16012 33210 16068 33212
rect 16092 33210 16148 33212
rect 15852 33158 15898 33210
rect 15898 33158 15908 33210
rect 15932 33158 15962 33210
rect 15962 33158 15974 33210
rect 15974 33158 15988 33210
rect 16012 33158 16026 33210
rect 16026 33158 16038 33210
rect 16038 33158 16068 33210
rect 16092 33158 16102 33210
rect 16102 33158 16148 33210
rect 15852 33156 15908 33158
rect 15932 33156 15988 33158
rect 16012 33156 16068 33158
rect 16092 33156 16148 33158
rect 15852 32122 15908 32124
rect 15932 32122 15988 32124
rect 16012 32122 16068 32124
rect 16092 32122 16148 32124
rect 15852 32070 15898 32122
rect 15898 32070 15908 32122
rect 15932 32070 15962 32122
rect 15962 32070 15974 32122
rect 15974 32070 15988 32122
rect 16012 32070 16026 32122
rect 16026 32070 16038 32122
rect 16038 32070 16068 32122
rect 16092 32070 16102 32122
rect 16102 32070 16148 32122
rect 15852 32068 15908 32070
rect 15932 32068 15988 32070
rect 16012 32068 16068 32070
rect 16092 32068 16148 32070
rect 14278 27512 14334 27568
rect 15852 31034 15908 31036
rect 15932 31034 15988 31036
rect 16012 31034 16068 31036
rect 16092 31034 16148 31036
rect 15852 30982 15898 31034
rect 15898 30982 15908 31034
rect 15932 30982 15962 31034
rect 15962 30982 15974 31034
rect 15974 30982 15988 31034
rect 16012 30982 16026 31034
rect 16026 30982 16038 31034
rect 16038 30982 16068 31034
rect 16092 30982 16102 31034
rect 16102 30982 16148 31034
rect 15852 30980 15908 30982
rect 15932 30980 15988 30982
rect 16012 30980 16068 30982
rect 16092 30980 16148 30982
rect 15852 29946 15908 29948
rect 15932 29946 15988 29948
rect 16012 29946 16068 29948
rect 16092 29946 16148 29948
rect 15852 29894 15898 29946
rect 15898 29894 15908 29946
rect 15932 29894 15962 29946
rect 15962 29894 15974 29946
rect 15974 29894 15988 29946
rect 16012 29894 16026 29946
rect 16026 29894 16038 29946
rect 16038 29894 16068 29946
rect 16092 29894 16102 29946
rect 16102 29894 16148 29946
rect 15852 29892 15908 29894
rect 15932 29892 15988 29894
rect 16012 29892 16068 29894
rect 16092 29892 16148 29894
rect 15852 28858 15908 28860
rect 15932 28858 15988 28860
rect 16012 28858 16068 28860
rect 16092 28858 16148 28860
rect 15852 28806 15898 28858
rect 15898 28806 15908 28858
rect 15932 28806 15962 28858
rect 15962 28806 15974 28858
rect 15974 28806 15988 28858
rect 16012 28806 16026 28858
rect 16026 28806 16038 28858
rect 16038 28806 16068 28858
rect 16092 28806 16102 28858
rect 16102 28806 16148 28858
rect 15852 28804 15908 28806
rect 15932 28804 15988 28806
rect 16012 28804 16068 28806
rect 16092 28804 16148 28806
rect 10886 18522 10942 18524
rect 10966 18522 11022 18524
rect 11046 18522 11102 18524
rect 11126 18522 11182 18524
rect 10886 18470 10932 18522
rect 10932 18470 10942 18522
rect 10966 18470 10996 18522
rect 10996 18470 11008 18522
rect 11008 18470 11022 18522
rect 11046 18470 11060 18522
rect 11060 18470 11072 18522
rect 11072 18470 11102 18522
rect 11126 18470 11136 18522
rect 11136 18470 11182 18522
rect 10886 18468 10942 18470
rect 10966 18468 11022 18470
rect 11046 18468 11102 18470
rect 11126 18468 11182 18470
rect 10886 17434 10942 17436
rect 10966 17434 11022 17436
rect 11046 17434 11102 17436
rect 11126 17434 11182 17436
rect 10886 17382 10932 17434
rect 10932 17382 10942 17434
rect 10966 17382 10996 17434
rect 10996 17382 11008 17434
rect 11008 17382 11022 17434
rect 11046 17382 11060 17434
rect 11060 17382 11072 17434
rect 11072 17382 11102 17434
rect 11126 17382 11136 17434
rect 11136 17382 11182 17434
rect 10886 17380 10942 17382
rect 10966 17380 11022 17382
rect 11046 17380 11102 17382
rect 11126 17380 11182 17382
rect 10886 16346 10942 16348
rect 10966 16346 11022 16348
rect 11046 16346 11102 16348
rect 11126 16346 11182 16348
rect 10886 16294 10932 16346
rect 10932 16294 10942 16346
rect 10966 16294 10996 16346
rect 10996 16294 11008 16346
rect 11008 16294 11022 16346
rect 11046 16294 11060 16346
rect 11060 16294 11072 16346
rect 11072 16294 11102 16346
rect 11126 16294 11136 16346
rect 11136 16294 11182 16346
rect 10886 16292 10942 16294
rect 10966 16292 11022 16294
rect 11046 16292 11102 16294
rect 11126 16292 11182 16294
rect 10690 16088 10746 16144
rect 10506 11736 10562 11792
rect 10506 8472 10562 8528
rect 10886 15258 10942 15260
rect 10966 15258 11022 15260
rect 11046 15258 11102 15260
rect 11126 15258 11182 15260
rect 10886 15206 10932 15258
rect 10932 15206 10942 15258
rect 10966 15206 10996 15258
rect 10996 15206 11008 15258
rect 11008 15206 11022 15258
rect 11046 15206 11060 15258
rect 11060 15206 11072 15258
rect 11072 15206 11102 15258
rect 11126 15206 11136 15258
rect 11136 15206 11182 15258
rect 10886 15204 10942 15206
rect 10966 15204 11022 15206
rect 11046 15204 11102 15206
rect 11126 15204 11182 15206
rect 11242 14320 11298 14376
rect 12346 14456 12402 14512
rect 10886 14170 10942 14172
rect 10966 14170 11022 14172
rect 11046 14170 11102 14172
rect 11126 14170 11182 14172
rect 10886 14118 10932 14170
rect 10932 14118 10942 14170
rect 10966 14118 10996 14170
rect 10996 14118 11008 14170
rect 11008 14118 11022 14170
rect 11046 14118 11060 14170
rect 11060 14118 11072 14170
rect 11072 14118 11102 14170
rect 11126 14118 11136 14170
rect 11136 14118 11182 14170
rect 10886 14116 10942 14118
rect 10966 14116 11022 14118
rect 11046 14116 11102 14118
rect 11126 14116 11182 14118
rect 11886 14320 11942 14376
rect 10886 13082 10942 13084
rect 10966 13082 11022 13084
rect 11046 13082 11102 13084
rect 11126 13082 11182 13084
rect 10886 13030 10932 13082
rect 10932 13030 10942 13082
rect 10966 13030 10996 13082
rect 10996 13030 11008 13082
rect 11008 13030 11022 13082
rect 11046 13030 11060 13082
rect 11060 13030 11072 13082
rect 11072 13030 11102 13082
rect 11126 13030 11136 13082
rect 11136 13030 11182 13082
rect 10886 13028 10942 13030
rect 10966 13028 11022 13030
rect 11046 13028 11102 13030
rect 11126 13028 11182 13030
rect 10886 11994 10942 11996
rect 10966 11994 11022 11996
rect 11046 11994 11102 11996
rect 11126 11994 11182 11996
rect 10886 11942 10932 11994
rect 10932 11942 10942 11994
rect 10966 11942 10996 11994
rect 10996 11942 11008 11994
rect 11008 11942 11022 11994
rect 11046 11942 11060 11994
rect 11060 11942 11072 11994
rect 11072 11942 11102 11994
rect 11126 11942 11136 11994
rect 11136 11942 11182 11994
rect 10886 11940 10942 11942
rect 10966 11940 11022 11942
rect 11046 11940 11102 11942
rect 11126 11940 11182 11942
rect 11978 11192 12034 11248
rect 10886 10906 10942 10908
rect 10966 10906 11022 10908
rect 11046 10906 11102 10908
rect 11126 10906 11182 10908
rect 10886 10854 10932 10906
rect 10932 10854 10942 10906
rect 10966 10854 10996 10906
rect 10996 10854 11008 10906
rect 11008 10854 11022 10906
rect 11046 10854 11060 10906
rect 11060 10854 11072 10906
rect 11072 10854 11102 10906
rect 11126 10854 11136 10906
rect 11136 10854 11182 10906
rect 10886 10852 10942 10854
rect 10966 10852 11022 10854
rect 11046 10852 11102 10854
rect 11126 10852 11182 10854
rect 10886 9818 10942 9820
rect 10966 9818 11022 9820
rect 11046 9818 11102 9820
rect 11126 9818 11182 9820
rect 10886 9766 10932 9818
rect 10932 9766 10942 9818
rect 10966 9766 10996 9818
rect 10996 9766 11008 9818
rect 11008 9766 11022 9818
rect 11046 9766 11060 9818
rect 11060 9766 11072 9818
rect 11072 9766 11102 9818
rect 11126 9766 11136 9818
rect 11136 9766 11182 9818
rect 10886 9764 10942 9766
rect 10966 9764 11022 9766
rect 11046 9764 11102 9766
rect 11126 9764 11182 9766
rect 10886 8730 10942 8732
rect 10966 8730 11022 8732
rect 11046 8730 11102 8732
rect 11126 8730 11182 8732
rect 10886 8678 10932 8730
rect 10932 8678 10942 8730
rect 10966 8678 10996 8730
rect 10996 8678 11008 8730
rect 11008 8678 11022 8730
rect 11046 8678 11060 8730
rect 11060 8678 11072 8730
rect 11072 8678 11102 8730
rect 11126 8678 11136 8730
rect 11136 8678 11182 8730
rect 10886 8676 10942 8678
rect 10966 8676 11022 8678
rect 11046 8676 11102 8678
rect 11126 8676 11182 8678
rect 10886 7642 10942 7644
rect 10966 7642 11022 7644
rect 11046 7642 11102 7644
rect 11126 7642 11182 7644
rect 10886 7590 10932 7642
rect 10932 7590 10942 7642
rect 10966 7590 10996 7642
rect 10996 7590 11008 7642
rect 11008 7590 11022 7642
rect 11046 7590 11060 7642
rect 11060 7590 11072 7642
rect 11072 7590 11102 7642
rect 11126 7590 11136 7642
rect 11136 7590 11182 7642
rect 10886 7588 10942 7590
rect 10966 7588 11022 7590
rect 11046 7588 11102 7590
rect 11126 7588 11182 7590
rect 11794 8508 11796 8528
rect 11796 8508 11848 8528
rect 11848 8508 11850 8528
rect 11794 8472 11850 8508
rect 10886 6554 10942 6556
rect 10966 6554 11022 6556
rect 11046 6554 11102 6556
rect 11126 6554 11182 6556
rect 10886 6502 10932 6554
rect 10932 6502 10942 6554
rect 10966 6502 10996 6554
rect 10996 6502 11008 6554
rect 11008 6502 11022 6554
rect 11046 6502 11060 6554
rect 11060 6502 11072 6554
rect 11072 6502 11102 6554
rect 11126 6502 11136 6554
rect 11136 6502 11182 6554
rect 10886 6500 10942 6502
rect 10966 6500 11022 6502
rect 11046 6500 11102 6502
rect 11126 6500 11182 6502
rect 10886 5466 10942 5468
rect 10966 5466 11022 5468
rect 11046 5466 11102 5468
rect 11126 5466 11182 5468
rect 10886 5414 10932 5466
rect 10932 5414 10942 5466
rect 10966 5414 10996 5466
rect 10996 5414 11008 5466
rect 11008 5414 11022 5466
rect 11046 5414 11060 5466
rect 11060 5414 11072 5466
rect 11072 5414 11102 5466
rect 11126 5414 11136 5466
rect 11136 5414 11182 5466
rect 10886 5412 10942 5414
rect 10966 5412 11022 5414
rect 11046 5412 11102 5414
rect 11126 5412 11182 5414
rect 10886 4378 10942 4380
rect 10966 4378 11022 4380
rect 11046 4378 11102 4380
rect 11126 4378 11182 4380
rect 10886 4326 10932 4378
rect 10932 4326 10942 4378
rect 10966 4326 10996 4378
rect 10996 4326 11008 4378
rect 11008 4326 11022 4378
rect 11046 4326 11060 4378
rect 11060 4326 11072 4378
rect 11072 4326 11102 4378
rect 11126 4326 11136 4378
rect 11136 4326 11182 4378
rect 10886 4324 10942 4326
rect 10966 4324 11022 4326
rect 11046 4324 11102 4326
rect 11126 4324 11182 4326
rect 10886 3290 10942 3292
rect 10966 3290 11022 3292
rect 11046 3290 11102 3292
rect 11126 3290 11182 3292
rect 10886 3238 10932 3290
rect 10932 3238 10942 3290
rect 10966 3238 10996 3290
rect 10996 3238 11008 3290
rect 11008 3238 11022 3290
rect 11046 3238 11060 3290
rect 11060 3238 11072 3290
rect 11072 3238 11102 3290
rect 11126 3238 11136 3290
rect 11136 3238 11182 3290
rect 10886 3236 10942 3238
rect 10966 3236 11022 3238
rect 11046 3236 11102 3238
rect 11126 3236 11182 3238
rect 12806 11328 12862 11384
rect 11886 3984 11942 4040
rect 11978 3476 11980 3496
rect 11980 3476 12032 3496
rect 12032 3476 12034 3496
rect 11978 3440 12034 3476
rect 10886 2202 10942 2204
rect 10966 2202 11022 2204
rect 11046 2202 11102 2204
rect 11126 2202 11182 2204
rect 10886 2150 10932 2202
rect 10932 2150 10942 2202
rect 10966 2150 10996 2202
rect 10996 2150 11008 2202
rect 11008 2150 11022 2202
rect 11046 2150 11060 2202
rect 11060 2150 11072 2202
rect 11072 2150 11102 2202
rect 11126 2150 11136 2202
rect 11136 2150 11182 2202
rect 10886 2148 10942 2150
rect 10966 2148 11022 2150
rect 11046 2148 11102 2150
rect 11126 2148 11182 2150
rect 2870 312 2926 368
rect 13726 13932 13782 13968
rect 13726 13912 13728 13932
rect 13728 13912 13780 13932
rect 13780 13912 13782 13932
rect 15852 27770 15908 27772
rect 15932 27770 15988 27772
rect 16012 27770 16068 27772
rect 16092 27770 16148 27772
rect 15852 27718 15898 27770
rect 15898 27718 15908 27770
rect 15932 27718 15962 27770
rect 15962 27718 15974 27770
rect 15974 27718 15988 27770
rect 16012 27718 16026 27770
rect 16026 27718 16038 27770
rect 16038 27718 16068 27770
rect 16092 27718 16102 27770
rect 16102 27718 16148 27770
rect 15852 27716 15908 27718
rect 15932 27716 15988 27718
rect 16012 27716 16068 27718
rect 16092 27716 16148 27718
rect 15852 26682 15908 26684
rect 15932 26682 15988 26684
rect 16012 26682 16068 26684
rect 16092 26682 16148 26684
rect 15852 26630 15898 26682
rect 15898 26630 15908 26682
rect 15932 26630 15962 26682
rect 15962 26630 15974 26682
rect 15974 26630 15988 26682
rect 16012 26630 16026 26682
rect 16026 26630 16038 26682
rect 16038 26630 16068 26682
rect 16092 26630 16102 26682
rect 16102 26630 16148 26682
rect 15852 26628 15908 26630
rect 15932 26628 15988 26630
rect 16012 26628 16068 26630
rect 16092 26628 16148 26630
rect 15852 25594 15908 25596
rect 15932 25594 15988 25596
rect 16012 25594 16068 25596
rect 16092 25594 16148 25596
rect 15852 25542 15898 25594
rect 15898 25542 15908 25594
rect 15932 25542 15962 25594
rect 15962 25542 15974 25594
rect 15974 25542 15988 25594
rect 16012 25542 16026 25594
rect 16026 25542 16038 25594
rect 16038 25542 16068 25594
rect 16092 25542 16102 25594
rect 16102 25542 16148 25594
rect 15852 25540 15908 25542
rect 15932 25540 15988 25542
rect 16012 25540 16068 25542
rect 16092 25540 16148 25542
rect 15852 24506 15908 24508
rect 15932 24506 15988 24508
rect 16012 24506 16068 24508
rect 16092 24506 16148 24508
rect 15852 24454 15898 24506
rect 15898 24454 15908 24506
rect 15932 24454 15962 24506
rect 15962 24454 15974 24506
rect 15974 24454 15988 24506
rect 16012 24454 16026 24506
rect 16026 24454 16038 24506
rect 16038 24454 16068 24506
rect 16092 24454 16102 24506
rect 16102 24454 16148 24506
rect 15852 24452 15908 24454
rect 15932 24452 15988 24454
rect 16012 24452 16068 24454
rect 16092 24452 16148 24454
rect 15852 23418 15908 23420
rect 15932 23418 15988 23420
rect 16012 23418 16068 23420
rect 16092 23418 16148 23420
rect 15852 23366 15898 23418
rect 15898 23366 15908 23418
rect 15932 23366 15962 23418
rect 15962 23366 15974 23418
rect 15974 23366 15988 23418
rect 16012 23366 16026 23418
rect 16026 23366 16038 23418
rect 16038 23366 16068 23418
rect 16092 23366 16102 23418
rect 16102 23366 16148 23418
rect 15852 23364 15908 23366
rect 15932 23364 15988 23366
rect 16012 23364 16068 23366
rect 16092 23364 16148 23366
rect 15852 22330 15908 22332
rect 15932 22330 15988 22332
rect 16012 22330 16068 22332
rect 16092 22330 16148 22332
rect 15852 22278 15898 22330
rect 15898 22278 15908 22330
rect 15932 22278 15962 22330
rect 15962 22278 15974 22330
rect 15974 22278 15988 22330
rect 16012 22278 16026 22330
rect 16026 22278 16038 22330
rect 16038 22278 16068 22330
rect 16092 22278 16102 22330
rect 16102 22278 16148 22330
rect 15852 22276 15908 22278
rect 15932 22276 15988 22278
rect 16012 22276 16068 22278
rect 16092 22276 16148 22278
rect 15750 22072 15806 22128
rect 16210 21936 16266 21992
rect 15852 21242 15908 21244
rect 15932 21242 15988 21244
rect 16012 21242 16068 21244
rect 16092 21242 16148 21244
rect 15852 21190 15898 21242
rect 15898 21190 15908 21242
rect 15932 21190 15962 21242
rect 15962 21190 15974 21242
rect 15974 21190 15988 21242
rect 16012 21190 16026 21242
rect 16026 21190 16038 21242
rect 16038 21190 16068 21242
rect 16092 21190 16102 21242
rect 16102 21190 16148 21242
rect 15852 21188 15908 21190
rect 15932 21188 15988 21190
rect 16012 21188 16068 21190
rect 16092 21188 16148 21190
rect 15852 20154 15908 20156
rect 15932 20154 15988 20156
rect 16012 20154 16068 20156
rect 16092 20154 16148 20156
rect 15852 20102 15898 20154
rect 15898 20102 15908 20154
rect 15932 20102 15962 20154
rect 15962 20102 15974 20154
rect 15974 20102 15988 20154
rect 16012 20102 16026 20154
rect 16026 20102 16038 20154
rect 16038 20102 16068 20154
rect 16092 20102 16102 20154
rect 16102 20102 16148 20154
rect 15852 20100 15908 20102
rect 15932 20100 15988 20102
rect 16012 20100 16068 20102
rect 16092 20100 16148 20102
rect 16578 22616 16634 22672
rect 15198 11328 15254 11384
rect 15852 19066 15908 19068
rect 15932 19066 15988 19068
rect 16012 19066 16068 19068
rect 16092 19066 16148 19068
rect 15852 19014 15898 19066
rect 15898 19014 15908 19066
rect 15932 19014 15962 19066
rect 15962 19014 15974 19066
rect 15974 19014 15988 19066
rect 16012 19014 16026 19066
rect 16026 19014 16038 19066
rect 16038 19014 16068 19066
rect 16092 19014 16102 19066
rect 16102 19014 16148 19066
rect 15852 19012 15908 19014
rect 15932 19012 15988 19014
rect 16012 19012 16068 19014
rect 16092 19012 16148 19014
rect 15852 17978 15908 17980
rect 15932 17978 15988 17980
rect 16012 17978 16068 17980
rect 16092 17978 16148 17980
rect 15852 17926 15898 17978
rect 15898 17926 15908 17978
rect 15932 17926 15962 17978
rect 15962 17926 15974 17978
rect 15974 17926 15988 17978
rect 16012 17926 16026 17978
rect 16026 17926 16038 17978
rect 16038 17926 16068 17978
rect 16092 17926 16102 17978
rect 16102 17926 16148 17978
rect 15852 17924 15908 17926
rect 15932 17924 15988 17926
rect 16012 17924 16068 17926
rect 16092 17924 16148 17926
rect 15852 16890 15908 16892
rect 15932 16890 15988 16892
rect 16012 16890 16068 16892
rect 16092 16890 16148 16892
rect 15852 16838 15898 16890
rect 15898 16838 15908 16890
rect 15932 16838 15962 16890
rect 15962 16838 15974 16890
rect 15974 16838 15988 16890
rect 16012 16838 16026 16890
rect 16026 16838 16038 16890
rect 16038 16838 16068 16890
rect 16092 16838 16102 16890
rect 16102 16838 16148 16890
rect 15852 16836 15908 16838
rect 15932 16836 15988 16838
rect 16012 16836 16068 16838
rect 16092 16836 16148 16838
rect 15852 15802 15908 15804
rect 15932 15802 15988 15804
rect 16012 15802 16068 15804
rect 16092 15802 16148 15804
rect 15852 15750 15898 15802
rect 15898 15750 15908 15802
rect 15932 15750 15962 15802
rect 15962 15750 15974 15802
rect 15974 15750 15988 15802
rect 16012 15750 16026 15802
rect 16026 15750 16038 15802
rect 16038 15750 16068 15802
rect 16092 15750 16102 15802
rect 16102 15750 16148 15802
rect 15852 15748 15908 15750
rect 15932 15748 15988 15750
rect 16012 15748 16068 15750
rect 16092 15748 16148 15750
rect 15852 14714 15908 14716
rect 15932 14714 15988 14716
rect 16012 14714 16068 14716
rect 16092 14714 16148 14716
rect 15852 14662 15898 14714
rect 15898 14662 15908 14714
rect 15932 14662 15962 14714
rect 15962 14662 15974 14714
rect 15974 14662 15988 14714
rect 16012 14662 16026 14714
rect 16026 14662 16038 14714
rect 16038 14662 16068 14714
rect 16092 14662 16102 14714
rect 16102 14662 16148 14714
rect 15852 14660 15908 14662
rect 15932 14660 15988 14662
rect 16012 14660 16068 14662
rect 16092 14660 16148 14662
rect 16302 14456 16358 14512
rect 15852 13626 15908 13628
rect 15932 13626 15988 13628
rect 16012 13626 16068 13628
rect 16092 13626 16148 13628
rect 15852 13574 15898 13626
rect 15898 13574 15908 13626
rect 15932 13574 15962 13626
rect 15962 13574 15974 13626
rect 15974 13574 15988 13626
rect 16012 13574 16026 13626
rect 16026 13574 16038 13626
rect 16038 13574 16068 13626
rect 16092 13574 16102 13626
rect 16102 13574 16148 13626
rect 15852 13572 15908 13574
rect 15932 13572 15988 13574
rect 16012 13572 16068 13574
rect 16092 13572 16148 13574
rect 15852 12538 15908 12540
rect 15932 12538 15988 12540
rect 16012 12538 16068 12540
rect 16092 12538 16148 12540
rect 15852 12486 15898 12538
rect 15898 12486 15908 12538
rect 15932 12486 15962 12538
rect 15962 12486 15974 12538
rect 15974 12486 15988 12538
rect 16012 12486 16026 12538
rect 16026 12486 16038 12538
rect 16038 12486 16068 12538
rect 16092 12486 16102 12538
rect 16102 12486 16148 12538
rect 15852 12484 15908 12486
rect 15932 12484 15988 12486
rect 16012 12484 16068 12486
rect 16092 12484 16148 12486
rect 15852 11450 15908 11452
rect 15932 11450 15988 11452
rect 16012 11450 16068 11452
rect 16092 11450 16148 11452
rect 15852 11398 15898 11450
rect 15898 11398 15908 11450
rect 15932 11398 15962 11450
rect 15962 11398 15974 11450
rect 15974 11398 15988 11450
rect 16012 11398 16026 11450
rect 16026 11398 16038 11450
rect 16038 11398 16068 11450
rect 16092 11398 16102 11450
rect 16102 11398 16148 11450
rect 15852 11396 15908 11398
rect 15932 11396 15988 11398
rect 16012 11396 16068 11398
rect 16092 11396 16148 11398
rect 15852 10362 15908 10364
rect 15932 10362 15988 10364
rect 16012 10362 16068 10364
rect 16092 10362 16148 10364
rect 15852 10310 15898 10362
rect 15898 10310 15908 10362
rect 15932 10310 15962 10362
rect 15962 10310 15974 10362
rect 15974 10310 15988 10362
rect 16012 10310 16026 10362
rect 16026 10310 16038 10362
rect 16038 10310 16068 10362
rect 16092 10310 16102 10362
rect 16102 10310 16148 10362
rect 15852 10308 15908 10310
rect 15932 10308 15988 10310
rect 16012 10308 16068 10310
rect 16092 10308 16148 10310
rect 15658 9596 15660 9616
rect 15660 9596 15712 9616
rect 15712 9596 15714 9616
rect 15658 9560 15714 9596
rect 15852 9274 15908 9276
rect 15932 9274 15988 9276
rect 16012 9274 16068 9276
rect 16092 9274 16148 9276
rect 15852 9222 15898 9274
rect 15898 9222 15908 9274
rect 15932 9222 15962 9274
rect 15962 9222 15974 9274
rect 15974 9222 15988 9274
rect 16012 9222 16026 9274
rect 16026 9222 16038 9274
rect 16038 9222 16068 9274
rect 16092 9222 16102 9274
rect 16102 9222 16148 9274
rect 15852 9220 15908 9222
rect 15932 9220 15988 9222
rect 16012 9220 16068 9222
rect 16092 9220 16148 9222
rect 15852 8186 15908 8188
rect 15932 8186 15988 8188
rect 16012 8186 16068 8188
rect 16092 8186 16148 8188
rect 15852 8134 15898 8186
rect 15898 8134 15908 8186
rect 15932 8134 15962 8186
rect 15962 8134 15974 8186
rect 15974 8134 15988 8186
rect 16012 8134 16026 8186
rect 16026 8134 16038 8186
rect 16038 8134 16068 8186
rect 16092 8134 16102 8186
rect 16102 8134 16148 8186
rect 15852 8132 15908 8134
rect 15932 8132 15988 8134
rect 16012 8132 16068 8134
rect 16092 8132 16148 8134
rect 15852 7098 15908 7100
rect 15932 7098 15988 7100
rect 16012 7098 16068 7100
rect 16092 7098 16148 7100
rect 15852 7046 15898 7098
rect 15898 7046 15908 7098
rect 15932 7046 15962 7098
rect 15962 7046 15974 7098
rect 15974 7046 15988 7098
rect 16012 7046 16026 7098
rect 16026 7046 16038 7098
rect 16038 7046 16068 7098
rect 16092 7046 16102 7098
rect 16102 7046 16148 7098
rect 15852 7044 15908 7046
rect 15932 7044 15988 7046
rect 16012 7044 16068 7046
rect 16092 7044 16148 7046
rect 15852 6010 15908 6012
rect 15932 6010 15988 6012
rect 16012 6010 16068 6012
rect 16092 6010 16148 6012
rect 15852 5958 15898 6010
rect 15898 5958 15908 6010
rect 15932 5958 15962 6010
rect 15962 5958 15974 6010
rect 15974 5958 15988 6010
rect 16012 5958 16026 6010
rect 16026 5958 16038 6010
rect 16038 5958 16068 6010
rect 16092 5958 16102 6010
rect 16102 5958 16148 6010
rect 15852 5956 15908 5958
rect 15932 5956 15988 5958
rect 16012 5956 16068 5958
rect 16092 5956 16148 5958
rect 16762 22752 16818 22808
rect 16578 19760 16634 19816
rect 17130 21664 17186 21720
rect 16670 16224 16726 16280
rect 16946 15816 17002 15872
rect 18050 29996 18052 30016
rect 18052 29996 18104 30016
rect 18104 29996 18106 30016
rect 18050 29960 18106 29996
rect 30102 43968 30158 44024
rect 25782 43002 25838 43004
rect 25862 43002 25918 43004
rect 25942 43002 25998 43004
rect 26022 43002 26078 43004
rect 25782 42950 25828 43002
rect 25828 42950 25838 43002
rect 25862 42950 25892 43002
rect 25892 42950 25904 43002
rect 25904 42950 25918 43002
rect 25942 42950 25956 43002
rect 25956 42950 25968 43002
rect 25968 42950 25998 43002
rect 26022 42950 26032 43002
rect 26032 42950 26078 43002
rect 25782 42948 25838 42950
rect 25862 42948 25918 42950
rect 25942 42948 25998 42950
rect 26022 42948 26078 42950
rect 20817 42458 20873 42460
rect 20897 42458 20953 42460
rect 20977 42458 21033 42460
rect 21057 42458 21113 42460
rect 20817 42406 20863 42458
rect 20863 42406 20873 42458
rect 20897 42406 20927 42458
rect 20927 42406 20939 42458
rect 20939 42406 20953 42458
rect 20977 42406 20991 42458
rect 20991 42406 21003 42458
rect 21003 42406 21033 42458
rect 21057 42406 21067 42458
rect 21067 42406 21113 42458
rect 20817 42404 20873 42406
rect 20897 42404 20953 42406
rect 20977 42404 21033 42406
rect 21057 42404 21113 42406
rect 25782 41914 25838 41916
rect 25862 41914 25918 41916
rect 25942 41914 25998 41916
rect 26022 41914 26078 41916
rect 25782 41862 25828 41914
rect 25828 41862 25838 41914
rect 25862 41862 25892 41914
rect 25892 41862 25904 41914
rect 25904 41862 25918 41914
rect 25942 41862 25956 41914
rect 25956 41862 25968 41914
rect 25968 41862 25998 41914
rect 26022 41862 26032 41914
rect 26032 41862 26078 41914
rect 25782 41860 25838 41862
rect 25862 41860 25918 41862
rect 25942 41860 25998 41862
rect 26022 41860 26078 41862
rect 30102 42472 30158 42528
rect 20817 41370 20873 41372
rect 20897 41370 20953 41372
rect 20977 41370 21033 41372
rect 21057 41370 21113 41372
rect 20817 41318 20863 41370
rect 20863 41318 20873 41370
rect 20897 41318 20927 41370
rect 20927 41318 20939 41370
rect 20939 41318 20953 41370
rect 20977 41318 20991 41370
rect 20991 41318 21003 41370
rect 21003 41318 21033 41370
rect 21057 41318 21067 41370
rect 21067 41318 21113 41370
rect 20817 41316 20873 41318
rect 20897 41316 20953 41318
rect 20977 41316 21033 41318
rect 21057 41316 21113 41318
rect 20817 40282 20873 40284
rect 20897 40282 20953 40284
rect 20977 40282 21033 40284
rect 21057 40282 21113 40284
rect 20817 40230 20863 40282
rect 20863 40230 20873 40282
rect 20897 40230 20927 40282
rect 20927 40230 20939 40282
rect 20939 40230 20953 40282
rect 20977 40230 20991 40282
rect 20991 40230 21003 40282
rect 21003 40230 21033 40282
rect 21057 40230 21067 40282
rect 21067 40230 21113 40282
rect 20817 40228 20873 40230
rect 20897 40228 20953 40230
rect 20977 40228 21033 40230
rect 21057 40228 21113 40230
rect 30102 40976 30158 41032
rect 25782 40826 25838 40828
rect 25862 40826 25918 40828
rect 25942 40826 25998 40828
rect 26022 40826 26078 40828
rect 25782 40774 25828 40826
rect 25828 40774 25838 40826
rect 25862 40774 25892 40826
rect 25892 40774 25904 40826
rect 25904 40774 25918 40826
rect 25942 40774 25956 40826
rect 25956 40774 25968 40826
rect 25968 40774 25998 40826
rect 26022 40774 26032 40826
rect 26032 40774 26078 40826
rect 25782 40772 25838 40774
rect 25862 40772 25918 40774
rect 25942 40772 25998 40774
rect 26022 40772 26078 40774
rect 25782 39738 25838 39740
rect 25862 39738 25918 39740
rect 25942 39738 25998 39740
rect 26022 39738 26078 39740
rect 25782 39686 25828 39738
rect 25828 39686 25838 39738
rect 25862 39686 25892 39738
rect 25892 39686 25904 39738
rect 25904 39686 25918 39738
rect 25942 39686 25956 39738
rect 25956 39686 25968 39738
rect 25968 39686 25998 39738
rect 26022 39686 26032 39738
rect 26032 39686 26078 39738
rect 25782 39684 25838 39686
rect 25862 39684 25918 39686
rect 25942 39684 25998 39686
rect 26022 39684 26078 39686
rect 20817 39194 20873 39196
rect 20897 39194 20953 39196
rect 20977 39194 21033 39196
rect 21057 39194 21113 39196
rect 20817 39142 20863 39194
rect 20863 39142 20873 39194
rect 20897 39142 20927 39194
rect 20927 39142 20939 39194
rect 20939 39142 20953 39194
rect 20977 39142 20991 39194
rect 20991 39142 21003 39194
rect 21003 39142 21033 39194
rect 21057 39142 21067 39194
rect 21067 39142 21113 39194
rect 20817 39140 20873 39142
rect 20897 39140 20953 39142
rect 20977 39140 21033 39142
rect 21057 39140 21113 39142
rect 17314 19760 17370 19816
rect 17590 21664 17646 21720
rect 17682 15952 17738 16008
rect 18050 23060 18052 23080
rect 18052 23060 18104 23080
rect 18104 23060 18106 23080
rect 18050 23024 18106 23060
rect 18050 16108 18106 16144
rect 18050 16088 18052 16108
rect 18052 16088 18104 16108
rect 18104 16088 18106 16108
rect 17038 13640 17094 13696
rect 17958 13932 18014 13968
rect 17958 13912 17960 13932
rect 17960 13912 18012 13932
rect 18012 13912 18014 13932
rect 15852 4922 15908 4924
rect 15932 4922 15988 4924
rect 16012 4922 16068 4924
rect 16092 4922 16148 4924
rect 15852 4870 15898 4922
rect 15898 4870 15908 4922
rect 15932 4870 15962 4922
rect 15962 4870 15974 4922
rect 15974 4870 15988 4922
rect 16012 4870 16026 4922
rect 16026 4870 16038 4922
rect 16038 4870 16068 4922
rect 16092 4870 16102 4922
rect 16102 4870 16148 4922
rect 15852 4868 15908 4870
rect 15932 4868 15988 4870
rect 16012 4868 16068 4870
rect 16092 4868 16148 4870
rect 15852 3834 15908 3836
rect 15932 3834 15988 3836
rect 16012 3834 16068 3836
rect 16092 3834 16148 3836
rect 15852 3782 15898 3834
rect 15898 3782 15908 3834
rect 15932 3782 15962 3834
rect 15962 3782 15974 3834
rect 15974 3782 15988 3834
rect 16012 3782 16026 3834
rect 16026 3782 16038 3834
rect 16038 3782 16068 3834
rect 16092 3782 16102 3834
rect 16102 3782 16148 3834
rect 15852 3780 15908 3782
rect 15932 3780 15988 3782
rect 16012 3780 16068 3782
rect 16092 3780 16148 3782
rect 18326 14356 18328 14376
rect 18328 14356 18380 14376
rect 18380 14356 18382 14376
rect 18326 14320 18382 14356
rect 18326 13676 18328 13696
rect 18328 13676 18380 13696
rect 18380 13676 18382 13696
rect 18326 13640 18382 13676
rect 18602 21664 18658 21720
rect 19062 23024 19118 23080
rect 20817 38106 20873 38108
rect 20897 38106 20953 38108
rect 20977 38106 21033 38108
rect 21057 38106 21113 38108
rect 20817 38054 20863 38106
rect 20863 38054 20873 38106
rect 20897 38054 20927 38106
rect 20927 38054 20939 38106
rect 20939 38054 20953 38106
rect 20977 38054 20991 38106
rect 20991 38054 21003 38106
rect 21003 38054 21033 38106
rect 21057 38054 21067 38106
rect 21067 38054 21113 38106
rect 20817 38052 20873 38054
rect 20897 38052 20953 38054
rect 20977 38052 21033 38054
rect 21057 38052 21113 38054
rect 19982 25744 20038 25800
rect 19246 21664 19302 21720
rect 18694 16244 18750 16280
rect 18694 16224 18696 16244
rect 18696 16224 18748 16244
rect 18748 16224 18750 16244
rect 18602 15952 18658 16008
rect 19062 15816 19118 15872
rect 16486 3068 16488 3088
rect 16488 3068 16540 3088
rect 16540 3068 16542 3088
rect 16486 3032 16542 3068
rect 17222 3440 17278 3496
rect 15852 2746 15908 2748
rect 15932 2746 15988 2748
rect 16012 2746 16068 2748
rect 16092 2746 16148 2748
rect 15852 2694 15898 2746
rect 15898 2694 15908 2746
rect 15932 2694 15962 2746
rect 15962 2694 15974 2746
rect 15974 2694 15988 2746
rect 16012 2694 16026 2746
rect 16026 2694 16038 2746
rect 16038 2694 16068 2746
rect 16092 2694 16102 2746
rect 16102 2694 16148 2746
rect 15852 2692 15908 2694
rect 15932 2692 15988 2694
rect 16012 2692 16068 2694
rect 16092 2692 16148 2694
rect 17866 3032 17922 3088
rect 20817 37018 20873 37020
rect 20897 37018 20953 37020
rect 20977 37018 21033 37020
rect 21057 37018 21113 37020
rect 20817 36966 20863 37018
rect 20863 36966 20873 37018
rect 20897 36966 20927 37018
rect 20927 36966 20939 37018
rect 20939 36966 20953 37018
rect 20977 36966 20991 37018
rect 20991 36966 21003 37018
rect 21003 36966 21033 37018
rect 21057 36966 21067 37018
rect 21067 36966 21113 37018
rect 20817 36964 20873 36966
rect 20897 36964 20953 36966
rect 20977 36964 21033 36966
rect 21057 36964 21113 36966
rect 20817 35930 20873 35932
rect 20897 35930 20953 35932
rect 20977 35930 21033 35932
rect 21057 35930 21113 35932
rect 20817 35878 20863 35930
rect 20863 35878 20873 35930
rect 20897 35878 20927 35930
rect 20927 35878 20939 35930
rect 20939 35878 20953 35930
rect 20977 35878 20991 35930
rect 20991 35878 21003 35930
rect 21003 35878 21033 35930
rect 21057 35878 21067 35930
rect 21067 35878 21113 35930
rect 20817 35876 20873 35878
rect 20897 35876 20953 35878
rect 20977 35876 21033 35878
rect 21057 35876 21113 35878
rect 20817 34842 20873 34844
rect 20897 34842 20953 34844
rect 20977 34842 21033 34844
rect 21057 34842 21113 34844
rect 20817 34790 20863 34842
rect 20863 34790 20873 34842
rect 20897 34790 20927 34842
rect 20927 34790 20939 34842
rect 20939 34790 20953 34842
rect 20977 34790 20991 34842
rect 20991 34790 21003 34842
rect 21003 34790 21033 34842
rect 21057 34790 21067 34842
rect 21067 34790 21113 34842
rect 20817 34788 20873 34790
rect 20897 34788 20953 34790
rect 20977 34788 21033 34790
rect 21057 34788 21113 34790
rect 20817 33754 20873 33756
rect 20897 33754 20953 33756
rect 20977 33754 21033 33756
rect 21057 33754 21113 33756
rect 20817 33702 20863 33754
rect 20863 33702 20873 33754
rect 20897 33702 20927 33754
rect 20927 33702 20939 33754
rect 20939 33702 20953 33754
rect 20977 33702 20991 33754
rect 20991 33702 21003 33754
rect 21003 33702 21033 33754
rect 21057 33702 21067 33754
rect 21067 33702 21113 33754
rect 20817 33700 20873 33702
rect 20897 33700 20953 33702
rect 20977 33700 21033 33702
rect 21057 33700 21113 33702
rect 20817 32666 20873 32668
rect 20897 32666 20953 32668
rect 20977 32666 21033 32668
rect 21057 32666 21113 32668
rect 20817 32614 20863 32666
rect 20863 32614 20873 32666
rect 20897 32614 20927 32666
rect 20927 32614 20939 32666
rect 20939 32614 20953 32666
rect 20977 32614 20991 32666
rect 20991 32614 21003 32666
rect 21003 32614 21033 32666
rect 21057 32614 21067 32666
rect 21067 32614 21113 32666
rect 20817 32612 20873 32614
rect 20897 32612 20953 32614
rect 20977 32612 21033 32614
rect 21057 32612 21113 32614
rect 20817 31578 20873 31580
rect 20897 31578 20953 31580
rect 20977 31578 21033 31580
rect 21057 31578 21113 31580
rect 20817 31526 20863 31578
rect 20863 31526 20873 31578
rect 20897 31526 20927 31578
rect 20927 31526 20939 31578
rect 20939 31526 20953 31578
rect 20977 31526 20991 31578
rect 20991 31526 21003 31578
rect 21003 31526 21033 31578
rect 21057 31526 21067 31578
rect 21067 31526 21113 31578
rect 20817 31524 20873 31526
rect 20897 31524 20953 31526
rect 20977 31524 21033 31526
rect 21057 31524 21113 31526
rect 20817 30490 20873 30492
rect 20897 30490 20953 30492
rect 20977 30490 21033 30492
rect 21057 30490 21113 30492
rect 20817 30438 20863 30490
rect 20863 30438 20873 30490
rect 20897 30438 20927 30490
rect 20927 30438 20939 30490
rect 20939 30438 20953 30490
rect 20977 30438 20991 30490
rect 20991 30438 21003 30490
rect 21003 30438 21033 30490
rect 21057 30438 21067 30490
rect 21067 30438 21113 30490
rect 20817 30436 20873 30438
rect 20897 30436 20953 30438
rect 20977 30436 21033 30438
rect 21057 30436 21113 30438
rect 20817 29402 20873 29404
rect 20897 29402 20953 29404
rect 20977 29402 21033 29404
rect 21057 29402 21113 29404
rect 20817 29350 20863 29402
rect 20863 29350 20873 29402
rect 20897 29350 20927 29402
rect 20927 29350 20939 29402
rect 20939 29350 20953 29402
rect 20977 29350 20991 29402
rect 20991 29350 21003 29402
rect 21003 29350 21033 29402
rect 21057 29350 21067 29402
rect 21067 29350 21113 29402
rect 20817 29348 20873 29350
rect 20897 29348 20953 29350
rect 20977 29348 21033 29350
rect 21057 29348 21113 29350
rect 20817 28314 20873 28316
rect 20897 28314 20953 28316
rect 20977 28314 21033 28316
rect 21057 28314 21113 28316
rect 20817 28262 20863 28314
rect 20863 28262 20873 28314
rect 20897 28262 20927 28314
rect 20927 28262 20939 28314
rect 20939 28262 20953 28314
rect 20977 28262 20991 28314
rect 20991 28262 21003 28314
rect 21003 28262 21033 28314
rect 21057 28262 21067 28314
rect 21067 28262 21113 28314
rect 20817 28260 20873 28262
rect 20897 28260 20953 28262
rect 20977 28260 21033 28262
rect 21057 28260 21113 28262
rect 20817 27226 20873 27228
rect 20897 27226 20953 27228
rect 20977 27226 21033 27228
rect 21057 27226 21113 27228
rect 20817 27174 20863 27226
rect 20863 27174 20873 27226
rect 20897 27174 20927 27226
rect 20927 27174 20939 27226
rect 20939 27174 20953 27226
rect 20977 27174 20991 27226
rect 20991 27174 21003 27226
rect 21003 27174 21033 27226
rect 21057 27174 21067 27226
rect 21067 27174 21113 27226
rect 20817 27172 20873 27174
rect 20897 27172 20953 27174
rect 20977 27172 21033 27174
rect 21057 27172 21113 27174
rect 20718 26288 20774 26344
rect 20534 25744 20590 25800
rect 20817 26138 20873 26140
rect 20897 26138 20953 26140
rect 20977 26138 21033 26140
rect 21057 26138 21113 26140
rect 20817 26086 20863 26138
rect 20863 26086 20873 26138
rect 20897 26086 20927 26138
rect 20927 26086 20939 26138
rect 20939 26086 20953 26138
rect 20977 26086 20991 26138
rect 20991 26086 21003 26138
rect 21003 26086 21033 26138
rect 21057 26086 21067 26138
rect 21067 26086 21113 26138
rect 20817 26084 20873 26086
rect 20897 26084 20953 26086
rect 20977 26084 21033 26086
rect 21057 26084 21113 26086
rect 20810 25900 20866 25936
rect 20810 25880 20812 25900
rect 20812 25880 20864 25900
rect 20864 25880 20866 25900
rect 20817 25050 20873 25052
rect 20897 25050 20953 25052
rect 20977 25050 21033 25052
rect 21057 25050 21113 25052
rect 20817 24998 20863 25050
rect 20863 24998 20873 25050
rect 20897 24998 20927 25050
rect 20927 24998 20939 25050
rect 20939 24998 20953 25050
rect 20977 24998 20991 25050
rect 20991 24998 21003 25050
rect 21003 24998 21033 25050
rect 21057 24998 21067 25050
rect 21067 24998 21113 25050
rect 20817 24996 20873 24998
rect 20897 24996 20953 24998
rect 20977 24996 21033 24998
rect 21057 24996 21113 24998
rect 20817 23962 20873 23964
rect 20897 23962 20953 23964
rect 20977 23962 21033 23964
rect 21057 23962 21113 23964
rect 20817 23910 20863 23962
rect 20863 23910 20873 23962
rect 20897 23910 20927 23962
rect 20927 23910 20939 23962
rect 20939 23910 20953 23962
rect 20977 23910 20991 23962
rect 20991 23910 21003 23962
rect 21003 23910 21033 23962
rect 21057 23910 21067 23962
rect 21067 23910 21113 23962
rect 20817 23908 20873 23910
rect 20897 23908 20953 23910
rect 20977 23908 21033 23910
rect 21057 23908 21113 23910
rect 20817 22874 20873 22876
rect 20897 22874 20953 22876
rect 20977 22874 21033 22876
rect 21057 22874 21113 22876
rect 20817 22822 20863 22874
rect 20863 22822 20873 22874
rect 20897 22822 20927 22874
rect 20927 22822 20939 22874
rect 20939 22822 20953 22874
rect 20977 22822 20991 22874
rect 20991 22822 21003 22874
rect 21003 22822 21033 22874
rect 21057 22822 21067 22874
rect 21067 22822 21113 22874
rect 20817 22820 20873 22822
rect 20897 22820 20953 22822
rect 20977 22820 21033 22822
rect 21057 22820 21113 22822
rect 20817 21786 20873 21788
rect 20897 21786 20953 21788
rect 20977 21786 21033 21788
rect 21057 21786 21113 21788
rect 20817 21734 20863 21786
rect 20863 21734 20873 21786
rect 20897 21734 20927 21786
rect 20927 21734 20939 21786
rect 20939 21734 20953 21786
rect 20977 21734 20991 21786
rect 20991 21734 21003 21786
rect 21003 21734 21033 21786
rect 21057 21734 21067 21786
rect 21067 21734 21113 21786
rect 20817 21732 20873 21734
rect 20897 21732 20953 21734
rect 20977 21732 21033 21734
rect 21057 21732 21113 21734
rect 20817 20698 20873 20700
rect 20897 20698 20953 20700
rect 20977 20698 21033 20700
rect 21057 20698 21113 20700
rect 20817 20646 20863 20698
rect 20863 20646 20873 20698
rect 20897 20646 20927 20698
rect 20927 20646 20939 20698
rect 20939 20646 20953 20698
rect 20977 20646 20991 20698
rect 20991 20646 21003 20698
rect 21003 20646 21033 20698
rect 21057 20646 21067 20698
rect 21067 20646 21113 20698
rect 20817 20644 20873 20646
rect 20897 20644 20953 20646
rect 20977 20644 21033 20646
rect 21057 20644 21113 20646
rect 20817 19610 20873 19612
rect 20897 19610 20953 19612
rect 20977 19610 21033 19612
rect 21057 19610 21113 19612
rect 20817 19558 20863 19610
rect 20863 19558 20873 19610
rect 20897 19558 20927 19610
rect 20927 19558 20939 19610
rect 20939 19558 20953 19610
rect 20977 19558 20991 19610
rect 20991 19558 21003 19610
rect 21003 19558 21033 19610
rect 21057 19558 21067 19610
rect 21067 19558 21113 19610
rect 20817 19556 20873 19558
rect 20897 19556 20953 19558
rect 20977 19556 21033 19558
rect 21057 19556 21113 19558
rect 20817 18522 20873 18524
rect 20897 18522 20953 18524
rect 20977 18522 21033 18524
rect 21057 18522 21113 18524
rect 20817 18470 20863 18522
rect 20863 18470 20873 18522
rect 20897 18470 20927 18522
rect 20927 18470 20939 18522
rect 20939 18470 20953 18522
rect 20977 18470 20991 18522
rect 20991 18470 21003 18522
rect 21003 18470 21033 18522
rect 21057 18470 21067 18522
rect 21067 18470 21113 18522
rect 20817 18468 20873 18470
rect 20897 18468 20953 18470
rect 20977 18468 21033 18470
rect 21057 18468 21113 18470
rect 20817 17434 20873 17436
rect 20897 17434 20953 17436
rect 20977 17434 21033 17436
rect 21057 17434 21113 17436
rect 20817 17382 20863 17434
rect 20863 17382 20873 17434
rect 20897 17382 20927 17434
rect 20927 17382 20939 17434
rect 20939 17382 20953 17434
rect 20977 17382 20991 17434
rect 20991 17382 21003 17434
rect 21003 17382 21033 17434
rect 21057 17382 21067 17434
rect 21067 17382 21113 17434
rect 20817 17380 20873 17382
rect 20897 17380 20953 17382
rect 20977 17380 21033 17382
rect 21057 17380 21113 17382
rect 20817 16346 20873 16348
rect 20897 16346 20953 16348
rect 20977 16346 21033 16348
rect 21057 16346 21113 16348
rect 20817 16294 20863 16346
rect 20863 16294 20873 16346
rect 20897 16294 20927 16346
rect 20927 16294 20939 16346
rect 20939 16294 20953 16346
rect 20977 16294 20991 16346
rect 20991 16294 21003 16346
rect 21003 16294 21033 16346
rect 21057 16294 21067 16346
rect 21067 16294 21113 16346
rect 20817 16292 20873 16294
rect 20897 16292 20953 16294
rect 20977 16292 21033 16294
rect 21057 16292 21113 16294
rect 20817 15258 20873 15260
rect 20897 15258 20953 15260
rect 20977 15258 21033 15260
rect 21057 15258 21113 15260
rect 20817 15206 20863 15258
rect 20863 15206 20873 15258
rect 20897 15206 20927 15258
rect 20927 15206 20939 15258
rect 20939 15206 20953 15258
rect 20977 15206 20991 15258
rect 20991 15206 21003 15258
rect 21003 15206 21033 15258
rect 21057 15206 21067 15258
rect 21067 15206 21113 15258
rect 20817 15204 20873 15206
rect 20897 15204 20953 15206
rect 20977 15204 21033 15206
rect 21057 15204 21113 15206
rect 30102 39380 30104 39400
rect 30104 39380 30156 39400
rect 30156 39380 30158 39400
rect 30102 39344 30158 39380
rect 25782 38650 25838 38652
rect 25862 38650 25918 38652
rect 25942 38650 25998 38652
rect 26022 38650 26078 38652
rect 25782 38598 25828 38650
rect 25828 38598 25838 38650
rect 25862 38598 25892 38650
rect 25892 38598 25904 38650
rect 25904 38598 25918 38650
rect 25942 38598 25956 38650
rect 25956 38598 25968 38650
rect 25968 38598 25998 38650
rect 26022 38598 26032 38650
rect 26032 38598 26078 38650
rect 25782 38596 25838 38598
rect 25862 38596 25918 38598
rect 25942 38596 25998 38598
rect 26022 38596 26078 38598
rect 30102 37848 30158 37904
rect 25782 37562 25838 37564
rect 25862 37562 25918 37564
rect 25942 37562 25998 37564
rect 26022 37562 26078 37564
rect 25782 37510 25828 37562
rect 25828 37510 25838 37562
rect 25862 37510 25892 37562
rect 25892 37510 25904 37562
rect 25904 37510 25918 37562
rect 25942 37510 25956 37562
rect 25956 37510 25968 37562
rect 25968 37510 25998 37562
rect 26022 37510 26032 37562
rect 26032 37510 26078 37562
rect 25782 37508 25838 37510
rect 25862 37508 25918 37510
rect 25942 37508 25998 37510
rect 26022 37508 26078 37510
rect 25782 36474 25838 36476
rect 25862 36474 25918 36476
rect 25942 36474 25998 36476
rect 26022 36474 26078 36476
rect 25782 36422 25828 36474
rect 25828 36422 25838 36474
rect 25862 36422 25892 36474
rect 25892 36422 25904 36474
rect 25904 36422 25918 36474
rect 25942 36422 25956 36474
rect 25956 36422 25968 36474
rect 25968 36422 25998 36474
rect 26022 36422 26032 36474
rect 26032 36422 26078 36474
rect 25782 36420 25838 36422
rect 25862 36420 25918 36422
rect 25942 36420 25998 36422
rect 26022 36420 26078 36422
rect 30102 36216 30158 36272
rect 25782 35386 25838 35388
rect 25862 35386 25918 35388
rect 25942 35386 25998 35388
rect 26022 35386 26078 35388
rect 25782 35334 25828 35386
rect 25828 35334 25838 35386
rect 25862 35334 25892 35386
rect 25892 35334 25904 35386
rect 25904 35334 25918 35386
rect 25942 35334 25956 35386
rect 25956 35334 25968 35386
rect 25968 35334 25998 35386
rect 26022 35334 26032 35386
rect 26032 35334 26078 35386
rect 25782 35332 25838 35334
rect 25862 35332 25918 35334
rect 25942 35332 25998 35334
rect 26022 35332 26078 35334
rect 30102 34720 30158 34776
rect 25782 34298 25838 34300
rect 25862 34298 25918 34300
rect 25942 34298 25998 34300
rect 26022 34298 26078 34300
rect 25782 34246 25828 34298
rect 25828 34246 25838 34298
rect 25862 34246 25892 34298
rect 25892 34246 25904 34298
rect 25904 34246 25918 34298
rect 25942 34246 25956 34298
rect 25956 34246 25968 34298
rect 25968 34246 25998 34298
rect 26022 34246 26032 34298
rect 26032 34246 26078 34298
rect 25782 34244 25838 34246
rect 25862 34244 25918 34246
rect 25942 34244 25998 34246
rect 26022 34244 26078 34246
rect 30010 33260 30012 33280
rect 30012 33260 30064 33280
rect 30064 33260 30066 33280
rect 30010 33224 30066 33260
rect 25782 33210 25838 33212
rect 25862 33210 25918 33212
rect 25942 33210 25998 33212
rect 26022 33210 26078 33212
rect 25782 33158 25828 33210
rect 25828 33158 25838 33210
rect 25862 33158 25892 33210
rect 25892 33158 25904 33210
rect 25904 33158 25918 33210
rect 25942 33158 25956 33210
rect 25956 33158 25968 33210
rect 25968 33158 25998 33210
rect 26022 33158 26032 33210
rect 26032 33158 26078 33210
rect 25782 33156 25838 33158
rect 25862 33156 25918 33158
rect 25942 33156 25998 33158
rect 26022 33156 26078 33158
rect 25782 32122 25838 32124
rect 25862 32122 25918 32124
rect 25942 32122 25998 32124
rect 26022 32122 26078 32124
rect 25782 32070 25828 32122
rect 25828 32070 25838 32122
rect 25862 32070 25892 32122
rect 25892 32070 25904 32122
rect 25904 32070 25918 32122
rect 25942 32070 25956 32122
rect 25956 32070 25968 32122
rect 25968 32070 25998 32122
rect 26022 32070 26032 32122
rect 26032 32070 26078 32122
rect 25782 32068 25838 32070
rect 25862 32068 25918 32070
rect 25942 32068 25998 32070
rect 26022 32068 26078 32070
rect 25782 31034 25838 31036
rect 25862 31034 25918 31036
rect 25942 31034 25998 31036
rect 26022 31034 26078 31036
rect 25782 30982 25828 31034
rect 25828 30982 25838 31034
rect 25862 30982 25892 31034
rect 25892 30982 25904 31034
rect 25904 30982 25918 31034
rect 25942 30982 25956 31034
rect 25956 30982 25968 31034
rect 25968 30982 25998 31034
rect 26022 30982 26032 31034
rect 26032 30982 26078 31034
rect 25782 30980 25838 30982
rect 25862 30980 25918 30982
rect 25942 30980 25998 30982
rect 26022 30980 26078 30982
rect 30010 31628 30012 31648
rect 30012 31628 30064 31648
rect 30064 31628 30066 31648
rect 30010 31592 30066 31628
rect 25782 29946 25838 29948
rect 25862 29946 25918 29948
rect 25942 29946 25998 29948
rect 26022 29946 26078 29948
rect 25782 29894 25828 29946
rect 25828 29894 25838 29946
rect 25862 29894 25892 29946
rect 25892 29894 25904 29946
rect 25904 29894 25918 29946
rect 25942 29894 25956 29946
rect 25956 29894 25968 29946
rect 25968 29894 25998 29946
rect 26022 29894 26032 29946
rect 26032 29894 26078 29946
rect 25782 29892 25838 29894
rect 25862 29892 25918 29894
rect 25942 29892 25998 29894
rect 26022 29892 26078 29894
rect 25782 28858 25838 28860
rect 25862 28858 25918 28860
rect 25942 28858 25998 28860
rect 26022 28858 26078 28860
rect 25782 28806 25828 28858
rect 25828 28806 25838 28858
rect 25862 28806 25892 28858
rect 25892 28806 25904 28858
rect 25904 28806 25918 28858
rect 25942 28806 25956 28858
rect 25956 28806 25968 28858
rect 25968 28806 25998 28858
rect 26022 28806 26032 28858
rect 26032 28806 26078 28858
rect 25782 28804 25838 28806
rect 25862 28804 25918 28806
rect 25942 28804 25998 28806
rect 26022 28804 26078 28806
rect 25782 27770 25838 27772
rect 25862 27770 25918 27772
rect 25942 27770 25998 27772
rect 26022 27770 26078 27772
rect 25782 27718 25828 27770
rect 25828 27718 25838 27770
rect 25862 27718 25892 27770
rect 25892 27718 25904 27770
rect 25904 27718 25918 27770
rect 25942 27718 25956 27770
rect 25956 27718 25968 27770
rect 25968 27718 25998 27770
rect 26022 27718 26032 27770
rect 26032 27718 26078 27770
rect 25782 27716 25838 27718
rect 25862 27716 25918 27718
rect 25942 27716 25998 27718
rect 26022 27716 26078 27718
rect 25782 26682 25838 26684
rect 25862 26682 25918 26684
rect 25942 26682 25998 26684
rect 26022 26682 26078 26684
rect 25782 26630 25828 26682
rect 25828 26630 25838 26682
rect 25862 26630 25892 26682
rect 25892 26630 25904 26682
rect 25904 26630 25918 26682
rect 25942 26630 25956 26682
rect 25956 26630 25968 26682
rect 25968 26630 25998 26682
rect 26022 26630 26032 26682
rect 26032 26630 26078 26682
rect 25782 26628 25838 26630
rect 25862 26628 25918 26630
rect 25942 26628 25998 26630
rect 26022 26628 26078 26630
rect 25782 25594 25838 25596
rect 25862 25594 25918 25596
rect 25942 25594 25998 25596
rect 26022 25594 26078 25596
rect 25782 25542 25828 25594
rect 25828 25542 25838 25594
rect 25862 25542 25892 25594
rect 25892 25542 25904 25594
rect 25904 25542 25918 25594
rect 25942 25542 25956 25594
rect 25956 25542 25968 25594
rect 25968 25542 25998 25594
rect 26022 25542 26032 25594
rect 26032 25542 26078 25594
rect 25782 25540 25838 25542
rect 25862 25540 25918 25542
rect 25942 25540 25998 25542
rect 26022 25540 26078 25542
rect 25782 24506 25838 24508
rect 25862 24506 25918 24508
rect 25942 24506 25998 24508
rect 26022 24506 26078 24508
rect 25782 24454 25828 24506
rect 25828 24454 25838 24506
rect 25862 24454 25892 24506
rect 25892 24454 25904 24506
rect 25904 24454 25918 24506
rect 25942 24454 25956 24506
rect 25956 24454 25968 24506
rect 25968 24454 25998 24506
rect 26022 24454 26032 24506
rect 26032 24454 26078 24506
rect 25782 24452 25838 24454
rect 25862 24452 25918 24454
rect 25942 24452 25998 24454
rect 26022 24452 26078 24454
rect 25782 23418 25838 23420
rect 25862 23418 25918 23420
rect 25942 23418 25998 23420
rect 26022 23418 26078 23420
rect 25782 23366 25828 23418
rect 25828 23366 25838 23418
rect 25862 23366 25892 23418
rect 25892 23366 25904 23418
rect 25904 23366 25918 23418
rect 25942 23366 25956 23418
rect 25956 23366 25968 23418
rect 25968 23366 25998 23418
rect 26022 23366 26032 23418
rect 26032 23366 26078 23418
rect 25782 23364 25838 23366
rect 25862 23364 25918 23366
rect 25942 23364 25998 23366
rect 26022 23364 26078 23366
rect 20817 14170 20873 14172
rect 20897 14170 20953 14172
rect 20977 14170 21033 14172
rect 21057 14170 21113 14172
rect 20817 14118 20863 14170
rect 20863 14118 20873 14170
rect 20897 14118 20927 14170
rect 20927 14118 20939 14170
rect 20939 14118 20953 14170
rect 20977 14118 20991 14170
rect 20991 14118 21003 14170
rect 21003 14118 21033 14170
rect 21057 14118 21067 14170
rect 21067 14118 21113 14170
rect 20817 14116 20873 14118
rect 20897 14116 20953 14118
rect 20977 14116 21033 14118
rect 21057 14116 21113 14118
rect 25782 22330 25838 22332
rect 25862 22330 25918 22332
rect 25942 22330 25998 22332
rect 26022 22330 26078 22332
rect 25782 22278 25828 22330
rect 25828 22278 25838 22330
rect 25862 22278 25892 22330
rect 25892 22278 25904 22330
rect 25904 22278 25918 22330
rect 25942 22278 25956 22330
rect 25956 22278 25968 22330
rect 25968 22278 25998 22330
rect 26022 22278 26032 22330
rect 26032 22278 26078 22330
rect 25782 22276 25838 22278
rect 25862 22276 25918 22278
rect 25942 22276 25998 22278
rect 26022 22276 26078 22278
rect 25782 21242 25838 21244
rect 25862 21242 25918 21244
rect 25942 21242 25998 21244
rect 26022 21242 26078 21244
rect 25782 21190 25828 21242
rect 25828 21190 25838 21242
rect 25862 21190 25892 21242
rect 25892 21190 25904 21242
rect 25904 21190 25918 21242
rect 25942 21190 25956 21242
rect 25956 21190 25968 21242
rect 25968 21190 25998 21242
rect 26022 21190 26032 21242
rect 26032 21190 26078 21242
rect 25782 21188 25838 21190
rect 25862 21188 25918 21190
rect 25942 21188 25998 21190
rect 26022 21188 26078 21190
rect 25782 20154 25838 20156
rect 25862 20154 25918 20156
rect 25942 20154 25998 20156
rect 26022 20154 26078 20156
rect 25782 20102 25828 20154
rect 25828 20102 25838 20154
rect 25862 20102 25892 20154
rect 25892 20102 25904 20154
rect 25904 20102 25918 20154
rect 25942 20102 25956 20154
rect 25956 20102 25968 20154
rect 25968 20102 25998 20154
rect 26022 20102 26032 20154
rect 26032 20102 26078 20154
rect 25782 20100 25838 20102
rect 25862 20100 25918 20102
rect 25942 20100 25998 20102
rect 26022 20100 26078 20102
rect 25782 19066 25838 19068
rect 25862 19066 25918 19068
rect 25942 19066 25998 19068
rect 26022 19066 26078 19068
rect 25782 19014 25828 19066
rect 25828 19014 25838 19066
rect 25862 19014 25892 19066
rect 25892 19014 25904 19066
rect 25904 19014 25918 19066
rect 25942 19014 25956 19066
rect 25956 19014 25968 19066
rect 25968 19014 25998 19066
rect 26022 19014 26032 19066
rect 26032 19014 26078 19066
rect 25782 19012 25838 19014
rect 25862 19012 25918 19014
rect 25942 19012 25998 19014
rect 26022 19012 26078 19014
rect 25782 17978 25838 17980
rect 25862 17978 25918 17980
rect 25942 17978 25998 17980
rect 26022 17978 26078 17980
rect 25782 17926 25828 17978
rect 25828 17926 25838 17978
rect 25862 17926 25892 17978
rect 25892 17926 25904 17978
rect 25904 17926 25918 17978
rect 25942 17926 25956 17978
rect 25956 17926 25968 17978
rect 25968 17926 25998 17978
rect 26022 17926 26032 17978
rect 26032 17926 26078 17978
rect 25782 17924 25838 17926
rect 25862 17924 25918 17926
rect 25942 17924 25998 17926
rect 26022 17924 26078 17926
rect 25782 16890 25838 16892
rect 25862 16890 25918 16892
rect 25942 16890 25998 16892
rect 26022 16890 26078 16892
rect 25782 16838 25828 16890
rect 25828 16838 25838 16890
rect 25862 16838 25892 16890
rect 25892 16838 25904 16890
rect 25904 16838 25918 16890
rect 25942 16838 25956 16890
rect 25956 16838 25968 16890
rect 25968 16838 25998 16890
rect 26022 16838 26032 16890
rect 26032 16838 26078 16890
rect 25782 16836 25838 16838
rect 25862 16836 25918 16838
rect 25942 16836 25998 16838
rect 26022 16836 26078 16838
rect 25782 15802 25838 15804
rect 25862 15802 25918 15804
rect 25942 15802 25998 15804
rect 26022 15802 26078 15804
rect 25782 15750 25828 15802
rect 25828 15750 25838 15802
rect 25862 15750 25892 15802
rect 25892 15750 25904 15802
rect 25904 15750 25918 15802
rect 25942 15750 25956 15802
rect 25956 15750 25968 15802
rect 25968 15750 25998 15802
rect 26022 15750 26032 15802
rect 26032 15750 26078 15802
rect 25782 15748 25838 15750
rect 25862 15748 25918 15750
rect 25942 15748 25998 15750
rect 26022 15748 26078 15750
rect 20817 13082 20873 13084
rect 20897 13082 20953 13084
rect 20977 13082 21033 13084
rect 21057 13082 21113 13084
rect 20817 13030 20863 13082
rect 20863 13030 20873 13082
rect 20897 13030 20927 13082
rect 20927 13030 20939 13082
rect 20939 13030 20953 13082
rect 20977 13030 20991 13082
rect 20991 13030 21003 13082
rect 21003 13030 21033 13082
rect 21057 13030 21067 13082
rect 21067 13030 21113 13082
rect 20817 13028 20873 13030
rect 20897 13028 20953 13030
rect 20977 13028 21033 13030
rect 21057 13028 21113 13030
rect 20817 11994 20873 11996
rect 20897 11994 20953 11996
rect 20977 11994 21033 11996
rect 21057 11994 21113 11996
rect 20817 11942 20863 11994
rect 20863 11942 20873 11994
rect 20897 11942 20927 11994
rect 20927 11942 20939 11994
rect 20939 11942 20953 11994
rect 20977 11942 20991 11994
rect 20991 11942 21003 11994
rect 21003 11942 21033 11994
rect 21057 11942 21067 11994
rect 21067 11942 21113 11994
rect 20817 11940 20873 11942
rect 20897 11940 20953 11942
rect 20977 11940 21033 11942
rect 21057 11940 21113 11942
rect 25782 14714 25838 14716
rect 25862 14714 25918 14716
rect 25942 14714 25998 14716
rect 26022 14714 26078 14716
rect 25782 14662 25828 14714
rect 25828 14662 25838 14714
rect 25862 14662 25892 14714
rect 25892 14662 25904 14714
rect 25904 14662 25918 14714
rect 25942 14662 25956 14714
rect 25956 14662 25968 14714
rect 25968 14662 25998 14714
rect 26022 14662 26032 14714
rect 26032 14662 26078 14714
rect 25782 14660 25838 14662
rect 25862 14660 25918 14662
rect 25942 14660 25998 14662
rect 26022 14660 26078 14662
rect 25782 13626 25838 13628
rect 25862 13626 25918 13628
rect 25942 13626 25998 13628
rect 26022 13626 26078 13628
rect 25782 13574 25828 13626
rect 25828 13574 25838 13626
rect 25862 13574 25892 13626
rect 25892 13574 25904 13626
rect 25904 13574 25918 13626
rect 25942 13574 25956 13626
rect 25956 13574 25968 13626
rect 25968 13574 25998 13626
rect 26022 13574 26032 13626
rect 26032 13574 26078 13626
rect 25782 13572 25838 13574
rect 25862 13572 25918 13574
rect 25942 13572 25998 13574
rect 26022 13572 26078 13574
rect 25782 12538 25838 12540
rect 25862 12538 25918 12540
rect 25942 12538 25998 12540
rect 26022 12538 26078 12540
rect 25782 12486 25828 12538
rect 25828 12486 25838 12538
rect 25862 12486 25892 12538
rect 25892 12486 25904 12538
rect 25904 12486 25918 12538
rect 25942 12486 25956 12538
rect 25956 12486 25968 12538
rect 25968 12486 25998 12538
rect 26022 12486 26032 12538
rect 26032 12486 26078 12538
rect 25782 12484 25838 12486
rect 25862 12484 25918 12486
rect 25942 12484 25998 12486
rect 26022 12484 26078 12486
rect 20817 10906 20873 10908
rect 20897 10906 20953 10908
rect 20977 10906 21033 10908
rect 21057 10906 21113 10908
rect 20817 10854 20863 10906
rect 20863 10854 20873 10906
rect 20897 10854 20927 10906
rect 20927 10854 20939 10906
rect 20939 10854 20953 10906
rect 20977 10854 20991 10906
rect 20991 10854 21003 10906
rect 21003 10854 21033 10906
rect 21057 10854 21067 10906
rect 21067 10854 21113 10906
rect 20817 10852 20873 10854
rect 20897 10852 20953 10854
rect 20977 10852 21033 10854
rect 21057 10852 21113 10854
rect 20817 9818 20873 9820
rect 20897 9818 20953 9820
rect 20977 9818 21033 9820
rect 21057 9818 21113 9820
rect 20817 9766 20863 9818
rect 20863 9766 20873 9818
rect 20897 9766 20927 9818
rect 20927 9766 20939 9818
rect 20939 9766 20953 9818
rect 20977 9766 20991 9818
rect 20991 9766 21003 9818
rect 21003 9766 21033 9818
rect 21057 9766 21067 9818
rect 21067 9766 21113 9818
rect 20817 9764 20873 9766
rect 20897 9764 20953 9766
rect 20977 9764 21033 9766
rect 21057 9764 21113 9766
rect 20817 8730 20873 8732
rect 20897 8730 20953 8732
rect 20977 8730 21033 8732
rect 21057 8730 21113 8732
rect 20817 8678 20863 8730
rect 20863 8678 20873 8730
rect 20897 8678 20927 8730
rect 20927 8678 20939 8730
rect 20939 8678 20953 8730
rect 20977 8678 20991 8730
rect 20991 8678 21003 8730
rect 21003 8678 21033 8730
rect 21057 8678 21067 8730
rect 21067 8678 21113 8730
rect 20817 8676 20873 8678
rect 20897 8676 20953 8678
rect 20977 8676 21033 8678
rect 21057 8676 21113 8678
rect 20817 7642 20873 7644
rect 20897 7642 20953 7644
rect 20977 7642 21033 7644
rect 21057 7642 21113 7644
rect 20817 7590 20863 7642
rect 20863 7590 20873 7642
rect 20897 7590 20927 7642
rect 20927 7590 20939 7642
rect 20939 7590 20953 7642
rect 20977 7590 20991 7642
rect 20991 7590 21003 7642
rect 21003 7590 21033 7642
rect 21057 7590 21067 7642
rect 21067 7590 21113 7642
rect 20817 7588 20873 7590
rect 20897 7588 20953 7590
rect 20977 7588 21033 7590
rect 21057 7588 21113 7590
rect 20817 6554 20873 6556
rect 20897 6554 20953 6556
rect 20977 6554 21033 6556
rect 21057 6554 21113 6556
rect 20817 6502 20863 6554
rect 20863 6502 20873 6554
rect 20897 6502 20927 6554
rect 20927 6502 20939 6554
rect 20939 6502 20953 6554
rect 20977 6502 20991 6554
rect 20991 6502 21003 6554
rect 21003 6502 21033 6554
rect 21057 6502 21067 6554
rect 21067 6502 21113 6554
rect 20817 6500 20873 6502
rect 20897 6500 20953 6502
rect 20977 6500 21033 6502
rect 21057 6500 21113 6502
rect 20817 5466 20873 5468
rect 20897 5466 20953 5468
rect 20977 5466 21033 5468
rect 21057 5466 21113 5468
rect 20817 5414 20863 5466
rect 20863 5414 20873 5466
rect 20897 5414 20927 5466
rect 20927 5414 20939 5466
rect 20939 5414 20953 5466
rect 20977 5414 20991 5466
rect 20991 5414 21003 5466
rect 21003 5414 21033 5466
rect 21057 5414 21067 5466
rect 21067 5414 21113 5466
rect 20817 5412 20873 5414
rect 20897 5412 20953 5414
rect 20977 5412 21033 5414
rect 21057 5412 21113 5414
rect 20817 4378 20873 4380
rect 20897 4378 20953 4380
rect 20977 4378 21033 4380
rect 21057 4378 21113 4380
rect 20817 4326 20863 4378
rect 20863 4326 20873 4378
rect 20897 4326 20927 4378
rect 20927 4326 20939 4378
rect 20939 4326 20953 4378
rect 20977 4326 20991 4378
rect 20991 4326 21003 4378
rect 21003 4326 21033 4378
rect 21057 4326 21067 4378
rect 21067 4326 21113 4378
rect 20817 4324 20873 4326
rect 20897 4324 20953 4326
rect 20977 4324 21033 4326
rect 21057 4324 21113 4326
rect 20166 3052 20222 3088
rect 20166 3032 20168 3052
rect 20168 3032 20220 3052
rect 20220 3032 20222 3052
rect 20817 3290 20873 3292
rect 20897 3290 20953 3292
rect 20977 3290 21033 3292
rect 21057 3290 21113 3292
rect 20817 3238 20863 3290
rect 20863 3238 20873 3290
rect 20897 3238 20927 3290
rect 20927 3238 20939 3290
rect 20939 3238 20953 3290
rect 20977 3238 20991 3290
rect 20991 3238 21003 3290
rect 21003 3238 21033 3290
rect 21057 3238 21067 3290
rect 21067 3238 21113 3290
rect 20817 3236 20873 3238
rect 20897 3236 20953 3238
rect 20977 3236 21033 3238
rect 21057 3236 21113 3238
rect 20817 2202 20873 2204
rect 20897 2202 20953 2204
rect 20977 2202 21033 2204
rect 21057 2202 21113 2204
rect 20817 2150 20863 2202
rect 20863 2150 20873 2202
rect 20897 2150 20927 2202
rect 20927 2150 20939 2202
rect 20939 2150 20953 2202
rect 20977 2150 20991 2202
rect 20991 2150 21003 2202
rect 21003 2150 21033 2202
rect 21057 2150 21067 2202
rect 21067 2150 21113 2202
rect 20817 2148 20873 2150
rect 20897 2148 20953 2150
rect 20977 2148 21033 2150
rect 21057 2148 21113 2150
rect 25782 11450 25838 11452
rect 25862 11450 25918 11452
rect 25942 11450 25998 11452
rect 26022 11450 26078 11452
rect 25782 11398 25828 11450
rect 25828 11398 25838 11450
rect 25862 11398 25892 11450
rect 25892 11398 25904 11450
rect 25904 11398 25918 11450
rect 25942 11398 25956 11450
rect 25956 11398 25968 11450
rect 25968 11398 25998 11450
rect 26022 11398 26032 11450
rect 26032 11398 26078 11450
rect 25782 11396 25838 11398
rect 25862 11396 25918 11398
rect 25942 11396 25998 11398
rect 26022 11396 26078 11398
rect 25782 10362 25838 10364
rect 25862 10362 25918 10364
rect 25942 10362 25998 10364
rect 26022 10362 26078 10364
rect 25782 10310 25828 10362
rect 25828 10310 25838 10362
rect 25862 10310 25892 10362
rect 25892 10310 25904 10362
rect 25904 10310 25918 10362
rect 25942 10310 25956 10362
rect 25956 10310 25968 10362
rect 25968 10310 25998 10362
rect 26022 10310 26032 10362
rect 26032 10310 26078 10362
rect 25782 10308 25838 10310
rect 25862 10308 25918 10310
rect 25942 10308 25998 10310
rect 26022 10308 26078 10310
rect 25782 9274 25838 9276
rect 25862 9274 25918 9276
rect 25942 9274 25998 9276
rect 26022 9274 26078 9276
rect 25782 9222 25828 9274
rect 25828 9222 25838 9274
rect 25862 9222 25892 9274
rect 25892 9222 25904 9274
rect 25904 9222 25918 9274
rect 25942 9222 25956 9274
rect 25956 9222 25968 9274
rect 25968 9222 25998 9274
rect 26022 9222 26032 9274
rect 26032 9222 26078 9274
rect 25782 9220 25838 9222
rect 25862 9220 25918 9222
rect 25942 9220 25998 9222
rect 26022 9220 26078 9222
rect 25782 8186 25838 8188
rect 25862 8186 25918 8188
rect 25942 8186 25998 8188
rect 26022 8186 26078 8188
rect 25782 8134 25828 8186
rect 25828 8134 25838 8186
rect 25862 8134 25892 8186
rect 25892 8134 25904 8186
rect 25904 8134 25918 8186
rect 25942 8134 25956 8186
rect 25956 8134 25968 8186
rect 25968 8134 25998 8186
rect 26022 8134 26032 8186
rect 26032 8134 26078 8186
rect 25782 8132 25838 8134
rect 25862 8132 25918 8134
rect 25942 8132 25998 8134
rect 26022 8132 26078 8134
rect 25782 7098 25838 7100
rect 25862 7098 25918 7100
rect 25942 7098 25998 7100
rect 26022 7098 26078 7100
rect 25782 7046 25828 7098
rect 25828 7046 25838 7098
rect 25862 7046 25892 7098
rect 25892 7046 25904 7098
rect 25904 7046 25918 7098
rect 25942 7046 25956 7098
rect 25956 7046 25968 7098
rect 25968 7046 25998 7098
rect 26022 7046 26032 7098
rect 26032 7046 26078 7098
rect 25782 7044 25838 7046
rect 25862 7044 25918 7046
rect 25942 7044 25998 7046
rect 26022 7044 26078 7046
rect 25782 6010 25838 6012
rect 25862 6010 25918 6012
rect 25942 6010 25998 6012
rect 26022 6010 26078 6012
rect 25782 5958 25828 6010
rect 25828 5958 25838 6010
rect 25862 5958 25892 6010
rect 25892 5958 25904 6010
rect 25904 5958 25918 6010
rect 25942 5958 25956 6010
rect 25956 5958 25968 6010
rect 25968 5958 25998 6010
rect 26022 5958 26032 6010
rect 26032 5958 26078 6010
rect 25782 5956 25838 5958
rect 25862 5956 25918 5958
rect 25942 5956 25998 5958
rect 26022 5956 26078 5958
rect 25782 4922 25838 4924
rect 25862 4922 25918 4924
rect 25942 4922 25998 4924
rect 26022 4922 26078 4924
rect 25782 4870 25828 4922
rect 25828 4870 25838 4922
rect 25862 4870 25892 4922
rect 25892 4870 25904 4922
rect 25904 4870 25918 4922
rect 25942 4870 25956 4922
rect 25956 4870 25968 4922
rect 25968 4870 25998 4922
rect 26022 4870 26032 4922
rect 26032 4870 26078 4922
rect 25782 4868 25838 4870
rect 25862 4868 25918 4870
rect 25942 4868 25998 4870
rect 26022 4868 26078 4870
rect 25782 3834 25838 3836
rect 25862 3834 25918 3836
rect 25942 3834 25998 3836
rect 26022 3834 26078 3836
rect 25782 3782 25828 3834
rect 25828 3782 25838 3834
rect 25862 3782 25892 3834
rect 25892 3782 25904 3834
rect 25904 3782 25918 3834
rect 25942 3782 25956 3834
rect 25956 3782 25968 3834
rect 25968 3782 25998 3834
rect 26022 3782 26032 3834
rect 26032 3782 26078 3834
rect 25782 3780 25838 3782
rect 25862 3780 25918 3782
rect 25942 3780 25998 3782
rect 26022 3780 26078 3782
rect 22926 3032 22982 3088
rect 25782 2746 25838 2748
rect 25862 2746 25918 2748
rect 25942 2746 25998 2748
rect 26022 2746 26078 2748
rect 25782 2694 25828 2746
rect 25828 2694 25838 2746
rect 25862 2694 25892 2746
rect 25892 2694 25904 2746
rect 25904 2694 25918 2746
rect 25942 2694 25956 2746
rect 25956 2694 25968 2746
rect 25968 2694 25998 2746
rect 26022 2694 26032 2746
rect 26032 2694 26078 2746
rect 25782 2692 25838 2694
rect 25862 2692 25918 2694
rect 25942 2692 25998 2694
rect 26022 2692 26078 2694
rect 30010 30116 30066 30152
rect 30010 30096 30012 30116
rect 30012 30096 30064 30116
rect 30064 30096 30066 30116
rect 30010 28464 30066 28520
rect 30010 26968 30066 27024
rect 30010 25472 30066 25528
rect 30010 23840 30066 23896
rect 30010 22380 30012 22400
rect 30012 22380 30064 22400
rect 30064 22380 30066 22400
rect 30010 22344 30066 22380
rect 30010 20848 30066 20904
rect 30010 19216 30066 19272
rect 30010 17720 30066 17776
rect 30010 16088 30066 16144
rect 30010 14592 30066 14648
rect 30010 13132 30012 13152
rect 30012 13132 30064 13152
rect 30064 13132 30066 13152
rect 30010 13096 30066 13132
rect 30010 11500 30012 11520
rect 30012 11500 30064 11520
rect 30064 11500 30066 11520
rect 30010 11464 30066 11500
rect 30010 9968 30066 10024
rect 30010 8356 30066 8392
rect 30010 8336 30012 8356
rect 30012 8336 30064 8356
rect 30064 8336 30066 8356
rect 30010 6840 30066 6896
rect 30010 5364 30066 5400
rect 30010 5344 30012 5364
rect 30012 5344 30064 5364
rect 30064 5344 30066 5364
rect 30010 3712 30066 3768
rect 30010 2252 30012 2272
rect 30012 2252 30064 2272
rect 30064 2252 30066 2272
rect 30010 2216 30066 2252
rect 28906 720 28962 776
<< metal3 >>
rect 0 47562 800 47592
rect 2773 47562 2839 47565
rect 0 47560 2839 47562
rect 0 47504 2778 47560
rect 2834 47504 2839 47560
rect 0 47502 2839 47504
rect 0 47472 800 47502
rect 2773 47499 2839 47502
rect 30189 47154 30255 47157
rect 31200 47154 32000 47184
rect 30189 47152 32000 47154
rect 30189 47096 30194 47152
rect 30250 47096 32000 47152
rect 30189 47094 32000 47096
rect 30189 47091 30255 47094
rect 31200 47064 32000 47094
rect 0 46882 800 46912
rect 2865 46882 2931 46885
rect 0 46880 2931 46882
rect 0 46824 2870 46880
rect 2926 46824 2931 46880
rect 0 46822 2931 46824
rect 0 46792 800 46822
rect 2865 46819 2931 46822
rect 0 46066 800 46096
rect 2957 46066 3023 46069
rect 0 46064 3023 46066
rect 0 46008 2962 46064
rect 3018 46008 3023 46064
rect 0 46006 3023 46008
rect 0 45976 800 46006
rect 2957 46003 3023 46006
rect 10874 45728 11194 45729
rect 10874 45664 10882 45728
rect 10946 45664 10962 45728
rect 11026 45664 11042 45728
rect 11106 45664 11122 45728
rect 11186 45664 11194 45728
rect 10874 45663 11194 45664
rect 20805 45728 21125 45729
rect 20805 45664 20813 45728
rect 20877 45664 20893 45728
rect 20957 45664 20973 45728
rect 21037 45664 21053 45728
rect 21117 45664 21125 45728
rect 20805 45663 21125 45664
rect 30097 45658 30163 45661
rect 31200 45658 32000 45688
rect 30097 45656 32000 45658
rect 30097 45600 30102 45656
rect 30158 45600 32000 45656
rect 30097 45598 32000 45600
rect 30097 45595 30163 45598
rect 31200 45568 32000 45598
rect 0 45386 800 45416
rect 2221 45386 2287 45389
rect 0 45384 2287 45386
rect 0 45328 2226 45384
rect 2282 45328 2287 45384
rect 0 45326 2287 45328
rect 0 45296 800 45326
rect 2221 45323 2287 45326
rect 5909 45184 6229 45185
rect 5909 45120 5917 45184
rect 5981 45120 5997 45184
rect 6061 45120 6077 45184
rect 6141 45120 6157 45184
rect 6221 45120 6229 45184
rect 5909 45119 6229 45120
rect 15840 45184 16160 45185
rect 15840 45120 15848 45184
rect 15912 45120 15928 45184
rect 15992 45120 16008 45184
rect 16072 45120 16088 45184
rect 16152 45120 16160 45184
rect 15840 45119 16160 45120
rect 25770 45184 26090 45185
rect 25770 45120 25778 45184
rect 25842 45120 25858 45184
rect 25922 45120 25938 45184
rect 26002 45120 26018 45184
rect 26082 45120 26090 45184
rect 25770 45119 26090 45120
rect 10874 44640 11194 44641
rect 0 44570 800 44600
rect 10874 44576 10882 44640
rect 10946 44576 10962 44640
rect 11026 44576 11042 44640
rect 11106 44576 11122 44640
rect 11186 44576 11194 44640
rect 10874 44575 11194 44576
rect 20805 44640 21125 44641
rect 20805 44576 20813 44640
rect 20877 44576 20893 44640
rect 20957 44576 20973 44640
rect 21037 44576 21053 44640
rect 21117 44576 21125 44640
rect 20805 44575 21125 44576
rect 1485 44570 1551 44573
rect 0 44568 1551 44570
rect 0 44512 1490 44568
rect 1546 44512 1551 44568
rect 0 44510 1551 44512
rect 0 44480 800 44510
rect 1485 44507 1551 44510
rect 5909 44096 6229 44097
rect 5909 44032 5917 44096
rect 5981 44032 5997 44096
rect 6061 44032 6077 44096
rect 6141 44032 6157 44096
rect 6221 44032 6229 44096
rect 5909 44031 6229 44032
rect 15840 44096 16160 44097
rect 15840 44032 15848 44096
rect 15912 44032 15928 44096
rect 15992 44032 16008 44096
rect 16072 44032 16088 44096
rect 16152 44032 16160 44096
rect 15840 44031 16160 44032
rect 25770 44096 26090 44097
rect 25770 44032 25778 44096
rect 25842 44032 25858 44096
rect 25922 44032 25938 44096
rect 26002 44032 26018 44096
rect 26082 44032 26090 44096
rect 25770 44031 26090 44032
rect 30097 44026 30163 44029
rect 31200 44026 32000 44056
rect 30097 44024 32000 44026
rect 30097 43968 30102 44024
rect 30158 43968 32000 44024
rect 30097 43966 32000 43968
rect 30097 43963 30163 43966
rect 31200 43936 32000 43966
rect 0 43890 800 43920
rect 1485 43890 1551 43893
rect 0 43888 1551 43890
rect 0 43832 1490 43888
rect 1546 43832 1551 43888
rect 0 43830 1551 43832
rect 0 43800 800 43830
rect 1485 43827 1551 43830
rect 10874 43552 11194 43553
rect 10874 43488 10882 43552
rect 10946 43488 10962 43552
rect 11026 43488 11042 43552
rect 11106 43488 11122 43552
rect 11186 43488 11194 43552
rect 10874 43487 11194 43488
rect 20805 43552 21125 43553
rect 20805 43488 20813 43552
rect 20877 43488 20893 43552
rect 20957 43488 20973 43552
rect 21037 43488 21053 43552
rect 21117 43488 21125 43552
rect 20805 43487 21125 43488
rect 0 43074 800 43104
rect 1485 43074 1551 43077
rect 0 43072 1551 43074
rect 0 43016 1490 43072
rect 1546 43016 1551 43072
rect 0 43014 1551 43016
rect 0 42984 800 43014
rect 1485 43011 1551 43014
rect 5909 43008 6229 43009
rect 5909 42944 5917 43008
rect 5981 42944 5997 43008
rect 6061 42944 6077 43008
rect 6141 42944 6157 43008
rect 6221 42944 6229 43008
rect 5909 42943 6229 42944
rect 15840 43008 16160 43009
rect 15840 42944 15848 43008
rect 15912 42944 15928 43008
rect 15992 42944 16008 43008
rect 16072 42944 16088 43008
rect 16152 42944 16160 43008
rect 15840 42943 16160 42944
rect 25770 43008 26090 43009
rect 25770 42944 25778 43008
rect 25842 42944 25858 43008
rect 25922 42944 25938 43008
rect 26002 42944 26018 43008
rect 26082 42944 26090 43008
rect 25770 42943 26090 42944
rect 30097 42530 30163 42533
rect 31200 42530 32000 42560
rect 30097 42528 32000 42530
rect 30097 42472 30102 42528
rect 30158 42472 32000 42528
rect 30097 42470 32000 42472
rect 30097 42467 30163 42470
rect 10874 42464 11194 42465
rect 0 42394 800 42424
rect 10874 42400 10882 42464
rect 10946 42400 10962 42464
rect 11026 42400 11042 42464
rect 11106 42400 11122 42464
rect 11186 42400 11194 42464
rect 10874 42399 11194 42400
rect 20805 42464 21125 42465
rect 20805 42400 20813 42464
rect 20877 42400 20893 42464
rect 20957 42400 20973 42464
rect 21037 42400 21053 42464
rect 21117 42400 21125 42464
rect 31200 42440 32000 42470
rect 20805 42399 21125 42400
rect 1485 42394 1551 42397
rect 0 42392 1551 42394
rect 0 42336 1490 42392
rect 1546 42336 1551 42392
rect 0 42334 1551 42336
rect 0 42304 800 42334
rect 1485 42331 1551 42334
rect 5909 41920 6229 41921
rect 5909 41856 5917 41920
rect 5981 41856 5997 41920
rect 6061 41856 6077 41920
rect 6141 41856 6157 41920
rect 6221 41856 6229 41920
rect 5909 41855 6229 41856
rect 15840 41920 16160 41921
rect 15840 41856 15848 41920
rect 15912 41856 15928 41920
rect 15992 41856 16008 41920
rect 16072 41856 16088 41920
rect 16152 41856 16160 41920
rect 15840 41855 16160 41856
rect 25770 41920 26090 41921
rect 25770 41856 25778 41920
rect 25842 41856 25858 41920
rect 25922 41856 25938 41920
rect 26002 41856 26018 41920
rect 26082 41856 26090 41920
rect 25770 41855 26090 41856
rect 0 41714 800 41744
rect 1485 41714 1551 41717
rect 0 41712 1551 41714
rect 0 41656 1490 41712
rect 1546 41656 1551 41712
rect 0 41654 1551 41656
rect 0 41624 800 41654
rect 1485 41651 1551 41654
rect 10874 41376 11194 41377
rect 10874 41312 10882 41376
rect 10946 41312 10962 41376
rect 11026 41312 11042 41376
rect 11106 41312 11122 41376
rect 11186 41312 11194 41376
rect 10874 41311 11194 41312
rect 20805 41376 21125 41377
rect 20805 41312 20813 41376
rect 20877 41312 20893 41376
rect 20957 41312 20973 41376
rect 21037 41312 21053 41376
rect 21117 41312 21125 41376
rect 20805 41311 21125 41312
rect 30097 41034 30163 41037
rect 31200 41034 32000 41064
rect 30097 41032 32000 41034
rect 30097 40976 30102 41032
rect 30158 40976 32000 41032
rect 30097 40974 32000 40976
rect 30097 40971 30163 40974
rect 31200 40944 32000 40974
rect 0 40898 800 40928
rect 1485 40898 1551 40901
rect 0 40896 1551 40898
rect 0 40840 1490 40896
rect 1546 40840 1551 40896
rect 0 40838 1551 40840
rect 0 40808 800 40838
rect 1485 40835 1551 40838
rect 5909 40832 6229 40833
rect 5909 40768 5917 40832
rect 5981 40768 5997 40832
rect 6061 40768 6077 40832
rect 6141 40768 6157 40832
rect 6221 40768 6229 40832
rect 5909 40767 6229 40768
rect 15840 40832 16160 40833
rect 15840 40768 15848 40832
rect 15912 40768 15928 40832
rect 15992 40768 16008 40832
rect 16072 40768 16088 40832
rect 16152 40768 16160 40832
rect 15840 40767 16160 40768
rect 25770 40832 26090 40833
rect 25770 40768 25778 40832
rect 25842 40768 25858 40832
rect 25922 40768 25938 40832
rect 26002 40768 26018 40832
rect 26082 40768 26090 40832
rect 25770 40767 26090 40768
rect 10874 40288 11194 40289
rect 0 40218 800 40248
rect 10874 40224 10882 40288
rect 10946 40224 10962 40288
rect 11026 40224 11042 40288
rect 11106 40224 11122 40288
rect 11186 40224 11194 40288
rect 10874 40223 11194 40224
rect 20805 40288 21125 40289
rect 20805 40224 20813 40288
rect 20877 40224 20893 40288
rect 20957 40224 20973 40288
rect 21037 40224 21053 40288
rect 21117 40224 21125 40288
rect 20805 40223 21125 40224
rect 1485 40218 1551 40221
rect 0 40216 1551 40218
rect 0 40160 1490 40216
rect 1546 40160 1551 40216
rect 0 40158 1551 40160
rect 0 40128 800 40158
rect 1485 40155 1551 40158
rect 5909 39744 6229 39745
rect 5909 39680 5917 39744
rect 5981 39680 5997 39744
rect 6061 39680 6077 39744
rect 6141 39680 6157 39744
rect 6221 39680 6229 39744
rect 5909 39679 6229 39680
rect 15840 39744 16160 39745
rect 15840 39680 15848 39744
rect 15912 39680 15928 39744
rect 15992 39680 16008 39744
rect 16072 39680 16088 39744
rect 16152 39680 16160 39744
rect 15840 39679 16160 39680
rect 25770 39744 26090 39745
rect 25770 39680 25778 39744
rect 25842 39680 25858 39744
rect 25922 39680 25938 39744
rect 26002 39680 26018 39744
rect 26082 39680 26090 39744
rect 25770 39679 26090 39680
rect 0 39402 800 39432
rect 2221 39402 2287 39405
rect 0 39400 2287 39402
rect 0 39344 2226 39400
rect 2282 39344 2287 39400
rect 0 39342 2287 39344
rect 0 39312 800 39342
rect 2221 39339 2287 39342
rect 30097 39402 30163 39405
rect 31200 39402 32000 39432
rect 30097 39400 32000 39402
rect 30097 39344 30102 39400
rect 30158 39344 32000 39400
rect 30097 39342 32000 39344
rect 30097 39339 30163 39342
rect 31200 39312 32000 39342
rect 10874 39200 11194 39201
rect 10874 39136 10882 39200
rect 10946 39136 10962 39200
rect 11026 39136 11042 39200
rect 11106 39136 11122 39200
rect 11186 39136 11194 39200
rect 10874 39135 11194 39136
rect 20805 39200 21125 39201
rect 20805 39136 20813 39200
rect 20877 39136 20893 39200
rect 20957 39136 20973 39200
rect 21037 39136 21053 39200
rect 21117 39136 21125 39200
rect 20805 39135 21125 39136
rect 0 38722 800 38752
rect 3049 38722 3115 38725
rect 0 38720 3115 38722
rect 0 38664 3054 38720
rect 3110 38664 3115 38720
rect 0 38662 3115 38664
rect 0 38632 800 38662
rect 3049 38659 3115 38662
rect 5909 38656 6229 38657
rect 5909 38592 5917 38656
rect 5981 38592 5997 38656
rect 6061 38592 6077 38656
rect 6141 38592 6157 38656
rect 6221 38592 6229 38656
rect 5909 38591 6229 38592
rect 15840 38656 16160 38657
rect 15840 38592 15848 38656
rect 15912 38592 15928 38656
rect 15992 38592 16008 38656
rect 16072 38592 16088 38656
rect 16152 38592 16160 38656
rect 15840 38591 16160 38592
rect 25770 38656 26090 38657
rect 25770 38592 25778 38656
rect 25842 38592 25858 38656
rect 25922 38592 25938 38656
rect 26002 38592 26018 38656
rect 26082 38592 26090 38656
rect 25770 38591 26090 38592
rect 10874 38112 11194 38113
rect 10874 38048 10882 38112
rect 10946 38048 10962 38112
rect 11026 38048 11042 38112
rect 11106 38048 11122 38112
rect 11186 38048 11194 38112
rect 10874 38047 11194 38048
rect 20805 38112 21125 38113
rect 20805 38048 20813 38112
rect 20877 38048 20893 38112
rect 20957 38048 20973 38112
rect 21037 38048 21053 38112
rect 21117 38048 21125 38112
rect 20805 38047 21125 38048
rect 0 37906 800 37936
rect 1485 37906 1551 37909
rect 0 37904 1551 37906
rect 0 37848 1490 37904
rect 1546 37848 1551 37904
rect 0 37846 1551 37848
rect 0 37816 800 37846
rect 1485 37843 1551 37846
rect 30097 37906 30163 37909
rect 31200 37906 32000 37936
rect 30097 37904 32000 37906
rect 30097 37848 30102 37904
rect 30158 37848 32000 37904
rect 30097 37846 32000 37848
rect 30097 37843 30163 37846
rect 31200 37816 32000 37846
rect 5909 37568 6229 37569
rect 5909 37504 5917 37568
rect 5981 37504 5997 37568
rect 6061 37504 6077 37568
rect 6141 37504 6157 37568
rect 6221 37504 6229 37568
rect 5909 37503 6229 37504
rect 15840 37568 16160 37569
rect 15840 37504 15848 37568
rect 15912 37504 15928 37568
rect 15992 37504 16008 37568
rect 16072 37504 16088 37568
rect 16152 37504 16160 37568
rect 15840 37503 16160 37504
rect 25770 37568 26090 37569
rect 25770 37504 25778 37568
rect 25842 37504 25858 37568
rect 25922 37504 25938 37568
rect 26002 37504 26018 37568
rect 26082 37504 26090 37568
rect 25770 37503 26090 37504
rect 0 37226 800 37256
rect 3049 37226 3115 37229
rect 0 37224 3115 37226
rect 0 37168 3054 37224
rect 3110 37168 3115 37224
rect 0 37166 3115 37168
rect 0 37136 800 37166
rect 3049 37163 3115 37166
rect 10874 37024 11194 37025
rect 10874 36960 10882 37024
rect 10946 36960 10962 37024
rect 11026 36960 11042 37024
rect 11106 36960 11122 37024
rect 11186 36960 11194 37024
rect 10874 36959 11194 36960
rect 20805 37024 21125 37025
rect 20805 36960 20813 37024
rect 20877 36960 20893 37024
rect 20957 36960 20973 37024
rect 21037 36960 21053 37024
rect 21117 36960 21125 37024
rect 20805 36959 21125 36960
rect 0 36546 800 36576
rect 2313 36546 2379 36549
rect 0 36544 2379 36546
rect 0 36488 2318 36544
rect 2374 36488 2379 36544
rect 0 36486 2379 36488
rect 0 36456 800 36486
rect 2313 36483 2379 36486
rect 5909 36480 6229 36481
rect 5909 36416 5917 36480
rect 5981 36416 5997 36480
rect 6061 36416 6077 36480
rect 6141 36416 6157 36480
rect 6221 36416 6229 36480
rect 5909 36415 6229 36416
rect 15840 36480 16160 36481
rect 15840 36416 15848 36480
rect 15912 36416 15928 36480
rect 15992 36416 16008 36480
rect 16072 36416 16088 36480
rect 16152 36416 16160 36480
rect 15840 36415 16160 36416
rect 25770 36480 26090 36481
rect 25770 36416 25778 36480
rect 25842 36416 25858 36480
rect 25922 36416 25938 36480
rect 26002 36416 26018 36480
rect 26082 36416 26090 36480
rect 25770 36415 26090 36416
rect 10041 36274 10107 36277
rect 11513 36274 11579 36277
rect 10041 36272 11579 36274
rect 10041 36216 10046 36272
rect 10102 36216 11518 36272
rect 11574 36216 11579 36272
rect 10041 36214 11579 36216
rect 10041 36211 10107 36214
rect 11513 36211 11579 36214
rect 30097 36274 30163 36277
rect 31200 36274 32000 36304
rect 30097 36272 32000 36274
rect 30097 36216 30102 36272
rect 30158 36216 32000 36272
rect 30097 36214 32000 36216
rect 30097 36211 30163 36214
rect 31200 36184 32000 36214
rect 9673 36138 9739 36141
rect 11513 36138 11579 36141
rect 9673 36136 11579 36138
rect 9673 36080 9678 36136
rect 9734 36080 11518 36136
rect 11574 36080 11579 36136
rect 9673 36078 11579 36080
rect 9673 36075 9739 36078
rect 11513 36075 11579 36078
rect 10874 35936 11194 35937
rect 10874 35872 10882 35936
rect 10946 35872 10962 35936
rect 11026 35872 11042 35936
rect 11106 35872 11122 35936
rect 11186 35872 11194 35936
rect 10874 35871 11194 35872
rect 20805 35936 21125 35937
rect 20805 35872 20813 35936
rect 20877 35872 20893 35936
rect 20957 35872 20973 35936
rect 21037 35872 21053 35936
rect 21117 35872 21125 35936
rect 20805 35871 21125 35872
rect 0 35730 800 35760
rect 1393 35730 1459 35733
rect 0 35728 1459 35730
rect 0 35672 1398 35728
rect 1454 35672 1459 35728
rect 0 35670 1459 35672
rect 0 35640 800 35670
rect 1393 35667 1459 35670
rect 5909 35392 6229 35393
rect 5909 35328 5917 35392
rect 5981 35328 5997 35392
rect 6061 35328 6077 35392
rect 6141 35328 6157 35392
rect 6221 35328 6229 35392
rect 5909 35327 6229 35328
rect 15840 35392 16160 35393
rect 15840 35328 15848 35392
rect 15912 35328 15928 35392
rect 15992 35328 16008 35392
rect 16072 35328 16088 35392
rect 16152 35328 16160 35392
rect 15840 35327 16160 35328
rect 25770 35392 26090 35393
rect 25770 35328 25778 35392
rect 25842 35328 25858 35392
rect 25922 35328 25938 35392
rect 26002 35328 26018 35392
rect 26082 35328 26090 35392
rect 25770 35327 26090 35328
rect 0 35050 800 35080
rect 1485 35050 1551 35053
rect 0 35048 1551 35050
rect 0 34992 1490 35048
rect 1546 34992 1551 35048
rect 0 34990 1551 34992
rect 0 34960 800 34990
rect 1485 34987 1551 34990
rect 10874 34848 11194 34849
rect 10874 34784 10882 34848
rect 10946 34784 10962 34848
rect 11026 34784 11042 34848
rect 11106 34784 11122 34848
rect 11186 34784 11194 34848
rect 10874 34783 11194 34784
rect 20805 34848 21125 34849
rect 20805 34784 20813 34848
rect 20877 34784 20893 34848
rect 20957 34784 20973 34848
rect 21037 34784 21053 34848
rect 21117 34784 21125 34848
rect 20805 34783 21125 34784
rect 30097 34778 30163 34781
rect 31200 34778 32000 34808
rect 30097 34776 32000 34778
rect 30097 34720 30102 34776
rect 30158 34720 32000 34776
rect 30097 34718 32000 34720
rect 30097 34715 30163 34718
rect 31200 34688 32000 34718
rect 5909 34304 6229 34305
rect 0 34234 800 34264
rect 5909 34240 5917 34304
rect 5981 34240 5997 34304
rect 6061 34240 6077 34304
rect 6141 34240 6157 34304
rect 6221 34240 6229 34304
rect 5909 34239 6229 34240
rect 15840 34304 16160 34305
rect 15840 34240 15848 34304
rect 15912 34240 15928 34304
rect 15992 34240 16008 34304
rect 16072 34240 16088 34304
rect 16152 34240 16160 34304
rect 15840 34239 16160 34240
rect 25770 34304 26090 34305
rect 25770 34240 25778 34304
rect 25842 34240 25858 34304
rect 25922 34240 25938 34304
rect 26002 34240 26018 34304
rect 26082 34240 26090 34304
rect 25770 34239 26090 34240
rect 2957 34234 3023 34237
rect 0 34232 3023 34234
rect 0 34176 2962 34232
rect 3018 34176 3023 34232
rect 0 34174 3023 34176
rect 0 34144 800 34174
rect 2957 34171 3023 34174
rect 10874 33760 11194 33761
rect 10874 33696 10882 33760
rect 10946 33696 10962 33760
rect 11026 33696 11042 33760
rect 11106 33696 11122 33760
rect 11186 33696 11194 33760
rect 10874 33695 11194 33696
rect 20805 33760 21125 33761
rect 20805 33696 20813 33760
rect 20877 33696 20893 33760
rect 20957 33696 20973 33760
rect 21037 33696 21053 33760
rect 21117 33696 21125 33760
rect 20805 33695 21125 33696
rect 0 33554 800 33584
rect 2957 33554 3023 33557
rect 0 33552 3023 33554
rect 0 33496 2962 33552
rect 3018 33496 3023 33552
rect 0 33494 3023 33496
rect 0 33464 800 33494
rect 2957 33491 3023 33494
rect 30005 33282 30071 33285
rect 31200 33282 32000 33312
rect 30005 33280 32000 33282
rect 30005 33224 30010 33280
rect 30066 33224 32000 33280
rect 30005 33222 32000 33224
rect 30005 33219 30071 33222
rect 5909 33216 6229 33217
rect 5909 33152 5917 33216
rect 5981 33152 5997 33216
rect 6061 33152 6077 33216
rect 6141 33152 6157 33216
rect 6221 33152 6229 33216
rect 5909 33151 6229 33152
rect 15840 33216 16160 33217
rect 15840 33152 15848 33216
rect 15912 33152 15928 33216
rect 15992 33152 16008 33216
rect 16072 33152 16088 33216
rect 16152 33152 16160 33216
rect 15840 33151 16160 33152
rect 25770 33216 26090 33217
rect 25770 33152 25778 33216
rect 25842 33152 25858 33216
rect 25922 33152 25938 33216
rect 26002 33152 26018 33216
rect 26082 33152 26090 33216
rect 31200 33192 32000 33222
rect 25770 33151 26090 33152
rect 0 32738 800 32768
rect 1485 32738 1551 32741
rect 0 32736 1551 32738
rect 0 32680 1490 32736
rect 1546 32680 1551 32736
rect 0 32678 1551 32680
rect 0 32648 800 32678
rect 1485 32675 1551 32678
rect 10874 32672 11194 32673
rect 10874 32608 10882 32672
rect 10946 32608 10962 32672
rect 11026 32608 11042 32672
rect 11106 32608 11122 32672
rect 11186 32608 11194 32672
rect 10874 32607 11194 32608
rect 20805 32672 21125 32673
rect 20805 32608 20813 32672
rect 20877 32608 20893 32672
rect 20957 32608 20973 32672
rect 21037 32608 21053 32672
rect 21117 32608 21125 32672
rect 20805 32607 21125 32608
rect 5909 32128 6229 32129
rect 0 32058 800 32088
rect 5909 32064 5917 32128
rect 5981 32064 5997 32128
rect 6061 32064 6077 32128
rect 6141 32064 6157 32128
rect 6221 32064 6229 32128
rect 5909 32063 6229 32064
rect 15840 32128 16160 32129
rect 15840 32064 15848 32128
rect 15912 32064 15928 32128
rect 15992 32064 16008 32128
rect 16072 32064 16088 32128
rect 16152 32064 16160 32128
rect 15840 32063 16160 32064
rect 25770 32128 26090 32129
rect 25770 32064 25778 32128
rect 25842 32064 25858 32128
rect 25922 32064 25938 32128
rect 26002 32064 26018 32128
rect 26082 32064 26090 32128
rect 25770 32063 26090 32064
rect 2221 32058 2287 32061
rect 0 32056 2287 32058
rect 0 32000 2226 32056
rect 2282 32000 2287 32056
rect 0 31998 2287 32000
rect 0 31968 800 31998
rect 2221 31995 2287 31998
rect 30005 31650 30071 31653
rect 31200 31650 32000 31680
rect 30005 31648 32000 31650
rect 30005 31592 30010 31648
rect 30066 31592 32000 31648
rect 30005 31590 32000 31592
rect 30005 31587 30071 31590
rect 10874 31584 11194 31585
rect 10874 31520 10882 31584
rect 10946 31520 10962 31584
rect 11026 31520 11042 31584
rect 11106 31520 11122 31584
rect 11186 31520 11194 31584
rect 10874 31519 11194 31520
rect 20805 31584 21125 31585
rect 20805 31520 20813 31584
rect 20877 31520 20893 31584
rect 20957 31520 20973 31584
rect 21037 31520 21053 31584
rect 21117 31520 21125 31584
rect 31200 31560 32000 31590
rect 20805 31519 21125 31520
rect 0 31378 800 31408
rect 1485 31378 1551 31381
rect 0 31376 1551 31378
rect 0 31320 1490 31376
rect 1546 31320 1551 31376
rect 0 31318 1551 31320
rect 0 31288 800 31318
rect 1485 31315 1551 31318
rect 5909 31040 6229 31041
rect 5909 30976 5917 31040
rect 5981 30976 5997 31040
rect 6061 30976 6077 31040
rect 6141 30976 6157 31040
rect 6221 30976 6229 31040
rect 5909 30975 6229 30976
rect 15840 31040 16160 31041
rect 15840 30976 15848 31040
rect 15912 30976 15928 31040
rect 15992 30976 16008 31040
rect 16072 30976 16088 31040
rect 16152 30976 16160 31040
rect 15840 30975 16160 30976
rect 25770 31040 26090 31041
rect 25770 30976 25778 31040
rect 25842 30976 25858 31040
rect 25922 30976 25938 31040
rect 26002 30976 26018 31040
rect 26082 30976 26090 31040
rect 25770 30975 26090 30976
rect 0 30562 800 30592
rect 3141 30562 3207 30565
rect 0 30560 3207 30562
rect 0 30504 3146 30560
rect 3202 30504 3207 30560
rect 0 30502 3207 30504
rect 0 30472 800 30502
rect 3141 30499 3207 30502
rect 10874 30496 11194 30497
rect 10874 30432 10882 30496
rect 10946 30432 10962 30496
rect 11026 30432 11042 30496
rect 11106 30432 11122 30496
rect 11186 30432 11194 30496
rect 10874 30431 11194 30432
rect 20805 30496 21125 30497
rect 20805 30432 20813 30496
rect 20877 30432 20893 30496
rect 20957 30432 20973 30496
rect 21037 30432 21053 30496
rect 21117 30432 21125 30496
rect 20805 30431 21125 30432
rect 9029 30428 9095 30429
rect 9029 30426 9076 30428
rect 8984 30424 9076 30426
rect 8984 30368 9034 30424
rect 8984 30366 9076 30368
rect 9029 30364 9076 30366
rect 9140 30364 9146 30428
rect 9029 30363 9095 30364
rect 30005 30154 30071 30157
rect 31200 30154 32000 30184
rect 30005 30152 32000 30154
rect 30005 30096 30010 30152
rect 30066 30096 32000 30152
rect 30005 30094 32000 30096
rect 30005 30091 30071 30094
rect 31200 30064 32000 30094
rect 18045 30018 18111 30021
rect 18270 30018 18276 30020
rect 18045 30016 18276 30018
rect 18045 29960 18050 30016
rect 18106 29960 18276 30016
rect 18045 29958 18276 29960
rect 18045 29955 18111 29958
rect 18270 29956 18276 29958
rect 18340 29956 18346 30020
rect 5909 29952 6229 29953
rect 0 29882 800 29912
rect 5909 29888 5917 29952
rect 5981 29888 5997 29952
rect 6061 29888 6077 29952
rect 6141 29888 6157 29952
rect 6221 29888 6229 29952
rect 5909 29887 6229 29888
rect 15840 29952 16160 29953
rect 15840 29888 15848 29952
rect 15912 29888 15928 29952
rect 15992 29888 16008 29952
rect 16072 29888 16088 29952
rect 16152 29888 16160 29952
rect 15840 29887 16160 29888
rect 25770 29952 26090 29953
rect 25770 29888 25778 29952
rect 25842 29888 25858 29952
rect 25922 29888 25938 29952
rect 26002 29888 26018 29952
rect 26082 29888 26090 29952
rect 25770 29887 26090 29888
rect 1485 29882 1551 29885
rect 0 29880 1551 29882
rect 0 29824 1490 29880
rect 1546 29824 1551 29880
rect 0 29822 1551 29824
rect 0 29792 800 29822
rect 1485 29819 1551 29822
rect 10874 29408 11194 29409
rect 10874 29344 10882 29408
rect 10946 29344 10962 29408
rect 11026 29344 11042 29408
rect 11106 29344 11122 29408
rect 11186 29344 11194 29408
rect 10874 29343 11194 29344
rect 20805 29408 21125 29409
rect 20805 29344 20813 29408
rect 20877 29344 20893 29408
rect 20957 29344 20973 29408
rect 21037 29344 21053 29408
rect 21117 29344 21125 29408
rect 20805 29343 21125 29344
rect 0 29066 800 29096
rect 1485 29066 1551 29069
rect 0 29064 1551 29066
rect 0 29008 1490 29064
rect 1546 29008 1551 29064
rect 0 29006 1551 29008
rect 0 28976 800 29006
rect 1485 29003 1551 29006
rect 5909 28864 6229 28865
rect 5909 28800 5917 28864
rect 5981 28800 5997 28864
rect 6061 28800 6077 28864
rect 6141 28800 6157 28864
rect 6221 28800 6229 28864
rect 5909 28799 6229 28800
rect 15840 28864 16160 28865
rect 15840 28800 15848 28864
rect 15912 28800 15928 28864
rect 15992 28800 16008 28864
rect 16072 28800 16088 28864
rect 16152 28800 16160 28864
rect 15840 28799 16160 28800
rect 25770 28864 26090 28865
rect 25770 28800 25778 28864
rect 25842 28800 25858 28864
rect 25922 28800 25938 28864
rect 26002 28800 26018 28864
rect 26082 28800 26090 28864
rect 25770 28799 26090 28800
rect 30005 28522 30071 28525
rect 31200 28522 32000 28552
rect 30005 28520 32000 28522
rect 30005 28464 30010 28520
rect 30066 28464 32000 28520
rect 30005 28462 32000 28464
rect 30005 28459 30071 28462
rect 31200 28432 32000 28462
rect 0 28386 800 28416
rect 1485 28386 1551 28389
rect 0 28384 1551 28386
rect 0 28328 1490 28384
rect 1546 28328 1551 28384
rect 0 28326 1551 28328
rect 0 28296 800 28326
rect 1485 28323 1551 28326
rect 10874 28320 11194 28321
rect 10874 28256 10882 28320
rect 10946 28256 10962 28320
rect 11026 28256 11042 28320
rect 11106 28256 11122 28320
rect 11186 28256 11194 28320
rect 10874 28255 11194 28256
rect 20805 28320 21125 28321
rect 20805 28256 20813 28320
rect 20877 28256 20893 28320
rect 20957 28256 20973 28320
rect 21037 28256 21053 28320
rect 21117 28256 21125 28320
rect 20805 28255 21125 28256
rect 5909 27776 6229 27777
rect 5909 27712 5917 27776
rect 5981 27712 5997 27776
rect 6061 27712 6077 27776
rect 6141 27712 6157 27776
rect 6221 27712 6229 27776
rect 5909 27711 6229 27712
rect 15840 27776 16160 27777
rect 15840 27712 15848 27776
rect 15912 27712 15928 27776
rect 15992 27712 16008 27776
rect 16072 27712 16088 27776
rect 16152 27712 16160 27776
rect 15840 27711 16160 27712
rect 25770 27776 26090 27777
rect 25770 27712 25778 27776
rect 25842 27712 25858 27776
rect 25922 27712 25938 27776
rect 26002 27712 26018 27776
rect 26082 27712 26090 27776
rect 25770 27711 26090 27712
rect 6361 27706 6427 27709
rect 6729 27706 6795 27709
rect 9489 27706 9555 27709
rect 6361 27704 9555 27706
rect 6361 27648 6366 27704
rect 6422 27648 6734 27704
rect 6790 27648 9494 27704
rect 9550 27648 9555 27704
rect 6361 27646 9555 27648
rect 6361 27643 6427 27646
rect 6729 27643 6795 27646
rect 9489 27643 9555 27646
rect 0 27570 800 27600
rect 1485 27570 1551 27573
rect 0 27568 1551 27570
rect 0 27512 1490 27568
rect 1546 27512 1551 27568
rect 0 27510 1551 27512
rect 0 27480 800 27510
rect 1485 27507 1551 27510
rect 9029 27570 9095 27573
rect 9305 27570 9371 27573
rect 14273 27570 14339 27573
rect 9029 27568 9371 27570
rect 9029 27512 9034 27568
rect 9090 27512 9310 27568
rect 9366 27512 9371 27568
rect 9029 27510 9371 27512
rect 9029 27507 9095 27510
rect 9305 27507 9371 27510
rect 10366 27568 14339 27570
rect 10366 27512 14278 27568
rect 14334 27512 14339 27568
rect 10366 27510 14339 27512
rect 10366 27437 10426 27510
rect 14273 27507 14339 27510
rect 8385 27436 8451 27437
rect 8334 27372 8340 27436
rect 8404 27434 8451 27436
rect 8404 27432 8496 27434
rect 8446 27376 8496 27432
rect 8404 27374 8496 27376
rect 10317 27432 10426 27437
rect 10777 27434 10843 27437
rect 10317 27376 10322 27432
rect 10378 27376 10426 27432
rect 10317 27374 10426 27376
rect 10734 27432 10843 27434
rect 10734 27376 10782 27432
rect 10838 27376 10843 27432
rect 8404 27372 8451 27374
rect 8385 27371 8451 27372
rect 10317 27371 10383 27374
rect 10734 27371 10843 27376
rect 7465 27162 7531 27165
rect 9581 27162 9647 27165
rect 7465 27160 9647 27162
rect 7465 27104 7470 27160
rect 7526 27104 9586 27160
rect 9642 27104 9647 27160
rect 7465 27102 9647 27104
rect 7465 27099 7531 27102
rect 9581 27099 9647 27102
rect 10225 27026 10291 27029
rect 10225 27024 10426 27026
rect 10225 26968 10230 27024
rect 10286 26968 10426 27024
rect 10225 26966 10426 26968
rect 10225 26963 10291 26966
rect 0 26890 800 26920
rect 1485 26890 1551 26893
rect 0 26888 1551 26890
rect 0 26832 1490 26888
rect 1546 26832 1551 26888
rect 0 26830 1551 26832
rect 0 26800 800 26830
rect 1485 26827 1551 26830
rect 10366 26754 10426 26966
rect 10501 26890 10567 26893
rect 10734 26890 10794 27371
rect 10874 27232 11194 27233
rect 10874 27168 10882 27232
rect 10946 27168 10962 27232
rect 11026 27168 11042 27232
rect 11106 27168 11122 27232
rect 11186 27168 11194 27232
rect 10874 27167 11194 27168
rect 20805 27232 21125 27233
rect 20805 27168 20813 27232
rect 20877 27168 20893 27232
rect 20957 27168 20973 27232
rect 21037 27168 21053 27232
rect 21117 27168 21125 27232
rect 20805 27167 21125 27168
rect 30005 27026 30071 27029
rect 31200 27026 32000 27056
rect 30005 27024 32000 27026
rect 30005 26968 30010 27024
rect 30066 26968 32000 27024
rect 30005 26966 32000 26968
rect 30005 26963 30071 26966
rect 31200 26936 32000 26966
rect 10501 26888 10794 26890
rect 10501 26832 10506 26888
rect 10562 26832 10794 26888
rect 10501 26830 10794 26832
rect 10501 26827 10567 26830
rect 11605 26754 11671 26757
rect 10366 26752 11671 26754
rect 10366 26696 11610 26752
rect 11666 26696 11671 26752
rect 10366 26694 11671 26696
rect 11605 26691 11671 26694
rect 5909 26688 6229 26689
rect 5909 26624 5917 26688
rect 5981 26624 5997 26688
rect 6061 26624 6077 26688
rect 6141 26624 6157 26688
rect 6221 26624 6229 26688
rect 5909 26623 6229 26624
rect 15840 26688 16160 26689
rect 15840 26624 15848 26688
rect 15912 26624 15928 26688
rect 15992 26624 16008 26688
rect 16072 26624 16088 26688
rect 16152 26624 16160 26688
rect 15840 26623 16160 26624
rect 25770 26688 26090 26689
rect 25770 26624 25778 26688
rect 25842 26624 25858 26688
rect 25922 26624 25938 26688
rect 26002 26624 26018 26688
rect 26082 26624 26090 26688
rect 25770 26623 26090 26624
rect 3785 26482 3851 26485
rect 5717 26482 5783 26485
rect 5901 26482 5967 26485
rect 3785 26480 5967 26482
rect 3785 26424 3790 26480
rect 3846 26424 5722 26480
rect 5778 26424 5906 26480
rect 5962 26424 5967 26480
rect 3785 26422 5967 26424
rect 3785 26419 3851 26422
rect 5717 26419 5783 26422
rect 5901 26419 5967 26422
rect 8334 26284 8340 26348
rect 8404 26346 8410 26348
rect 9581 26346 9647 26349
rect 20713 26346 20779 26349
rect 8404 26344 9647 26346
rect 8404 26288 9586 26344
rect 9642 26288 9647 26344
rect 8404 26286 9647 26288
rect 8404 26284 8410 26286
rect 9581 26283 9647 26286
rect 20670 26344 20779 26346
rect 20670 26288 20718 26344
rect 20774 26288 20779 26344
rect 20670 26283 20779 26288
rect 0 26210 800 26240
rect 1485 26210 1551 26213
rect 0 26208 1551 26210
rect 0 26152 1490 26208
rect 1546 26152 1551 26208
rect 0 26150 1551 26152
rect 0 26120 800 26150
rect 1485 26147 1551 26150
rect 10874 26144 11194 26145
rect 10874 26080 10882 26144
rect 10946 26080 10962 26144
rect 11026 26080 11042 26144
rect 11106 26080 11122 26144
rect 11186 26080 11194 26144
rect 10874 26079 11194 26080
rect 5073 26074 5139 26077
rect 6085 26074 6151 26077
rect 5073 26072 6151 26074
rect 5073 26016 5078 26072
rect 5134 26016 6090 26072
rect 6146 26016 6151 26072
rect 5073 26014 6151 26016
rect 5073 26011 5139 26014
rect 6085 26011 6151 26014
rect 4889 25938 4955 25941
rect 6729 25938 6795 25941
rect 4889 25936 6795 25938
rect 4889 25880 4894 25936
rect 4950 25880 6734 25936
rect 6790 25880 6795 25936
rect 4889 25878 6795 25880
rect 4889 25875 4955 25878
rect 6729 25875 6795 25878
rect 7649 25938 7715 25941
rect 8569 25938 8635 25941
rect 7649 25936 8635 25938
rect 7649 25880 7654 25936
rect 7710 25880 8574 25936
rect 8630 25880 8635 25936
rect 7649 25878 8635 25880
rect 20670 25938 20730 26283
rect 20805 26144 21125 26145
rect 20805 26080 20813 26144
rect 20877 26080 20893 26144
rect 20957 26080 20973 26144
rect 21037 26080 21053 26144
rect 21117 26080 21125 26144
rect 20805 26079 21125 26080
rect 20805 25938 20871 25941
rect 20670 25936 20871 25938
rect 20670 25880 20810 25936
rect 20866 25880 20871 25936
rect 20670 25878 20871 25880
rect 7649 25875 7715 25878
rect 8569 25875 8635 25878
rect 20805 25875 20871 25878
rect 4797 25802 4863 25805
rect 9397 25802 9463 25805
rect 4797 25800 9463 25802
rect 4797 25744 4802 25800
rect 4858 25744 9402 25800
rect 9458 25744 9463 25800
rect 4797 25742 9463 25744
rect 4797 25739 4863 25742
rect 9397 25739 9463 25742
rect 19977 25802 20043 25805
rect 20529 25802 20595 25805
rect 19977 25800 20595 25802
rect 19977 25744 19982 25800
rect 20038 25744 20534 25800
rect 20590 25744 20595 25800
rect 19977 25742 20595 25744
rect 19977 25739 20043 25742
rect 20529 25739 20595 25742
rect 5909 25600 6229 25601
rect 5909 25536 5917 25600
rect 5981 25536 5997 25600
rect 6061 25536 6077 25600
rect 6141 25536 6157 25600
rect 6221 25536 6229 25600
rect 5909 25535 6229 25536
rect 15840 25600 16160 25601
rect 15840 25536 15848 25600
rect 15912 25536 15928 25600
rect 15992 25536 16008 25600
rect 16072 25536 16088 25600
rect 16152 25536 16160 25600
rect 15840 25535 16160 25536
rect 25770 25600 26090 25601
rect 25770 25536 25778 25600
rect 25842 25536 25858 25600
rect 25922 25536 25938 25600
rect 26002 25536 26018 25600
rect 26082 25536 26090 25600
rect 25770 25535 26090 25536
rect 30005 25530 30071 25533
rect 31200 25530 32000 25560
rect 30005 25528 32000 25530
rect 30005 25472 30010 25528
rect 30066 25472 32000 25528
rect 30005 25470 32000 25472
rect 30005 25467 30071 25470
rect 31200 25440 32000 25470
rect 0 25394 800 25424
rect 1485 25394 1551 25397
rect 0 25392 1551 25394
rect 0 25336 1490 25392
rect 1546 25336 1551 25392
rect 0 25334 1551 25336
rect 0 25304 800 25334
rect 1485 25331 1551 25334
rect 7925 25258 7991 25261
rect 9305 25258 9371 25261
rect 7925 25256 9371 25258
rect 7925 25200 7930 25256
rect 7986 25200 9310 25256
rect 9366 25200 9371 25256
rect 7925 25198 9371 25200
rect 7925 25195 7991 25198
rect 9305 25195 9371 25198
rect 10874 25056 11194 25057
rect 10874 24992 10882 25056
rect 10946 24992 10962 25056
rect 11026 24992 11042 25056
rect 11106 24992 11122 25056
rect 11186 24992 11194 25056
rect 10874 24991 11194 24992
rect 20805 25056 21125 25057
rect 20805 24992 20813 25056
rect 20877 24992 20893 25056
rect 20957 24992 20973 25056
rect 21037 24992 21053 25056
rect 21117 24992 21125 25056
rect 20805 24991 21125 24992
rect 5809 24850 5875 24853
rect 8109 24850 8175 24853
rect 5809 24848 8175 24850
rect 5809 24792 5814 24848
rect 5870 24792 8114 24848
rect 8170 24792 8175 24848
rect 5809 24790 8175 24792
rect 5809 24787 5875 24790
rect 8109 24787 8175 24790
rect 0 24714 800 24744
rect 1485 24714 1551 24717
rect 0 24712 1551 24714
rect 0 24656 1490 24712
rect 1546 24656 1551 24712
rect 0 24654 1551 24656
rect 0 24624 800 24654
rect 1485 24651 1551 24654
rect 5909 24512 6229 24513
rect 5909 24448 5917 24512
rect 5981 24448 5997 24512
rect 6061 24448 6077 24512
rect 6141 24448 6157 24512
rect 6221 24448 6229 24512
rect 5909 24447 6229 24448
rect 15840 24512 16160 24513
rect 15840 24448 15848 24512
rect 15912 24448 15928 24512
rect 15992 24448 16008 24512
rect 16072 24448 16088 24512
rect 16152 24448 16160 24512
rect 15840 24447 16160 24448
rect 25770 24512 26090 24513
rect 25770 24448 25778 24512
rect 25842 24448 25858 24512
rect 25922 24448 25938 24512
rect 26002 24448 26018 24512
rect 26082 24448 26090 24512
rect 25770 24447 26090 24448
rect 5073 24306 5139 24309
rect 6177 24306 6243 24309
rect 5073 24304 6243 24306
rect 5073 24248 5078 24304
rect 5134 24248 6182 24304
rect 6238 24248 6243 24304
rect 5073 24246 6243 24248
rect 5073 24243 5139 24246
rect 6177 24243 6243 24246
rect 9765 24170 9831 24173
rect 10685 24170 10751 24173
rect 9765 24168 10751 24170
rect 9765 24112 9770 24168
rect 9826 24112 10690 24168
rect 10746 24112 10751 24168
rect 9765 24110 10751 24112
rect 9765 24107 9831 24110
rect 10685 24107 10751 24110
rect 10874 23968 11194 23969
rect 0 23898 800 23928
rect 10874 23904 10882 23968
rect 10946 23904 10962 23968
rect 11026 23904 11042 23968
rect 11106 23904 11122 23968
rect 11186 23904 11194 23968
rect 10874 23903 11194 23904
rect 20805 23968 21125 23969
rect 20805 23904 20813 23968
rect 20877 23904 20893 23968
rect 20957 23904 20973 23968
rect 21037 23904 21053 23968
rect 21117 23904 21125 23968
rect 20805 23903 21125 23904
rect 1485 23898 1551 23901
rect 0 23896 1551 23898
rect 0 23840 1490 23896
rect 1546 23840 1551 23896
rect 0 23838 1551 23840
rect 0 23808 800 23838
rect 1485 23835 1551 23838
rect 30005 23898 30071 23901
rect 31200 23898 32000 23928
rect 30005 23896 32000 23898
rect 30005 23840 30010 23896
rect 30066 23840 32000 23896
rect 30005 23838 32000 23840
rect 30005 23835 30071 23838
rect 31200 23808 32000 23838
rect 8109 23626 8175 23629
rect 8937 23626 9003 23629
rect 8109 23624 9003 23626
rect 8109 23568 8114 23624
rect 8170 23568 8942 23624
rect 8998 23568 9003 23624
rect 8109 23566 9003 23568
rect 8109 23563 8175 23566
rect 8937 23563 9003 23566
rect 5909 23424 6229 23425
rect 5909 23360 5917 23424
rect 5981 23360 5997 23424
rect 6061 23360 6077 23424
rect 6141 23360 6157 23424
rect 6221 23360 6229 23424
rect 5909 23359 6229 23360
rect 15840 23424 16160 23425
rect 15840 23360 15848 23424
rect 15912 23360 15928 23424
rect 15992 23360 16008 23424
rect 16072 23360 16088 23424
rect 16152 23360 16160 23424
rect 15840 23359 16160 23360
rect 25770 23424 26090 23425
rect 25770 23360 25778 23424
rect 25842 23360 25858 23424
rect 25922 23360 25938 23424
rect 26002 23360 26018 23424
rect 26082 23360 26090 23424
rect 25770 23359 26090 23360
rect 0 23218 800 23248
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 800 23158
rect 1393 23155 1459 23158
rect 18045 23082 18111 23085
rect 19057 23082 19123 23085
rect 18045 23080 19123 23082
rect 18045 23024 18050 23080
rect 18106 23024 19062 23080
rect 19118 23024 19123 23080
rect 18045 23022 19123 23024
rect 18045 23019 18111 23022
rect 19057 23019 19123 23022
rect 10874 22880 11194 22881
rect 10874 22816 10882 22880
rect 10946 22816 10962 22880
rect 11026 22816 11042 22880
rect 11106 22816 11122 22880
rect 11186 22816 11194 22880
rect 10874 22815 11194 22816
rect 20805 22880 21125 22881
rect 20805 22816 20813 22880
rect 20877 22816 20893 22880
rect 20957 22816 20973 22880
rect 21037 22816 21053 22880
rect 21117 22816 21125 22880
rect 20805 22815 21125 22816
rect 16757 22810 16823 22813
rect 16576 22808 16823 22810
rect 16576 22752 16762 22808
rect 16818 22752 16823 22808
rect 16576 22750 16823 22752
rect 16576 22677 16636 22750
rect 16757 22747 16823 22750
rect 16573 22672 16639 22677
rect 16573 22616 16578 22672
rect 16634 22616 16639 22672
rect 16573 22611 16639 22616
rect 0 22402 800 22432
rect 2773 22402 2839 22405
rect 0 22400 2839 22402
rect 0 22344 2778 22400
rect 2834 22344 2839 22400
rect 0 22342 2839 22344
rect 0 22312 800 22342
rect 2773 22339 2839 22342
rect 30005 22402 30071 22405
rect 31200 22402 32000 22432
rect 30005 22400 32000 22402
rect 30005 22344 30010 22400
rect 30066 22344 32000 22400
rect 30005 22342 32000 22344
rect 30005 22339 30071 22342
rect 5909 22336 6229 22337
rect 5909 22272 5917 22336
rect 5981 22272 5997 22336
rect 6061 22272 6077 22336
rect 6141 22272 6157 22336
rect 6221 22272 6229 22336
rect 5909 22271 6229 22272
rect 15840 22336 16160 22337
rect 15840 22272 15848 22336
rect 15912 22272 15928 22336
rect 15992 22272 16008 22336
rect 16072 22272 16088 22336
rect 16152 22272 16160 22336
rect 15840 22271 16160 22272
rect 25770 22336 26090 22337
rect 25770 22272 25778 22336
rect 25842 22272 25858 22336
rect 25922 22272 25938 22336
rect 26002 22272 26018 22336
rect 26082 22272 26090 22336
rect 31200 22312 32000 22342
rect 25770 22271 26090 22272
rect 15745 22130 15811 22133
rect 15745 22128 15946 22130
rect 15745 22072 15750 22128
rect 15806 22072 15946 22128
rect 15745 22070 15946 22072
rect 15745 22067 15811 22070
rect 8201 21994 8267 21997
rect 8334 21994 8340 21996
rect 8201 21992 8340 21994
rect 8201 21936 8206 21992
rect 8262 21936 8340 21992
rect 8201 21934 8340 21936
rect 8201 21931 8267 21934
rect 8334 21932 8340 21934
rect 8404 21932 8410 21996
rect 15886 21994 15946 22070
rect 16205 21994 16271 21997
rect 15886 21992 16271 21994
rect 15886 21936 16210 21992
rect 16266 21936 16271 21992
rect 15886 21934 16271 21936
rect 16205 21931 16271 21934
rect 10874 21792 11194 21793
rect 0 21722 800 21752
rect 10874 21728 10882 21792
rect 10946 21728 10962 21792
rect 11026 21728 11042 21792
rect 11106 21728 11122 21792
rect 11186 21728 11194 21792
rect 10874 21727 11194 21728
rect 20805 21792 21125 21793
rect 20805 21728 20813 21792
rect 20877 21728 20893 21792
rect 20957 21728 20973 21792
rect 21037 21728 21053 21792
rect 21117 21728 21125 21792
rect 20805 21727 21125 21728
rect 2037 21722 2103 21725
rect 0 21720 2103 21722
rect 0 21664 2042 21720
rect 2098 21664 2103 21720
rect 0 21662 2103 21664
rect 0 21632 800 21662
rect 2037 21659 2103 21662
rect 17125 21722 17191 21725
rect 17585 21722 17651 21725
rect 17125 21720 17651 21722
rect 17125 21664 17130 21720
rect 17186 21664 17590 21720
rect 17646 21664 17651 21720
rect 17125 21662 17651 21664
rect 17125 21659 17191 21662
rect 17585 21659 17651 21662
rect 18597 21722 18663 21725
rect 19241 21722 19307 21725
rect 18597 21720 19307 21722
rect 18597 21664 18602 21720
rect 18658 21664 19246 21720
rect 19302 21664 19307 21720
rect 18597 21662 19307 21664
rect 18597 21659 18663 21662
rect 19241 21659 19307 21662
rect 5909 21248 6229 21249
rect 5909 21184 5917 21248
rect 5981 21184 5997 21248
rect 6061 21184 6077 21248
rect 6141 21184 6157 21248
rect 6221 21184 6229 21248
rect 5909 21183 6229 21184
rect 15840 21248 16160 21249
rect 15840 21184 15848 21248
rect 15912 21184 15928 21248
rect 15992 21184 16008 21248
rect 16072 21184 16088 21248
rect 16152 21184 16160 21248
rect 15840 21183 16160 21184
rect 25770 21248 26090 21249
rect 25770 21184 25778 21248
rect 25842 21184 25858 21248
rect 25922 21184 25938 21248
rect 26002 21184 26018 21248
rect 26082 21184 26090 21248
rect 25770 21183 26090 21184
rect 0 21042 800 21072
rect 1393 21042 1459 21045
rect 0 21040 1459 21042
rect 0 20984 1398 21040
rect 1454 20984 1459 21040
rect 0 20982 1459 20984
rect 0 20952 800 20982
rect 1393 20979 1459 20982
rect 30005 20906 30071 20909
rect 31200 20906 32000 20936
rect 30005 20904 32000 20906
rect 30005 20848 30010 20904
rect 30066 20848 32000 20904
rect 30005 20846 32000 20848
rect 30005 20843 30071 20846
rect 31200 20816 32000 20846
rect 10874 20704 11194 20705
rect 10874 20640 10882 20704
rect 10946 20640 10962 20704
rect 11026 20640 11042 20704
rect 11106 20640 11122 20704
rect 11186 20640 11194 20704
rect 10874 20639 11194 20640
rect 20805 20704 21125 20705
rect 20805 20640 20813 20704
rect 20877 20640 20893 20704
rect 20957 20640 20973 20704
rect 21037 20640 21053 20704
rect 21117 20640 21125 20704
rect 20805 20639 21125 20640
rect 0 20226 800 20256
rect 4061 20226 4127 20229
rect 0 20224 4127 20226
rect 0 20168 4066 20224
rect 4122 20168 4127 20224
rect 0 20166 4127 20168
rect 0 20136 800 20166
rect 4061 20163 4127 20166
rect 5909 20160 6229 20161
rect 5909 20096 5917 20160
rect 5981 20096 5997 20160
rect 6061 20096 6077 20160
rect 6141 20096 6157 20160
rect 6221 20096 6229 20160
rect 5909 20095 6229 20096
rect 15840 20160 16160 20161
rect 15840 20096 15848 20160
rect 15912 20096 15928 20160
rect 15992 20096 16008 20160
rect 16072 20096 16088 20160
rect 16152 20096 16160 20160
rect 15840 20095 16160 20096
rect 25770 20160 26090 20161
rect 25770 20096 25778 20160
rect 25842 20096 25858 20160
rect 25922 20096 25938 20160
rect 26002 20096 26018 20160
rect 26082 20096 26090 20160
rect 25770 20095 26090 20096
rect 3141 19954 3207 19957
rect 8017 19954 8083 19957
rect 3141 19952 8083 19954
rect 3141 19896 3146 19952
rect 3202 19896 8022 19952
rect 8078 19896 8083 19952
rect 3141 19894 8083 19896
rect 3141 19891 3207 19894
rect 8017 19891 8083 19894
rect 5809 19818 5875 19821
rect 6913 19818 6979 19821
rect 5809 19816 6979 19818
rect 5809 19760 5814 19816
rect 5870 19760 6918 19816
rect 6974 19760 6979 19816
rect 5809 19758 6979 19760
rect 5809 19755 5875 19758
rect 6913 19755 6979 19758
rect 16573 19818 16639 19821
rect 17309 19818 17375 19821
rect 16573 19816 17375 19818
rect 16573 19760 16578 19816
rect 16634 19760 17314 19816
rect 17370 19760 17375 19816
rect 16573 19758 17375 19760
rect 16573 19755 16639 19758
rect 17309 19755 17375 19758
rect 10874 19616 11194 19617
rect 0 19546 800 19576
rect 10874 19552 10882 19616
rect 10946 19552 10962 19616
rect 11026 19552 11042 19616
rect 11106 19552 11122 19616
rect 11186 19552 11194 19616
rect 10874 19551 11194 19552
rect 20805 19616 21125 19617
rect 20805 19552 20813 19616
rect 20877 19552 20893 19616
rect 20957 19552 20973 19616
rect 21037 19552 21053 19616
rect 21117 19552 21125 19616
rect 20805 19551 21125 19552
rect 3233 19546 3299 19549
rect 0 19544 3299 19546
rect 0 19488 3238 19544
rect 3294 19488 3299 19544
rect 0 19486 3299 19488
rect 0 19456 800 19486
rect 3233 19483 3299 19486
rect 30005 19274 30071 19277
rect 31200 19274 32000 19304
rect 30005 19272 32000 19274
rect 30005 19216 30010 19272
rect 30066 19216 32000 19272
rect 30005 19214 32000 19216
rect 30005 19211 30071 19214
rect 31200 19184 32000 19214
rect 5909 19072 6229 19073
rect 5909 19008 5917 19072
rect 5981 19008 5997 19072
rect 6061 19008 6077 19072
rect 6141 19008 6157 19072
rect 6221 19008 6229 19072
rect 5909 19007 6229 19008
rect 15840 19072 16160 19073
rect 15840 19008 15848 19072
rect 15912 19008 15928 19072
rect 15992 19008 16008 19072
rect 16072 19008 16088 19072
rect 16152 19008 16160 19072
rect 15840 19007 16160 19008
rect 25770 19072 26090 19073
rect 25770 19008 25778 19072
rect 25842 19008 25858 19072
rect 25922 19008 25938 19072
rect 26002 19008 26018 19072
rect 26082 19008 26090 19072
rect 25770 19007 26090 19008
rect 0 18730 800 18760
rect 2957 18730 3023 18733
rect 0 18728 3023 18730
rect 0 18672 2962 18728
rect 3018 18672 3023 18728
rect 0 18670 3023 18672
rect 0 18640 800 18670
rect 2957 18667 3023 18670
rect 10874 18528 11194 18529
rect 10874 18464 10882 18528
rect 10946 18464 10962 18528
rect 11026 18464 11042 18528
rect 11106 18464 11122 18528
rect 11186 18464 11194 18528
rect 10874 18463 11194 18464
rect 20805 18528 21125 18529
rect 20805 18464 20813 18528
rect 20877 18464 20893 18528
rect 20957 18464 20973 18528
rect 21037 18464 21053 18528
rect 21117 18464 21125 18528
rect 20805 18463 21125 18464
rect 6637 18322 6703 18325
rect 9489 18322 9555 18325
rect 6637 18320 6746 18322
rect 6637 18264 6642 18320
rect 6698 18264 6746 18320
rect 6637 18259 6746 18264
rect 0 18050 800 18080
rect 6686 18053 6746 18259
rect 9446 18320 9555 18322
rect 9446 18264 9494 18320
rect 9550 18264 9555 18320
rect 9446 18259 9555 18264
rect 3049 18050 3115 18053
rect 0 18048 3115 18050
rect 0 17992 3054 18048
rect 3110 17992 3115 18048
rect 0 17990 3115 17992
rect 0 17960 800 17990
rect 3049 17987 3115 17990
rect 6637 18048 6746 18053
rect 6637 17992 6642 18048
rect 6698 17992 6746 18048
rect 6637 17990 6746 17992
rect 9305 18050 9371 18053
rect 9446 18050 9506 18259
rect 9305 18048 9506 18050
rect 9305 17992 9310 18048
rect 9366 17992 9506 18048
rect 9305 17990 9506 17992
rect 6637 17987 6703 17990
rect 9305 17987 9371 17990
rect 5909 17984 6229 17985
rect 5909 17920 5917 17984
rect 5981 17920 5997 17984
rect 6061 17920 6077 17984
rect 6141 17920 6157 17984
rect 6221 17920 6229 17984
rect 5909 17919 6229 17920
rect 15840 17984 16160 17985
rect 15840 17920 15848 17984
rect 15912 17920 15928 17984
rect 15992 17920 16008 17984
rect 16072 17920 16088 17984
rect 16152 17920 16160 17984
rect 15840 17919 16160 17920
rect 25770 17984 26090 17985
rect 25770 17920 25778 17984
rect 25842 17920 25858 17984
rect 25922 17920 25938 17984
rect 26002 17920 26018 17984
rect 26082 17920 26090 17984
rect 25770 17919 26090 17920
rect 30005 17778 30071 17781
rect 31200 17778 32000 17808
rect 30005 17776 32000 17778
rect 30005 17720 30010 17776
rect 30066 17720 32000 17776
rect 30005 17718 32000 17720
rect 30005 17715 30071 17718
rect 31200 17688 32000 17718
rect 10874 17440 11194 17441
rect 10874 17376 10882 17440
rect 10946 17376 10962 17440
rect 11026 17376 11042 17440
rect 11106 17376 11122 17440
rect 11186 17376 11194 17440
rect 10874 17375 11194 17376
rect 20805 17440 21125 17441
rect 20805 17376 20813 17440
rect 20877 17376 20893 17440
rect 20957 17376 20973 17440
rect 21037 17376 21053 17440
rect 21117 17376 21125 17440
rect 20805 17375 21125 17376
rect 0 17234 800 17264
rect 2773 17234 2839 17237
rect 0 17232 2839 17234
rect 0 17176 2778 17232
rect 2834 17176 2839 17232
rect 0 17174 2839 17176
rect 0 17144 800 17174
rect 2773 17171 2839 17174
rect 5909 16896 6229 16897
rect 5909 16832 5917 16896
rect 5981 16832 5997 16896
rect 6061 16832 6077 16896
rect 6141 16832 6157 16896
rect 6221 16832 6229 16896
rect 5909 16831 6229 16832
rect 15840 16896 16160 16897
rect 15840 16832 15848 16896
rect 15912 16832 15928 16896
rect 15992 16832 16008 16896
rect 16072 16832 16088 16896
rect 16152 16832 16160 16896
rect 15840 16831 16160 16832
rect 25770 16896 26090 16897
rect 25770 16832 25778 16896
rect 25842 16832 25858 16896
rect 25922 16832 25938 16896
rect 26002 16832 26018 16896
rect 26082 16832 26090 16896
rect 25770 16831 26090 16832
rect 0 16554 800 16584
rect 3233 16554 3299 16557
rect 0 16552 3299 16554
rect 0 16496 3238 16552
rect 3294 16496 3299 16552
rect 0 16494 3299 16496
rect 0 16464 800 16494
rect 3233 16491 3299 16494
rect 10874 16352 11194 16353
rect 10874 16288 10882 16352
rect 10946 16288 10962 16352
rect 11026 16288 11042 16352
rect 11106 16288 11122 16352
rect 11186 16288 11194 16352
rect 10874 16287 11194 16288
rect 20805 16352 21125 16353
rect 20805 16288 20813 16352
rect 20877 16288 20893 16352
rect 20957 16288 20973 16352
rect 21037 16288 21053 16352
rect 21117 16288 21125 16352
rect 20805 16287 21125 16288
rect 16665 16282 16731 16285
rect 18689 16282 18755 16285
rect 16665 16280 18755 16282
rect 16665 16224 16670 16280
rect 16726 16224 18694 16280
rect 18750 16224 18755 16280
rect 16665 16222 18755 16224
rect 16665 16219 16731 16222
rect 18689 16219 18755 16222
rect 7465 16146 7531 16149
rect 10685 16146 10751 16149
rect 7465 16144 10751 16146
rect 7465 16088 7470 16144
rect 7526 16088 10690 16144
rect 10746 16088 10751 16144
rect 7465 16086 10751 16088
rect 7465 16083 7531 16086
rect 10685 16083 10751 16086
rect 18045 16146 18111 16149
rect 18270 16146 18276 16148
rect 18045 16144 18276 16146
rect 18045 16088 18050 16144
rect 18106 16088 18276 16144
rect 18045 16086 18276 16088
rect 18045 16083 18111 16086
rect 18270 16084 18276 16086
rect 18340 16084 18346 16148
rect 30005 16146 30071 16149
rect 31200 16146 32000 16176
rect 30005 16144 32000 16146
rect 30005 16088 30010 16144
rect 30066 16088 32000 16144
rect 30005 16086 32000 16088
rect 30005 16083 30071 16086
rect 31200 16056 32000 16086
rect 5758 15948 5764 16012
rect 5828 16010 5834 16012
rect 6269 16010 6335 16013
rect 5828 16008 6335 16010
rect 5828 15952 6274 16008
rect 6330 15952 6335 16008
rect 5828 15950 6335 15952
rect 5828 15948 5834 15950
rect 6269 15947 6335 15950
rect 17677 16010 17743 16013
rect 18597 16010 18663 16013
rect 17677 16008 18663 16010
rect 17677 15952 17682 16008
rect 17738 15952 18602 16008
rect 18658 15952 18663 16008
rect 17677 15950 18663 15952
rect 17677 15947 17743 15950
rect 18597 15947 18663 15950
rect 0 15874 800 15904
rect 1393 15874 1459 15877
rect 0 15872 1459 15874
rect 0 15816 1398 15872
rect 1454 15816 1459 15872
rect 0 15814 1459 15816
rect 0 15784 800 15814
rect 1393 15811 1459 15814
rect 16941 15874 17007 15877
rect 19057 15874 19123 15877
rect 16941 15872 19123 15874
rect 16941 15816 16946 15872
rect 17002 15816 19062 15872
rect 19118 15816 19123 15872
rect 16941 15814 19123 15816
rect 16941 15811 17007 15814
rect 19057 15811 19123 15814
rect 5909 15808 6229 15809
rect 5909 15744 5917 15808
rect 5981 15744 5997 15808
rect 6061 15744 6077 15808
rect 6141 15744 6157 15808
rect 6221 15744 6229 15808
rect 5909 15743 6229 15744
rect 15840 15808 16160 15809
rect 15840 15744 15848 15808
rect 15912 15744 15928 15808
rect 15992 15744 16008 15808
rect 16072 15744 16088 15808
rect 16152 15744 16160 15808
rect 15840 15743 16160 15744
rect 25770 15808 26090 15809
rect 25770 15744 25778 15808
rect 25842 15744 25858 15808
rect 25922 15744 25938 15808
rect 26002 15744 26018 15808
rect 26082 15744 26090 15808
rect 25770 15743 26090 15744
rect 10874 15264 11194 15265
rect 10874 15200 10882 15264
rect 10946 15200 10962 15264
rect 11026 15200 11042 15264
rect 11106 15200 11122 15264
rect 11186 15200 11194 15264
rect 10874 15199 11194 15200
rect 20805 15264 21125 15265
rect 20805 15200 20813 15264
rect 20877 15200 20893 15264
rect 20957 15200 20973 15264
rect 21037 15200 21053 15264
rect 21117 15200 21125 15264
rect 20805 15199 21125 15200
rect 0 15058 800 15088
rect 1209 15058 1275 15061
rect 0 15056 1275 15058
rect 0 15000 1214 15056
rect 1270 15000 1275 15056
rect 0 14998 1275 15000
rect 0 14968 800 14998
rect 1209 14995 1275 14998
rect 5909 14720 6229 14721
rect 5909 14656 5917 14720
rect 5981 14656 5997 14720
rect 6061 14656 6077 14720
rect 6141 14656 6157 14720
rect 6221 14656 6229 14720
rect 5909 14655 6229 14656
rect 15840 14720 16160 14721
rect 15840 14656 15848 14720
rect 15912 14656 15928 14720
rect 15992 14656 16008 14720
rect 16072 14656 16088 14720
rect 16152 14656 16160 14720
rect 15840 14655 16160 14656
rect 25770 14720 26090 14721
rect 25770 14656 25778 14720
rect 25842 14656 25858 14720
rect 25922 14656 25938 14720
rect 26002 14656 26018 14720
rect 26082 14656 26090 14720
rect 25770 14655 26090 14656
rect 30005 14650 30071 14653
rect 31200 14650 32000 14680
rect 30005 14648 32000 14650
rect 30005 14592 30010 14648
rect 30066 14592 32000 14648
rect 30005 14590 32000 14592
rect 30005 14587 30071 14590
rect 31200 14560 32000 14590
rect 1393 14514 1459 14517
rect 798 14512 1459 14514
rect 798 14456 1398 14512
rect 1454 14456 1459 14512
rect 798 14454 1459 14456
rect 798 14408 858 14454
rect 1393 14451 1459 14454
rect 12341 14514 12407 14517
rect 16297 14514 16363 14517
rect 12341 14512 16363 14514
rect 12341 14456 12346 14512
rect 12402 14456 16302 14512
rect 16358 14456 16363 14512
rect 12341 14454 16363 14456
rect 12341 14451 12407 14454
rect 16297 14451 16363 14454
rect 0 14318 858 14408
rect 6177 14378 6243 14381
rect 11237 14378 11303 14381
rect 6177 14376 11303 14378
rect 6177 14320 6182 14376
rect 6238 14320 11242 14376
rect 11298 14320 11303 14376
rect 6177 14318 11303 14320
rect 0 14288 800 14318
rect 6177 14315 6243 14318
rect 11237 14315 11303 14318
rect 11881 14378 11947 14381
rect 18321 14378 18387 14381
rect 11881 14376 18387 14378
rect 11881 14320 11886 14376
rect 11942 14320 18326 14376
rect 18382 14320 18387 14376
rect 11881 14318 18387 14320
rect 11881 14315 11947 14318
rect 18321 14315 18387 14318
rect 10874 14176 11194 14177
rect 10874 14112 10882 14176
rect 10946 14112 10962 14176
rect 11026 14112 11042 14176
rect 11106 14112 11122 14176
rect 11186 14112 11194 14176
rect 10874 14111 11194 14112
rect 20805 14176 21125 14177
rect 20805 14112 20813 14176
rect 20877 14112 20893 14176
rect 20957 14112 20973 14176
rect 21037 14112 21053 14176
rect 21117 14112 21125 14176
rect 20805 14111 21125 14112
rect 7557 14106 7623 14109
rect 9581 14106 9647 14109
rect 7557 14104 9647 14106
rect 7557 14048 7562 14104
rect 7618 14048 9586 14104
rect 9642 14048 9647 14104
rect 7557 14046 9647 14048
rect 7557 14043 7623 14046
rect 9581 14043 9647 14046
rect 8017 13970 8083 13973
rect 9121 13970 9187 13973
rect 8017 13968 9187 13970
rect 8017 13912 8022 13968
rect 8078 13912 9126 13968
rect 9182 13912 9187 13968
rect 8017 13910 9187 13912
rect 8017 13907 8083 13910
rect 9121 13907 9187 13910
rect 13721 13970 13787 13973
rect 17953 13970 18019 13973
rect 13721 13968 18019 13970
rect 13721 13912 13726 13968
rect 13782 13912 17958 13968
rect 18014 13912 18019 13968
rect 13721 13910 18019 13912
rect 13721 13907 13787 13910
rect 17953 13907 18019 13910
rect 17033 13698 17099 13701
rect 18321 13698 18387 13701
rect 17033 13696 18387 13698
rect 17033 13640 17038 13696
rect 17094 13640 18326 13696
rect 18382 13640 18387 13696
rect 17033 13638 18387 13640
rect 17033 13635 17099 13638
rect 18321 13635 18387 13638
rect 5909 13632 6229 13633
rect 0 13562 800 13592
rect 5909 13568 5917 13632
rect 5981 13568 5997 13632
rect 6061 13568 6077 13632
rect 6141 13568 6157 13632
rect 6221 13568 6229 13632
rect 5909 13567 6229 13568
rect 15840 13632 16160 13633
rect 15840 13568 15848 13632
rect 15912 13568 15928 13632
rect 15992 13568 16008 13632
rect 16072 13568 16088 13632
rect 16152 13568 16160 13632
rect 15840 13567 16160 13568
rect 25770 13632 26090 13633
rect 25770 13568 25778 13632
rect 25842 13568 25858 13632
rect 25922 13568 25938 13632
rect 26002 13568 26018 13632
rect 26082 13568 26090 13632
rect 25770 13567 26090 13568
rect 2773 13562 2839 13565
rect 0 13560 2839 13562
rect 0 13504 2778 13560
rect 2834 13504 2839 13560
rect 0 13502 2839 13504
rect 0 13472 800 13502
rect 2773 13499 2839 13502
rect 30005 13154 30071 13157
rect 31200 13154 32000 13184
rect 30005 13152 32000 13154
rect 30005 13096 30010 13152
rect 30066 13096 32000 13152
rect 30005 13094 32000 13096
rect 30005 13091 30071 13094
rect 10874 13088 11194 13089
rect 10874 13024 10882 13088
rect 10946 13024 10962 13088
rect 11026 13024 11042 13088
rect 11106 13024 11122 13088
rect 11186 13024 11194 13088
rect 10874 13023 11194 13024
rect 20805 13088 21125 13089
rect 20805 13024 20813 13088
rect 20877 13024 20893 13088
rect 20957 13024 20973 13088
rect 21037 13024 21053 13088
rect 21117 13024 21125 13088
rect 31200 13064 32000 13094
rect 20805 13023 21125 13024
rect 0 12882 800 12912
rect 1209 12882 1275 12885
rect 0 12880 1275 12882
rect 0 12824 1214 12880
rect 1270 12824 1275 12880
rect 0 12822 1275 12824
rect 0 12792 800 12822
rect 1209 12819 1275 12822
rect 5909 12544 6229 12545
rect 5909 12480 5917 12544
rect 5981 12480 5997 12544
rect 6061 12480 6077 12544
rect 6141 12480 6157 12544
rect 6221 12480 6229 12544
rect 5909 12479 6229 12480
rect 15840 12544 16160 12545
rect 15840 12480 15848 12544
rect 15912 12480 15928 12544
rect 15992 12480 16008 12544
rect 16072 12480 16088 12544
rect 16152 12480 16160 12544
rect 15840 12479 16160 12480
rect 25770 12544 26090 12545
rect 25770 12480 25778 12544
rect 25842 12480 25858 12544
rect 25922 12480 25938 12544
rect 26002 12480 26018 12544
rect 26082 12480 26090 12544
rect 25770 12479 26090 12480
rect 0 12066 800 12096
rect 2773 12066 2839 12069
rect 0 12064 2839 12066
rect 0 12008 2778 12064
rect 2834 12008 2839 12064
rect 0 12006 2839 12008
rect 0 11976 800 12006
rect 2773 12003 2839 12006
rect 10874 12000 11194 12001
rect 10874 11936 10882 12000
rect 10946 11936 10962 12000
rect 11026 11936 11042 12000
rect 11106 11936 11122 12000
rect 11186 11936 11194 12000
rect 10874 11935 11194 11936
rect 20805 12000 21125 12001
rect 20805 11936 20813 12000
rect 20877 11936 20893 12000
rect 20957 11936 20973 12000
rect 21037 11936 21053 12000
rect 21117 11936 21125 12000
rect 20805 11935 21125 11936
rect 10225 11794 10291 11797
rect 10501 11794 10567 11797
rect 10225 11792 10567 11794
rect 10225 11736 10230 11792
rect 10286 11736 10506 11792
rect 10562 11736 10567 11792
rect 10225 11734 10567 11736
rect 10225 11731 10291 11734
rect 10501 11731 10567 11734
rect 30005 11522 30071 11525
rect 31200 11522 32000 11552
rect 30005 11520 32000 11522
rect 30005 11464 30010 11520
rect 30066 11464 32000 11520
rect 30005 11462 32000 11464
rect 30005 11459 30071 11462
rect 5909 11456 6229 11457
rect 0 11386 800 11416
rect 5909 11392 5917 11456
rect 5981 11392 5997 11456
rect 6061 11392 6077 11456
rect 6141 11392 6157 11456
rect 6221 11392 6229 11456
rect 5909 11391 6229 11392
rect 15840 11456 16160 11457
rect 15840 11392 15848 11456
rect 15912 11392 15928 11456
rect 15992 11392 16008 11456
rect 16072 11392 16088 11456
rect 16152 11392 16160 11456
rect 15840 11391 16160 11392
rect 25770 11456 26090 11457
rect 25770 11392 25778 11456
rect 25842 11392 25858 11456
rect 25922 11392 25938 11456
rect 26002 11392 26018 11456
rect 26082 11392 26090 11456
rect 31200 11432 32000 11462
rect 25770 11391 26090 11392
rect 1393 11386 1459 11389
rect 0 11384 1459 11386
rect 0 11328 1398 11384
rect 1454 11328 1459 11384
rect 0 11326 1459 11328
rect 0 11296 800 11326
rect 1393 11323 1459 11326
rect 12801 11386 12867 11389
rect 15193 11386 15259 11389
rect 12801 11384 15259 11386
rect 12801 11328 12806 11384
rect 12862 11328 15198 11384
rect 15254 11328 15259 11384
rect 12801 11326 15259 11328
rect 12801 11323 12867 11326
rect 15193 11323 15259 11326
rect 10317 11250 10383 11253
rect 11973 11250 12039 11253
rect 10317 11248 12039 11250
rect 10317 11192 10322 11248
rect 10378 11192 11978 11248
rect 12034 11192 12039 11248
rect 10317 11190 12039 11192
rect 10317 11187 10383 11190
rect 11973 11187 12039 11190
rect 10874 10912 11194 10913
rect 10874 10848 10882 10912
rect 10946 10848 10962 10912
rect 11026 10848 11042 10912
rect 11106 10848 11122 10912
rect 11186 10848 11194 10912
rect 10874 10847 11194 10848
rect 20805 10912 21125 10913
rect 20805 10848 20813 10912
rect 20877 10848 20893 10912
rect 20957 10848 20973 10912
rect 21037 10848 21053 10912
rect 21117 10848 21125 10912
rect 20805 10847 21125 10848
rect 0 10706 800 10736
rect 1393 10706 1459 10709
rect 0 10704 1459 10706
rect 0 10648 1398 10704
rect 1454 10648 1459 10704
rect 0 10646 1459 10648
rect 0 10616 800 10646
rect 1393 10643 1459 10646
rect 5909 10368 6229 10369
rect 5909 10304 5917 10368
rect 5981 10304 5997 10368
rect 6061 10304 6077 10368
rect 6141 10304 6157 10368
rect 6221 10304 6229 10368
rect 5909 10303 6229 10304
rect 15840 10368 16160 10369
rect 15840 10304 15848 10368
rect 15912 10304 15928 10368
rect 15992 10304 16008 10368
rect 16072 10304 16088 10368
rect 16152 10304 16160 10368
rect 15840 10303 16160 10304
rect 25770 10368 26090 10369
rect 25770 10304 25778 10368
rect 25842 10304 25858 10368
rect 25922 10304 25938 10368
rect 26002 10304 26018 10368
rect 26082 10304 26090 10368
rect 25770 10303 26090 10304
rect 30005 10026 30071 10029
rect 31200 10026 32000 10056
rect 30005 10024 32000 10026
rect 30005 9968 30010 10024
rect 30066 9968 32000 10024
rect 30005 9966 32000 9968
rect 30005 9963 30071 9966
rect 31200 9936 32000 9966
rect 0 9890 800 9920
rect 2773 9890 2839 9893
rect 0 9888 2839 9890
rect 0 9832 2778 9888
rect 2834 9832 2839 9888
rect 0 9830 2839 9832
rect 0 9800 800 9830
rect 2773 9827 2839 9830
rect 10874 9824 11194 9825
rect 10874 9760 10882 9824
rect 10946 9760 10962 9824
rect 11026 9760 11042 9824
rect 11106 9760 11122 9824
rect 11186 9760 11194 9824
rect 10874 9759 11194 9760
rect 20805 9824 21125 9825
rect 20805 9760 20813 9824
rect 20877 9760 20893 9824
rect 20957 9760 20973 9824
rect 21037 9760 21053 9824
rect 21117 9760 21125 9824
rect 20805 9759 21125 9760
rect 10041 9618 10107 9621
rect 15653 9618 15719 9621
rect 10041 9616 15719 9618
rect 10041 9560 10046 9616
rect 10102 9560 15658 9616
rect 15714 9560 15719 9616
rect 10041 9558 15719 9560
rect 10041 9555 10107 9558
rect 15653 9555 15719 9558
rect 5909 9280 6229 9281
rect 0 9210 800 9240
rect 5909 9216 5917 9280
rect 5981 9216 5997 9280
rect 6061 9216 6077 9280
rect 6141 9216 6157 9280
rect 6221 9216 6229 9280
rect 5909 9215 6229 9216
rect 15840 9280 16160 9281
rect 15840 9216 15848 9280
rect 15912 9216 15928 9280
rect 15992 9216 16008 9280
rect 16072 9216 16088 9280
rect 16152 9216 16160 9280
rect 15840 9215 16160 9216
rect 25770 9280 26090 9281
rect 25770 9216 25778 9280
rect 25842 9216 25858 9280
rect 25922 9216 25938 9280
rect 26002 9216 26018 9280
rect 26082 9216 26090 9280
rect 25770 9215 26090 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 5257 9074 5323 9077
rect 5758 9074 5764 9076
rect 5257 9072 5764 9074
rect 5257 9016 5262 9072
rect 5318 9016 5764 9072
rect 5257 9014 5764 9016
rect 5257 9011 5323 9014
rect 5758 9012 5764 9014
rect 5828 9012 5834 9076
rect 10874 8736 11194 8737
rect 10874 8672 10882 8736
rect 10946 8672 10962 8736
rect 11026 8672 11042 8736
rect 11106 8672 11122 8736
rect 11186 8672 11194 8736
rect 10874 8671 11194 8672
rect 20805 8736 21125 8737
rect 20805 8672 20813 8736
rect 20877 8672 20893 8736
rect 20957 8672 20973 8736
rect 21037 8672 21053 8736
rect 21117 8672 21125 8736
rect 20805 8671 21125 8672
rect 10501 8530 10567 8533
rect 11789 8530 11855 8533
rect 10501 8528 11855 8530
rect 10501 8472 10506 8528
rect 10562 8472 11794 8528
rect 11850 8472 11855 8528
rect 10501 8470 11855 8472
rect 10501 8467 10567 8470
rect 11789 8467 11855 8470
rect 0 8394 800 8424
rect 1393 8394 1459 8397
rect 0 8392 1459 8394
rect 0 8336 1398 8392
rect 1454 8336 1459 8392
rect 0 8334 1459 8336
rect 0 8304 800 8334
rect 1393 8331 1459 8334
rect 30005 8394 30071 8397
rect 31200 8394 32000 8424
rect 30005 8392 32000 8394
rect 30005 8336 30010 8392
rect 30066 8336 32000 8392
rect 30005 8334 32000 8336
rect 30005 8331 30071 8334
rect 31200 8304 32000 8334
rect 5909 8192 6229 8193
rect 5909 8128 5917 8192
rect 5981 8128 5997 8192
rect 6061 8128 6077 8192
rect 6141 8128 6157 8192
rect 6221 8128 6229 8192
rect 5909 8127 6229 8128
rect 15840 8192 16160 8193
rect 15840 8128 15848 8192
rect 15912 8128 15928 8192
rect 15992 8128 16008 8192
rect 16072 8128 16088 8192
rect 16152 8128 16160 8192
rect 15840 8127 16160 8128
rect 25770 8192 26090 8193
rect 25770 8128 25778 8192
rect 25842 8128 25858 8192
rect 25922 8128 25938 8192
rect 26002 8128 26018 8192
rect 26082 8128 26090 8192
rect 25770 8127 26090 8128
rect 0 7714 800 7744
rect 1393 7714 1459 7717
rect 0 7712 1459 7714
rect 0 7656 1398 7712
rect 1454 7656 1459 7712
rect 0 7654 1459 7656
rect 0 7624 800 7654
rect 1393 7651 1459 7654
rect 10874 7648 11194 7649
rect 10874 7584 10882 7648
rect 10946 7584 10962 7648
rect 11026 7584 11042 7648
rect 11106 7584 11122 7648
rect 11186 7584 11194 7648
rect 10874 7583 11194 7584
rect 20805 7648 21125 7649
rect 20805 7584 20813 7648
rect 20877 7584 20893 7648
rect 20957 7584 20973 7648
rect 21037 7584 21053 7648
rect 21117 7584 21125 7648
rect 20805 7583 21125 7584
rect 5909 7104 6229 7105
rect 5909 7040 5917 7104
rect 5981 7040 5997 7104
rect 6061 7040 6077 7104
rect 6141 7040 6157 7104
rect 6221 7040 6229 7104
rect 5909 7039 6229 7040
rect 15840 7104 16160 7105
rect 15840 7040 15848 7104
rect 15912 7040 15928 7104
rect 15992 7040 16008 7104
rect 16072 7040 16088 7104
rect 16152 7040 16160 7104
rect 15840 7039 16160 7040
rect 25770 7104 26090 7105
rect 25770 7040 25778 7104
rect 25842 7040 25858 7104
rect 25922 7040 25938 7104
rect 26002 7040 26018 7104
rect 26082 7040 26090 7104
rect 25770 7039 26090 7040
rect 0 6898 800 6928
rect 3969 6898 4035 6901
rect 0 6896 4035 6898
rect 0 6840 3974 6896
rect 4030 6840 4035 6896
rect 0 6838 4035 6840
rect 0 6808 800 6838
rect 3969 6835 4035 6838
rect 30005 6898 30071 6901
rect 31200 6898 32000 6928
rect 30005 6896 32000 6898
rect 30005 6840 30010 6896
rect 30066 6840 32000 6896
rect 30005 6838 32000 6840
rect 30005 6835 30071 6838
rect 31200 6808 32000 6838
rect 10874 6560 11194 6561
rect 10874 6496 10882 6560
rect 10946 6496 10962 6560
rect 11026 6496 11042 6560
rect 11106 6496 11122 6560
rect 11186 6496 11194 6560
rect 10874 6495 11194 6496
rect 20805 6560 21125 6561
rect 20805 6496 20813 6560
rect 20877 6496 20893 6560
rect 20957 6496 20973 6560
rect 21037 6496 21053 6560
rect 21117 6496 21125 6560
rect 20805 6495 21125 6496
rect 0 6218 800 6248
rect 2773 6218 2839 6221
rect 0 6216 2839 6218
rect 0 6160 2778 6216
rect 2834 6160 2839 6216
rect 0 6158 2839 6160
rect 0 6128 800 6158
rect 2773 6155 2839 6158
rect 5909 6016 6229 6017
rect 5909 5952 5917 6016
rect 5981 5952 5997 6016
rect 6061 5952 6077 6016
rect 6141 5952 6157 6016
rect 6221 5952 6229 6016
rect 5909 5951 6229 5952
rect 15840 6016 16160 6017
rect 15840 5952 15848 6016
rect 15912 5952 15928 6016
rect 15992 5952 16008 6016
rect 16072 5952 16088 6016
rect 16152 5952 16160 6016
rect 15840 5951 16160 5952
rect 25770 6016 26090 6017
rect 25770 5952 25778 6016
rect 25842 5952 25858 6016
rect 25922 5952 25938 6016
rect 26002 5952 26018 6016
rect 26082 5952 26090 6016
rect 25770 5951 26090 5952
rect 0 5538 800 5568
rect 1209 5538 1275 5541
rect 0 5536 1275 5538
rect 0 5480 1214 5536
rect 1270 5480 1275 5536
rect 0 5478 1275 5480
rect 0 5448 800 5478
rect 1209 5475 1275 5478
rect 10874 5472 11194 5473
rect 10874 5408 10882 5472
rect 10946 5408 10962 5472
rect 11026 5408 11042 5472
rect 11106 5408 11122 5472
rect 11186 5408 11194 5472
rect 10874 5407 11194 5408
rect 20805 5472 21125 5473
rect 20805 5408 20813 5472
rect 20877 5408 20893 5472
rect 20957 5408 20973 5472
rect 21037 5408 21053 5472
rect 21117 5408 21125 5472
rect 20805 5407 21125 5408
rect 30005 5402 30071 5405
rect 31200 5402 32000 5432
rect 30005 5400 32000 5402
rect 30005 5344 30010 5400
rect 30066 5344 32000 5400
rect 30005 5342 32000 5344
rect 30005 5339 30071 5342
rect 31200 5312 32000 5342
rect 5909 4928 6229 4929
rect 5909 4864 5917 4928
rect 5981 4864 5997 4928
rect 6061 4864 6077 4928
rect 6141 4864 6157 4928
rect 6221 4864 6229 4928
rect 5909 4863 6229 4864
rect 15840 4928 16160 4929
rect 15840 4864 15848 4928
rect 15912 4864 15928 4928
rect 15992 4864 16008 4928
rect 16072 4864 16088 4928
rect 16152 4864 16160 4928
rect 15840 4863 16160 4864
rect 25770 4928 26090 4929
rect 25770 4864 25778 4928
rect 25842 4864 25858 4928
rect 25922 4864 25938 4928
rect 26002 4864 26018 4928
rect 26082 4864 26090 4928
rect 25770 4863 26090 4864
rect 0 4722 800 4752
rect 1393 4722 1459 4725
rect 0 4720 1459 4722
rect 0 4664 1398 4720
rect 1454 4664 1459 4720
rect 0 4662 1459 4664
rect 0 4632 800 4662
rect 1393 4659 1459 4662
rect 10874 4384 11194 4385
rect 10874 4320 10882 4384
rect 10946 4320 10962 4384
rect 11026 4320 11042 4384
rect 11106 4320 11122 4384
rect 11186 4320 11194 4384
rect 10874 4319 11194 4320
rect 20805 4384 21125 4385
rect 20805 4320 20813 4384
rect 20877 4320 20893 4384
rect 20957 4320 20973 4384
rect 21037 4320 21053 4384
rect 21117 4320 21125 4384
rect 20805 4319 21125 4320
rect 0 4042 800 4072
rect 2773 4042 2839 4045
rect 0 4040 2839 4042
rect 0 3984 2778 4040
rect 2834 3984 2839 4040
rect 0 3982 2839 3984
rect 0 3952 800 3982
rect 2773 3979 2839 3982
rect 9070 3980 9076 4044
rect 9140 4042 9146 4044
rect 11881 4042 11947 4045
rect 9140 4040 11947 4042
rect 9140 3984 11886 4040
rect 11942 3984 11947 4040
rect 9140 3982 11947 3984
rect 9140 3980 9146 3982
rect 11881 3979 11947 3982
rect 5909 3840 6229 3841
rect 5909 3776 5917 3840
rect 5981 3776 5997 3840
rect 6061 3776 6077 3840
rect 6141 3776 6157 3840
rect 6221 3776 6229 3840
rect 5909 3775 6229 3776
rect 15840 3840 16160 3841
rect 15840 3776 15848 3840
rect 15912 3776 15928 3840
rect 15992 3776 16008 3840
rect 16072 3776 16088 3840
rect 16152 3776 16160 3840
rect 15840 3775 16160 3776
rect 25770 3840 26090 3841
rect 25770 3776 25778 3840
rect 25842 3776 25858 3840
rect 25922 3776 25938 3840
rect 26002 3776 26018 3840
rect 26082 3776 26090 3840
rect 25770 3775 26090 3776
rect 30005 3770 30071 3773
rect 31200 3770 32000 3800
rect 30005 3768 32000 3770
rect 30005 3712 30010 3768
rect 30066 3712 32000 3768
rect 30005 3710 32000 3712
rect 30005 3707 30071 3710
rect 31200 3680 32000 3710
rect 11973 3498 12039 3501
rect 17217 3498 17283 3501
rect 11973 3496 17283 3498
rect 11973 3440 11978 3496
rect 12034 3440 17222 3496
rect 17278 3440 17283 3496
rect 11973 3438 17283 3440
rect 11973 3435 12039 3438
rect 17217 3435 17283 3438
rect 10874 3296 11194 3297
rect 0 3226 800 3256
rect 10874 3232 10882 3296
rect 10946 3232 10962 3296
rect 11026 3232 11042 3296
rect 11106 3232 11122 3296
rect 11186 3232 11194 3296
rect 10874 3231 11194 3232
rect 20805 3296 21125 3297
rect 20805 3232 20813 3296
rect 20877 3232 20893 3296
rect 20957 3232 20973 3296
rect 21037 3232 21053 3296
rect 21117 3232 21125 3296
rect 20805 3231 21125 3232
rect 2773 3226 2839 3229
rect 0 3224 2839 3226
rect 0 3168 2778 3224
rect 2834 3168 2839 3224
rect 0 3166 2839 3168
rect 0 3136 800 3166
rect 2773 3163 2839 3166
rect 16481 3090 16547 3093
rect 17861 3090 17927 3093
rect 16481 3088 17927 3090
rect 16481 3032 16486 3088
rect 16542 3032 17866 3088
rect 17922 3032 17927 3088
rect 16481 3030 17927 3032
rect 16481 3027 16547 3030
rect 17861 3027 17927 3030
rect 20161 3090 20227 3093
rect 22921 3090 22987 3093
rect 20161 3088 22987 3090
rect 20161 3032 20166 3088
rect 20222 3032 22926 3088
rect 22982 3032 22987 3088
rect 20161 3030 22987 3032
rect 20161 3027 20227 3030
rect 22921 3027 22987 3030
rect 5909 2752 6229 2753
rect 5909 2688 5917 2752
rect 5981 2688 5997 2752
rect 6061 2688 6077 2752
rect 6141 2688 6157 2752
rect 6221 2688 6229 2752
rect 5909 2687 6229 2688
rect 15840 2752 16160 2753
rect 15840 2688 15848 2752
rect 15912 2688 15928 2752
rect 15992 2688 16008 2752
rect 16072 2688 16088 2752
rect 16152 2688 16160 2752
rect 15840 2687 16160 2688
rect 25770 2752 26090 2753
rect 25770 2688 25778 2752
rect 25842 2688 25858 2752
rect 25922 2688 25938 2752
rect 26002 2688 26018 2752
rect 26082 2688 26090 2752
rect 25770 2687 26090 2688
rect 0 2546 800 2576
rect 1853 2546 1919 2549
rect 0 2544 1919 2546
rect 0 2488 1858 2544
rect 1914 2488 1919 2544
rect 0 2486 1919 2488
rect 0 2456 800 2486
rect 1853 2483 1919 2486
rect 30005 2274 30071 2277
rect 31200 2274 32000 2304
rect 30005 2272 32000 2274
rect 30005 2216 30010 2272
rect 30066 2216 32000 2272
rect 30005 2214 32000 2216
rect 30005 2211 30071 2214
rect 10874 2208 11194 2209
rect 10874 2144 10882 2208
rect 10946 2144 10962 2208
rect 11026 2144 11042 2208
rect 11106 2144 11122 2208
rect 11186 2144 11194 2208
rect 10874 2143 11194 2144
rect 20805 2208 21125 2209
rect 20805 2144 20813 2208
rect 20877 2144 20893 2208
rect 20957 2144 20973 2208
rect 21037 2144 21053 2208
rect 21117 2144 21125 2208
rect 31200 2184 32000 2214
rect 20805 2143 21125 2144
rect 0 1730 800 1760
rect 2773 1730 2839 1733
rect 0 1728 2839 1730
rect 0 1672 2778 1728
rect 2834 1672 2839 1728
rect 0 1670 2839 1672
rect 0 1640 800 1670
rect 2773 1667 2839 1670
rect 0 1050 800 1080
rect 2957 1050 3023 1053
rect 0 1048 3023 1050
rect 0 992 2962 1048
rect 3018 992 3023 1048
rect 0 990 3023 992
rect 0 960 800 990
rect 2957 987 3023 990
rect 28901 778 28967 781
rect 31200 778 32000 808
rect 28901 776 32000 778
rect 28901 720 28906 776
rect 28962 720 32000 776
rect 28901 718 32000 720
rect 28901 715 28967 718
rect 31200 688 32000 718
rect 0 370 800 400
rect 2865 370 2931 373
rect 0 368 2931 370
rect 0 312 2870 368
rect 2926 312 2931 368
rect 0 310 2931 312
rect 0 280 800 310
rect 2865 307 2931 310
<< via3 >>
rect 10882 45724 10946 45728
rect 10882 45668 10886 45724
rect 10886 45668 10942 45724
rect 10942 45668 10946 45724
rect 10882 45664 10946 45668
rect 10962 45724 11026 45728
rect 10962 45668 10966 45724
rect 10966 45668 11022 45724
rect 11022 45668 11026 45724
rect 10962 45664 11026 45668
rect 11042 45724 11106 45728
rect 11042 45668 11046 45724
rect 11046 45668 11102 45724
rect 11102 45668 11106 45724
rect 11042 45664 11106 45668
rect 11122 45724 11186 45728
rect 11122 45668 11126 45724
rect 11126 45668 11182 45724
rect 11182 45668 11186 45724
rect 11122 45664 11186 45668
rect 20813 45724 20877 45728
rect 20813 45668 20817 45724
rect 20817 45668 20873 45724
rect 20873 45668 20877 45724
rect 20813 45664 20877 45668
rect 20893 45724 20957 45728
rect 20893 45668 20897 45724
rect 20897 45668 20953 45724
rect 20953 45668 20957 45724
rect 20893 45664 20957 45668
rect 20973 45724 21037 45728
rect 20973 45668 20977 45724
rect 20977 45668 21033 45724
rect 21033 45668 21037 45724
rect 20973 45664 21037 45668
rect 21053 45724 21117 45728
rect 21053 45668 21057 45724
rect 21057 45668 21113 45724
rect 21113 45668 21117 45724
rect 21053 45664 21117 45668
rect 5917 45180 5981 45184
rect 5917 45124 5921 45180
rect 5921 45124 5977 45180
rect 5977 45124 5981 45180
rect 5917 45120 5981 45124
rect 5997 45180 6061 45184
rect 5997 45124 6001 45180
rect 6001 45124 6057 45180
rect 6057 45124 6061 45180
rect 5997 45120 6061 45124
rect 6077 45180 6141 45184
rect 6077 45124 6081 45180
rect 6081 45124 6137 45180
rect 6137 45124 6141 45180
rect 6077 45120 6141 45124
rect 6157 45180 6221 45184
rect 6157 45124 6161 45180
rect 6161 45124 6217 45180
rect 6217 45124 6221 45180
rect 6157 45120 6221 45124
rect 15848 45180 15912 45184
rect 15848 45124 15852 45180
rect 15852 45124 15908 45180
rect 15908 45124 15912 45180
rect 15848 45120 15912 45124
rect 15928 45180 15992 45184
rect 15928 45124 15932 45180
rect 15932 45124 15988 45180
rect 15988 45124 15992 45180
rect 15928 45120 15992 45124
rect 16008 45180 16072 45184
rect 16008 45124 16012 45180
rect 16012 45124 16068 45180
rect 16068 45124 16072 45180
rect 16008 45120 16072 45124
rect 16088 45180 16152 45184
rect 16088 45124 16092 45180
rect 16092 45124 16148 45180
rect 16148 45124 16152 45180
rect 16088 45120 16152 45124
rect 25778 45180 25842 45184
rect 25778 45124 25782 45180
rect 25782 45124 25838 45180
rect 25838 45124 25842 45180
rect 25778 45120 25842 45124
rect 25858 45180 25922 45184
rect 25858 45124 25862 45180
rect 25862 45124 25918 45180
rect 25918 45124 25922 45180
rect 25858 45120 25922 45124
rect 25938 45180 26002 45184
rect 25938 45124 25942 45180
rect 25942 45124 25998 45180
rect 25998 45124 26002 45180
rect 25938 45120 26002 45124
rect 26018 45180 26082 45184
rect 26018 45124 26022 45180
rect 26022 45124 26078 45180
rect 26078 45124 26082 45180
rect 26018 45120 26082 45124
rect 10882 44636 10946 44640
rect 10882 44580 10886 44636
rect 10886 44580 10942 44636
rect 10942 44580 10946 44636
rect 10882 44576 10946 44580
rect 10962 44636 11026 44640
rect 10962 44580 10966 44636
rect 10966 44580 11022 44636
rect 11022 44580 11026 44636
rect 10962 44576 11026 44580
rect 11042 44636 11106 44640
rect 11042 44580 11046 44636
rect 11046 44580 11102 44636
rect 11102 44580 11106 44636
rect 11042 44576 11106 44580
rect 11122 44636 11186 44640
rect 11122 44580 11126 44636
rect 11126 44580 11182 44636
rect 11182 44580 11186 44636
rect 11122 44576 11186 44580
rect 20813 44636 20877 44640
rect 20813 44580 20817 44636
rect 20817 44580 20873 44636
rect 20873 44580 20877 44636
rect 20813 44576 20877 44580
rect 20893 44636 20957 44640
rect 20893 44580 20897 44636
rect 20897 44580 20953 44636
rect 20953 44580 20957 44636
rect 20893 44576 20957 44580
rect 20973 44636 21037 44640
rect 20973 44580 20977 44636
rect 20977 44580 21033 44636
rect 21033 44580 21037 44636
rect 20973 44576 21037 44580
rect 21053 44636 21117 44640
rect 21053 44580 21057 44636
rect 21057 44580 21113 44636
rect 21113 44580 21117 44636
rect 21053 44576 21117 44580
rect 5917 44092 5981 44096
rect 5917 44036 5921 44092
rect 5921 44036 5977 44092
rect 5977 44036 5981 44092
rect 5917 44032 5981 44036
rect 5997 44092 6061 44096
rect 5997 44036 6001 44092
rect 6001 44036 6057 44092
rect 6057 44036 6061 44092
rect 5997 44032 6061 44036
rect 6077 44092 6141 44096
rect 6077 44036 6081 44092
rect 6081 44036 6137 44092
rect 6137 44036 6141 44092
rect 6077 44032 6141 44036
rect 6157 44092 6221 44096
rect 6157 44036 6161 44092
rect 6161 44036 6217 44092
rect 6217 44036 6221 44092
rect 6157 44032 6221 44036
rect 15848 44092 15912 44096
rect 15848 44036 15852 44092
rect 15852 44036 15908 44092
rect 15908 44036 15912 44092
rect 15848 44032 15912 44036
rect 15928 44092 15992 44096
rect 15928 44036 15932 44092
rect 15932 44036 15988 44092
rect 15988 44036 15992 44092
rect 15928 44032 15992 44036
rect 16008 44092 16072 44096
rect 16008 44036 16012 44092
rect 16012 44036 16068 44092
rect 16068 44036 16072 44092
rect 16008 44032 16072 44036
rect 16088 44092 16152 44096
rect 16088 44036 16092 44092
rect 16092 44036 16148 44092
rect 16148 44036 16152 44092
rect 16088 44032 16152 44036
rect 25778 44092 25842 44096
rect 25778 44036 25782 44092
rect 25782 44036 25838 44092
rect 25838 44036 25842 44092
rect 25778 44032 25842 44036
rect 25858 44092 25922 44096
rect 25858 44036 25862 44092
rect 25862 44036 25918 44092
rect 25918 44036 25922 44092
rect 25858 44032 25922 44036
rect 25938 44092 26002 44096
rect 25938 44036 25942 44092
rect 25942 44036 25998 44092
rect 25998 44036 26002 44092
rect 25938 44032 26002 44036
rect 26018 44092 26082 44096
rect 26018 44036 26022 44092
rect 26022 44036 26078 44092
rect 26078 44036 26082 44092
rect 26018 44032 26082 44036
rect 10882 43548 10946 43552
rect 10882 43492 10886 43548
rect 10886 43492 10942 43548
rect 10942 43492 10946 43548
rect 10882 43488 10946 43492
rect 10962 43548 11026 43552
rect 10962 43492 10966 43548
rect 10966 43492 11022 43548
rect 11022 43492 11026 43548
rect 10962 43488 11026 43492
rect 11042 43548 11106 43552
rect 11042 43492 11046 43548
rect 11046 43492 11102 43548
rect 11102 43492 11106 43548
rect 11042 43488 11106 43492
rect 11122 43548 11186 43552
rect 11122 43492 11126 43548
rect 11126 43492 11182 43548
rect 11182 43492 11186 43548
rect 11122 43488 11186 43492
rect 20813 43548 20877 43552
rect 20813 43492 20817 43548
rect 20817 43492 20873 43548
rect 20873 43492 20877 43548
rect 20813 43488 20877 43492
rect 20893 43548 20957 43552
rect 20893 43492 20897 43548
rect 20897 43492 20953 43548
rect 20953 43492 20957 43548
rect 20893 43488 20957 43492
rect 20973 43548 21037 43552
rect 20973 43492 20977 43548
rect 20977 43492 21033 43548
rect 21033 43492 21037 43548
rect 20973 43488 21037 43492
rect 21053 43548 21117 43552
rect 21053 43492 21057 43548
rect 21057 43492 21113 43548
rect 21113 43492 21117 43548
rect 21053 43488 21117 43492
rect 5917 43004 5981 43008
rect 5917 42948 5921 43004
rect 5921 42948 5977 43004
rect 5977 42948 5981 43004
rect 5917 42944 5981 42948
rect 5997 43004 6061 43008
rect 5997 42948 6001 43004
rect 6001 42948 6057 43004
rect 6057 42948 6061 43004
rect 5997 42944 6061 42948
rect 6077 43004 6141 43008
rect 6077 42948 6081 43004
rect 6081 42948 6137 43004
rect 6137 42948 6141 43004
rect 6077 42944 6141 42948
rect 6157 43004 6221 43008
rect 6157 42948 6161 43004
rect 6161 42948 6217 43004
rect 6217 42948 6221 43004
rect 6157 42944 6221 42948
rect 15848 43004 15912 43008
rect 15848 42948 15852 43004
rect 15852 42948 15908 43004
rect 15908 42948 15912 43004
rect 15848 42944 15912 42948
rect 15928 43004 15992 43008
rect 15928 42948 15932 43004
rect 15932 42948 15988 43004
rect 15988 42948 15992 43004
rect 15928 42944 15992 42948
rect 16008 43004 16072 43008
rect 16008 42948 16012 43004
rect 16012 42948 16068 43004
rect 16068 42948 16072 43004
rect 16008 42944 16072 42948
rect 16088 43004 16152 43008
rect 16088 42948 16092 43004
rect 16092 42948 16148 43004
rect 16148 42948 16152 43004
rect 16088 42944 16152 42948
rect 25778 43004 25842 43008
rect 25778 42948 25782 43004
rect 25782 42948 25838 43004
rect 25838 42948 25842 43004
rect 25778 42944 25842 42948
rect 25858 43004 25922 43008
rect 25858 42948 25862 43004
rect 25862 42948 25918 43004
rect 25918 42948 25922 43004
rect 25858 42944 25922 42948
rect 25938 43004 26002 43008
rect 25938 42948 25942 43004
rect 25942 42948 25998 43004
rect 25998 42948 26002 43004
rect 25938 42944 26002 42948
rect 26018 43004 26082 43008
rect 26018 42948 26022 43004
rect 26022 42948 26078 43004
rect 26078 42948 26082 43004
rect 26018 42944 26082 42948
rect 10882 42460 10946 42464
rect 10882 42404 10886 42460
rect 10886 42404 10942 42460
rect 10942 42404 10946 42460
rect 10882 42400 10946 42404
rect 10962 42460 11026 42464
rect 10962 42404 10966 42460
rect 10966 42404 11022 42460
rect 11022 42404 11026 42460
rect 10962 42400 11026 42404
rect 11042 42460 11106 42464
rect 11042 42404 11046 42460
rect 11046 42404 11102 42460
rect 11102 42404 11106 42460
rect 11042 42400 11106 42404
rect 11122 42460 11186 42464
rect 11122 42404 11126 42460
rect 11126 42404 11182 42460
rect 11182 42404 11186 42460
rect 11122 42400 11186 42404
rect 20813 42460 20877 42464
rect 20813 42404 20817 42460
rect 20817 42404 20873 42460
rect 20873 42404 20877 42460
rect 20813 42400 20877 42404
rect 20893 42460 20957 42464
rect 20893 42404 20897 42460
rect 20897 42404 20953 42460
rect 20953 42404 20957 42460
rect 20893 42400 20957 42404
rect 20973 42460 21037 42464
rect 20973 42404 20977 42460
rect 20977 42404 21033 42460
rect 21033 42404 21037 42460
rect 20973 42400 21037 42404
rect 21053 42460 21117 42464
rect 21053 42404 21057 42460
rect 21057 42404 21113 42460
rect 21113 42404 21117 42460
rect 21053 42400 21117 42404
rect 5917 41916 5981 41920
rect 5917 41860 5921 41916
rect 5921 41860 5977 41916
rect 5977 41860 5981 41916
rect 5917 41856 5981 41860
rect 5997 41916 6061 41920
rect 5997 41860 6001 41916
rect 6001 41860 6057 41916
rect 6057 41860 6061 41916
rect 5997 41856 6061 41860
rect 6077 41916 6141 41920
rect 6077 41860 6081 41916
rect 6081 41860 6137 41916
rect 6137 41860 6141 41916
rect 6077 41856 6141 41860
rect 6157 41916 6221 41920
rect 6157 41860 6161 41916
rect 6161 41860 6217 41916
rect 6217 41860 6221 41916
rect 6157 41856 6221 41860
rect 15848 41916 15912 41920
rect 15848 41860 15852 41916
rect 15852 41860 15908 41916
rect 15908 41860 15912 41916
rect 15848 41856 15912 41860
rect 15928 41916 15992 41920
rect 15928 41860 15932 41916
rect 15932 41860 15988 41916
rect 15988 41860 15992 41916
rect 15928 41856 15992 41860
rect 16008 41916 16072 41920
rect 16008 41860 16012 41916
rect 16012 41860 16068 41916
rect 16068 41860 16072 41916
rect 16008 41856 16072 41860
rect 16088 41916 16152 41920
rect 16088 41860 16092 41916
rect 16092 41860 16148 41916
rect 16148 41860 16152 41916
rect 16088 41856 16152 41860
rect 25778 41916 25842 41920
rect 25778 41860 25782 41916
rect 25782 41860 25838 41916
rect 25838 41860 25842 41916
rect 25778 41856 25842 41860
rect 25858 41916 25922 41920
rect 25858 41860 25862 41916
rect 25862 41860 25918 41916
rect 25918 41860 25922 41916
rect 25858 41856 25922 41860
rect 25938 41916 26002 41920
rect 25938 41860 25942 41916
rect 25942 41860 25998 41916
rect 25998 41860 26002 41916
rect 25938 41856 26002 41860
rect 26018 41916 26082 41920
rect 26018 41860 26022 41916
rect 26022 41860 26078 41916
rect 26078 41860 26082 41916
rect 26018 41856 26082 41860
rect 10882 41372 10946 41376
rect 10882 41316 10886 41372
rect 10886 41316 10942 41372
rect 10942 41316 10946 41372
rect 10882 41312 10946 41316
rect 10962 41372 11026 41376
rect 10962 41316 10966 41372
rect 10966 41316 11022 41372
rect 11022 41316 11026 41372
rect 10962 41312 11026 41316
rect 11042 41372 11106 41376
rect 11042 41316 11046 41372
rect 11046 41316 11102 41372
rect 11102 41316 11106 41372
rect 11042 41312 11106 41316
rect 11122 41372 11186 41376
rect 11122 41316 11126 41372
rect 11126 41316 11182 41372
rect 11182 41316 11186 41372
rect 11122 41312 11186 41316
rect 20813 41372 20877 41376
rect 20813 41316 20817 41372
rect 20817 41316 20873 41372
rect 20873 41316 20877 41372
rect 20813 41312 20877 41316
rect 20893 41372 20957 41376
rect 20893 41316 20897 41372
rect 20897 41316 20953 41372
rect 20953 41316 20957 41372
rect 20893 41312 20957 41316
rect 20973 41372 21037 41376
rect 20973 41316 20977 41372
rect 20977 41316 21033 41372
rect 21033 41316 21037 41372
rect 20973 41312 21037 41316
rect 21053 41372 21117 41376
rect 21053 41316 21057 41372
rect 21057 41316 21113 41372
rect 21113 41316 21117 41372
rect 21053 41312 21117 41316
rect 5917 40828 5981 40832
rect 5917 40772 5921 40828
rect 5921 40772 5977 40828
rect 5977 40772 5981 40828
rect 5917 40768 5981 40772
rect 5997 40828 6061 40832
rect 5997 40772 6001 40828
rect 6001 40772 6057 40828
rect 6057 40772 6061 40828
rect 5997 40768 6061 40772
rect 6077 40828 6141 40832
rect 6077 40772 6081 40828
rect 6081 40772 6137 40828
rect 6137 40772 6141 40828
rect 6077 40768 6141 40772
rect 6157 40828 6221 40832
rect 6157 40772 6161 40828
rect 6161 40772 6217 40828
rect 6217 40772 6221 40828
rect 6157 40768 6221 40772
rect 15848 40828 15912 40832
rect 15848 40772 15852 40828
rect 15852 40772 15908 40828
rect 15908 40772 15912 40828
rect 15848 40768 15912 40772
rect 15928 40828 15992 40832
rect 15928 40772 15932 40828
rect 15932 40772 15988 40828
rect 15988 40772 15992 40828
rect 15928 40768 15992 40772
rect 16008 40828 16072 40832
rect 16008 40772 16012 40828
rect 16012 40772 16068 40828
rect 16068 40772 16072 40828
rect 16008 40768 16072 40772
rect 16088 40828 16152 40832
rect 16088 40772 16092 40828
rect 16092 40772 16148 40828
rect 16148 40772 16152 40828
rect 16088 40768 16152 40772
rect 25778 40828 25842 40832
rect 25778 40772 25782 40828
rect 25782 40772 25838 40828
rect 25838 40772 25842 40828
rect 25778 40768 25842 40772
rect 25858 40828 25922 40832
rect 25858 40772 25862 40828
rect 25862 40772 25918 40828
rect 25918 40772 25922 40828
rect 25858 40768 25922 40772
rect 25938 40828 26002 40832
rect 25938 40772 25942 40828
rect 25942 40772 25998 40828
rect 25998 40772 26002 40828
rect 25938 40768 26002 40772
rect 26018 40828 26082 40832
rect 26018 40772 26022 40828
rect 26022 40772 26078 40828
rect 26078 40772 26082 40828
rect 26018 40768 26082 40772
rect 10882 40284 10946 40288
rect 10882 40228 10886 40284
rect 10886 40228 10942 40284
rect 10942 40228 10946 40284
rect 10882 40224 10946 40228
rect 10962 40284 11026 40288
rect 10962 40228 10966 40284
rect 10966 40228 11022 40284
rect 11022 40228 11026 40284
rect 10962 40224 11026 40228
rect 11042 40284 11106 40288
rect 11042 40228 11046 40284
rect 11046 40228 11102 40284
rect 11102 40228 11106 40284
rect 11042 40224 11106 40228
rect 11122 40284 11186 40288
rect 11122 40228 11126 40284
rect 11126 40228 11182 40284
rect 11182 40228 11186 40284
rect 11122 40224 11186 40228
rect 20813 40284 20877 40288
rect 20813 40228 20817 40284
rect 20817 40228 20873 40284
rect 20873 40228 20877 40284
rect 20813 40224 20877 40228
rect 20893 40284 20957 40288
rect 20893 40228 20897 40284
rect 20897 40228 20953 40284
rect 20953 40228 20957 40284
rect 20893 40224 20957 40228
rect 20973 40284 21037 40288
rect 20973 40228 20977 40284
rect 20977 40228 21033 40284
rect 21033 40228 21037 40284
rect 20973 40224 21037 40228
rect 21053 40284 21117 40288
rect 21053 40228 21057 40284
rect 21057 40228 21113 40284
rect 21113 40228 21117 40284
rect 21053 40224 21117 40228
rect 5917 39740 5981 39744
rect 5917 39684 5921 39740
rect 5921 39684 5977 39740
rect 5977 39684 5981 39740
rect 5917 39680 5981 39684
rect 5997 39740 6061 39744
rect 5997 39684 6001 39740
rect 6001 39684 6057 39740
rect 6057 39684 6061 39740
rect 5997 39680 6061 39684
rect 6077 39740 6141 39744
rect 6077 39684 6081 39740
rect 6081 39684 6137 39740
rect 6137 39684 6141 39740
rect 6077 39680 6141 39684
rect 6157 39740 6221 39744
rect 6157 39684 6161 39740
rect 6161 39684 6217 39740
rect 6217 39684 6221 39740
rect 6157 39680 6221 39684
rect 15848 39740 15912 39744
rect 15848 39684 15852 39740
rect 15852 39684 15908 39740
rect 15908 39684 15912 39740
rect 15848 39680 15912 39684
rect 15928 39740 15992 39744
rect 15928 39684 15932 39740
rect 15932 39684 15988 39740
rect 15988 39684 15992 39740
rect 15928 39680 15992 39684
rect 16008 39740 16072 39744
rect 16008 39684 16012 39740
rect 16012 39684 16068 39740
rect 16068 39684 16072 39740
rect 16008 39680 16072 39684
rect 16088 39740 16152 39744
rect 16088 39684 16092 39740
rect 16092 39684 16148 39740
rect 16148 39684 16152 39740
rect 16088 39680 16152 39684
rect 25778 39740 25842 39744
rect 25778 39684 25782 39740
rect 25782 39684 25838 39740
rect 25838 39684 25842 39740
rect 25778 39680 25842 39684
rect 25858 39740 25922 39744
rect 25858 39684 25862 39740
rect 25862 39684 25918 39740
rect 25918 39684 25922 39740
rect 25858 39680 25922 39684
rect 25938 39740 26002 39744
rect 25938 39684 25942 39740
rect 25942 39684 25998 39740
rect 25998 39684 26002 39740
rect 25938 39680 26002 39684
rect 26018 39740 26082 39744
rect 26018 39684 26022 39740
rect 26022 39684 26078 39740
rect 26078 39684 26082 39740
rect 26018 39680 26082 39684
rect 10882 39196 10946 39200
rect 10882 39140 10886 39196
rect 10886 39140 10942 39196
rect 10942 39140 10946 39196
rect 10882 39136 10946 39140
rect 10962 39196 11026 39200
rect 10962 39140 10966 39196
rect 10966 39140 11022 39196
rect 11022 39140 11026 39196
rect 10962 39136 11026 39140
rect 11042 39196 11106 39200
rect 11042 39140 11046 39196
rect 11046 39140 11102 39196
rect 11102 39140 11106 39196
rect 11042 39136 11106 39140
rect 11122 39196 11186 39200
rect 11122 39140 11126 39196
rect 11126 39140 11182 39196
rect 11182 39140 11186 39196
rect 11122 39136 11186 39140
rect 20813 39196 20877 39200
rect 20813 39140 20817 39196
rect 20817 39140 20873 39196
rect 20873 39140 20877 39196
rect 20813 39136 20877 39140
rect 20893 39196 20957 39200
rect 20893 39140 20897 39196
rect 20897 39140 20953 39196
rect 20953 39140 20957 39196
rect 20893 39136 20957 39140
rect 20973 39196 21037 39200
rect 20973 39140 20977 39196
rect 20977 39140 21033 39196
rect 21033 39140 21037 39196
rect 20973 39136 21037 39140
rect 21053 39196 21117 39200
rect 21053 39140 21057 39196
rect 21057 39140 21113 39196
rect 21113 39140 21117 39196
rect 21053 39136 21117 39140
rect 5917 38652 5981 38656
rect 5917 38596 5921 38652
rect 5921 38596 5977 38652
rect 5977 38596 5981 38652
rect 5917 38592 5981 38596
rect 5997 38652 6061 38656
rect 5997 38596 6001 38652
rect 6001 38596 6057 38652
rect 6057 38596 6061 38652
rect 5997 38592 6061 38596
rect 6077 38652 6141 38656
rect 6077 38596 6081 38652
rect 6081 38596 6137 38652
rect 6137 38596 6141 38652
rect 6077 38592 6141 38596
rect 6157 38652 6221 38656
rect 6157 38596 6161 38652
rect 6161 38596 6217 38652
rect 6217 38596 6221 38652
rect 6157 38592 6221 38596
rect 15848 38652 15912 38656
rect 15848 38596 15852 38652
rect 15852 38596 15908 38652
rect 15908 38596 15912 38652
rect 15848 38592 15912 38596
rect 15928 38652 15992 38656
rect 15928 38596 15932 38652
rect 15932 38596 15988 38652
rect 15988 38596 15992 38652
rect 15928 38592 15992 38596
rect 16008 38652 16072 38656
rect 16008 38596 16012 38652
rect 16012 38596 16068 38652
rect 16068 38596 16072 38652
rect 16008 38592 16072 38596
rect 16088 38652 16152 38656
rect 16088 38596 16092 38652
rect 16092 38596 16148 38652
rect 16148 38596 16152 38652
rect 16088 38592 16152 38596
rect 25778 38652 25842 38656
rect 25778 38596 25782 38652
rect 25782 38596 25838 38652
rect 25838 38596 25842 38652
rect 25778 38592 25842 38596
rect 25858 38652 25922 38656
rect 25858 38596 25862 38652
rect 25862 38596 25918 38652
rect 25918 38596 25922 38652
rect 25858 38592 25922 38596
rect 25938 38652 26002 38656
rect 25938 38596 25942 38652
rect 25942 38596 25998 38652
rect 25998 38596 26002 38652
rect 25938 38592 26002 38596
rect 26018 38652 26082 38656
rect 26018 38596 26022 38652
rect 26022 38596 26078 38652
rect 26078 38596 26082 38652
rect 26018 38592 26082 38596
rect 10882 38108 10946 38112
rect 10882 38052 10886 38108
rect 10886 38052 10942 38108
rect 10942 38052 10946 38108
rect 10882 38048 10946 38052
rect 10962 38108 11026 38112
rect 10962 38052 10966 38108
rect 10966 38052 11022 38108
rect 11022 38052 11026 38108
rect 10962 38048 11026 38052
rect 11042 38108 11106 38112
rect 11042 38052 11046 38108
rect 11046 38052 11102 38108
rect 11102 38052 11106 38108
rect 11042 38048 11106 38052
rect 11122 38108 11186 38112
rect 11122 38052 11126 38108
rect 11126 38052 11182 38108
rect 11182 38052 11186 38108
rect 11122 38048 11186 38052
rect 20813 38108 20877 38112
rect 20813 38052 20817 38108
rect 20817 38052 20873 38108
rect 20873 38052 20877 38108
rect 20813 38048 20877 38052
rect 20893 38108 20957 38112
rect 20893 38052 20897 38108
rect 20897 38052 20953 38108
rect 20953 38052 20957 38108
rect 20893 38048 20957 38052
rect 20973 38108 21037 38112
rect 20973 38052 20977 38108
rect 20977 38052 21033 38108
rect 21033 38052 21037 38108
rect 20973 38048 21037 38052
rect 21053 38108 21117 38112
rect 21053 38052 21057 38108
rect 21057 38052 21113 38108
rect 21113 38052 21117 38108
rect 21053 38048 21117 38052
rect 5917 37564 5981 37568
rect 5917 37508 5921 37564
rect 5921 37508 5977 37564
rect 5977 37508 5981 37564
rect 5917 37504 5981 37508
rect 5997 37564 6061 37568
rect 5997 37508 6001 37564
rect 6001 37508 6057 37564
rect 6057 37508 6061 37564
rect 5997 37504 6061 37508
rect 6077 37564 6141 37568
rect 6077 37508 6081 37564
rect 6081 37508 6137 37564
rect 6137 37508 6141 37564
rect 6077 37504 6141 37508
rect 6157 37564 6221 37568
rect 6157 37508 6161 37564
rect 6161 37508 6217 37564
rect 6217 37508 6221 37564
rect 6157 37504 6221 37508
rect 15848 37564 15912 37568
rect 15848 37508 15852 37564
rect 15852 37508 15908 37564
rect 15908 37508 15912 37564
rect 15848 37504 15912 37508
rect 15928 37564 15992 37568
rect 15928 37508 15932 37564
rect 15932 37508 15988 37564
rect 15988 37508 15992 37564
rect 15928 37504 15992 37508
rect 16008 37564 16072 37568
rect 16008 37508 16012 37564
rect 16012 37508 16068 37564
rect 16068 37508 16072 37564
rect 16008 37504 16072 37508
rect 16088 37564 16152 37568
rect 16088 37508 16092 37564
rect 16092 37508 16148 37564
rect 16148 37508 16152 37564
rect 16088 37504 16152 37508
rect 25778 37564 25842 37568
rect 25778 37508 25782 37564
rect 25782 37508 25838 37564
rect 25838 37508 25842 37564
rect 25778 37504 25842 37508
rect 25858 37564 25922 37568
rect 25858 37508 25862 37564
rect 25862 37508 25918 37564
rect 25918 37508 25922 37564
rect 25858 37504 25922 37508
rect 25938 37564 26002 37568
rect 25938 37508 25942 37564
rect 25942 37508 25998 37564
rect 25998 37508 26002 37564
rect 25938 37504 26002 37508
rect 26018 37564 26082 37568
rect 26018 37508 26022 37564
rect 26022 37508 26078 37564
rect 26078 37508 26082 37564
rect 26018 37504 26082 37508
rect 10882 37020 10946 37024
rect 10882 36964 10886 37020
rect 10886 36964 10942 37020
rect 10942 36964 10946 37020
rect 10882 36960 10946 36964
rect 10962 37020 11026 37024
rect 10962 36964 10966 37020
rect 10966 36964 11022 37020
rect 11022 36964 11026 37020
rect 10962 36960 11026 36964
rect 11042 37020 11106 37024
rect 11042 36964 11046 37020
rect 11046 36964 11102 37020
rect 11102 36964 11106 37020
rect 11042 36960 11106 36964
rect 11122 37020 11186 37024
rect 11122 36964 11126 37020
rect 11126 36964 11182 37020
rect 11182 36964 11186 37020
rect 11122 36960 11186 36964
rect 20813 37020 20877 37024
rect 20813 36964 20817 37020
rect 20817 36964 20873 37020
rect 20873 36964 20877 37020
rect 20813 36960 20877 36964
rect 20893 37020 20957 37024
rect 20893 36964 20897 37020
rect 20897 36964 20953 37020
rect 20953 36964 20957 37020
rect 20893 36960 20957 36964
rect 20973 37020 21037 37024
rect 20973 36964 20977 37020
rect 20977 36964 21033 37020
rect 21033 36964 21037 37020
rect 20973 36960 21037 36964
rect 21053 37020 21117 37024
rect 21053 36964 21057 37020
rect 21057 36964 21113 37020
rect 21113 36964 21117 37020
rect 21053 36960 21117 36964
rect 5917 36476 5981 36480
rect 5917 36420 5921 36476
rect 5921 36420 5977 36476
rect 5977 36420 5981 36476
rect 5917 36416 5981 36420
rect 5997 36476 6061 36480
rect 5997 36420 6001 36476
rect 6001 36420 6057 36476
rect 6057 36420 6061 36476
rect 5997 36416 6061 36420
rect 6077 36476 6141 36480
rect 6077 36420 6081 36476
rect 6081 36420 6137 36476
rect 6137 36420 6141 36476
rect 6077 36416 6141 36420
rect 6157 36476 6221 36480
rect 6157 36420 6161 36476
rect 6161 36420 6217 36476
rect 6217 36420 6221 36476
rect 6157 36416 6221 36420
rect 15848 36476 15912 36480
rect 15848 36420 15852 36476
rect 15852 36420 15908 36476
rect 15908 36420 15912 36476
rect 15848 36416 15912 36420
rect 15928 36476 15992 36480
rect 15928 36420 15932 36476
rect 15932 36420 15988 36476
rect 15988 36420 15992 36476
rect 15928 36416 15992 36420
rect 16008 36476 16072 36480
rect 16008 36420 16012 36476
rect 16012 36420 16068 36476
rect 16068 36420 16072 36476
rect 16008 36416 16072 36420
rect 16088 36476 16152 36480
rect 16088 36420 16092 36476
rect 16092 36420 16148 36476
rect 16148 36420 16152 36476
rect 16088 36416 16152 36420
rect 25778 36476 25842 36480
rect 25778 36420 25782 36476
rect 25782 36420 25838 36476
rect 25838 36420 25842 36476
rect 25778 36416 25842 36420
rect 25858 36476 25922 36480
rect 25858 36420 25862 36476
rect 25862 36420 25918 36476
rect 25918 36420 25922 36476
rect 25858 36416 25922 36420
rect 25938 36476 26002 36480
rect 25938 36420 25942 36476
rect 25942 36420 25998 36476
rect 25998 36420 26002 36476
rect 25938 36416 26002 36420
rect 26018 36476 26082 36480
rect 26018 36420 26022 36476
rect 26022 36420 26078 36476
rect 26078 36420 26082 36476
rect 26018 36416 26082 36420
rect 10882 35932 10946 35936
rect 10882 35876 10886 35932
rect 10886 35876 10942 35932
rect 10942 35876 10946 35932
rect 10882 35872 10946 35876
rect 10962 35932 11026 35936
rect 10962 35876 10966 35932
rect 10966 35876 11022 35932
rect 11022 35876 11026 35932
rect 10962 35872 11026 35876
rect 11042 35932 11106 35936
rect 11042 35876 11046 35932
rect 11046 35876 11102 35932
rect 11102 35876 11106 35932
rect 11042 35872 11106 35876
rect 11122 35932 11186 35936
rect 11122 35876 11126 35932
rect 11126 35876 11182 35932
rect 11182 35876 11186 35932
rect 11122 35872 11186 35876
rect 20813 35932 20877 35936
rect 20813 35876 20817 35932
rect 20817 35876 20873 35932
rect 20873 35876 20877 35932
rect 20813 35872 20877 35876
rect 20893 35932 20957 35936
rect 20893 35876 20897 35932
rect 20897 35876 20953 35932
rect 20953 35876 20957 35932
rect 20893 35872 20957 35876
rect 20973 35932 21037 35936
rect 20973 35876 20977 35932
rect 20977 35876 21033 35932
rect 21033 35876 21037 35932
rect 20973 35872 21037 35876
rect 21053 35932 21117 35936
rect 21053 35876 21057 35932
rect 21057 35876 21113 35932
rect 21113 35876 21117 35932
rect 21053 35872 21117 35876
rect 5917 35388 5981 35392
rect 5917 35332 5921 35388
rect 5921 35332 5977 35388
rect 5977 35332 5981 35388
rect 5917 35328 5981 35332
rect 5997 35388 6061 35392
rect 5997 35332 6001 35388
rect 6001 35332 6057 35388
rect 6057 35332 6061 35388
rect 5997 35328 6061 35332
rect 6077 35388 6141 35392
rect 6077 35332 6081 35388
rect 6081 35332 6137 35388
rect 6137 35332 6141 35388
rect 6077 35328 6141 35332
rect 6157 35388 6221 35392
rect 6157 35332 6161 35388
rect 6161 35332 6217 35388
rect 6217 35332 6221 35388
rect 6157 35328 6221 35332
rect 15848 35388 15912 35392
rect 15848 35332 15852 35388
rect 15852 35332 15908 35388
rect 15908 35332 15912 35388
rect 15848 35328 15912 35332
rect 15928 35388 15992 35392
rect 15928 35332 15932 35388
rect 15932 35332 15988 35388
rect 15988 35332 15992 35388
rect 15928 35328 15992 35332
rect 16008 35388 16072 35392
rect 16008 35332 16012 35388
rect 16012 35332 16068 35388
rect 16068 35332 16072 35388
rect 16008 35328 16072 35332
rect 16088 35388 16152 35392
rect 16088 35332 16092 35388
rect 16092 35332 16148 35388
rect 16148 35332 16152 35388
rect 16088 35328 16152 35332
rect 25778 35388 25842 35392
rect 25778 35332 25782 35388
rect 25782 35332 25838 35388
rect 25838 35332 25842 35388
rect 25778 35328 25842 35332
rect 25858 35388 25922 35392
rect 25858 35332 25862 35388
rect 25862 35332 25918 35388
rect 25918 35332 25922 35388
rect 25858 35328 25922 35332
rect 25938 35388 26002 35392
rect 25938 35332 25942 35388
rect 25942 35332 25998 35388
rect 25998 35332 26002 35388
rect 25938 35328 26002 35332
rect 26018 35388 26082 35392
rect 26018 35332 26022 35388
rect 26022 35332 26078 35388
rect 26078 35332 26082 35388
rect 26018 35328 26082 35332
rect 10882 34844 10946 34848
rect 10882 34788 10886 34844
rect 10886 34788 10942 34844
rect 10942 34788 10946 34844
rect 10882 34784 10946 34788
rect 10962 34844 11026 34848
rect 10962 34788 10966 34844
rect 10966 34788 11022 34844
rect 11022 34788 11026 34844
rect 10962 34784 11026 34788
rect 11042 34844 11106 34848
rect 11042 34788 11046 34844
rect 11046 34788 11102 34844
rect 11102 34788 11106 34844
rect 11042 34784 11106 34788
rect 11122 34844 11186 34848
rect 11122 34788 11126 34844
rect 11126 34788 11182 34844
rect 11182 34788 11186 34844
rect 11122 34784 11186 34788
rect 20813 34844 20877 34848
rect 20813 34788 20817 34844
rect 20817 34788 20873 34844
rect 20873 34788 20877 34844
rect 20813 34784 20877 34788
rect 20893 34844 20957 34848
rect 20893 34788 20897 34844
rect 20897 34788 20953 34844
rect 20953 34788 20957 34844
rect 20893 34784 20957 34788
rect 20973 34844 21037 34848
rect 20973 34788 20977 34844
rect 20977 34788 21033 34844
rect 21033 34788 21037 34844
rect 20973 34784 21037 34788
rect 21053 34844 21117 34848
rect 21053 34788 21057 34844
rect 21057 34788 21113 34844
rect 21113 34788 21117 34844
rect 21053 34784 21117 34788
rect 5917 34300 5981 34304
rect 5917 34244 5921 34300
rect 5921 34244 5977 34300
rect 5977 34244 5981 34300
rect 5917 34240 5981 34244
rect 5997 34300 6061 34304
rect 5997 34244 6001 34300
rect 6001 34244 6057 34300
rect 6057 34244 6061 34300
rect 5997 34240 6061 34244
rect 6077 34300 6141 34304
rect 6077 34244 6081 34300
rect 6081 34244 6137 34300
rect 6137 34244 6141 34300
rect 6077 34240 6141 34244
rect 6157 34300 6221 34304
rect 6157 34244 6161 34300
rect 6161 34244 6217 34300
rect 6217 34244 6221 34300
rect 6157 34240 6221 34244
rect 15848 34300 15912 34304
rect 15848 34244 15852 34300
rect 15852 34244 15908 34300
rect 15908 34244 15912 34300
rect 15848 34240 15912 34244
rect 15928 34300 15992 34304
rect 15928 34244 15932 34300
rect 15932 34244 15988 34300
rect 15988 34244 15992 34300
rect 15928 34240 15992 34244
rect 16008 34300 16072 34304
rect 16008 34244 16012 34300
rect 16012 34244 16068 34300
rect 16068 34244 16072 34300
rect 16008 34240 16072 34244
rect 16088 34300 16152 34304
rect 16088 34244 16092 34300
rect 16092 34244 16148 34300
rect 16148 34244 16152 34300
rect 16088 34240 16152 34244
rect 25778 34300 25842 34304
rect 25778 34244 25782 34300
rect 25782 34244 25838 34300
rect 25838 34244 25842 34300
rect 25778 34240 25842 34244
rect 25858 34300 25922 34304
rect 25858 34244 25862 34300
rect 25862 34244 25918 34300
rect 25918 34244 25922 34300
rect 25858 34240 25922 34244
rect 25938 34300 26002 34304
rect 25938 34244 25942 34300
rect 25942 34244 25998 34300
rect 25998 34244 26002 34300
rect 25938 34240 26002 34244
rect 26018 34300 26082 34304
rect 26018 34244 26022 34300
rect 26022 34244 26078 34300
rect 26078 34244 26082 34300
rect 26018 34240 26082 34244
rect 10882 33756 10946 33760
rect 10882 33700 10886 33756
rect 10886 33700 10942 33756
rect 10942 33700 10946 33756
rect 10882 33696 10946 33700
rect 10962 33756 11026 33760
rect 10962 33700 10966 33756
rect 10966 33700 11022 33756
rect 11022 33700 11026 33756
rect 10962 33696 11026 33700
rect 11042 33756 11106 33760
rect 11042 33700 11046 33756
rect 11046 33700 11102 33756
rect 11102 33700 11106 33756
rect 11042 33696 11106 33700
rect 11122 33756 11186 33760
rect 11122 33700 11126 33756
rect 11126 33700 11182 33756
rect 11182 33700 11186 33756
rect 11122 33696 11186 33700
rect 20813 33756 20877 33760
rect 20813 33700 20817 33756
rect 20817 33700 20873 33756
rect 20873 33700 20877 33756
rect 20813 33696 20877 33700
rect 20893 33756 20957 33760
rect 20893 33700 20897 33756
rect 20897 33700 20953 33756
rect 20953 33700 20957 33756
rect 20893 33696 20957 33700
rect 20973 33756 21037 33760
rect 20973 33700 20977 33756
rect 20977 33700 21033 33756
rect 21033 33700 21037 33756
rect 20973 33696 21037 33700
rect 21053 33756 21117 33760
rect 21053 33700 21057 33756
rect 21057 33700 21113 33756
rect 21113 33700 21117 33756
rect 21053 33696 21117 33700
rect 5917 33212 5981 33216
rect 5917 33156 5921 33212
rect 5921 33156 5977 33212
rect 5977 33156 5981 33212
rect 5917 33152 5981 33156
rect 5997 33212 6061 33216
rect 5997 33156 6001 33212
rect 6001 33156 6057 33212
rect 6057 33156 6061 33212
rect 5997 33152 6061 33156
rect 6077 33212 6141 33216
rect 6077 33156 6081 33212
rect 6081 33156 6137 33212
rect 6137 33156 6141 33212
rect 6077 33152 6141 33156
rect 6157 33212 6221 33216
rect 6157 33156 6161 33212
rect 6161 33156 6217 33212
rect 6217 33156 6221 33212
rect 6157 33152 6221 33156
rect 15848 33212 15912 33216
rect 15848 33156 15852 33212
rect 15852 33156 15908 33212
rect 15908 33156 15912 33212
rect 15848 33152 15912 33156
rect 15928 33212 15992 33216
rect 15928 33156 15932 33212
rect 15932 33156 15988 33212
rect 15988 33156 15992 33212
rect 15928 33152 15992 33156
rect 16008 33212 16072 33216
rect 16008 33156 16012 33212
rect 16012 33156 16068 33212
rect 16068 33156 16072 33212
rect 16008 33152 16072 33156
rect 16088 33212 16152 33216
rect 16088 33156 16092 33212
rect 16092 33156 16148 33212
rect 16148 33156 16152 33212
rect 16088 33152 16152 33156
rect 25778 33212 25842 33216
rect 25778 33156 25782 33212
rect 25782 33156 25838 33212
rect 25838 33156 25842 33212
rect 25778 33152 25842 33156
rect 25858 33212 25922 33216
rect 25858 33156 25862 33212
rect 25862 33156 25918 33212
rect 25918 33156 25922 33212
rect 25858 33152 25922 33156
rect 25938 33212 26002 33216
rect 25938 33156 25942 33212
rect 25942 33156 25998 33212
rect 25998 33156 26002 33212
rect 25938 33152 26002 33156
rect 26018 33212 26082 33216
rect 26018 33156 26022 33212
rect 26022 33156 26078 33212
rect 26078 33156 26082 33212
rect 26018 33152 26082 33156
rect 10882 32668 10946 32672
rect 10882 32612 10886 32668
rect 10886 32612 10942 32668
rect 10942 32612 10946 32668
rect 10882 32608 10946 32612
rect 10962 32668 11026 32672
rect 10962 32612 10966 32668
rect 10966 32612 11022 32668
rect 11022 32612 11026 32668
rect 10962 32608 11026 32612
rect 11042 32668 11106 32672
rect 11042 32612 11046 32668
rect 11046 32612 11102 32668
rect 11102 32612 11106 32668
rect 11042 32608 11106 32612
rect 11122 32668 11186 32672
rect 11122 32612 11126 32668
rect 11126 32612 11182 32668
rect 11182 32612 11186 32668
rect 11122 32608 11186 32612
rect 20813 32668 20877 32672
rect 20813 32612 20817 32668
rect 20817 32612 20873 32668
rect 20873 32612 20877 32668
rect 20813 32608 20877 32612
rect 20893 32668 20957 32672
rect 20893 32612 20897 32668
rect 20897 32612 20953 32668
rect 20953 32612 20957 32668
rect 20893 32608 20957 32612
rect 20973 32668 21037 32672
rect 20973 32612 20977 32668
rect 20977 32612 21033 32668
rect 21033 32612 21037 32668
rect 20973 32608 21037 32612
rect 21053 32668 21117 32672
rect 21053 32612 21057 32668
rect 21057 32612 21113 32668
rect 21113 32612 21117 32668
rect 21053 32608 21117 32612
rect 5917 32124 5981 32128
rect 5917 32068 5921 32124
rect 5921 32068 5977 32124
rect 5977 32068 5981 32124
rect 5917 32064 5981 32068
rect 5997 32124 6061 32128
rect 5997 32068 6001 32124
rect 6001 32068 6057 32124
rect 6057 32068 6061 32124
rect 5997 32064 6061 32068
rect 6077 32124 6141 32128
rect 6077 32068 6081 32124
rect 6081 32068 6137 32124
rect 6137 32068 6141 32124
rect 6077 32064 6141 32068
rect 6157 32124 6221 32128
rect 6157 32068 6161 32124
rect 6161 32068 6217 32124
rect 6217 32068 6221 32124
rect 6157 32064 6221 32068
rect 15848 32124 15912 32128
rect 15848 32068 15852 32124
rect 15852 32068 15908 32124
rect 15908 32068 15912 32124
rect 15848 32064 15912 32068
rect 15928 32124 15992 32128
rect 15928 32068 15932 32124
rect 15932 32068 15988 32124
rect 15988 32068 15992 32124
rect 15928 32064 15992 32068
rect 16008 32124 16072 32128
rect 16008 32068 16012 32124
rect 16012 32068 16068 32124
rect 16068 32068 16072 32124
rect 16008 32064 16072 32068
rect 16088 32124 16152 32128
rect 16088 32068 16092 32124
rect 16092 32068 16148 32124
rect 16148 32068 16152 32124
rect 16088 32064 16152 32068
rect 25778 32124 25842 32128
rect 25778 32068 25782 32124
rect 25782 32068 25838 32124
rect 25838 32068 25842 32124
rect 25778 32064 25842 32068
rect 25858 32124 25922 32128
rect 25858 32068 25862 32124
rect 25862 32068 25918 32124
rect 25918 32068 25922 32124
rect 25858 32064 25922 32068
rect 25938 32124 26002 32128
rect 25938 32068 25942 32124
rect 25942 32068 25998 32124
rect 25998 32068 26002 32124
rect 25938 32064 26002 32068
rect 26018 32124 26082 32128
rect 26018 32068 26022 32124
rect 26022 32068 26078 32124
rect 26078 32068 26082 32124
rect 26018 32064 26082 32068
rect 10882 31580 10946 31584
rect 10882 31524 10886 31580
rect 10886 31524 10942 31580
rect 10942 31524 10946 31580
rect 10882 31520 10946 31524
rect 10962 31580 11026 31584
rect 10962 31524 10966 31580
rect 10966 31524 11022 31580
rect 11022 31524 11026 31580
rect 10962 31520 11026 31524
rect 11042 31580 11106 31584
rect 11042 31524 11046 31580
rect 11046 31524 11102 31580
rect 11102 31524 11106 31580
rect 11042 31520 11106 31524
rect 11122 31580 11186 31584
rect 11122 31524 11126 31580
rect 11126 31524 11182 31580
rect 11182 31524 11186 31580
rect 11122 31520 11186 31524
rect 20813 31580 20877 31584
rect 20813 31524 20817 31580
rect 20817 31524 20873 31580
rect 20873 31524 20877 31580
rect 20813 31520 20877 31524
rect 20893 31580 20957 31584
rect 20893 31524 20897 31580
rect 20897 31524 20953 31580
rect 20953 31524 20957 31580
rect 20893 31520 20957 31524
rect 20973 31580 21037 31584
rect 20973 31524 20977 31580
rect 20977 31524 21033 31580
rect 21033 31524 21037 31580
rect 20973 31520 21037 31524
rect 21053 31580 21117 31584
rect 21053 31524 21057 31580
rect 21057 31524 21113 31580
rect 21113 31524 21117 31580
rect 21053 31520 21117 31524
rect 5917 31036 5981 31040
rect 5917 30980 5921 31036
rect 5921 30980 5977 31036
rect 5977 30980 5981 31036
rect 5917 30976 5981 30980
rect 5997 31036 6061 31040
rect 5997 30980 6001 31036
rect 6001 30980 6057 31036
rect 6057 30980 6061 31036
rect 5997 30976 6061 30980
rect 6077 31036 6141 31040
rect 6077 30980 6081 31036
rect 6081 30980 6137 31036
rect 6137 30980 6141 31036
rect 6077 30976 6141 30980
rect 6157 31036 6221 31040
rect 6157 30980 6161 31036
rect 6161 30980 6217 31036
rect 6217 30980 6221 31036
rect 6157 30976 6221 30980
rect 15848 31036 15912 31040
rect 15848 30980 15852 31036
rect 15852 30980 15908 31036
rect 15908 30980 15912 31036
rect 15848 30976 15912 30980
rect 15928 31036 15992 31040
rect 15928 30980 15932 31036
rect 15932 30980 15988 31036
rect 15988 30980 15992 31036
rect 15928 30976 15992 30980
rect 16008 31036 16072 31040
rect 16008 30980 16012 31036
rect 16012 30980 16068 31036
rect 16068 30980 16072 31036
rect 16008 30976 16072 30980
rect 16088 31036 16152 31040
rect 16088 30980 16092 31036
rect 16092 30980 16148 31036
rect 16148 30980 16152 31036
rect 16088 30976 16152 30980
rect 25778 31036 25842 31040
rect 25778 30980 25782 31036
rect 25782 30980 25838 31036
rect 25838 30980 25842 31036
rect 25778 30976 25842 30980
rect 25858 31036 25922 31040
rect 25858 30980 25862 31036
rect 25862 30980 25918 31036
rect 25918 30980 25922 31036
rect 25858 30976 25922 30980
rect 25938 31036 26002 31040
rect 25938 30980 25942 31036
rect 25942 30980 25998 31036
rect 25998 30980 26002 31036
rect 25938 30976 26002 30980
rect 26018 31036 26082 31040
rect 26018 30980 26022 31036
rect 26022 30980 26078 31036
rect 26078 30980 26082 31036
rect 26018 30976 26082 30980
rect 10882 30492 10946 30496
rect 10882 30436 10886 30492
rect 10886 30436 10942 30492
rect 10942 30436 10946 30492
rect 10882 30432 10946 30436
rect 10962 30492 11026 30496
rect 10962 30436 10966 30492
rect 10966 30436 11022 30492
rect 11022 30436 11026 30492
rect 10962 30432 11026 30436
rect 11042 30492 11106 30496
rect 11042 30436 11046 30492
rect 11046 30436 11102 30492
rect 11102 30436 11106 30492
rect 11042 30432 11106 30436
rect 11122 30492 11186 30496
rect 11122 30436 11126 30492
rect 11126 30436 11182 30492
rect 11182 30436 11186 30492
rect 11122 30432 11186 30436
rect 20813 30492 20877 30496
rect 20813 30436 20817 30492
rect 20817 30436 20873 30492
rect 20873 30436 20877 30492
rect 20813 30432 20877 30436
rect 20893 30492 20957 30496
rect 20893 30436 20897 30492
rect 20897 30436 20953 30492
rect 20953 30436 20957 30492
rect 20893 30432 20957 30436
rect 20973 30492 21037 30496
rect 20973 30436 20977 30492
rect 20977 30436 21033 30492
rect 21033 30436 21037 30492
rect 20973 30432 21037 30436
rect 21053 30492 21117 30496
rect 21053 30436 21057 30492
rect 21057 30436 21113 30492
rect 21113 30436 21117 30492
rect 21053 30432 21117 30436
rect 9076 30424 9140 30428
rect 9076 30368 9090 30424
rect 9090 30368 9140 30424
rect 9076 30364 9140 30368
rect 18276 29956 18340 30020
rect 5917 29948 5981 29952
rect 5917 29892 5921 29948
rect 5921 29892 5977 29948
rect 5977 29892 5981 29948
rect 5917 29888 5981 29892
rect 5997 29948 6061 29952
rect 5997 29892 6001 29948
rect 6001 29892 6057 29948
rect 6057 29892 6061 29948
rect 5997 29888 6061 29892
rect 6077 29948 6141 29952
rect 6077 29892 6081 29948
rect 6081 29892 6137 29948
rect 6137 29892 6141 29948
rect 6077 29888 6141 29892
rect 6157 29948 6221 29952
rect 6157 29892 6161 29948
rect 6161 29892 6217 29948
rect 6217 29892 6221 29948
rect 6157 29888 6221 29892
rect 15848 29948 15912 29952
rect 15848 29892 15852 29948
rect 15852 29892 15908 29948
rect 15908 29892 15912 29948
rect 15848 29888 15912 29892
rect 15928 29948 15992 29952
rect 15928 29892 15932 29948
rect 15932 29892 15988 29948
rect 15988 29892 15992 29948
rect 15928 29888 15992 29892
rect 16008 29948 16072 29952
rect 16008 29892 16012 29948
rect 16012 29892 16068 29948
rect 16068 29892 16072 29948
rect 16008 29888 16072 29892
rect 16088 29948 16152 29952
rect 16088 29892 16092 29948
rect 16092 29892 16148 29948
rect 16148 29892 16152 29948
rect 16088 29888 16152 29892
rect 25778 29948 25842 29952
rect 25778 29892 25782 29948
rect 25782 29892 25838 29948
rect 25838 29892 25842 29948
rect 25778 29888 25842 29892
rect 25858 29948 25922 29952
rect 25858 29892 25862 29948
rect 25862 29892 25918 29948
rect 25918 29892 25922 29948
rect 25858 29888 25922 29892
rect 25938 29948 26002 29952
rect 25938 29892 25942 29948
rect 25942 29892 25998 29948
rect 25998 29892 26002 29948
rect 25938 29888 26002 29892
rect 26018 29948 26082 29952
rect 26018 29892 26022 29948
rect 26022 29892 26078 29948
rect 26078 29892 26082 29948
rect 26018 29888 26082 29892
rect 10882 29404 10946 29408
rect 10882 29348 10886 29404
rect 10886 29348 10942 29404
rect 10942 29348 10946 29404
rect 10882 29344 10946 29348
rect 10962 29404 11026 29408
rect 10962 29348 10966 29404
rect 10966 29348 11022 29404
rect 11022 29348 11026 29404
rect 10962 29344 11026 29348
rect 11042 29404 11106 29408
rect 11042 29348 11046 29404
rect 11046 29348 11102 29404
rect 11102 29348 11106 29404
rect 11042 29344 11106 29348
rect 11122 29404 11186 29408
rect 11122 29348 11126 29404
rect 11126 29348 11182 29404
rect 11182 29348 11186 29404
rect 11122 29344 11186 29348
rect 20813 29404 20877 29408
rect 20813 29348 20817 29404
rect 20817 29348 20873 29404
rect 20873 29348 20877 29404
rect 20813 29344 20877 29348
rect 20893 29404 20957 29408
rect 20893 29348 20897 29404
rect 20897 29348 20953 29404
rect 20953 29348 20957 29404
rect 20893 29344 20957 29348
rect 20973 29404 21037 29408
rect 20973 29348 20977 29404
rect 20977 29348 21033 29404
rect 21033 29348 21037 29404
rect 20973 29344 21037 29348
rect 21053 29404 21117 29408
rect 21053 29348 21057 29404
rect 21057 29348 21113 29404
rect 21113 29348 21117 29404
rect 21053 29344 21117 29348
rect 5917 28860 5981 28864
rect 5917 28804 5921 28860
rect 5921 28804 5977 28860
rect 5977 28804 5981 28860
rect 5917 28800 5981 28804
rect 5997 28860 6061 28864
rect 5997 28804 6001 28860
rect 6001 28804 6057 28860
rect 6057 28804 6061 28860
rect 5997 28800 6061 28804
rect 6077 28860 6141 28864
rect 6077 28804 6081 28860
rect 6081 28804 6137 28860
rect 6137 28804 6141 28860
rect 6077 28800 6141 28804
rect 6157 28860 6221 28864
rect 6157 28804 6161 28860
rect 6161 28804 6217 28860
rect 6217 28804 6221 28860
rect 6157 28800 6221 28804
rect 15848 28860 15912 28864
rect 15848 28804 15852 28860
rect 15852 28804 15908 28860
rect 15908 28804 15912 28860
rect 15848 28800 15912 28804
rect 15928 28860 15992 28864
rect 15928 28804 15932 28860
rect 15932 28804 15988 28860
rect 15988 28804 15992 28860
rect 15928 28800 15992 28804
rect 16008 28860 16072 28864
rect 16008 28804 16012 28860
rect 16012 28804 16068 28860
rect 16068 28804 16072 28860
rect 16008 28800 16072 28804
rect 16088 28860 16152 28864
rect 16088 28804 16092 28860
rect 16092 28804 16148 28860
rect 16148 28804 16152 28860
rect 16088 28800 16152 28804
rect 25778 28860 25842 28864
rect 25778 28804 25782 28860
rect 25782 28804 25838 28860
rect 25838 28804 25842 28860
rect 25778 28800 25842 28804
rect 25858 28860 25922 28864
rect 25858 28804 25862 28860
rect 25862 28804 25918 28860
rect 25918 28804 25922 28860
rect 25858 28800 25922 28804
rect 25938 28860 26002 28864
rect 25938 28804 25942 28860
rect 25942 28804 25998 28860
rect 25998 28804 26002 28860
rect 25938 28800 26002 28804
rect 26018 28860 26082 28864
rect 26018 28804 26022 28860
rect 26022 28804 26078 28860
rect 26078 28804 26082 28860
rect 26018 28800 26082 28804
rect 10882 28316 10946 28320
rect 10882 28260 10886 28316
rect 10886 28260 10942 28316
rect 10942 28260 10946 28316
rect 10882 28256 10946 28260
rect 10962 28316 11026 28320
rect 10962 28260 10966 28316
rect 10966 28260 11022 28316
rect 11022 28260 11026 28316
rect 10962 28256 11026 28260
rect 11042 28316 11106 28320
rect 11042 28260 11046 28316
rect 11046 28260 11102 28316
rect 11102 28260 11106 28316
rect 11042 28256 11106 28260
rect 11122 28316 11186 28320
rect 11122 28260 11126 28316
rect 11126 28260 11182 28316
rect 11182 28260 11186 28316
rect 11122 28256 11186 28260
rect 20813 28316 20877 28320
rect 20813 28260 20817 28316
rect 20817 28260 20873 28316
rect 20873 28260 20877 28316
rect 20813 28256 20877 28260
rect 20893 28316 20957 28320
rect 20893 28260 20897 28316
rect 20897 28260 20953 28316
rect 20953 28260 20957 28316
rect 20893 28256 20957 28260
rect 20973 28316 21037 28320
rect 20973 28260 20977 28316
rect 20977 28260 21033 28316
rect 21033 28260 21037 28316
rect 20973 28256 21037 28260
rect 21053 28316 21117 28320
rect 21053 28260 21057 28316
rect 21057 28260 21113 28316
rect 21113 28260 21117 28316
rect 21053 28256 21117 28260
rect 5917 27772 5981 27776
rect 5917 27716 5921 27772
rect 5921 27716 5977 27772
rect 5977 27716 5981 27772
rect 5917 27712 5981 27716
rect 5997 27772 6061 27776
rect 5997 27716 6001 27772
rect 6001 27716 6057 27772
rect 6057 27716 6061 27772
rect 5997 27712 6061 27716
rect 6077 27772 6141 27776
rect 6077 27716 6081 27772
rect 6081 27716 6137 27772
rect 6137 27716 6141 27772
rect 6077 27712 6141 27716
rect 6157 27772 6221 27776
rect 6157 27716 6161 27772
rect 6161 27716 6217 27772
rect 6217 27716 6221 27772
rect 6157 27712 6221 27716
rect 15848 27772 15912 27776
rect 15848 27716 15852 27772
rect 15852 27716 15908 27772
rect 15908 27716 15912 27772
rect 15848 27712 15912 27716
rect 15928 27772 15992 27776
rect 15928 27716 15932 27772
rect 15932 27716 15988 27772
rect 15988 27716 15992 27772
rect 15928 27712 15992 27716
rect 16008 27772 16072 27776
rect 16008 27716 16012 27772
rect 16012 27716 16068 27772
rect 16068 27716 16072 27772
rect 16008 27712 16072 27716
rect 16088 27772 16152 27776
rect 16088 27716 16092 27772
rect 16092 27716 16148 27772
rect 16148 27716 16152 27772
rect 16088 27712 16152 27716
rect 25778 27772 25842 27776
rect 25778 27716 25782 27772
rect 25782 27716 25838 27772
rect 25838 27716 25842 27772
rect 25778 27712 25842 27716
rect 25858 27772 25922 27776
rect 25858 27716 25862 27772
rect 25862 27716 25918 27772
rect 25918 27716 25922 27772
rect 25858 27712 25922 27716
rect 25938 27772 26002 27776
rect 25938 27716 25942 27772
rect 25942 27716 25998 27772
rect 25998 27716 26002 27772
rect 25938 27712 26002 27716
rect 26018 27772 26082 27776
rect 26018 27716 26022 27772
rect 26022 27716 26078 27772
rect 26078 27716 26082 27772
rect 26018 27712 26082 27716
rect 8340 27432 8404 27436
rect 8340 27376 8390 27432
rect 8390 27376 8404 27432
rect 8340 27372 8404 27376
rect 10882 27228 10946 27232
rect 10882 27172 10886 27228
rect 10886 27172 10942 27228
rect 10942 27172 10946 27228
rect 10882 27168 10946 27172
rect 10962 27228 11026 27232
rect 10962 27172 10966 27228
rect 10966 27172 11022 27228
rect 11022 27172 11026 27228
rect 10962 27168 11026 27172
rect 11042 27228 11106 27232
rect 11042 27172 11046 27228
rect 11046 27172 11102 27228
rect 11102 27172 11106 27228
rect 11042 27168 11106 27172
rect 11122 27228 11186 27232
rect 11122 27172 11126 27228
rect 11126 27172 11182 27228
rect 11182 27172 11186 27228
rect 11122 27168 11186 27172
rect 20813 27228 20877 27232
rect 20813 27172 20817 27228
rect 20817 27172 20873 27228
rect 20873 27172 20877 27228
rect 20813 27168 20877 27172
rect 20893 27228 20957 27232
rect 20893 27172 20897 27228
rect 20897 27172 20953 27228
rect 20953 27172 20957 27228
rect 20893 27168 20957 27172
rect 20973 27228 21037 27232
rect 20973 27172 20977 27228
rect 20977 27172 21033 27228
rect 21033 27172 21037 27228
rect 20973 27168 21037 27172
rect 21053 27228 21117 27232
rect 21053 27172 21057 27228
rect 21057 27172 21113 27228
rect 21113 27172 21117 27228
rect 21053 27168 21117 27172
rect 5917 26684 5981 26688
rect 5917 26628 5921 26684
rect 5921 26628 5977 26684
rect 5977 26628 5981 26684
rect 5917 26624 5981 26628
rect 5997 26684 6061 26688
rect 5997 26628 6001 26684
rect 6001 26628 6057 26684
rect 6057 26628 6061 26684
rect 5997 26624 6061 26628
rect 6077 26684 6141 26688
rect 6077 26628 6081 26684
rect 6081 26628 6137 26684
rect 6137 26628 6141 26684
rect 6077 26624 6141 26628
rect 6157 26684 6221 26688
rect 6157 26628 6161 26684
rect 6161 26628 6217 26684
rect 6217 26628 6221 26684
rect 6157 26624 6221 26628
rect 15848 26684 15912 26688
rect 15848 26628 15852 26684
rect 15852 26628 15908 26684
rect 15908 26628 15912 26684
rect 15848 26624 15912 26628
rect 15928 26684 15992 26688
rect 15928 26628 15932 26684
rect 15932 26628 15988 26684
rect 15988 26628 15992 26684
rect 15928 26624 15992 26628
rect 16008 26684 16072 26688
rect 16008 26628 16012 26684
rect 16012 26628 16068 26684
rect 16068 26628 16072 26684
rect 16008 26624 16072 26628
rect 16088 26684 16152 26688
rect 16088 26628 16092 26684
rect 16092 26628 16148 26684
rect 16148 26628 16152 26684
rect 16088 26624 16152 26628
rect 25778 26684 25842 26688
rect 25778 26628 25782 26684
rect 25782 26628 25838 26684
rect 25838 26628 25842 26684
rect 25778 26624 25842 26628
rect 25858 26684 25922 26688
rect 25858 26628 25862 26684
rect 25862 26628 25918 26684
rect 25918 26628 25922 26684
rect 25858 26624 25922 26628
rect 25938 26684 26002 26688
rect 25938 26628 25942 26684
rect 25942 26628 25998 26684
rect 25998 26628 26002 26684
rect 25938 26624 26002 26628
rect 26018 26684 26082 26688
rect 26018 26628 26022 26684
rect 26022 26628 26078 26684
rect 26078 26628 26082 26684
rect 26018 26624 26082 26628
rect 8340 26284 8404 26348
rect 10882 26140 10946 26144
rect 10882 26084 10886 26140
rect 10886 26084 10942 26140
rect 10942 26084 10946 26140
rect 10882 26080 10946 26084
rect 10962 26140 11026 26144
rect 10962 26084 10966 26140
rect 10966 26084 11022 26140
rect 11022 26084 11026 26140
rect 10962 26080 11026 26084
rect 11042 26140 11106 26144
rect 11042 26084 11046 26140
rect 11046 26084 11102 26140
rect 11102 26084 11106 26140
rect 11042 26080 11106 26084
rect 11122 26140 11186 26144
rect 11122 26084 11126 26140
rect 11126 26084 11182 26140
rect 11182 26084 11186 26140
rect 11122 26080 11186 26084
rect 20813 26140 20877 26144
rect 20813 26084 20817 26140
rect 20817 26084 20873 26140
rect 20873 26084 20877 26140
rect 20813 26080 20877 26084
rect 20893 26140 20957 26144
rect 20893 26084 20897 26140
rect 20897 26084 20953 26140
rect 20953 26084 20957 26140
rect 20893 26080 20957 26084
rect 20973 26140 21037 26144
rect 20973 26084 20977 26140
rect 20977 26084 21033 26140
rect 21033 26084 21037 26140
rect 20973 26080 21037 26084
rect 21053 26140 21117 26144
rect 21053 26084 21057 26140
rect 21057 26084 21113 26140
rect 21113 26084 21117 26140
rect 21053 26080 21117 26084
rect 5917 25596 5981 25600
rect 5917 25540 5921 25596
rect 5921 25540 5977 25596
rect 5977 25540 5981 25596
rect 5917 25536 5981 25540
rect 5997 25596 6061 25600
rect 5997 25540 6001 25596
rect 6001 25540 6057 25596
rect 6057 25540 6061 25596
rect 5997 25536 6061 25540
rect 6077 25596 6141 25600
rect 6077 25540 6081 25596
rect 6081 25540 6137 25596
rect 6137 25540 6141 25596
rect 6077 25536 6141 25540
rect 6157 25596 6221 25600
rect 6157 25540 6161 25596
rect 6161 25540 6217 25596
rect 6217 25540 6221 25596
rect 6157 25536 6221 25540
rect 15848 25596 15912 25600
rect 15848 25540 15852 25596
rect 15852 25540 15908 25596
rect 15908 25540 15912 25596
rect 15848 25536 15912 25540
rect 15928 25596 15992 25600
rect 15928 25540 15932 25596
rect 15932 25540 15988 25596
rect 15988 25540 15992 25596
rect 15928 25536 15992 25540
rect 16008 25596 16072 25600
rect 16008 25540 16012 25596
rect 16012 25540 16068 25596
rect 16068 25540 16072 25596
rect 16008 25536 16072 25540
rect 16088 25596 16152 25600
rect 16088 25540 16092 25596
rect 16092 25540 16148 25596
rect 16148 25540 16152 25596
rect 16088 25536 16152 25540
rect 25778 25596 25842 25600
rect 25778 25540 25782 25596
rect 25782 25540 25838 25596
rect 25838 25540 25842 25596
rect 25778 25536 25842 25540
rect 25858 25596 25922 25600
rect 25858 25540 25862 25596
rect 25862 25540 25918 25596
rect 25918 25540 25922 25596
rect 25858 25536 25922 25540
rect 25938 25596 26002 25600
rect 25938 25540 25942 25596
rect 25942 25540 25998 25596
rect 25998 25540 26002 25596
rect 25938 25536 26002 25540
rect 26018 25596 26082 25600
rect 26018 25540 26022 25596
rect 26022 25540 26078 25596
rect 26078 25540 26082 25596
rect 26018 25536 26082 25540
rect 10882 25052 10946 25056
rect 10882 24996 10886 25052
rect 10886 24996 10942 25052
rect 10942 24996 10946 25052
rect 10882 24992 10946 24996
rect 10962 25052 11026 25056
rect 10962 24996 10966 25052
rect 10966 24996 11022 25052
rect 11022 24996 11026 25052
rect 10962 24992 11026 24996
rect 11042 25052 11106 25056
rect 11042 24996 11046 25052
rect 11046 24996 11102 25052
rect 11102 24996 11106 25052
rect 11042 24992 11106 24996
rect 11122 25052 11186 25056
rect 11122 24996 11126 25052
rect 11126 24996 11182 25052
rect 11182 24996 11186 25052
rect 11122 24992 11186 24996
rect 20813 25052 20877 25056
rect 20813 24996 20817 25052
rect 20817 24996 20873 25052
rect 20873 24996 20877 25052
rect 20813 24992 20877 24996
rect 20893 25052 20957 25056
rect 20893 24996 20897 25052
rect 20897 24996 20953 25052
rect 20953 24996 20957 25052
rect 20893 24992 20957 24996
rect 20973 25052 21037 25056
rect 20973 24996 20977 25052
rect 20977 24996 21033 25052
rect 21033 24996 21037 25052
rect 20973 24992 21037 24996
rect 21053 25052 21117 25056
rect 21053 24996 21057 25052
rect 21057 24996 21113 25052
rect 21113 24996 21117 25052
rect 21053 24992 21117 24996
rect 5917 24508 5981 24512
rect 5917 24452 5921 24508
rect 5921 24452 5977 24508
rect 5977 24452 5981 24508
rect 5917 24448 5981 24452
rect 5997 24508 6061 24512
rect 5997 24452 6001 24508
rect 6001 24452 6057 24508
rect 6057 24452 6061 24508
rect 5997 24448 6061 24452
rect 6077 24508 6141 24512
rect 6077 24452 6081 24508
rect 6081 24452 6137 24508
rect 6137 24452 6141 24508
rect 6077 24448 6141 24452
rect 6157 24508 6221 24512
rect 6157 24452 6161 24508
rect 6161 24452 6217 24508
rect 6217 24452 6221 24508
rect 6157 24448 6221 24452
rect 15848 24508 15912 24512
rect 15848 24452 15852 24508
rect 15852 24452 15908 24508
rect 15908 24452 15912 24508
rect 15848 24448 15912 24452
rect 15928 24508 15992 24512
rect 15928 24452 15932 24508
rect 15932 24452 15988 24508
rect 15988 24452 15992 24508
rect 15928 24448 15992 24452
rect 16008 24508 16072 24512
rect 16008 24452 16012 24508
rect 16012 24452 16068 24508
rect 16068 24452 16072 24508
rect 16008 24448 16072 24452
rect 16088 24508 16152 24512
rect 16088 24452 16092 24508
rect 16092 24452 16148 24508
rect 16148 24452 16152 24508
rect 16088 24448 16152 24452
rect 25778 24508 25842 24512
rect 25778 24452 25782 24508
rect 25782 24452 25838 24508
rect 25838 24452 25842 24508
rect 25778 24448 25842 24452
rect 25858 24508 25922 24512
rect 25858 24452 25862 24508
rect 25862 24452 25918 24508
rect 25918 24452 25922 24508
rect 25858 24448 25922 24452
rect 25938 24508 26002 24512
rect 25938 24452 25942 24508
rect 25942 24452 25998 24508
rect 25998 24452 26002 24508
rect 25938 24448 26002 24452
rect 26018 24508 26082 24512
rect 26018 24452 26022 24508
rect 26022 24452 26078 24508
rect 26078 24452 26082 24508
rect 26018 24448 26082 24452
rect 10882 23964 10946 23968
rect 10882 23908 10886 23964
rect 10886 23908 10942 23964
rect 10942 23908 10946 23964
rect 10882 23904 10946 23908
rect 10962 23964 11026 23968
rect 10962 23908 10966 23964
rect 10966 23908 11022 23964
rect 11022 23908 11026 23964
rect 10962 23904 11026 23908
rect 11042 23964 11106 23968
rect 11042 23908 11046 23964
rect 11046 23908 11102 23964
rect 11102 23908 11106 23964
rect 11042 23904 11106 23908
rect 11122 23964 11186 23968
rect 11122 23908 11126 23964
rect 11126 23908 11182 23964
rect 11182 23908 11186 23964
rect 11122 23904 11186 23908
rect 20813 23964 20877 23968
rect 20813 23908 20817 23964
rect 20817 23908 20873 23964
rect 20873 23908 20877 23964
rect 20813 23904 20877 23908
rect 20893 23964 20957 23968
rect 20893 23908 20897 23964
rect 20897 23908 20953 23964
rect 20953 23908 20957 23964
rect 20893 23904 20957 23908
rect 20973 23964 21037 23968
rect 20973 23908 20977 23964
rect 20977 23908 21033 23964
rect 21033 23908 21037 23964
rect 20973 23904 21037 23908
rect 21053 23964 21117 23968
rect 21053 23908 21057 23964
rect 21057 23908 21113 23964
rect 21113 23908 21117 23964
rect 21053 23904 21117 23908
rect 5917 23420 5981 23424
rect 5917 23364 5921 23420
rect 5921 23364 5977 23420
rect 5977 23364 5981 23420
rect 5917 23360 5981 23364
rect 5997 23420 6061 23424
rect 5997 23364 6001 23420
rect 6001 23364 6057 23420
rect 6057 23364 6061 23420
rect 5997 23360 6061 23364
rect 6077 23420 6141 23424
rect 6077 23364 6081 23420
rect 6081 23364 6137 23420
rect 6137 23364 6141 23420
rect 6077 23360 6141 23364
rect 6157 23420 6221 23424
rect 6157 23364 6161 23420
rect 6161 23364 6217 23420
rect 6217 23364 6221 23420
rect 6157 23360 6221 23364
rect 15848 23420 15912 23424
rect 15848 23364 15852 23420
rect 15852 23364 15908 23420
rect 15908 23364 15912 23420
rect 15848 23360 15912 23364
rect 15928 23420 15992 23424
rect 15928 23364 15932 23420
rect 15932 23364 15988 23420
rect 15988 23364 15992 23420
rect 15928 23360 15992 23364
rect 16008 23420 16072 23424
rect 16008 23364 16012 23420
rect 16012 23364 16068 23420
rect 16068 23364 16072 23420
rect 16008 23360 16072 23364
rect 16088 23420 16152 23424
rect 16088 23364 16092 23420
rect 16092 23364 16148 23420
rect 16148 23364 16152 23420
rect 16088 23360 16152 23364
rect 25778 23420 25842 23424
rect 25778 23364 25782 23420
rect 25782 23364 25838 23420
rect 25838 23364 25842 23420
rect 25778 23360 25842 23364
rect 25858 23420 25922 23424
rect 25858 23364 25862 23420
rect 25862 23364 25918 23420
rect 25918 23364 25922 23420
rect 25858 23360 25922 23364
rect 25938 23420 26002 23424
rect 25938 23364 25942 23420
rect 25942 23364 25998 23420
rect 25998 23364 26002 23420
rect 25938 23360 26002 23364
rect 26018 23420 26082 23424
rect 26018 23364 26022 23420
rect 26022 23364 26078 23420
rect 26078 23364 26082 23420
rect 26018 23360 26082 23364
rect 10882 22876 10946 22880
rect 10882 22820 10886 22876
rect 10886 22820 10942 22876
rect 10942 22820 10946 22876
rect 10882 22816 10946 22820
rect 10962 22876 11026 22880
rect 10962 22820 10966 22876
rect 10966 22820 11022 22876
rect 11022 22820 11026 22876
rect 10962 22816 11026 22820
rect 11042 22876 11106 22880
rect 11042 22820 11046 22876
rect 11046 22820 11102 22876
rect 11102 22820 11106 22876
rect 11042 22816 11106 22820
rect 11122 22876 11186 22880
rect 11122 22820 11126 22876
rect 11126 22820 11182 22876
rect 11182 22820 11186 22876
rect 11122 22816 11186 22820
rect 20813 22876 20877 22880
rect 20813 22820 20817 22876
rect 20817 22820 20873 22876
rect 20873 22820 20877 22876
rect 20813 22816 20877 22820
rect 20893 22876 20957 22880
rect 20893 22820 20897 22876
rect 20897 22820 20953 22876
rect 20953 22820 20957 22876
rect 20893 22816 20957 22820
rect 20973 22876 21037 22880
rect 20973 22820 20977 22876
rect 20977 22820 21033 22876
rect 21033 22820 21037 22876
rect 20973 22816 21037 22820
rect 21053 22876 21117 22880
rect 21053 22820 21057 22876
rect 21057 22820 21113 22876
rect 21113 22820 21117 22876
rect 21053 22816 21117 22820
rect 5917 22332 5981 22336
rect 5917 22276 5921 22332
rect 5921 22276 5977 22332
rect 5977 22276 5981 22332
rect 5917 22272 5981 22276
rect 5997 22332 6061 22336
rect 5997 22276 6001 22332
rect 6001 22276 6057 22332
rect 6057 22276 6061 22332
rect 5997 22272 6061 22276
rect 6077 22332 6141 22336
rect 6077 22276 6081 22332
rect 6081 22276 6137 22332
rect 6137 22276 6141 22332
rect 6077 22272 6141 22276
rect 6157 22332 6221 22336
rect 6157 22276 6161 22332
rect 6161 22276 6217 22332
rect 6217 22276 6221 22332
rect 6157 22272 6221 22276
rect 15848 22332 15912 22336
rect 15848 22276 15852 22332
rect 15852 22276 15908 22332
rect 15908 22276 15912 22332
rect 15848 22272 15912 22276
rect 15928 22332 15992 22336
rect 15928 22276 15932 22332
rect 15932 22276 15988 22332
rect 15988 22276 15992 22332
rect 15928 22272 15992 22276
rect 16008 22332 16072 22336
rect 16008 22276 16012 22332
rect 16012 22276 16068 22332
rect 16068 22276 16072 22332
rect 16008 22272 16072 22276
rect 16088 22332 16152 22336
rect 16088 22276 16092 22332
rect 16092 22276 16148 22332
rect 16148 22276 16152 22332
rect 16088 22272 16152 22276
rect 25778 22332 25842 22336
rect 25778 22276 25782 22332
rect 25782 22276 25838 22332
rect 25838 22276 25842 22332
rect 25778 22272 25842 22276
rect 25858 22332 25922 22336
rect 25858 22276 25862 22332
rect 25862 22276 25918 22332
rect 25918 22276 25922 22332
rect 25858 22272 25922 22276
rect 25938 22332 26002 22336
rect 25938 22276 25942 22332
rect 25942 22276 25998 22332
rect 25998 22276 26002 22332
rect 25938 22272 26002 22276
rect 26018 22332 26082 22336
rect 26018 22276 26022 22332
rect 26022 22276 26078 22332
rect 26078 22276 26082 22332
rect 26018 22272 26082 22276
rect 8340 21932 8404 21996
rect 10882 21788 10946 21792
rect 10882 21732 10886 21788
rect 10886 21732 10942 21788
rect 10942 21732 10946 21788
rect 10882 21728 10946 21732
rect 10962 21788 11026 21792
rect 10962 21732 10966 21788
rect 10966 21732 11022 21788
rect 11022 21732 11026 21788
rect 10962 21728 11026 21732
rect 11042 21788 11106 21792
rect 11042 21732 11046 21788
rect 11046 21732 11102 21788
rect 11102 21732 11106 21788
rect 11042 21728 11106 21732
rect 11122 21788 11186 21792
rect 11122 21732 11126 21788
rect 11126 21732 11182 21788
rect 11182 21732 11186 21788
rect 11122 21728 11186 21732
rect 20813 21788 20877 21792
rect 20813 21732 20817 21788
rect 20817 21732 20873 21788
rect 20873 21732 20877 21788
rect 20813 21728 20877 21732
rect 20893 21788 20957 21792
rect 20893 21732 20897 21788
rect 20897 21732 20953 21788
rect 20953 21732 20957 21788
rect 20893 21728 20957 21732
rect 20973 21788 21037 21792
rect 20973 21732 20977 21788
rect 20977 21732 21033 21788
rect 21033 21732 21037 21788
rect 20973 21728 21037 21732
rect 21053 21788 21117 21792
rect 21053 21732 21057 21788
rect 21057 21732 21113 21788
rect 21113 21732 21117 21788
rect 21053 21728 21117 21732
rect 5917 21244 5981 21248
rect 5917 21188 5921 21244
rect 5921 21188 5977 21244
rect 5977 21188 5981 21244
rect 5917 21184 5981 21188
rect 5997 21244 6061 21248
rect 5997 21188 6001 21244
rect 6001 21188 6057 21244
rect 6057 21188 6061 21244
rect 5997 21184 6061 21188
rect 6077 21244 6141 21248
rect 6077 21188 6081 21244
rect 6081 21188 6137 21244
rect 6137 21188 6141 21244
rect 6077 21184 6141 21188
rect 6157 21244 6221 21248
rect 6157 21188 6161 21244
rect 6161 21188 6217 21244
rect 6217 21188 6221 21244
rect 6157 21184 6221 21188
rect 15848 21244 15912 21248
rect 15848 21188 15852 21244
rect 15852 21188 15908 21244
rect 15908 21188 15912 21244
rect 15848 21184 15912 21188
rect 15928 21244 15992 21248
rect 15928 21188 15932 21244
rect 15932 21188 15988 21244
rect 15988 21188 15992 21244
rect 15928 21184 15992 21188
rect 16008 21244 16072 21248
rect 16008 21188 16012 21244
rect 16012 21188 16068 21244
rect 16068 21188 16072 21244
rect 16008 21184 16072 21188
rect 16088 21244 16152 21248
rect 16088 21188 16092 21244
rect 16092 21188 16148 21244
rect 16148 21188 16152 21244
rect 16088 21184 16152 21188
rect 25778 21244 25842 21248
rect 25778 21188 25782 21244
rect 25782 21188 25838 21244
rect 25838 21188 25842 21244
rect 25778 21184 25842 21188
rect 25858 21244 25922 21248
rect 25858 21188 25862 21244
rect 25862 21188 25918 21244
rect 25918 21188 25922 21244
rect 25858 21184 25922 21188
rect 25938 21244 26002 21248
rect 25938 21188 25942 21244
rect 25942 21188 25998 21244
rect 25998 21188 26002 21244
rect 25938 21184 26002 21188
rect 26018 21244 26082 21248
rect 26018 21188 26022 21244
rect 26022 21188 26078 21244
rect 26078 21188 26082 21244
rect 26018 21184 26082 21188
rect 10882 20700 10946 20704
rect 10882 20644 10886 20700
rect 10886 20644 10942 20700
rect 10942 20644 10946 20700
rect 10882 20640 10946 20644
rect 10962 20700 11026 20704
rect 10962 20644 10966 20700
rect 10966 20644 11022 20700
rect 11022 20644 11026 20700
rect 10962 20640 11026 20644
rect 11042 20700 11106 20704
rect 11042 20644 11046 20700
rect 11046 20644 11102 20700
rect 11102 20644 11106 20700
rect 11042 20640 11106 20644
rect 11122 20700 11186 20704
rect 11122 20644 11126 20700
rect 11126 20644 11182 20700
rect 11182 20644 11186 20700
rect 11122 20640 11186 20644
rect 20813 20700 20877 20704
rect 20813 20644 20817 20700
rect 20817 20644 20873 20700
rect 20873 20644 20877 20700
rect 20813 20640 20877 20644
rect 20893 20700 20957 20704
rect 20893 20644 20897 20700
rect 20897 20644 20953 20700
rect 20953 20644 20957 20700
rect 20893 20640 20957 20644
rect 20973 20700 21037 20704
rect 20973 20644 20977 20700
rect 20977 20644 21033 20700
rect 21033 20644 21037 20700
rect 20973 20640 21037 20644
rect 21053 20700 21117 20704
rect 21053 20644 21057 20700
rect 21057 20644 21113 20700
rect 21113 20644 21117 20700
rect 21053 20640 21117 20644
rect 5917 20156 5981 20160
rect 5917 20100 5921 20156
rect 5921 20100 5977 20156
rect 5977 20100 5981 20156
rect 5917 20096 5981 20100
rect 5997 20156 6061 20160
rect 5997 20100 6001 20156
rect 6001 20100 6057 20156
rect 6057 20100 6061 20156
rect 5997 20096 6061 20100
rect 6077 20156 6141 20160
rect 6077 20100 6081 20156
rect 6081 20100 6137 20156
rect 6137 20100 6141 20156
rect 6077 20096 6141 20100
rect 6157 20156 6221 20160
rect 6157 20100 6161 20156
rect 6161 20100 6217 20156
rect 6217 20100 6221 20156
rect 6157 20096 6221 20100
rect 15848 20156 15912 20160
rect 15848 20100 15852 20156
rect 15852 20100 15908 20156
rect 15908 20100 15912 20156
rect 15848 20096 15912 20100
rect 15928 20156 15992 20160
rect 15928 20100 15932 20156
rect 15932 20100 15988 20156
rect 15988 20100 15992 20156
rect 15928 20096 15992 20100
rect 16008 20156 16072 20160
rect 16008 20100 16012 20156
rect 16012 20100 16068 20156
rect 16068 20100 16072 20156
rect 16008 20096 16072 20100
rect 16088 20156 16152 20160
rect 16088 20100 16092 20156
rect 16092 20100 16148 20156
rect 16148 20100 16152 20156
rect 16088 20096 16152 20100
rect 25778 20156 25842 20160
rect 25778 20100 25782 20156
rect 25782 20100 25838 20156
rect 25838 20100 25842 20156
rect 25778 20096 25842 20100
rect 25858 20156 25922 20160
rect 25858 20100 25862 20156
rect 25862 20100 25918 20156
rect 25918 20100 25922 20156
rect 25858 20096 25922 20100
rect 25938 20156 26002 20160
rect 25938 20100 25942 20156
rect 25942 20100 25998 20156
rect 25998 20100 26002 20156
rect 25938 20096 26002 20100
rect 26018 20156 26082 20160
rect 26018 20100 26022 20156
rect 26022 20100 26078 20156
rect 26078 20100 26082 20156
rect 26018 20096 26082 20100
rect 10882 19612 10946 19616
rect 10882 19556 10886 19612
rect 10886 19556 10942 19612
rect 10942 19556 10946 19612
rect 10882 19552 10946 19556
rect 10962 19612 11026 19616
rect 10962 19556 10966 19612
rect 10966 19556 11022 19612
rect 11022 19556 11026 19612
rect 10962 19552 11026 19556
rect 11042 19612 11106 19616
rect 11042 19556 11046 19612
rect 11046 19556 11102 19612
rect 11102 19556 11106 19612
rect 11042 19552 11106 19556
rect 11122 19612 11186 19616
rect 11122 19556 11126 19612
rect 11126 19556 11182 19612
rect 11182 19556 11186 19612
rect 11122 19552 11186 19556
rect 20813 19612 20877 19616
rect 20813 19556 20817 19612
rect 20817 19556 20873 19612
rect 20873 19556 20877 19612
rect 20813 19552 20877 19556
rect 20893 19612 20957 19616
rect 20893 19556 20897 19612
rect 20897 19556 20953 19612
rect 20953 19556 20957 19612
rect 20893 19552 20957 19556
rect 20973 19612 21037 19616
rect 20973 19556 20977 19612
rect 20977 19556 21033 19612
rect 21033 19556 21037 19612
rect 20973 19552 21037 19556
rect 21053 19612 21117 19616
rect 21053 19556 21057 19612
rect 21057 19556 21113 19612
rect 21113 19556 21117 19612
rect 21053 19552 21117 19556
rect 5917 19068 5981 19072
rect 5917 19012 5921 19068
rect 5921 19012 5977 19068
rect 5977 19012 5981 19068
rect 5917 19008 5981 19012
rect 5997 19068 6061 19072
rect 5997 19012 6001 19068
rect 6001 19012 6057 19068
rect 6057 19012 6061 19068
rect 5997 19008 6061 19012
rect 6077 19068 6141 19072
rect 6077 19012 6081 19068
rect 6081 19012 6137 19068
rect 6137 19012 6141 19068
rect 6077 19008 6141 19012
rect 6157 19068 6221 19072
rect 6157 19012 6161 19068
rect 6161 19012 6217 19068
rect 6217 19012 6221 19068
rect 6157 19008 6221 19012
rect 15848 19068 15912 19072
rect 15848 19012 15852 19068
rect 15852 19012 15908 19068
rect 15908 19012 15912 19068
rect 15848 19008 15912 19012
rect 15928 19068 15992 19072
rect 15928 19012 15932 19068
rect 15932 19012 15988 19068
rect 15988 19012 15992 19068
rect 15928 19008 15992 19012
rect 16008 19068 16072 19072
rect 16008 19012 16012 19068
rect 16012 19012 16068 19068
rect 16068 19012 16072 19068
rect 16008 19008 16072 19012
rect 16088 19068 16152 19072
rect 16088 19012 16092 19068
rect 16092 19012 16148 19068
rect 16148 19012 16152 19068
rect 16088 19008 16152 19012
rect 25778 19068 25842 19072
rect 25778 19012 25782 19068
rect 25782 19012 25838 19068
rect 25838 19012 25842 19068
rect 25778 19008 25842 19012
rect 25858 19068 25922 19072
rect 25858 19012 25862 19068
rect 25862 19012 25918 19068
rect 25918 19012 25922 19068
rect 25858 19008 25922 19012
rect 25938 19068 26002 19072
rect 25938 19012 25942 19068
rect 25942 19012 25998 19068
rect 25998 19012 26002 19068
rect 25938 19008 26002 19012
rect 26018 19068 26082 19072
rect 26018 19012 26022 19068
rect 26022 19012 26078 19068
rect 26078 19012 26082 19068
rect 26018 19008 26082 19012
rect 10882 18524 10946 18528
rect 10882 18468 10886 18524
rect 10886 18468 10942 18524
rect 10942 18468 10946 18524
rect 10882 18464 10946 18468
rect 10962 18524 11026 18528
rect 10962 18468 10966 18524
rect 10966 18468 11022 18524
rect 11022 18468 11026 18524
rect 10962 18464 11026 18468
rect 11042 18524 11106 18528
rect 11042 18468 11046 18524
rect 11046 18468 11102 18524
rect 11102 18468 11106 18524
rect 11042 18464 11106 18468
rect 11122 18524 11186 18528
rect 11122 18468 11126 18524
rect 11126 18468 11182 18524
rect 11182 18468 11186 18524
rect 11122 18464 11186 18468
rect 20813 18524 20877 18528
rect 20813 18468 20817 18524
rect 20817 18468 20873 18524
rect 20873 18468 20877 18524
rect 20813 18464 20877 18468
rect 20893 18524 20957 18528
rect 20893 18468 20897 18524
rect 20897 18468 20953 18524
rect 20953 18468 20957 18524
rect 20893 18464 20957 18468
rect 20973 18524 21037 18528
rect 20973 18468 20977 18524
rect 20977 18468 21033 18524
rect 21033 18468 21037 18524
rect 20973 18464 21037 18468
rect 21053 18524 21117 18528
rect 21053 18468 21057 18524
rect 21057 18468 21113 18524
rect 21113 18468 21117 18524
rect 21053 18464 21117 18468
rect 5917 17980 5981 17984
rect 5917 17924 5921 17980
rect 5921 17924 5977 17980
rect 5977 17924 5981 17980
rect 5917 17920 5981 17924
rect 5997 17980 6061 17984
rect 5997 17924 6001 17980
rect 6001 17924 6057 17980
rect 6057 17924 6061 17980
rect 5997 17920 6061 17924
rect 6077 17980 6141 17984
rect 6077 17924 6081 17980
rect 6081 17924 6137 17980
rect 6137 17924 6141 17980
rect 6077 17920 6141 17924
rect 6157 17980 6221 17984
rect 6157 17924 6161 17980
rect 6161 17924 6217 17980
rect 6217 17924 6221 17980
rect 6157 17920 6221 17924
rect 15848 17980 15912 17984
rect 15848 17924 15852 17980
rect 15852 17924 15908 17980
rect 15908 17924 15912 17980
rect 15848 17920 15912 17924
rect 15928 17980 15992 17984
rect 15928 17924 15932 17980
rect 15932 17924 15988 17980
rect 15988 17924 15992 17980
rect 15928 17920 15992 17924
rect 16008 17980 16072 17984
rect 16008 17924 16012 17980
rect 16012 17924 16068 17980
rect 16068 17924 16072 17980
rect 16008 17920 16072 17924
rect 16088 17980 16152 17984
rect 16088 17924 16092 17980
rect 16092 17924 16148 17980
rect 16148 17924 16152 17980
rect 16088 17920 16152 17924
rect 25778 17980 25842 17984
rect 25778 17924 25782 17980
rect 25782 17924 25838 17980
rect 25838 17924 25842 17980
rect 25778 17920 25842 17924
rect 25858 17980 25922 17984
rect 25858 17924 25862 17980
rect 25862 17924 25918 17980
rect 25918 17924 25922 17980
rect 25858 17920 25922 17924
rect 25938 17980 26002 17984
rect 25938 17924 25942 17980
rect 25942 17924 25998 17980
rect 25998 17924 26002 17980
rect 25938 17920 26002 17924
rect 26018 17980 26082 17984
rect 26018 17924 26022 17980
rect 26022 17924 26078 17980
rect 26078 17924 26082 17980
rect 26018 17920 26082 17924
rect 10882 17436 10946 17440
rect 10882 17380 10886 17436
rect 10886 17380 10942 17436
rect 10942 17380 10946 17436
rect 10882 17376 10946 17380
rect 10962 17436 11026 17440
rect 10962 17380 10966 17436
rect 10966 17380 11022 17436
rect 11022 17380 11026 17436
rect 10962 17376 11026 17380
rect 11042 17436 11106 17440
rect 11042 17380 11046 17436
rect 11046 17380 11102 17436
rect 11102 17380 11106 17436
rect 11042 17376 11106 17380
rect 11122 17436 11186 17440
rect 11122 17380 11126 17436
rect 11126 17380 11182 17436
rect 11182 17380 11186 17436
rect 11122 17376 11186 17380
rect 20813 17436 20877 17440
rect 20813 17380 20817 17436
rect 20817 17380 20873 17436
rect 20873 17380 20877 17436
rect 20813 17376 20877 17380
rect 20893 17436 20957 17440
rect 20893 17380 20897 17436
rect 20897 17380 20953 17436
rect 20953 17380 20957 17436
rect 20893 17376 20957 17380
rect 20973 17436 21037 17440
rect 20973 17380 20977 17436
rect 20977 17380 21033 17436
rect 21033 17380 21037 17436
rect 20973 17376 21037 17380
rect 21053 17436 21117 17440
rect 21053 17380 21057 17436
rect 21057 17380 21113 17436
rect 21113 17380 21117 17436
rect 21053 17376 21117 17380
rect 5917 16892 5981 16896
rect 5917 16836 5921 16892
rect 5921 16836 5977 16892
rect 5977 16836 5981 16892
rect 5917 16832 5981 16836
rect 5997 16892 6061 16896
rect 5997 16836 6001 16892
rect 6001 16836 6057 16892
rect 6057 16836 6061 16892
rect 5997 16832 6061 16836
rect 6077 16892 6141 16896
rect 6077 16836 6081 16892
rect 6081 16836 6137 16892
rect 6137 16836 6141 16892
rect 6077 16832 6141 16836
rect 6157 16892 6221 16896
rect 6157 16836 6161 16892
rect 6161 16836 6217 16892
rect 6217 16836 6221 16892
rect 6157 16832 6221 16836
rect 15848 16892 15912 16896
rect 15848 16836 15852 16892
rect 15852 16836 15908 16892
rect 15908 16836 15912 16892
rect 15848 16832 15912 16836
rect 15928 16892 15992 16896
rect 15928 16836 15932 16892
rect 15932 16836 15988 16892
rect 15988 16836 15992 16892
rect 15928 16832 15992 16836
rect 16008 16892 16072 16896
rect 16008 16836 16012 16892
rect 16012 16836 16068 16892
rect 16068 16836 16072 16892
rect 16008 16832 16072 16836
rect 16088 16892 16152 16896
rect 16088 16836 16092 16892
rect 16092 16836 16148 16892
rect 16148 16836 16152 16892
rect 16088 16832 16152 16836
rect 25778 16892 25842 16896
rect 25778 16836 25782 16892
rect 25782 16836 25838 16892
rect 25838 16836 25842 16892
rect 25778 16832 25842 16836
rect 25858 16892 25922 16896
rect 25858 16836 25862 16892
rect 25862 16836 25918 16892
rect 25918 16836 25922 16892
rect 25858 16832 25922 16836
rect 25938 16892 26002 16896
rect 25938 16836 25942 16892
rect 25942 16836 25998 16892
rect 25998 16836 26002 16892
rect 25938 16832 26002 16836
rect 26018 16892 26082 16896
rect 26018 16836 26022 16892
rect 26022 16836 26078 16892
rect 26078 16836 26082 16892
rect 26018 16832 26082 16836
rect 10882 16348 10946 16352
rect 10882 16292 10886 16348
rect 10886 16292 10942 16348
rect 10942 16292 10946 16348
rect 10882 16288 10946 16292
rect 10962 16348 11026 16352
rect 10962 16292 10966 16348
rect 10966 16292 11022 16348
rect 11022 16292 11026 16348
rect 10962 16288 11026 16292
rect 11042 16348 11106 16352
rect 11042 16292 11046 16348
rect 11046 16292 11102 16348
rect 11102 16292 11106 16348
rect 11042 16288 11106 16292
rect 11122 16348 11186 16352
rect 11122 16292 11126 16348
rect 11126 16292 11182 16348
rect 11182 16292 11186 16348
rect 11122 16288 11186 16292
rect 20813 16348 20877 16352
rect 20813 16292 20817 16348
rect 20817 16292 20873 16348
rect 20873 16292 20877 16348
rect 20813 16288 20877 16292
rect 20893 16348 20957 16352
rect 20893 16292 20897 16348
rect 20897 16292 20953 16348
rect 20953 16292 20957 16348
rect 20893 16288 20957 16292
rect 20973 16348 21037 16352
rect 20973 16292 20977 16348
rect 20977 16292 21033 16348
rect 21033 16292 21037 16348
rect 20973 16288 21037 16292
rect 21053 16348 21117 16352
rect 21053 16292 21057 16348
rect 21057 16292 21113 16348
rect 21113 16292 21117 16348
rect 21053 16288 21117 16292
rect 18276 16084 18340 16148
rect 5764 15948 5828 16012
rect 5917 15804 5981 15808
rect 5917 15748 5921 15804
rect 5921 15748 5977 15804
rect 5977 15748 5981 15804
rect 5917 15744 5981 15748
rect 5997 15804 6061 15808
rect 5997 15748 6001 15804
rect 6001 15748 6057 15804
rect 6057 15748 6061 15804
rect 5997 15744 6061 15748
rect 6077 15804 6141 15808
rect 6077 15748 6081 15804
rect 6081 15748 6137 15804
rect 6137 15748 6141 15804
rect 6077 15744 6141 15748
rect 6157 15804 6221 15808
rect 6157 15748 6161 15804
rect 6161 15748 6217 15804
rect 6217 15748 6221 15804
rect 6157 15744 6221 15748
rect 15848 15804 15912 15808
rect 15848 15748 15852 15804
rect 15852 15748 15908 15804
rect 15908 15748 15912 15804
rect 15848 15744 15912 15748
rect 15928 15804 15992 15808
rect 15928 15748 15932 15804
rect 15932 15748 15988 15804
rect 15988 15748 15992 15804
rect 15928 15744 15992 15748
rect 16008 15804 16072 15808
rect 16008 15748 16012 15804
rect 16012 15748 16068 15804
rect 16068 15748 16072 15804
rect 16008 15744 16072 15748
rect 16088 15804 16152 15808
rect 16088 15748 16092 15804
rect 16092 15748 16148 15804
rect 16148 15748 16152 15804
rect 16088 15744 16152 15748
rect 25778 15804 25842 15808
rect 25778 15748 25782 15804
rect 25782 15748 25838 15804
rect 25838 15748 25842 15804
rect 25778 15744 25842 15748
rect 25858 15804 25922 15808
rect 25858 15748 25862 15804
rect 25862 15748 25918 15804
rect 25918 15748 25922 15804
rect 25858 15744 25922 15748
rect 25938 15804 26002 15808
rect 25938 15748 25942 15804
rect 25942 15748 25998 15804
rect 25998 15748 26002 15804
rect 25938 15744 26002 15748
rect 26018 15804 26082 15808
rect 26018 15748 26022 15804
rect 26022 15748 26078 15804
rect 26078 15748 26082 15804
rect 26018 15744 26082 15748
rect 10882 15260 10946 15264
rect 10882 15204 10886 15260
rect 10886 15204 10942 15260
rect 10942 15204 10946 15260
rect 10882 15200 10946 15204
rect 10962 15260 11026 15264
rect 10962 15204 10966 15260
rect 10966 15204 11022 15260
rect 11022 15204 11026 15260
rect 10962 15200 11026 15204
rect 11042 15260 11106 15264
rect 11042 15204 11046 15260
rect 11046 15204 11102 15260
rect 11102 15204 11106 15260
rect 11042 15200 11106 15204
rect 11122 15260 11186 15264
rect 11122 15204 11126 15260
rect 11126 15204 11182 15260
rect 11182 15204 11186 15260
rect 11122 15200 11186 15204
rect 20813 15260 20877 15264
rect 20813 15204 20817 15260
rect 20817 15204 20873 15260
rect 20873 15204 20877 15260
rect 20813 15200 20877 15204
rect 20893 15260 20957 15264
rect 20893 15204 20897 15260
rect 20897 15204 20953 15260
rect 20953 15204 20957 15260
rect 20893 15200 20957 15204
rect 20973 15260 21037 15264
rect 20973 15204 20977 15260
rect 20977 15204 21033 15260
rect 21033 15204 21037 15260
rect 20973 15200 21037 15204
rect 21053 15260 21117 15264
rect 21053 15204 21057 15260
rect 21057 15204 21113 15260
rect 21113 15204 21117 15260
rect 21053 15200 21117 15204
rect 5917 14716 5981 14720
rect 5917 14660 5921 14716
rect 5921 14660 5977 14716
rect 5977 14660 5981 14716
rect 5917 14656 5981 14660
rect 5997 14716 6061 14720
rect 5997 14660 6001 14716
rect 6001 14660 6057 14716
rect 6057 14660 6061 14716
rect 5997 14656 6061 14660
rect 6077 14716 6141 14720
rect 6077 14660 6081 14716
rect 6081 14660 6137 14716
rect 6137 14660 6141 14716
rect 6077 14656 6141 14660
rect 6157 14716 6221 14720
rect 6157 14660 6161 14716
rect 6161 14660 6217 14716
rect 6217 14660 6221 14716
rect 6157 14656 6221 14660
rect 15848 14716 15912 14720
rect 15848 14660 15852 14716
rect 15852 14660 15908 14716
rect 15908 14660 15912 14716
rect 15848 14656 15912 14660
rect 15928 14716 15992 14720
rect 15928 14660 15932 14716
rect 15932 14660 15988 14716
rect 15988 14660 15992 14716
rect 15928 14656 15992 14660
rect 16008 14716 16072 14720
rect 16008 14660 16012 14716
rect 16012 14660 16068 14716
rect 16068 14660 16072 14716
rect 16008 14656 16072 14660
rect 16088 14716 16152 14720
rect 16088 14660 16092 14716
rect 16092 14660 16148 14716
rect 16148 14660 16152 14716
rect 16088 14656 16152 14660
rect 25778 14716 25842 14720
rect 25778 14660 25782 14716
rect 25782 14660 25838 14716
rect 25838 14660 25842 14716
rect 25778 14656 25842 14660
rect 25858 14716 25922 14720
rect 25858 14660 25862 14716
rect 25862 14660 25918 14716
rect 25918 14660 25922 14716
rect 25858 14656 25922 14660
rect 25938 14716 26002 14720
rect 25938 14660 25942 14716
rect 25942 14660 25998 14716
rect 25998 14660 26002 14716
rect 25938 14656 26002 14660
rect 26018 14716 26082 14720
rect 26018 14660 26022 14716
rect 26022 14660 26078 14716
rect 26078 14660 26082 14716
rect 26018 14656 26082 14660
rect 10882 14172 10946 14176
rect 10882 14116 10886 14172
rect 10886 14116 10942 14172
rect 10942 14116 10946 14172
rect 10882 14112 10946 14116
rect 10962 14172 11026 14176
rect 10962 14116 10966 14172
rect 10966 14116 11022 14172
rect 11022 14116 11026 14172
rect 10962 14112 11026 14116
rect 11042 14172 11106 14176
rect 11042 14116 11046 14172
rect 11046 14116 11102 14172
rect 11102 14116 11106 14172
rect 11042 14112 11106 14116
rect 11122 14172 11186 14176
rect 11122 14116 11126 14172
rect 11126 14116 11182 14172
rect 11182 14116 11186 14172
rect 11122 14112 11186 14116
rect 20813 14172 20877 14176
rect 20813 14116 20817 14172
rect 20817 14116 20873 14172
rect 20873 14116 20877 14172
rect 20813 14112 20877 14116
rect 20893 14172 20957 14176
rect 20893 14116 20897 14172
rect 20897 14116 20953 14172
rect 20953 14116 20957 14172
rect 20893 14112 20957 14116
rect 20973 14172 21037 14176
rect 20973 14116 20977 14172
rect 20977 14116 21033 14172
rect 21033 14116 21037 14172
rect 20973 14112 21037 14116
rect 21053 14172 21117 14176
rect 21053 14116 21057 14172
rect 21057 14116 21113 14172
rect 21113 14116 21117 14172
rect 21053 14112 21117 14116
rect 5917 13628 5981 13632
rect 5917 13572 5921 13628
rect 5921 13572 5977 13628
rect 5977 13572 5981 13628
rect 5917 13568 5981 13572
rect 5997 13628 6061 13632
rect 5997 13572 6001 13628
rect 6001 13572 6057 13628
rect 6057 13572 6061 13628
rect 5997 13568 6061 13572
rect 6077 13628 6141 13632
rect 6077 13572 6081 13628
rect 6081 13572 6137 13628
rect 6137 13572 6141 13628
rect 6077 13568 6141 13572
rect 6157 13628 6221 13632
rect 6157 13572 6161 13628
rect 6161 13572 6217 13628
rect 6217 13572 6221 13628
rect 6157 13568 6221 13572
rect 15848 13628 15912 13632
rect 15848 13572 15852 13628
rect 15852 13572 15908 13628
rect 15908 13572 15912 13628
rect 15848 13568 15912 13572
rect 15928 13628 15992 13632
rect 15928 13572 15932 13628
rect 15932 13572 15988 13628
rect 15988 13572 15992 13628
rect 15928 13568 15992 13572
rect 16008 13628 16072 13632
rect 16008 13572 16012 13628
rect 16012 13572 16068 13628
rect 16068 13572 16072 13628
rect 16008 13568 16072 13572
rect 16088 13628 16152 13632
rect 16088 13572 16092 13628
rect 16092 13572 16148 13628
rect 16148 13572 16152 13628
rect 16088 13568 16152 13572
rect 25778 13628 25842 13632
rect 25778 13572 25782 13628
rect 25782 13572 25838 13628
rect 25838 13572 25842 13628
rect 25778 13568 25842 13572
rect 25858 13628 25922 13632
rect 25858 13572 25862 13628
rect 25862 13572 25918 13628
rect 25918 13572 25922 13628
rect 25858 13568 25922 13572
rect 25938 13628 26002 13632
rect 25938 13572 25942 13628
rect 25942 13572 25998 13628
rect 25998 13572 26002 13628
rect 25938 13568 26002 13572
rect 26018 13628 26082 13632
rect 26018 13572 26022 13628
rect 26022 13572 26078 13628
rect 26078 13572 26082 13628
rect 26018 13568 26082 13572
rect 10882 13084 10946 13088
rect 10882 13028 10886 13084
rect 10886 13028 10942 13084
rect 10942 13028 10946 13084
rect 10882 13024 10946 13028
rect 10962 13084 11026 13088
rect 10962 13028 10966 13084
rect 10966 13028 11022 13084
rect 11022 13028 11026 13084
rect 10962 13024 11026 13028
rect 11042 13084 11106 13088
rect 11042 13028 11046 13084
rect 11046 13028 11102 13084
rect 11102 13028 11106 13084
rect 11042 13024 11106 13028
rect 11122 13084 11186 13088
rect 11122 13028 11126 13084
rect 11126 13028 11182 13084
rect 11182 13028 11186 13084
rect 11122 13024 11186 13028
rect 20813 13084 20877 13088
rect 20813 13028 20817 13084
rect 20817 13028 20873 13084
rect 20873 13028 20877 13084
rect 20813 13024 20877 13028
rect 20893 13084 20957 13088
rect 20893 13028 20897 13084
rect 20897 13028 20953 13084
rect 20953 13028 20957 13084
rect 20893 13024 20957 13028
rect 20973 13084 21037 13088
rect 20973 13028 20977 13084
rect 20977 13028 21033 13084
rect 21033 13028 21037 13084
rect 20973 13024 21037 13028
rect 21053 13084 21117 13088
rect 21053 13028 21057 13084
rect 21057 13028 21113 13084
rect 21113 13028 21117 13084
rect 21053 13024 21117 13028
rect 5917 12540 5981 12544
rect 5917 12484 5921 12540
rect 5921 12484 5977 12540
rect 5977 12484 5981 12540
rect 5917 12480 5981 12484
rect 5997 12540 6061 12544
rect 5997 12484 6001 12540
rect 6001 12484 6057 12540
rect 6057 12484 6061 12540
rect 5997 12480 6061 12484
rect 6077 12540 6141 12544
rect 6077 12484 6081 12540
rect 6081 12484 6137 12540
rect 6137 12484 6141 12540
rect 6077 12480 6141 12484
rect 6157 12540 6221 12544
rect 6157 12484 6161 12540
rect 6161 12484 6217 12540
rect 6217 12484 6221 12540
rect 6157 12480 6221 12484
rect 15848 12540 15912 12544
rect 15848 12484 15852 12540
rect 15852 12484 15908 12540
rect 15908 12484 15912 12540
rect 15848 12480 15912 12484
rect 15928 12540 15992 12544
rect 15928 12484 15932 12540
rect 15932 12484 15988 12540
rect 15988 12484 15992 12540
rect 15928 12480 15992 12484
rect 16008 12540 16072 12544
rect 16008 12484 16012 12540
rect 16012 12484 16068 12540
rect 16068 12484 16072 12540
rect 16008 12480 16072 12484
rect 16088 12540 16152 12544
rect 16088 12484 16092 12540
rect 16092 12484 16148 12540
rect 16148 12484 16152 12540
rect 16088 12480 16152 12484
rect 25778 12540 25842 12544
rect 25778 12484 25782 12540
rect 25782 12484 25838 12540
rect 25838 12484 25842 12540
rect 25778 12480 25842 12484
rect 25858 12540 25922 12544
rect 25858 12484 25862 12540
rect 25862 12484 25918 12540
rect 25918 12484 25922 12540
rect 25858 12480 25922 12484
rect 25938 12540 26002 12544
rect 25938 12484 25942 12540
rect 25942 12484 25998 12540
rect 25998 12484 26002 12540
rect 25938 12480 26002 12484
rect 26018 12540 26082 12544
rect 26018 12484 26022 12540
rect 26022 12484 26078 12540
rect 26078 12484 26082 12540
rect 26018 12480 26082 12484
rect 10882 11996 10946 12000
rect 10882 11940 10886 11996
rect 10886 11940 10942 11996
rect 10942 11940 10946 11996
rect 10882 11936 10946 11940
rect 10962 11996 11026 12000
rect 10962 11940 10966 11996
rect 10966 11940 11022 11996
rect 11022 11940 11026 11996
rect 10962 11936 11026 11940
rect 11042 11996 11106 12000
rect 11042 11940 11046 11996
rect 11046 11940 11102 11996
rect 11102 11940 11106 11996
rect 11042 11936 11106 11940
rect 11122 11996 11186 12000
rect 11122 11940 11126 11996
rect 11126 11940 11182 11996
rect 11182 11940 11186 11996
rect 11122 11936 11186 11940
rect 20813 11996 20877 12000
rect 20813 11940 20817 11996
rect 20817 11940 20873 11996
rect 20873 11940 20877 11996
rect 20813 11936 20877 11940
rect 20893 11996 20957 12000
rect 20893 11940 20897 11996
rect 20897 11940 20953 11996
rect 20953 11940 20957 11996
rect 20893 11936 20957 11940
rect 20973 11996 21037 12000
rect 20973 11940 20977 11996
rect 20977 11940 21033 11996
rect 21033 11940 21037 11996
rect 20973 11936 21037 11940
rect 21053 11996 21117 12000
rect 21053 11940 21057 11996
rect 21057 11940 21113 11996
rect 21113 11940 21117 11996
rect 21053 11936 21117 11940
rect 5917 11452 5981 11456
rect 5917 11396 5921 11452
rect 5921 11396 5977 11452
rect 5977 11396 5981 11452
rect 5917 11392 5981 11396
rect 5997 11452 6061 11456
rect 5997 11396 6001 11452
rect 6001 11396 6057 11452
rect 6057 11396 6061 11452
rect 5997 11392 6061 11396
rect 6077 11452 6141 11456
rect 6077 11396 6081 11452
rect 6081 11396 6137 11452
rect 6137 11396 6141 11452
rect 6077 11392 6141 11396
rect 6157 11452 6221 11456
rect 6157 11396 6161 11452
rect 6161 11396 6217 11452
rect 6217 11396 6221 11452
rect 6157 11392 6221 11396
rect 15848 11452 15912 11456
rect 15848 11396 15852 11452
rect 15852 11396 15908 11452
rect 15908 11396 15912 11452
rect 15848 11392 15912 11396
rect 15928 11452 15992 11456
rect 15928 11396 15932 11452
rect 15932 11396 15988 11452
rect 15988 11396 15992 11452
rect 15928 11392 15992 11396
rect 16008 11452 16072 11456
rect 16008 11396 16012 11452
rect 16012 11396 16068 11452
rect 16068 11396 16072 11452
rect 16008 11392 16072 11396
rect 16088 11452 16152 11456
rect 16088 11396 16092 11452
rect 16092 11396 16148 11452
rect 16148 11396 16152 11452
rect 16088 11392 16152 11396
rect 25778 11452 25842 11456
rect 25778 11396 25782 11452
rect 25782 11396 25838 11452
rect 25838 11396 25842 11452
rect 25778 11392 25842 11396
rect 25858 11452 25922 11456
rect 25858 11396 25862 11452
rect 25862 11396 25918 11452
rect 25918 11396 25922 11452
rect 25858 11392 25922 11396
rect 25938 11452 26002 11456
rect 25938 11396 25942 11452
rect 25942 11396 25998 11452
rect 25998 11396 26002 11452
rect 25938 11392 26002 11396
rect 26018 11452 26082 11456
rect 26018 11396 26022 11452
rect 26022 11396 26078 11452
rect 26078 11396 26082 11452
rect 26018 11392 26082 11396
rect 10882 10908 10946 10912
rect 10882 10852 10886 10908
rect 10886 10852 10942 10908
rect 10942 10852 10946 10908
rect 10882 10848 10946 10852
rect 10962 10908 11026 10912
rect 10962 10852 10966 10908
rect 10966 10852 11022 10908
rect 11022 10852 11026 10908
rect 10962 10848 11026 10852
rect 11042 10908 11106 10912
rect 11042 10852 11046 10908
rect 11046 10852 11102 10908
rect 11102 10852 11106 10908
rect 11042 10848 11106 10852
rect 11122 10908 11186 10912
rect 11122 10852 11126 10908
rect 11126 10852 11182 10908
rect 11182 10852 11186 10908
rect 11122 10848 11186 10852
rect 20813 10908 20877 10912
rect 20813 10852 20817 10908
rect 20817 10852 20873 10908
rect 20873 10852 20877 10908
rect 20813 10848 20877 10852
rect 20893 10908 20957 10912
rect 20893 10852 20897 10908
rect 20897 10852 20953 10908
rect 20953 10852 20957 10908
rect 20893 10848 20957 10852
rect 20973 10908 21037 10912
rect 20973 10852 20977 10908
rect 20977 10852 21033 10908
rect 21033 10852 21037 10908
rect 20973 10848 21037 10852
rect 21053 10908 21117 10912
rect 21053 10852 21057 10908
rect 21057 10852 21113 10908
rect 21113 10852 21117 10908
rect 21053 10848 21117 10852
rect 5917 10364 5981 10368
rect 5917 10308 5921 10364
rect 5921 10308 5977 10364
rect 5977 10308 5981 10364
rect 5917 10304 5981 10308
rect 5997 10364 6061 10368
rect 5997 10308 6001 10364
rect 6001 10308 6057 10364
rect 6057 10308 6061 10364
rect 5997 10304 6061 10308
rect 6077 10364 6141 10368
rect 6077 10308 6081 10364
rect 6081 10308 6137 10364
rect 6137 10308 6141 10364
rect 6077 10304 6141 10308
rect 6157 10364 6221 10368
rect 6157 10308 6161 10364
rect 6161 10308 6217 10364
rect 6217 10308 6221 10364
rect 6157 10304 6221 10308
rect 15848 10364 15912 10368
rect 15848 10308 15852 10364
rect 15852 10308 15908 10364
rect 15908 10308 15912 10364
rect 15848 10304 15912 10308
rect 15928 10364 15992 10368
rect 15928 10308 15932 10364
rect 15932 10308 15988 10364
rect 15988 10308 15992 10364
rect 15928 10304 15992 10308
rect 16008 10364 16072 10368
rect 16008 10308 16012 10364
rect 16012 10308 16068 10364
rect 16068 10308 16072 10364
rect 16008 10304 16072 10308
rect 16088 10364 16152 10368
rect 16088 10308 16092 10364
rect 16092 10308 16148 10364
rect 16148 10308 16152 10364
rect 16088 10304 16152 10308
rect 25778 10364 25842 10368
rect 25778 10308 25782 10364
rect 25782 10308 25838 10364
rect 25838 10308 25842 10364
rect 25778 10304 25842 10308
rect 25858 10364 25922 10368
rect 25858 10308 25862 10364
rect 25862 10308 25918 10364
rect 25918 10308 25922 10364
rect 25858 10304 25922 10308
rect 25938 10364 26002 10368
rect 25938 10308 25942 10364
rect 25942 10308 25998 10364
rect 25998 10308 26002 10364
rect 25938 10304 26002 10308
rect 26018 10364 26082 10368
rect 26018 10308 26022 10364
rect 26022 10308 26078 10364
rect 26078 10308 26082 10364
rect 26018 10304 26082 10308
rect 10882 9820 10946 9824
rect 10882 9764 10886 9820
rect 10886 9764 10942 9820
rect 10942 9764 10946 9820
rect 10882 9760 10946 9764
rect 10962 9820 11026 9824
rect 10962 9764 10966 9820
rect 10966 9764 11022 9820
rect 11022 9764 11026 9820
rect 10962 9760 11026 9764
rect 11042 9820 11106 9824
rect 11042 9764 11046 9820
rect 11046 9764 11102 9820
rect 11102 9764 11106 9820
rect 11042 9760 11106 9764
rect 11122 9820 11186 9824
rect 11122 9764 11126 9820
rect 11126 9764 11182 9820
rect 11182 9764 11186 9820
rect 11122 9760 11186 9764
rect 20813 9820 20877 9824
rect 20813 9764 20817 9820
rect 20817 9764 20873 9820
rect 20873 9764 20877 9820
rect 20813 9760 20877 9764
rect 20893 9820 20957 9824
rect 20893 9764 20897 9820
rect 20897 9764 20953 9820
rect 20953 9764 20957 9820
rect 20893 9760 20957 9764
rect 20973 9820 21037 9824
rect 20973 9764 20977 9820
rect 20977 9764 21033 9820
rect 21033 9764 21037 9820
rect 20973 9760 21037 9764
rect 21053 9820 21117 9824
rect 21053 9764 21057 9820
rect 21057 9764 21113 9820
rect 21113 9764 21117 9820
rect 21053 9760 21117 9764
rect 5917 9276 5981 9280
rect 5917 9220 5921 9276
rect 5921 9220 5977 9276
rect 5977 9220 5981 9276
rect 5917 9216 5981 9220
rect 5997 9276 6061 9280
rect 5997 9220 6001 9276
rect 6001 9220 6057 9276
rect 6057 9220 6061 9276
rect 5997 9216 6061 9220
rect 6077 9276 6141 9280
rect 6077 9220 6081 9276
rect 6081 9220 6137 9276
rect 6137 9220 6141 9276
rect 6077 9216 6141 9220
rect 6157 9276 6221 9280
rect 6157 9220 6161 9276
rect 6161 9220 6217 9276
rect 6217 9220 6221 9276
rect 6157 9216 6221 9220
rect 15848 9276 15912 9280
rect 15848 9220 15852 9276
rect 15852 9220 15908 9276
rect 15908 9220 15912 9276
rect 15848 9216 15912 9220
rect 15928 9276 15992 9280
rect 15928 9220 15932 9276
rect 15932 9220 15988 9276
rect 15988 9220 15992 9276
rect 15928 9216 15992 9220
rect 16008 9276 16072 9280
rect 16008 9220 16012 9276
rect 16012 9220 16068 9276
rect 16068 9220 16072 9276
rect 16008 9216 16072 9220
rect 16088 9276 16152 9280
rect 16088 9220 16092 9276
rect 16092 9220 16148 9276
rect 16148 9220 16152 9276
rect 16088 9216 16152 9220
rect 25778 9276 25842 9280
rect 25778 9220 25782 9276
rect 25782 9220 25838 9276
rect 25838 9220 25842 9276
rect 25778 9216 25842 9220
rect 25858 9276 25922 9280
rect 25858 9220 25862 9276
rect 25862 9220 25918 9276
rect 25918 9220 25922 9276
rect 25858 9216 25922 9220
rect 25938 9276 26002 9280
rect 25938 9220 25942 9276
rect 25942 9220 25998 9276
rect 25998 9220 26002 9276
rect 25938 9216 26002 9220
rect 26018 9276 26082 9280
rect 26018 9220 26022 9276
rect 26022 9220 26078 9276
rect 26078 9220 26082 9276
rect 26018 9216 26082 9220
rect 5764 9012 5828 9076
rect 10882 8732 10946 8736
rect 10882 8676 10886 8732
rect 10886 8676 10942 8732
rect 10942 8676 10946 8732
rect 10882 8672 10946 8676
rect 10962 8732 11026 8736
rect 10962 8676 10966 8732
rect 10966 8676 11022 8732
rect 11022 8676 11026 8732
rect 10962 8672 11026 8676
rect 11042 8732 11106 8736
rect 11042 8676 11046 8732
rect 11046 8676 11102 8732
rect 11102 8676 11106 8732
rect 11042 8672 11106 8676
rect 11122 8732 11186 8736
rect 11122 8676 11126 8732
rect 11126 8676 11182 8732
rect 11182 8676 11186 8732
rect 11122 8672 11186 8676
rect 20813 8732 20877 8736
rect 20813 8676 20817 8732
rect 20817 8676 20873 8732
rect 20873 8676 20877 8732
rect 20813 8672 20877 8676
rect 20893 8732 20957 8736
rect 20893 8676 20897 8732
rect 20897 8676 20953 8732
rect 20953 8676 20957 8732
rect 20893 8672 20957 8676
rect 20973 8732 21037 8736
rect 20973 8676 20977 8732
rect 20977 8676 21033 8732
rect 21033 8676 21037 8732
rect 20973 8672 21037 8676
rect 21053 8732 21117 8736
rect 21053 8676 21057 8732
rect 21057 8676 21113 8732
rect 21113 8676 21117 8732
rect 21053 8672 21117 8676
rect 5917 8188 5981 8192
rect 5917 8132 5921 8188
rect 5921 8132 5977 8188
rect 5977 8132 5981 8188
rect 5917 8128 5981 8132
rect 5997 8188 6061 8192
rect 5997 8132 6001 8188
rect 6001 8132 6057 8188
rect 6057 8132 6061 8188
rect 5997 8128 6061 8132
rect 6077 8188 6141 8192
rect 6077 8132 6081 8188
rect 6081 8132 6137 8188
rect 6137 8132 6141 8188
rect 6077 8128 6141 8132
rect 6157 8188 6221 8192
rect 6157 8132 6161 8188
rect 6161 8132 6217 8188
rect 6217 8132 6221 8188
rect 6157 8128 6221 8132
rect 15848 8188 15912 8192
rect 15848 8132 15852 8188
rect 15852 8132 15908 8188
rect 15908 8132 15912 8188
rect 15848 8128 15912 8132
rect 15928 8188 15992 8192
rect 15928 8132 15932 8188
rect 15932 8132 15988 8188
rect 15988 8132 15992 8188
rect 15928 8128 15992 8132
rect 16008 8188 16072 8192
rect 16008 8132 16012 8188
rect 16012 8132 16068 8188
rect 16068 8132 16072 8188
rect 16008 8128 16072 8132
rect 16088 8188 16152 8192
rect 16088 8132 16092 8188
rect 16092 8132 16148 8188
rect 16148 8132 16152 8188
rect 16088 8128 16152 8132
rect 25778 8188 25842 8192
rect 25778 8132 25782 8188
rect 25782 8132 25838 8188
rect 25838 8132 25842 8188
rect 25778 8128 25842 8132
rect 25858 8188 25922 8192
rect 25858 8132 25862 8188
rect 25862 8132 25918 8188
rect 25918 8132 25922 8188
rect 25858 8128 25922 8132
rect 25938 8188 26002 8192
rect 25938 8132 25942 8188
rect 25942 8132 25998 8188
rect 25998 8132 26002 8188
rect 25938 8128 26002 8132
rect 26018 8188 26082 8192
rect 26018 8132 26022 8188
rect 26022 8132 26078 8188
rect 26078 8132 26082 8188
rect 26018 8128 26082 8132
rect 10882 7644 10946 7648
rect 10882 7588 10886 7644
rect 10886 7588 10942 7644
rect 10942 7588 10946 7644
rect 10882 7584 10946 7588
rect 10962 7644 11026 7648
rect 10962 7588 10966 7644
rect 10966 7588 11022 7644
rect 11022 7588 11026 7644
rect 10962 7584 11026 7588
rect 11042 7644 11106 7648
rect 11042 7588 11046 7644
rect 11046 7588 11102 7644
rect 11102 7588 11106 7644
rect 11042 7584 11106 7588
rect 11122 7644 11186 7648
rect 11122 7588 11126 7644
rect 11126 7588 11182 7644
rect 11182 7588 11186 7644
rect 11122 7584 11186 7588
rect 20813 7644 20877 7648
rect 20813 7588 20817 7644
rect 20817 7588 20873 7644
rect 20873 7588 20877 7644
rect 20813 7584 20877 7588
rect 20893 7644 20957 7648
rect 20893 7588 20897 7644
rect 20897 7588 20953 7644
rect 20953 7588 20957 7644
rect 20893 7584 20957 7588
rect 20973 7644 21037 7648
rect 20973 7588 20977 7644
rect 20977 7588 21033 7644
rect 21033 7588 21037 7644
rect 20973 7584 21037 7588
rect 21053 7644 21117 7648
rect 21053 7588 21057 7644
rect 21057 7588 21113 7644
rect 21113 7588 21117 7644
rect 21053 7584 21117 7588
rect 5917 7100 5981 7104
rect 5917 7044 5921 7100
rect 5921 7044 5977 7100
rect 5977 7044 5981 7100
rect 5917 7040 5981 7044
rect 5997 7100 6061 7104
rect 5997 7044 6001 7100
rect 6001 7044 6057 7100
rect 6057 7044 6061 7100
rect 5997 7040 6061 7044
rect 6077 7100 6141 7104
rect 6077 7044 6081 7100
rect 6081 7044 6137 7100
rect 6137 7044 6141 7100
rect 6077 7040 6141 7044
rect 6157 7100 6221 7104
rect 6157 7044 6161 7100
rect 6161 7044 6217 7100
rect 6217 7044 6221 7100
rect 6157 7040 6221 7044
rect 15848 7100 15912 7104
rect 15848 7044 15852 7100
rect 15852 7044 15908 7100
rect 15908 7044 15912 7100
rect 15848 7040 15912 7044
rect 15928 7100 15992 7104
rect 15928 7044 15932 7100
rect 15932 7044 15988 7100
rect 15988 7044 15992 7100
rect 15928 7040 15992 7044
rect 16008 7100 16072 7104
rect 16008 7044 16012 7100
rect 16012 7044 16068 7100
rect 16068 7044 16072 7100
rect 16008 7040 16072 7044
rect 16088 7100 16152 7104
rect 16088 7044 16092 7100
rect 16092 7044 16148 7100
rect 16148 7044 16152 7100
rect 16088 7040 16152 7044
rect 25778 7100 25842 7104
rect 25778 7044 25782 7100
rect 25782 7044 25838 7100
rect 25838 7044 25842 7100
rect 25778 7040 25842 7044
rect 25858 7100 25922 7104
rect 25858 7044 25862 7100
rect 25862 7044 25918 7100
rect 25918 7044 25922 7100
rect 25858 7040 25922 7044
rect 25938 7100 26002 7104
rect 25938 7044 25942 7100
rect 25942 7044 25998 7100
rect 25998 7044 26002 7100
rect 25938 7040 26002 7044
rect 26018 7100 26082 7104
rect 26018 7044 26022 7100
rect 26022 7044 26078 7100
rect 26078 7044 26082 7100
rect 26018 7040 26082 7044
rect 10882 6556 10946 6560
rect 10882 6500 10886 6556
rect 10886 6500 10942 6556
rect 10942 6500 10946 6556
rect 10882 6496 10946 6500
rect 10962 6556 11026 6560
rect 10962 6500 10966 6556
rect 10966 6500 11022 6556
rect 11022 6500 11026 6556
rect 10962 6496 11026 6500
rect 11042 6556 11106 6560
rect 11042 6500 11046 6556
rect 11046 6500 11102 6556
rect 11102 6500 11106 6556
rect 11042 6496 11106 6500
rect 11122 6556 11186 6560
rect 11122 6500 11126 6556
rect 11126 6500 11182 6556
rect 11182 6500 11186 6556
rect 11122 6496 11186 6500
rect 20813 6556 20877 6560
rect 20813 6500 20817 6556
rect 20817 6500 20873 6556
rect 20873 6500 20877 6556
rect 20813 6496 20877 6500
rect 20893 6556 20957 6560
rect 20893 6500 20897 6556
rect 20897 6500 20953 6556
rect 20953 6500 20957 6556
rect 20893 6496 20957 6500
rect 20973 6556 21037 6560
rect 20973 6500 20977 6556
rect 20977 6500 21033 6556
rect 21033 6500 21037 6556
rect 20973 6496 21037 6500
rect 21053 6556 21117 6560
rect 21053 6500 21057 6556
rect 21057 6500 21113 6556
rect 21113 6500 21117 6556
rect 21053 6496 21117 6500
rect 5917 6012 5981 6016
rect 5917 5956 5921 6012
rect 5921 5956 5977 6012
rect 5977 5956 5981 6012
rect 5917 5952 5981 5956
rect 5997 6012 6061 6016
rect 5997 5956 6001 6012
rect 6001 5956 6057 6012
rect 6057 5956 6061 6012
rect 5997 5952 6061 5956
rect 6077 6012 6141 6016
rect 6077 5956 6081 6012
rect 6081 5956 6137 6012
rect 6137 5956 6141 6012
rect 6077 5952 6141 5956
rect 6157 6012 6221 6016
rect 6157 5956 6161 6012
rect 6161 5956 6217 6012
rect 6217 5956 6221 6012
rect 6157 5952 6221 5956
rect 15848 6012 15912 6016
rect 15848 5956 15852 6012
rect 15852 5956 15908 6012
rect 15908 5956 15912 6012
rect 15848 5952 15912 5956
rect 15928 6012 15992 6016
rect 15928 5956 15932 6012
rect 15932 5956 15988 6012
rect 15988 5956 15992 6012
rect 15928 5952 15992 5956
rect 16008 6012 16072 6016
rect 16008 5956 16012 6012
rect 16012 5956 16068 6012
rect 16068 5956 16072 6012
rect 16008 5952 16072 5956
rect 16088 6012 16152 6016
rect 16088 5956 16092 6012
rect 16092 5956 16148 6012
rect 16148 5956 16152 6012
rect 16088 5952 16152 5956
rect 25778 6012 25842 6016
rect 25778 5956 25782 6012
rect 25782 5956 25838 6012
rect 25838 5956 25842 6012
rect 25778 5952 25842 5956
rect 25858 6012 25922 6016
rect 25858 5956 25862 6012
rect 25862 5956 25918 6012
rect 25918 5956 25922 6012
rect 25858 5952 25922 5956
rect 25938 6012 26002 6016
rect 25938 5956 25942 6012
rect 25942 5956 25998 6012
rect 25998 5956 26002 6012
rect 25938 5952 26002 5956
rect 26018 6012 26082 6016
rect 26018 5956 26022 6012
rect 26022 5956 26078 6012
rect 26078 5956 26082 6012
rect 26018 5952 26082 5956
rect 10882 5468 10946 5472
rect 10882 5412 10886 5468
rect 10886 5412 10942 5468
rect 10942 5412 10946 5468
rect 10882 5408 10946 5412
rect 10962 5468 11026 5472
rect 10962 5412 10966 5468
rect 10966 5412 11022 5468
rect 11022 5412 11026 5468
rect 10962 5408 11026 5412
rect 11042 5468 11106 5472
rect 11042 5412 11046 5468
rect 11046 5412 11102 5468
rect 11102 5412 11106 5468
rect 11042 5408 11106 5412
rect 11122 5468 11186 5472
rect 11122 5412 11126 5468
rect 11126 5412 11182 5468
rect 11182 5412 11186 5468
rect 11122 5408 11186 5412
rect 20813 5468 20877 5472
rect 20813 5412 20817 5468
rect 20817 5412 20873 5468
rect 20873 5412 20877 5468
rect 20813 5408 20877 5412
rect 20893 5468 20957 5472
rect 20893 5412 20897 5468
rect 20897 5412 20953 5468
rect 20953 5412 20957 5468
rect 20893 5408 20957 5412
rect 20973 5468 21037 5472
rect 20973 5412 20977 5468
rect 20977 5412 21033 5468
rect 21033 5412 21037 5468
rect 20973 5408 21037 5412
rect 21053 5468 21117 5472
rect 21053 5412 21057 5468
rect 21057 5412 21113 5468
rect 21113 5412 21117 5468
rect 21053 5408 21117 5412
rect 5917 4924 5981 4928
rect 5917 4868 5921 4924
rect 5921 4868 5977 4924
rect 5977 4868 5981 4924
rect 5917 4864 5981 4868
rect 5997 4924 6061 4928
rect 5997 4868 6001 4924
rect 6001 4868 6057 4924
rect 6057 4868 6061 4924
rect 5997 4864 6061 4868
rect 6077 4924 6141 4928
rect 6077 4868 6081 4924
rect 6081 4868 6137 4924
rect 6137 4868 6141 4924
rect 6077 4864 6141 4868
rect 6157 4924 6221 4928
rect 6157 4868 6161 4924
rect 6161 4868 6217 4924
rect 6217 4868 6221 4924
rect 6157 4864 6221 4868
rect 15848 4924 15912 4928
rect 15848 4868 15852 4924
rect 15852 4868 15908 4924
rect 15908 4868 15912 4924
rect 15848 4864 15912 4868
rect 15928 4924 15992 4928
rect 15928 4868 15932 4924
rect 15932 4868 15988 4924
rect 15988 4868 15992 4924
rect 15928 4864 15992 4868
rect 16008 4924 16072 4928
rect 16008 4868 16012 4924
rect 16012 4868 16068 4924
rect 16068 4868 16072 4924
rect 16008 4864 16072 4868
rect 16088 4924 16152 4928
rect 16088 4868 16092 4924
rect 16092 4868 16148 4924
rect 16148 4868 16152 4924
rect 16088 4864 16152 4868
rect 25778 4924 25842 4928
rect 25778 4868 25782 4924
rect 25782 4868 25838 4924
rect 25838 4868 25842 4924
rect 25778 4864 25842 4868
rect 25858 4924 25922 4928
rect 25858 4868 25862 4924
rect 25862 4868 25918 4924
rect 25918 4868 25922 4924
rect 25858 4864 25922 4868
rect 25938 4924 26002 4928
rect 25938 4868 25942 4924
rect 25942 4868 25998 4924
rect 25998 4868 26002 4924
rect 25938 4864 26002 4868
rect 26018 4924 26082 4928
rect 26018 4868 26022 4924
rect 26022 4868 26078 4924
rect 26078 4868 26082 4924
rect 26018 4864 26082 4868
rect 10882 4380 10946 4384
rect 10882 4324 10886 4380
rect 10886 4324 10942 4380
rect 10942 4324 10946 4380
rect 10882 4320 10946 4324
rect 10962 4380 11026 4384
rect 10962 4324 10966 4380
rect 10966 4324 11022 4380
rect 11022 4324 11026 4380
rect 10962 4320 11026 4324
rect 11042 4380 11106 4384
rect 11042 4324 11046 4380
rect 11046 4324 11102 4380
rect 11102 4324 11106 4380
rect 11042 4320 11106 4324
rect 11122 4380 11186 4384
rect 11122 4324 11126 4380
rect 11126 4324 11182 4380
rect 11182 4324 11186 4380
rect 11122 4320 11186 4324
rect 20813 4380 20877 4384
rect 20813 4324 20817 4380
rect 20817 4324 20873 4380
rect 20873 4324 20877 4380
rect 20813 4320 20877 4324
rect 20893 4380 20957 4384
rect 20893 4324 20897 4380
rect 20897 4324 20953 4380
rect 20953 4324 20957 4380
rect 20893 4320 20957 4324
rect 20973 4380 21037 4384
rect 20973 4324 20977 4380
rect 20977 4324 21033 4380
rect 21033 4324 21037 4380
rect 20973 4320 21037 4324
rect 21053 4380 21117 4384
rect 21053 4324 21057 4380
rect 21057 4324 21113 4380
rect 21113 4324 21117 4380
rect 21053 4320 21117 4324
rect 9076 3980 9140 4044
rect 5917 3836 5981 3840
rect 5917 3780 5921 3836
rect 5921 3780 5977 3836
rect 5977 3780 5981 3836
rect 5917 3776 5981 3780
rect 5997 3836 6061 3840
rect 5997 3780 6001 3836
rect 6001 3780 6057 3836
rect 6057 3780 6061 3836
rect 5997 3776 6061 3780
rect 6077 3836 6141 3840
rect 6077 3780 6081 3836
rect 6081 3780 6137 3836
rect 6137 3780 6141 3836
rect 6077 3776 6141 3780
rect 6157 3836 6221 3840
rect 6157 3780 6161 3836
rect 6161 3780 6217 3836
rect 6217 3780 6221 3836
rect 6157 3776 6221 3780
rect 15848 3836 15912 3840
rect 15848 3780 15852 3836
rect 15852 3780 15908 3836
rect 15908 3780 15912 3836
rect 15848 3776 15912 3780
rect 15928 3836 15992 3840
rect 15928 3780 15932 3836
rect 15932 3780 15988 3836
rect 15988 3780 15992 3836
rect 15928 3776 15992 3780
rect 16008 3836 16072 3840
rect 16008 3780 16012 3836
rect 16012 3780 16068 3836
rect 16068 3780 16072 3836
rect 16008 3776 16072 3780
rect 16088 3836 16152 3840
rect 16088 3780 16092 3836
rect 16092 3780 16148 3836
rect 16148 3780 16152 3836
rect 16088 3776 16152 3780
rect 25778 3836 25842 3840
rect 25778 3780 25782 3836
rect 25782 3780 25838 3836
rect 25838 3780 25842 3836
rect 25778 3776 25842 3780
rect 25858 3836 25922 3840
rect 25858 3780 25862 3836
rect 25862 3780 25918 3836
rect 25918 3780 25922 3836
rect 25858 3776 25922 3780
rect 25938 3836 26002 3840
rect 25938 3780 25942 3836
rect 25942 3780 25998 3836
rect 25998 3780 26002 3836
rect 25938 3776 26002 3780
rect 26018 3836 26082 3840
rect 26018 3780 26022 3836
rect 26022 3780 26078 3836
rect 26078 3780 26082 3836
rect 26018 3776 26082 3780
rect 10882 3292 10946 3296
rect 10882 3236 10886 3292
rect 10886 3236 10942 3292
rect 10942 3236 10946 3292
rect 10882 3232 10946 3236
rect 10962 3292 11026 3296
rect 10962 3236 10966 3292
rect 10966 3236 11022 3292
rect 11022 3236 11026 3292
rect 10962 3232 11026 3236
rect 11042 3292 11106 3296
rect 11042 3236 11046 3292
rect 11046 3236 11102 3292
rect 11102 3236 11106 3292
rect 11042 3232 11106 3236
rect 11122 3292 11186 3296
rect 11122 3236 11126 3292
rect 11126 3236 11182 3292
rect 11182 3236 11186 3292
rect 11122 3232 11186 3236
rect 20813 3292 20877 3296
rect 20813 3236 20817 3292
rect 20817 3236 20873 3292
rect 20873 3236 20877 3292
rect 20813 3232 20877 3236
rect 20893 3292 20957 3296
rect 20893 3236 20897 3292
rect 20897 3236 20953 3292
rect 20953 3236 20957 3292
rect 20893 3232 20957 3236
rect 20973 3292 21037 3296
rect 20973 3236 20977 3292
rect 20977 3236 21033 3292
rect 21033 3236 21037 3292
rect 20973 3232 21037 3236
rect 21053 3292 21117 3296
rect 21053 3236 21057 3292
rect 21057 3236 21113 3292
rect 21113 3236 21117 3292
rect 21053 3232 21117 3236
rect 5917 2748 5981 2752
rect 5917 2692 5921 2748
rect 5921 2692 5977 2748
rect 5977 2692 5981 2748
rect 5917 2688 5981 2692
rect 5997 2748 6061 2752
rect 5997 2692 6001 2748
rect 6001 2692 6057 2748
rect 6057 2692 6061 2748
rect 5997 2688 6061 2692
rect 6077 2748 6141 2752
rect 6077 2692 6081 2748
rect 6081 2692 6137 2748
rect 6137 2692 6141 2748
rect 6077 2688 6141 2692
rect 6157 2748 6221 2752
rect 6157 2692 6161 2748
rect 6161 2692 6217 2748
rect 6217 2692 6221 2748
rect 6157 2688 6221 2692
rect 15848 2748 15912 2752
rect 15848 2692 15852 2748
rect 15852 2692 15908 2748
rect 15908 2692 15912 2748
rect 15848 2688 15912 2692
rect 15928 2748 15992 2752
rect 15928 2692 15932 2748
rect 15932 2692 15988 2748
rect 15988 2692 15992 2748
rect 15928 2688 15992 2692
rect 16008 2748 16072 2752
rect 16008 2692 16012 2748
rect 16012 2692 16068 2748
rect 16068 2692 16072 2748
rect 16008 2688 16072 2692
rect 16088 2748 16152 2752
rect 16088 2692 16092 2748
rect 16092 2692 16148 2748
rect 16148 2692 16152 2748
rect 16088 2688 16152 2692
rect 25778 2748 25842 2752
rect 25778 2692 25782 2748
rect 25782 2692 25838 2748
rect 25838 2692 25842 2748
rect 25778 2688 25842 2692
rect 25858 2748 25922 2752
rect 25858 2692 25862 2748
rect 25862 2692 25918 2748
rect 25918 2692 25922 2748
rect 25858 2688 25922 2692
rect 25938 2748 26002 2752
rect 25938 2692 25942 2748
rect 25942 2692 25998 2748
rect 25998 2692 26002 2748
rect 25938 2688 26002 2692
rect 26018 2748 26082 2752
rect 26018 2692 26022 2748
rect 26022 2692 26078 2748
rect 26078 2692 26082 2748
rect 26018 2688 26082 2692
rect 10882 2204 10946 2208
rect 10882 2148 10886 2204
rect 10886 2148 10942 2204
rect 10942 2148 10946 2204
rect 10882 2144 10946 2148
rect 10962 2204 11026 2208
rect 10962 2148 10966 2204
rect 10966 2148 11022 2204
rect 11022 2148 11026 2204
rect 10962 2144 11026 2148
rect 11042 2204 11106 2208
rect 11042 2148 11046 2204
rect 11046 2148 11102 2204
rect 11102 2148 11106 2204
rect 11042 2144 11106 2148
rect 11122 2204 11186 2208
rect 11122 2148 11126 2204
rect 11126 2148 11182 2204
rect 11182 2148 11186 2204
rect 11122 2144 11186 2148
rect 20813 2204 20877 2208
rect 20813 2148 20817 2204
rect 20817 2148 20873 2204
rect 20873 2148 20877 2204
rect 20813 2144 20877 2148
rect 20893 2204 20957 2208
rect 20893 2148 20897 2204
rect 20897 2148 20953 2204
rect 20953 2148 20957 2204
rect 20893 2144 20957 2148
rect 20973 2204 21037 2208
rect 20973 2148 20977 2204
rect 20977 2148 21033 2204
rect 21033 2148 21037 2204
rect 20973 2144 21037 2148
rect 21053 2204 21117 2208
rect 21053 2148 21057 2204
rect 21057 2148 21113 2204
rect 21113 2148 21117 2204
rect 21053 2144 21117 2148
<< metal4 >>
rect 5909 45184 6229 45744
rect 5909 45120 5917 45184
rect 5981 45120 5997 45184
rect 6061 45120 6077 45184
rect 6141 45120 6157 45184
rect 6221 45120 6229 45184
rect 5909 44096 6229 45120
rect 5909 44032 5917 44096
rect 5981 44032 5997 44096
rect 6061 44032 6077 44096
rect 6141 44032 6157 44096
rect 6221 44032 6229 44096
rect 5909 43008 6229 44032
rect 5909 42944 5917 43008
rect 5981 42944 5997 43008
rect 6061 42944 6077 43008
rect 6141 42944 6157 43008
rect 6221 42944 6229 43008
rect 5909 41920 6229 42944
rect 5909 41856 5917 41920
rect 5981 41856 5997 41920
rect 6061 41856 6077 41920
rect 6141 41856 6157 41920
rect 6221 41856 6229 41920
rect 5909 40832 6229 41856
rect 5909 40768 5917 40832
rect 5981 40768 5997 40832
rect 6061 40768 6077 40832
rect 6141 40768 6157 40832
rect 6221 40768 6229 40832
rect 5909 39744 6229 40768
rect 5909 39680 5917 39744
rect 5981 39680 5997 39744
rect 6061 39680 6077 39744
rect 6141 39680 6157 39744
rect 6221 39680 6229 39744
rect 5909 38656 6229 39680
rect 5909 38592 5917 38656
rect 5981 38592 5997 38656
rect 6061 38592 6077 38656
rect 6141 38592 6157 38656
rect 6221 38592 6229 38656
rect 5909 37568 6229 38592
rect 5909 37504 5917 37568
rect 5981 37504 5997 37568
rect 6061 37504 6077 37568
rect 6141 37504 6157 37568
rect 6221 37504 6229 37568
rect 5909 36480 6229 37504
rect 5909 36416 5917 36480
rect 5981 36416 5997 36480
rect 6061 36416 6077 36480
rect 6141 36416 6157 36480
rect 6221 36416 6229 36480
rect 5909 35392 6229 36416
rect 5909 35328 5917 35392
rect 5981 35328 5997 35392
rect 6061 35328 6077 35392
rect 6141 35328 6157 35392
rect 6221 35328 6229 35392
rect 5909 34304 6229 35328
rect 5909 34240 5917 34304
rect 5981 34240 5997 34304
rect 6061 34240 6077 34304
rect 6141 34240 6157 34304
rect 6221 34240 6229 34304
rect 5909 33216 6229 34240
rect 5909 33152 5917 33216
rect 5981 33152 5997 33216
rect 6061 33152 6077 33216
rect 6141 33152 6157 33216
rect 6221 33152 6229 33216
rect 5909 32128 6229 33152
rect 5909 32064 5917 32128
rect 5981 32064 5997 32128
rect 6061 32064 6077 32128
rect 6141 32064 6157 32128
rect 6221 32064 6229 32128
rect 5909 31040 6229 32064
rect 5909 30976 5917 31040
rect 5981 30976 5997 31040
rect 6061 30976 6077 31040
rect 6141 30976 6157 31040
rect 6221 30976 6229 31040
rect 5909 29952 6229 30976
rect 10874 45728 11194 45744
rect 10874 45664 10882 45728
rect 10946 45664 10962 45728
rect 11026 45664 11042 45728
rect 11106 45664 11122 45728
rect 11186 45664 11194 45728
rect 10874 44640 11194 45664
rect 10874 44576 10882 44640
rect 10946 44576 10962 44640
rect 11026 44576 11042 44640
rect 11106 44576 11122 44640
rect 11186 44576 11194 44640
rect 10874 43552 11194 44576
rect 10874 43488 10882 43552
rect 10946 43488 10962 43552
rect 11026 43488 11042 43552
rect 11106 43488 11122 43552
rect 11186 43488 11194 43552
rect 10874 42464 11194 43488
rect 10874 42400 10882 42464
rect 10946 42400 10962 42464
rect 11026 42400 11042 42464
rect 11106 42400 11122 42464
rect 11186 42400 11194 42464
rect 10874 41376 11194 42400
rect 10874 41312 10882 41376
rect 10946 41312 10962 41376
rect 11026 41312 11042 41376
rect 11106 41312 11122 41376
rect 11186 41312 11194 41376
rect 10874 40288 11194 41312
rect 10874 40224 10882 40288
rect 10946 40224 10962 40288
rect 11026 40224 11042 40288
rect 11106 40224 11122 40288
rect 11186 40224 11194 40288
rect 10874 39200 11194 40224
rect 10874 39136 10882 39200
rect 10946 39136 10962 39200
rect 11026 39136 11042 39200
rect 11106 39136 11122 39200
rect 11186 39136 11194 39200
rect 10874 38112 11194 39136
rect 10874 38048 10882 38112
rect 10946 38048 10962 38112
rect 11026 38048 11042 38112
rect 11106 38048 11122 38112
rect 11186 38048 11194 38112
rect 10874 37024 11194 38048
rect 10874 36960 10882 37024
rect 10946 36960 10962 37024
rect 11026 36960 11042 37024
rect 11106 36960 11122 37024
rect 11186 36960 11194 37024
rect 10874 35936 11194 36960
rect 10874 35872 10882 35936
rect 10946 35872 10962 35936
rect 11026 35872 11042 35936
rect 11106 35872 11122 35936
rect 11186 35872 11194 35936
rect 10874 34848 11194 35872
rect 10874 34784 10882 34848
rect 10946 34784 10962 34848
rect 11026 34784 11042 34848
rect 11106 34784 11122 34848
rect 11186 34784 11194 34848
rect 10874 33760 11194 34784
rect 10874 33696 10882 33760
rect 10946 33696 10962 33760
rect 11026 33696 11042 33760
rect 11106 33696 11122 33760
rect 11186 33696 11194 33760
rect 10874 32672 11194 33696
rect 10874 32608 10882 32672
rect 10946 32608 10962 32672
rect 11026 32608 11042 32672
rect 11106 32608 11122 32672
rect 11186 32608 11194 32672
rect 10874 31584 11194 32608
rect 10874 31520 10882 31584
rect 10946 31520 10962 31584
rect 11026 31520 11042 31584
rect 11106 31520 11122 31584
rect 11186 31520 11194 31584
rect 10874 30496 11194 31520
rect 10874 30432 10882 30496
rect 10946 30432 10962 30496
rect 11026 30432 11042 30496
rect 11106 30432 11122 30496
rect 11186 30432 11194 30496
rect 9075 30428 9141 30429
rect 9075 30364 9076 30428
rect 9140 30364 9141 30428
rect 9075 30363 9141 30364
rect 5909 29888 5917 29952
rect 5981 29888 5997 29952
rect 6061 29888 6077 29952
rect 6141 29888 6157 29952
rect 6221 29888 6229 29952
rect 5909 28864 6229 29888
rect 5909 28800 5917 28864
rect 5981 28800 5997 28864
rect 6061 28800 6077 28864
rect 6141 28800 6157 28864
rect 6221 28800 6229 28864
rect 5909 27776 6229 28800
rect 5909 27712 5917 27776
rect 5981 27712 5997 27776
rect 6061 27712 6077 27776
rect 6141 27712 6157 27776
rect 6221 27712 6229 27776
rect 5909 26688 6229 27712
rect 8339 27436 8405 27437
rect 8339 27372 8340 27436
rect 8404 27372 8405 27436
rect 8339 27371 8405 27372
rect 5909 26624 5917 26688
rect 5981 26624 5997 26688
rect 6061 26624 6077 26688
rect 6141 26624 6157 26688
rect 6221 26624 6229 26688
rect 5909 25600 6229 26624
rect 8342 26349 8402 27371
rect 8339 26348 8405 26349
rect 8339 26284 8340 26348
rect 8404 26284 8405 26348
rect 8339 26283 8405 26284
rect 5909 25536 5917 25600
rect 5981 25536 5997 25600
rect 6061 25536 6077 25600
rect 6141 25536 6157 25600
rect 6221 25536 6229 25600
rect 5909 24512 6229 25536
rect 5909 24448 5917 24512
rect 5981 24448 5997 24512
rect 6061 24448 6077 24512
rect 6141 24448 6157 24512
rect 6221 24448 6229 24512
rect 5909 23424 6229 24448
rect 5909 23360 5917 23424
rect 5981 23360 5997 23424
rect 6061 23360 6077 23424
rect 6141 23360 6157 23424
rect 6221 23360 6229 23424
rect 5909 22336 6229 23360
rect 5909 22272 5917 22336
rect 5981 22272 5997 22336
rect 6061 22272 6077 22336
rect 6141 22272 6157 22336
rect 6221 22272 6229 22336
rect 5909 21248 6229 22272
rect 8342 21997 8402 26283
rect 8339 21996 8405 21997
rect 8339 21932 8340 21996
rect 8404 21932 8405 21996
rect 8339 21931 8405 21932
rect 5909 21184 5917 21248
rect 5981 21184 5997 21248
rect 6061 21184 6077 21248
rect 6141 21184 6157 21248
rect 6221 21184 6229 21248
rect 5909 20160 6229 21184
rect 5909 20096 5917 20160
rect 5981 20096 5997 20160
rect 6061 20096 6077 20160
rect 6141 20096 6157 20160
rect 6221 20096 6229 20160
rect 5909 19072 6229 20096
rect 5909 19008 5917 19072
rect 5981 19008 5997 19072
rect 6061 19008 6077 19072
rect 6141 19008 6157 19072
rect 6221 19008 6229 19072
rect 5909 17984 6229 19008
rect 5909 17920 5917 17984
rect 5981 17920 5997 17984
rect 6061 17920 6077 17984
rect 6141 17920 6157 17984
rect 6221 17920 6229 17984
rect 5909 16896 6229 17920
rect 5909 16832 5917 16896
rect 5981 16832 5997 16896
rect 6061 16832 6077 16896
rect 6141 16832 6157 16896
rect 6221 16832 6229 16896
rect 5763 16012 5829 16013
rect 5763 15948 5764 16012
rect 5828 15948 5829 16012
rect 5763 15947 5829 15948
rect 5766 9077 5826 15947
rect 5909 15808 6229 16832
rect 5909 15744 5917 15808
rect 5981 15744 5997 15808
rect 6061 15744 6077 15808
rect 6141 15744 6157 15808
rect 6221 15744 6229 15808
rect 5909 14720 6229 15744
rect 5909 14656 5917 14720
rect 5981 14656 5997 14720
rect 6061 14656 6077 14720
rect 6141 14656 6157 14720
rect 6221 14656 6229 14720
rect 5909 13632 6229 14656
rect 5909 13568 5917 13632
rect 5981 13568 5997 13632
rect 6061 13568 6077 13632
rect 6141 13568 6157 13632
rect 6221 13568 6229 13632
rect 5909 12544 6229 13568
rect 5909 12480 5917 12544
rect 5981 12480 5997 12544
rect 6061 12480 6077 12544
rect 6141 12480 6157 12544
rect 6221 12480 6229 12544
rect 5909 11456 6229 12480
rect 5909 11392 5917 11456
rect 5981 11392 5997 11456
rect 6061 11392 6077 11456
rect 6141 11392 6157 11456
rect 6221 11392 6229 11456
rect 5909 10368 6229 11392
rect 5909 10304 5917 10368
rect 5981 10304 5997 10368
rect 6061 10304 6077 10368
rect 6141 10304 6157 10368
rect 6221 10304 6229 10368
rect 5909 9280 6229 10304
rect 5909 9216 5917 9280
rect 5981 9216 5997 9280
rect 6061 9216 6077 9280
rect 6141 9216 6157 9280
rect 6221 9216 6229 9280
rect 5763 9076 5829 9077
rect 5763 9012 5764 9076
rect 5828 9012 5829 9076
rect 5763 9011 5829 9012
rect 5909 8192 6229 9216
rect 5909 8128 5917 8192
rect 5981 8128 5997 8192
rect 6061 8128 6077 8192
rect 6141 8128 6157 8192
rect 6221 8128 6229 8192
rect 5909 7104 6229 8128
rect 5909 7040 5917 7104
rect 5981 7040 5997 7104
rect 6061 7040 6077 7104
rect 6141 7040 6157 7104
rect 6221 7040 6229 7104
rect 5909 6016 6229 7040
rect 5909 5952 5917 6016
rect 5981 5952 5997 6016
rect 6061 5952 6077 6016
rect 6141 5952 6157 6016
rect 6221 5952 6229 6016
rect 5909 4928 6229 5952
rect 5909 4864 5917 4928
rect 5981 4864 5997 4928
rect 6061 4864 6077 4928
rect 6141 4864 6157 4928
rect 6221 4864 6229 4928
rect 5909 3840 6229 4864
rect 9078 4045 9138 30363
rect 10874 29408 11194 30432
rect 10874 29344 10882 29408
rect 10946 29344 10962 29408
rect 11026 29344 11042 29408
rect 11106 29344 11122 29408
rect 11186 29344 11194 29408
rect 10874 28320 11194 29344
rect 10874 28256 10882 28320
rect 10946 28256 10962 28320
rect 11026 28256 11042 28320
rect 11106 28256 11122 28320
rect 11186 28256 11194 28320
rect 10874 27232 11194 28256
rect 10874 27168 10882 27232
rect 10946 27168 10962 27232
rect 11026 27168 11042 27232
rect 11106 27168 11122 27232
rect 11186 27168 11194 27232
rect 10874 26144 11194 27168
rect 10874 26080 10882 26144
rect 10946 26080 10962 26144
rect 11026 26080 11042 26144
rect 11106 26080 11122 26144
rect 11186 26080 11194 26144
rect 10874 25056 11194 26080
rect 10874 24992 10882 25056
rect 10946 24992 10962 25056
rect 11026 24992 11042 25056
rect 11106 24992 11122 25056
rect 11186 24992 11194 25056
rect 10874 23968 11194 24992
rect 10874 23904 10882 23968
rect 10946 23904 10962 23968
rect 11026 23904 11042 23968
rect 11106 23904 11122 23968
rect 11186 23904 11194 23968
rect 10874 22880 11194 23904
rect 10874 22816 10882 22880
rect 10946 22816 10962 22880
rect 11026 22816 11042 22880
rect 11106 22816 11122 22880
rect 11186 22816 11194 22880
rect 10874 21792 11194 22816
rect 10874 21728 10882 21792
rect 10946 21728 10962 21792
rect 11026 21728 11042 21792
rect 11106 21728 11122 21792
rect 11186 21728 11194 21792
rect 10874 20704 11194 21728
rect 10874 20640 10882 20704
rect 10946 20640 10962 20704
rect 11026 20640 11042 20704
rect 11106 20640 11122 20704
rect 11186 20640 11194 20704
rect 10874 19616 11194 20640
rect 10874 19552 10882 19616
rect 10946 19552 10962 19616
rect 11026 19552 11042 19616
rect 11106 19552 11122 19616
rect 11186 19552 11194 19616
rect 10874 18528 11194 19552
rect 10874 18464 10882 18528
rect 10946 18464 10962 18528
rect 11026 18464 11042 18528
rect 11106 18464 11122 18528
rect 11186 18464 11194 18528
rect 10874 17440 11194 18464
rect 10874 17376 10882 17440
rect 10946 17376 10962 17440
rect 11026 17376 11042 17440
rect 11106 17376 11122 17440
rect 11186 17376 11194 17440
rect 10874 16352 11194 17376
rect 10874 16288 10882 16352
rect 10946 16288 10962 16352
rect 11026 16288 11042 16352
rect 11106 16288 11122 16352
rect 11186 16288 11194 16352
rect 10874 15264 11194 16288
rect 10874 15200 10882 15264
rect 10946 15200 10962 15264
rect 11026 15200 11042 15264
rect 11106 15200 11122 15264
rect 11186 15200 11194 15264
rect 10874 14176 11194 15200
rect 10874 14112 10882 14176
rect 10946 14112 10962 14176
rect 11026 14112 11042 14176
rect 11106 14112 11122 14176
rect 11186 14112 11194 14176
rect 10874 13088 11194 14112
rect 10874 13024 10882 13088
rect 10946 13024 10962 13088
rect 11026 13024 11042 13088
rect 11106 13024 11122 13088
rect 11186 13024 11194 13088
rect 10874 12000 11194 13024
rect 10874 11936 10882 12000
rect 10946 11936 10962 12000
rect 11026 11936 11042 12000
rect 11106 11936 11122 12000
rect 11186 11936 11194 12000
rect 10874 10912 11194 11936
rect 10874 10848 10882 10912
rect 10946 10848 10962 10912
rect 11026 10848 11042 10912
rect 11106 10848 11122 10912
rect 11186 10848 11194 10912
rect 10874 9824 11194 10848
rect 10874 9760 10882 9824
rect 10946 9760 10962 9824
rect 11026 9760 11042 9824
rect 11106 9760 11122 9824
rect 11186 9760 11194 9824
rect 10874 8736 11194 9760
rect 10874 8672 10882 8736
rect 10946 8672 10962 8736
rect 11026 8672 11042 8736
rect 11106 8672 11122 8736
rect 11186 8672 11194 8736
rect 10874 7648 11194 8672
rect 10874 7584 10882 7648
rect 10946 7584 10962 7648
rect 11026 7584 11042 7648
rect 11106 7584 11122 7648
rect 11186 7584 11194 7648
rect 10874 6560 11194 7584
rect 10874 6496 10882 6560
rect 10946 6496 10962 6560
rect 11026 6496 11042 6560
rect 11106 6496 11122 6560
rect 11186 6496 11194 6560
rect 10874 5472 11194 6496
rect 10874 5408 10882 5472
rect 10946 5408 10962 5472
rect 11026 5408 11042 5472
rect 11106 5408 11122 5472
rect 11186 5408 11194 5472
rect 10874 4384 11194 5408
rect 10874 4320 10882 4384
rect 10946 4320 10962 4384
rect 11026 4320 11042 4384
rect 11106 4320 11122 4384
rect 11186 4320 11194 4384
rect 9075 4044 9141 4045
rect 9075 3980 9076 4044
rect 9140 3980 9141 4044
rect 9075 3979 9141 3980
rect 5909 3776 5917 3840
rect 5981 3776 5997 3840
rect 6061 3776 6077 3840
rect 6141 3776 6157 3840
rect 6221 3776 6229 3840
rect 5909 2752 6229 3776
rect 5909 2688 5917 2752
rect 5981 2688 5997 2752
rect 6061 2688 6077 2752
rect 6141 2688 6157 2752
rect 6221 2688 6229 2752
rect 5909 2128 6229 2688
rect 10874 3296 11194 4320
rect 10874 3232 10882 3296
rect 10946 3232 10962 3296
rect 11026 3232 11042 3296
rect 11106 3232 11122 3296
rect 11186 3232 11194 3296
rect 10874 2208 11194 3232
rect 10874 2144 10882 2208
rect 10946 2144 10962 2208
rect 11026 2144 11042 2208
rect 11106 2144 11122 2208
rect 11186 2144 11194 2208
rect 10874 2128 11194 2144
rect 15839 45184 16160 45744
rect 15839 45120 15848 45184
rect 15912 45120 15928 45184
rect 15992 45120 16008 45184
rect 16072 45120 16088 45184
rect 16152 45120 16160 45184
rect 15839 44096 16160 45120
rect 15839 44032 15848 44096
rect 15912 44032 15928 44096
rect 15992 44032 16008 44096
rect 16072 44032 16088 44096
rect 16152 44032 16160 44096
rect 15839 43008 16160 44032
rect 15839 42944 15848 43008
rect 15912 42944 15928 43008
rect 15992 42944 16008 43008
rect 16072 42944 16088 43008
rect 16152 42944 16160 43008
rect 15839 41920 16160 42944
rect 15839 41856 15848 41920
rect 15912 41856 15928 41920
rect 15992 41856 16008 41920
rect 16072 41856 16088 41920
rect 16152 41856 16160 41920
rect 15839 40832 16160 41856
rect 15839 40768 15848 40832
rect 15912 40768 15928 40832
rect 15992 40768 16008 40832
rect 16072 40768 16088 40832
rect 16152 40768 16160 40832
rect 15839 39744 16160 40768
rect 15839 39680 15848 39744
rect 15912 39680 15928 39744
rect 15992 39680 16008 39744
rect 16072 39680 16088 39744
rect 16152 39680 16160 39744
rect 15839 38656 16160 39680
rect 15839 38592 15848 38656
rect 15912 38592 15928 38656
rect 15992 38592 16008 38656
rect 16072 38592 16088 38656
rect 16152 38592 16160 38656
rect 15839 37568 16160 38592
rect 15839 37504 15848 37568
rect 15912 37504 15928 37568
rect 15992 37504 16008 37568
rect 16072 37504 16088 37568
rect 16152 37504 16160 37568
rect 15839 36480 16160 37504
rect 15839 36416 15848 36480
rect 15912 36416 15928 36480
rect 15992 36416 16008 36480
rect 16072 36416 16088 36480
rect 16152 36416 16160 36480
rect 15839 35392 16160 36416
rect 15839 35328 15848 35392
rect 15912 35328 15928 35392
rect 15992 35328 16008 35392
rect 16072 35328 16088 35392
rect 16152 35328 16160 35392
rect 15839 34304 16160 35328
rect 15839 34240 15848 34304
rect 15912 34240 15928 34304
rect 15992 34240 16008 34304
rect 16072 34240 16088 34304
rect 16152 34240 16160 34304
rect 15839 33216 16160 34240
rect 15839 33152 15848 33216
rect 15912 33152 15928 33216
rect 15992 33152 16008 33216
rect 16072 33152 16088 33216
rect 16152 33152 16160 33216
rect 15839 32128 16160 33152
rect 15839 32064 15848 32128
rect 15912 32064 15928 32128
rect 15992 32064 16008 32128
rect 16072 32064 16088 32128
rect 16152 32064 16160 32128
rect 15839 31040 16160 32064
rect 15839 30976 15848 31040
rect 15912 30976 15928 31040
rect 15992 30976 16008 31040
rect 16072 30976 16088 31040
rect 16152 30976 16160 31040
rect 15839 29952 16160 30976
rect 20805 45728 21125 45744
rect 20805 45664 20813 45728
rect 20877 45664 20893 45728
rect 20957 45664 20973 45728
rect 21037 45664 21053 45728
rect 21117 45664 21125 45728
rect 20805 44640 21125 45664
rect 20805 44576 20813 44640
rect 20877 44576 20893 44640
rect 20957 44576 20973 44640
rect 21037 44576 21053 44640
rect 21117 44576 21125 44640
rect 20805 43552 21125 44576
rect 20805 43488 20813 43552
rect 20877 43488 20893 43552
rect 20957 43488 20973 43552
rect 21037 43488 21053 43552
rect 21117 43488 21125 43552
rect 20805 42464 21125 43488
rect 20805 42400 20813 42464
rect 20877 42400 20893 42464
rect 20957 42400 20973 42464
rect 21037 42400 21053 42464
rect 21117 42400 21125 42464
rect 20805 41376 21125 42400
rect 20805 41312 20813 41376
rect 20877 41312 20893 41376
rect 20957 41312 20973 41376
rect 21037 41312 21053 41376
rect 21117 41312 21125 41376
rect 20805 40288 21125 41312
rect 20805 40224 20813 40288
rect 20877 40224 20893 40288
rect 20957 40224 20973 40288
rect 21037 40224 21053 40288
rect 21117 40224 21125 40288
rect 20805 39200 21125 40224
rect 20805 39136 20813 39200
rect 20877 39136 20893 39200
rect 20957 39136 20973 39200
rect 21037 39136 21053 39200
rect 21117 39136 21125 39200
rect 20805 38112 21125 39136
rect 20805 38048 20813 38112
rect 20877 38048 20893 38112
rect 20957 38048 20973 38112
rect 21037 38048 21053 38112
rect 21117 38048 21125 38112
rect 20805 37024 21125 38048
rect 20805 36960 20813 37024
rect 20877 36960 20893 37024
rect 20957 36960 20973 37024
rect 21037 36960 21053 37024
rect 21117 36960 21125 37024
rect 20805 35936 21125 36960
rect 20805 35872 20813 35936
rect 20877 35872 20893 35936
rect 20957 35872 20973 35936
rect 21037 35872 21053 35936
rect 21117 35872 21125 35936
rect 20805 34848 21125 35872
rect 20805 34784 20813 34848
rect 20877 34784 20893 34848
rect 20957 34784 20973 34848
rect 21037 34784 21053 34848
rect 21117 34784 21125 34848
rect 20805 33760 21125 34784
rect 20805 33696 20813 33760
rect 20877 33696 20893 33760
rect 20957 33696 20973 33760
rect 21037 33696 21053 33760
rect 21117 33696 21125 33760
rect 20805 32672 21125 33696
rect 20805 32608 20813 32672
rect 20877 32608 20893 32672
rect 20957 32608 20973 32672
rect 21037 32608 21053 32672
rect 21117 32608 21125 32672
rect 20805 31584 21125 32608
rect 20805 31520 20813 31584
rect 20877 31520 20893 31584
rect 20957 31520 20973 31584
rect 21037 31520 21053 31584
rect 21117 31520 21125 31584
rect 20805 30496 21125 31520
rect 20805 30432 20813 30496
rect 20877 30432 20893 30496
rect 20957 30432 20973 30496
rect 21037 30432 21053 30496
rect 21117 30432 21125 30496
rect 18275 30020 18341 30021
rect 18275 29956 18276 30020
rect 18340 29956 18341 30020
rect 18275 29955 18341 29956
rect 15839 29888 15848 29952
rect 15912 29888 15928 29952
rect 15992 29888 16008 29952
rect 16072 29888 16088 29952
rect 16152 29888 16160 29952
rect 15839 28864 16160 29888
rect 15839 28800 15848 28864
rect 15912 28800 15928 28864
rect 15992 28800 16008 28864
rect 16072 28800 16088 28864
rect 16152 28800 16160 28864
rect 15839 27776 16160 28800
rect 15839 27712 15848 27776
rect 15912 27712 15928 27776
rect 15992 27712 16008 27776
rect 16072 27712 16088 27776
rect 16152 27712 16160 27776
rect 15839 26688 16160 27712
rect 15839 26624 15848 26688
rect 15912 26624 15928 26688
rect 15992 26624 16008 26688
rect 16072 26624 16088 26688
rect 16152 26624 16160 26688
rect 15839 25600 16160 26624
rect 15839 25536 15848 25600
rect 15912 25536 15928 25600
rect 15992 25536 16008 25600
rect 16072 25536 16088 25600
rect 16152 25536 16160 25600
rect 15839 24512 16160 25536
rect 15839 24448 15848 24512
rect 15912 24448 15928 24512
rect 15992 24448 16008 24512
rect 16072 24448 16088 24512
rect 16152 24448 16160 24512
rect 15839 23424 16160 24448
rect 15839 23360 15848 23424
rect 15912 23360 15928 23424
rect 15992 23360 16008 23424
rect 16072 23360 16088 23424
rect 16152 23360 16160 23424
rect 15839 22336 16160 23360
rect 15839 22272 15848 22336
rect 15912 22272 15928 22336
rect 15992 22272 16008 22336
rect 16072 22272 16088 22336
rect 16152 22272 16160 22336
rect 15839 21248 16160 22272
rect 15839 21184 15848 21248
rect 15912 21184 15928 21248
rect 15992 21184 16008 21248
rect 16072 21184 16088 21248
rect 16152 21184 16160 21248
rect 15839 20160 16160 21184
rect 15839 20096 15848 20160
rect 15912 20096 15928 20160
rect 15992 20096 16008 20160
rect 16072 20096 16088 20160
rect 16152 20096 16160 20160
rect 15839 19072 16160 20096
rect 15839 19008 15848 19072
rect 15912 19008 15928 19072
rect 15992 19008 16008 19072
rect 16072 19008 16088 19072
rect 16152 19008 16160 19072
rect 15839 17984 16160 19008
rect 15839 17920 15848 17984
rect 15912 17920 15928 17984
rect 15992 17920 16008 17984
rect 16072 17920 16088 17984
rect 16152 17920 16160 17984
rect 15839 16896 16160 17920
rect 15839 16832 15848 16896
rect 15912 16832 15928 16896
rect 15992 16832 16008 16896
rect 16072 16832 16088 16896
rect 16152 16832 16160 16896
rect 15839 15808 16160 16832
rect 18278 16149 18338 29955
rect 20805 29408 21125 30432
rect 20805 29344 20813 29408
rect 20877 29344 20893 29408
rect 20957 29344 20973 29408
rect 21037 29344 21053 29408
rect 21117 29344 21125 29408
rect 20805 28320 21125 29344
rect 20805 28256 20813 28320
rect 20877 28256 20893 28320
rect 20957 28256 20973 28320
rect 21037 28256 21053 28320
rect 21117 28256 21125 28320
rect 20805 27232 21125 28256
rect 20805 27168 20813 27232
rect 20877 27168 20893 27232
rect 20957 27168 20973 27232
rect 21037 27168 21053 27232
rect 21117 27168 21125 27232
rect 20805 26144 21125 27168
rect 20805 26080 20813 26144
rect 20877 26080 20893 26144
rect 20957 26080 20973 26144
rect 21037 26080 21053 26144
rect 21117 26080 21125 26144
rect 20805 25056 21125 26080
rect 20805 24992 20813 25056
rect 20877 24992 20893 25056
rect 20957 24992 20973 25056
rect 21037 24992 21053 25056
rect 21117 24992 21125 25056
rect 20805 23968 21125 24992
rect 20805 23904 20813 23968
rect 20877 23904 20893 23968
rect 20957 23904 20973 23968
rect 21037 23904 21053 23968
rect 21117 23904 21125 23968
rect 20805 22880 21125 23904
rect 20805 22816 20813 22880
rect 20877 22816 20893 22880
rect 20957 22816 20973 22880
rect 21037 22816 21053 22880
rect 21117 22816 21125 22880
rect 20805 21792 21125 22816
rect 20805 21728 20813 21792
rect 20877 21728 20893 21792
rect 20957 21728 20973 21792
rect 21037 21728 21053 21792
rect 21117 21728 21125 21792
rect 20805 20704 21125 21728
rect 20805 20640 20813 20704
rect 20877 20640 20893 20704
rect 20957 20640 20973 20704
rect 21037 20640 21053 20704
rect 21117 20640 21125 20704
rect 20805 19616 21125 20640
rect 20805 19552 20813 19616
rect 20877 19552 20893 19616
rect 20957 19552 20973 19616
rect 21037 19552 21053 19616
rect 21117 19552 21125 19616
rect 20805 18528 21125 19552
rect 20805 18464 20813 18528
rect 20877 18464 20893 18528
rect 20957 18464 20973 18528
rect 21037 18464 21053 18528
rect 21117 18464 21125 18528
rect 20805 17440 21125 18464
rect 20805 17376 20813 17440
rect 20877 17376 20893 17440
rect 20957 17376 20973 17440
rect 21037 17376 21053 17440
rect 21117 17376 21125 17440
rect 20805 16352 21125 17376
rect 20805 16288 20813 16352
rect 20877 16288 20893 16352
rect 20957 16288 20973 16352
rect 21037 16288 21053 16352
rect 21117 16288 21125 16352
rect 18275 16148 18341 16149
rect 18275 16084 18276 16148
rect 18340 16084 18341 16148
rect 18275 16083 18341 16084
rect 15839 15744 15848 15808
rect 15912 15744 15928 15808
rect 15992 15744 16008 15808
rect 16072 15744 16088 15808
rect 16152 15744 16160 15808
rect 15839 14720 16160 15744
rect 15839 14656 15848 14720
rect 15912 14656 15928 14720
rect 15992 14656 16008 14720
rect 16072 14656 16088 14720
rect 16152 14656 16160 14720
rect 15839 13632 16160 14656
rect 15839 13568 15848 13632
rect 15912 13568 15928 13632
rect 15992 13568 16008 13632
rect 16072 13568 16088 13632
rect 16152 13568 16160 13632
rect 15839 12544 16160 13568
rect 15839 12480 15848 12544
rect 15912 12480 15928 12544
rect 15992 12480 16008 12544
rect 16072 12480 16088 12544
rect 16152 12480 16160 12544
rect 15839 11456 16160 12480
rect 15839 11392 15848 11456
rect 15912 11392 15928 11456
rect 15992 11392 16008 11456
rect 16072 11392 16088 11456
rect 16152 11392 16160 11456
rect 15839 10368 16160 11392
rect 15839 10304 15848 10368
rect 15912 10304 15928 10368
rect 15992 10304 16008 10368
rect 16072 10304 16088 10368
rect 16152 10304 16160 10368
rect 15839 9280 16160 10304
rect 15839 9216 15848 9280
rect 15912 9216 15928 9280
rect 15992 9216 16008 9280
rect 16072 9216 16088 9280
rect 16152 9216 16160 9280
rect 15839 8192 16160 9216
rect 15839 8128 15848 8192
rect 15912 8128 15928 8192
rect 15992 8128 16008 8192
rect 16072 8128 16088 8192
rect 16152 8128 16160 8192
rect 15839 7104 16160 8128
rect 15839 7040 15848 7104
rect 15912 7040 15928 7104
rect 15992 7040 16008 7104
rect 16072 7040 16088 7104
rect 16152 7040 16160 7104
rect 15839 6016 16160 7040
rect 15839 5952 15848 6016
rect 15912 5952 15928 6016
rect 15992 5952 16008 6016
rect 16072 5952 16088 6016
rect 16152 5952 16160 6016
rect 15839 4928 16160 5952
rect 15839 4864 15848 4928
rect 15912 4864 15928 4928
rect 15992 4864 16008 4928
rect 16072 4864 16088 4928
rect 16152 4864 16160 4928
rect 15839 3840 16160 4864
rect 15839 3776 15848 3840
rect 15912 3776 15928 3840
rect 15992 3776 16008 3840
rect 16072 3776 16088 3840
rect 16152 3776 16160 3840
rect 15839 2752 16160 3776
rect 15839 2688 15848 2752
rect 15912 2688 15928 2752
rect 15992 2688 16008 2752
rect 16072 2688 16088 2752
rect 16152 2688 16160 2752
rect 15839 2128 16160 2688
rect 20805 15264 21125 16288
rect 20805 15200 20813 15264
rect 20877 15200 20893 15264
rect 20957 15200 20973 15264
rect 21037 15200 21053 15264
rect 21117 15200 21125 15264
rect 20805 14176 21125 15200
rect 20805 14112 20813 14176
rect 20877 14112 20893 14176
rect 20957 14112 20973 14176
rect 21037 14112 21053 14176
rect 21117 14112 21125 14176
rect 20805 13088 21125 14112
rect 20805 13024 20813 13088
rect 20877 13024 20893 13088
rect 20957 13024 20973 13088
rect 21037 13024 21053 13088
rect 21117 13024 21125 13088
rect 20805 12000 21125 13024
rect 20805 11936 20813 12000
rect 20877 11936 20893 12000
rect 20957 11936 20973 12000
rect 21037 11936 21053 12000
rect 21117 11936 21125 12000
rect 20805 10912 21125 11936
rect 20805 10848 20813 10912
rect 20877 10848 20893 10912
rect 20957 10848 20973 10912
rect 21037 10848 21053 10912
rect 21117 10848 21125 10912
rect 20805 9824 21125 10848
rect 20805 9760 20813 9824
rect 20877 9760 20893 9824
rect 20957 9760 20973 9824
rect 21037 9760 21053 9824
rect 21117 9760 21125 9824
rect 20805 8736 21125 9760
rect 20805 8672 20813 8736
rect 20877 8672 20893 8736
rect 20957 8672 20973 8736
rect 21037 8672 21053 8736
rect 21117 8672 21125 8736
rect 20805 7648 21125 8672
rect 20805 7584 20813 7648
rect 20877 7584 20893 7648
rect 20957 7584 20973 7648
rect 21037 7584 21053 7648
rect 21117 7584 21125 7648
rect 20805 6560 21125 7584
rect 20805 6496 20813 6560
rect 20877 6496 20893 6560
rect 20957 6496 20973 6560
rect 21037 6496 21053 6560
rect 21117 6496 21125 6560
rect 20805 5472 21125 6496
rect 20805 5408 20813 5472
rect 20877 5408 20893 5472
rect 20957 5408 20973 5472
rect 21037 5408 21053 5472
rect 21117 5408 21125 5472
rect 20805 4384 21125 5408
rect 20805 4320 20813 4384
rect 20877 4320 20893 4384
rect 20957 4320 20973 4384
rect 21037 4320 21053 4384
rect 21117 4320 21125 4384
rect 20805 3296 21125 4320
rect 20805 3232 20813 3296
rect 20877 3232 20893 3296
rect 20957 3232 20973 3296
rect 21037 3232 21053 3296
rect 21117 3232 21125 3296
rect 20805 2208 21125 3232
rect 20805 2144 20813 2208
rect 20877 2144 20893 2208
rect 20957 2144 20973 2208
rect 21037 2144 21053 2208
rect 21117 2144 21125 2208
rect 20805 2128 21125 2144
rect 25770 45184 26090 45744
rect 25770 45120 25778 45184
rect 25842 45120 25858 45184
rect 25922 45120 25938 45184
rect 26002 45120 26018 45184
rect 26082 45120 26090 45184
rect 25770 44096 26090 45120
rect 25770 44032 25778 44096
rect 25842 44032 25858 44096
rect 25922 44032 25938 44096
rect 26002 44032 26018 44096
rect 26082 44032 26090 44096
rect 25770 43008 26090 44032
rect 25770 42944 25778 43008
rect 25842 42944 25858 43008
rect 25922 42944 25938 43008
rect 26002 42944 26018 43008
rect 26082 42944 26090 43008
rect 25770 41920 26090 42944
rect 25770 41856 25778 41920
rect 25842 41856 25858 41920
rect 25922 41856 25938 41920
rect 26002 41856 26018 41920
rect 26082 41856 26090 41920
rect 25770 40832 26090 41856
rect 25770 40768 25778 40832
rect 25842 40768 25858 40832
rect 25922 40768 25938 40832
rect 26002 40768 26018 40832
rect 26082 40768 26090 40832
rect 25770 39744 26090 40768
rect 25770 39680 25778 39744
rect 25842 39680 25858 39744
rect 25922 39680 25938 39744
rect 26002 39680 26018 39744
rect 26082 39680 26090 39744
rect 25770 38656 26090 39680
rect 25770 38592 25778 38656
rect 25842 38592 25858 38656
rect 25922 38592 25938 38656
rect 26002 38592 26018 38656
rect 26082 38592 26090 38656
rect 25770 37568 26090 38592
rect 25770 37504 25778 37568
rect 25842 37504 25858 37568
rect 25922 37504 25938 37568
rect 26002 37504 26018 37568
rect 26082 37504 26090 37568
rect 25770 36480 26090 37504
rect 25770 36416 25778 36480
rect 25842 36416 25858 36480
rect 25922 36416 25938 36480
rect 26002 36416 26018 36480
rect 26082 36416 26090 36480
rect 25770 35392 26090 36416
rect 25770 35328 25778 35392
rect 25842 35328 25858 35392
rect 25922 35328 25938 35392
rect 26002 35328 26018 35392
rect 26082 35328 26090 35392
rect 25770 34304 26090 35328
rect 25770 34240 25778 34304
rect 25842 34240 25858 34304
rect 25922 34240 25938 34304
rect 26002 34240 26018 34304
rect 26082 34240 26090 34304
rect 25770 33216 26090 34240
rect 25770 33152 25778 33216
rect 25842 33152 25858 33216
rect 25922 33152 25938 33216
rect 26002 33152 26018 33216
rect 26082 33152 26090 33216
rect 25770 32128 26090 33152
rect 25770 32064 25778 32128
rect 25842 32064 25858 32128
rect 25922 32064 25938 32128
rect 26002 32064 26018 32128
rect 26082 32064 26090 32128
rect 25770 31040 26090 32064
rect 25770 30976 25778 31040
rect 25842 30976 25858 31040
rect 25922 30976 25938 31040
rect 26002 30976 26018 31040
rect 26082 30976 26090 31040
rect 25770 29952 26090 30976
rect 25770 29888 25778 29952
rect 25842 29888 25858 29952
rect 25922 29888 25938 29952
rect 26002 29888 26018 29952
rect 26082 29888 26090 29952
rect 25770 28864 26090 29888
rect 25770 28800 25778 28864
rect 25842 28800 25858 28864
rect 25922 28800 25938 28864
rect 26002 28800 26018 28864
rect 26082 28800 26090 28864
rect 25770 27776 26090 28800
rect 25770 27712 25778 27776
rect 25842 27712 25858 27776
rect 25922 27712 25938 27776
rect 26002 27712 26018 27776
rect 26082 27712 26090 27776
rect 25770 26688 26090 27712
rect 25770 26624 25778 26688
rect 25842 26624 25858 26688
rect 25922 26624 25938 26688
rect 26002 26624 26018 26688
rect 26082 26624 26090 26688
rect 25770 25600 26090 26624
rect 25770 25536 25778 25600
rect 25842 25536 25858 25600
rect 25922 25536 25938 25600
rect 26002 25536 26018 25600
rect 26082 25536 26090 25600
rect 25770 24512 26090 25536
rect 25770 24448 25778 24512
rect 25842 24448 25858 24512
rect 25922 24448 25938 24512
rect 26002 24448 26018 24512
rect 26082 24448 26090 24512
rect 25770 23424 26090 24448
rect 25770 23360 25778 23424
rect 25842 23360 25858 23424
rect 25922 23360 25938 23424
rect 26002 23360 26018 23424
rect 26082 23360 26090 23424
rect 25770 22336 26090 23360
rect 25770 22272 25778 22336
rect 25842 22272 25858 22336
rect 25922 22272 25938 22336
rect 26002 22272 26018 22336
rect 26082 22272 26090 22336
rect 25770 21248 26090 22272
rect 25770 21184 25778 21248
rect 25842 21184 25858 21248
rect 25922 21184 25938 21248
rect 26002 21184 26018 21248
rect 26082 21184 26090 21248
rect 25770 20160 26090 21184
rect 25770 20096 25778 20160
rect 25842 20096 25858 20160
rect 25922 20096 25938 20160
rect 26002 20096 26018 20160
rect 26082 20096 26090 20160
rect 25770 19072 26090 20096
rect 25770 19008 25778 19072
rect 25842 19008 25858 19072
rect 25922 19008 25938 19072
rect 26002 19008 26018 19072
rect 26082 19008 26090 19072
rect 25770 17984 26090 19008
rect 25770 17920 25778 17984
rect 25842 17920 25858 17984
rect 25922 17920 25938 17984
rect 26002 17920 26018 17984
rect 26082 17920 26090 17984
rect 25770 16896 26090 17920
rect 25770 16832 25778 16896
rect 25842 16832 25858 16896
rect 25922 16832 25938 16896
rect 26002 16832 26018 16896
rect 26082 16832 26090 16896
rect 25770 15808 26090 16832
rect 25770 15744 25778 15808
rect 25842 15744 25858 15808
rect 25922 15744 25938 15808
rect 26002 15744 26018 15808
rect 26082 15744 26090 15808
rect 25770 14720 26090 15744
rect 25770 14656 25778 14720
rect 25842 14656 25858 14720
rect 25922 14656 25938 14720
rect 26002 14656 26018 14720
rect 26082 14656 26090 14720
rect 25770 13632 26090 14656
rect 25770 13568 25778 13632
rect 25842 13568 25858 13632
rect 25922 13568 25938 13632
rect 26002 13568 26018 13632
rect 26082 13568 26090 13632
rect 25770 12544 26090 13568
rect 25770 12480 25778 12544
rect 25842 12480 25858 12544
rect 25922 12480 25938 12544
rect 26002 12480 26018 12544
rect 26082 12480 26090 12544
rect 25770 11456 26090 12480
rect 25770 11392 25778 11456
rect 25842 11392 25858 11456
rect 25922 11392 25938 11456
rect 26002 11392 26018 11456
rect 26082 11392 26090 11456
rect 25770 10368 26090 11392
rect 25770 10304 25778 10368
rect 25842 10304 25858 10368
rect 25922 10304 25938 10368
rect 26002 10304 26018 10368
rect 26082 10304 26090 10368
rect 25770 9280 26090 10304
rect 25770 9216 25778 9280
rect 25842 9216 25858 9280
rect 25922 9216 25938 9280
rect 26002 9216 26018 9280
rect 26082 9216 26090 9280
rect 25770 8192 26090 9216
rect 25770 8128 25778 8192
rect 25842 8128 25858 8192
rect 25922 8128 25938 8192
rect 26002 8128 26018 8192
rect 26082 8128 26090 8192
rect 25770 7104 26090 8128
rect 25770 7040 25778 7104
rect 25842 7040 25858 7104
rect 25922 7040 25938 7104
rect 26002 7040 26018 7104
rect 26082 7040 26090 7104
rect 25770 6016 26090 7040
rect 25770 5952 25778 6016
rect 25842 5952 25858 6016
rect 25922 5952 25938 6016
rect 26002 5952 26018 6016
rect 26082 5952 26090 6016
rect 25770 4928 26090 5952
rect 25770 4864 25778 4928
rect 25842 4864 25858 4928
rect 25922 4864 25938 4928
rect 26002 4864 26018 4928
rect 26082 4864 26090 4928
rect 25770 3840 26090 4864
rect 25770 3776 25778 3840
rect 25842 3776 25858 3840
rect 25922 3776 25938 3840
rect 26002 3776 26018 3840
rect 26082 3776 26090 3840
rect 25770 2752 26090 3776
rect 25770 2688 25778 2752
rect 25842 2688 25858 2752
rect 25922 2688 25938 2752
rect 26002 2688 26018 2752
rect 26082 2688 26090 2752
rect 25770 2128 26090 2688
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1635444444
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input45 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1635444444
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input67
timestamp 1635444444
transform 1 0 2668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1635444444
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22
timestamp 1635444444
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp 1635444444
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1635444444
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3220 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1901_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3956 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 4968 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input82
timestamp 1635444444
transform 1 0 4048 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1635444444
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1635444444
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1635444444
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1635444444
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1635444444
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1635444444
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60
timestamp 1635444444
transform 1 0 6624 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1635444444
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1635444444
transform -1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1635444444
transform -1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_70
timestamp 1635444444
transform 1 0 7544 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66
timestamp 1635444444
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71
timestamp 1635444444
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635444444
transform -1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0881_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8372 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1635444444
transform 1 0 8280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1635444444
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1635444444
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1635444444
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1635444444
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102
timestamp 1635444444
transform 1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1635444444
transform 1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1635444444
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1956_
timestamp 1635444444
transform 1 0 9384 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1635444444
transform 1 0 9568 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1635444444
transform 1 0 11500 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 12052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1635444444
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1635444444
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_119
timestamp 1635444444
transform 1 0 12052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1635444444
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  input38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1015_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 13340 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_125
timestamp 1635444444
transform 1 0 12604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123
timestamp 1635444444
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1635444444
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 13800 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1635444444
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_137
timestamp 1635444444
transform 1 0 13708 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1635444444
transform 1 0 13340 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1635444444
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_147
timestamp 1635444444
transform 1 0 14628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_147
timestamp 1635444444
transform 1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1515_
timestamp 1635444444
transform -1 0 15548 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1258_
timestamp 1635444444
transform -1 0 15548 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_157
timestamp 1635444444
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_157
timestamp 1635444444
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1635444444
transform -1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1635444444
transform -1 0 16192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1635444444
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1635444444
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1635444444
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1516_
timestamp 1635444444
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1635444444
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1635444444
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_172
timestamp 1635444444
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1635444444
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1635444444
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_175
timestamp 1635444444
transform 1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1635444444
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1635444444
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _1259_
timestamp 1635444444
transform -1 0 17848 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1520_
timestamp 1635444444
transform 1 0 18216 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1759_
timestamp 1635444444
transform 1 0 17572 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1760_
timestamp 1635444444
transform 1 0 18768 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_200
timestamp 1635444444
transform 1 0 19504 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_214
timestamp 1635444444
transform 1 0 20792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_201
timestamp 1635444444
transform 1 0 19596 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215
timestamp 1635444444
transform 1 0 20884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1009_
timestamp 1635444444
transform 1 0 20240 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 20148 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1635444444
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 22264 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1008_
timestamp 1635444444
transform -1 0 22540 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1635444444
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1635444444
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1635444444
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1635444444
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1635444444
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_233
timestamp 1635444444
transform 1 0 22540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1635444444
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1635444444
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1635444444
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1635444444
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1635444444
transform 1 0 24196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1635444444
transform 1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1635444444
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1635444444
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244
timestamp 1635444444
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1635444444
transform 1 0 25024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1635444444
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1635444444
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_256
timestamp 1635444444
transform 1 0 24656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_254 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 24472 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1635444444
transform 1 0 25668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_270
timestamp 1635444444
transform 1 0 25944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_263
timestamp 1635444444
transform 1 0 25300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1635444444
transform -1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1635444444
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1635444444
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp 1635444444
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1635444444
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1635444444
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_266
timestamp 1635444444
transform 1 0 25576 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1635444444
transform 1 0 27600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 1635444444
transform -1 0 27784 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_290
timestamp 1635444444
transform 1 0 27784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_291
timestamp 1635444444
transform 1 0 27876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_284
timestamp 1635444444
transform 1 0 27232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1635444444
transform 1 0 28704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1012_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 28152 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_1_299
timestamp 1635444444
transform 1 0 28612 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_299
timestamp 1635444444
transform 1 0 28612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1635444444
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_309
timestamp 1635444444
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_316
timestamp 1635444444
transform 1 0 30176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_316
timestamp 1635444444
transform 1 0 30176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635444444
transform -1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635444444
transform -1 0 30820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1635444444
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__or4bb_1  _1010_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 30176 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1635444444
transform 1 0 29808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1635444444
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1635444444
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635444444
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1635444444
transform 1 0 1748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1635444444
transform 1 0 2668 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1635444444
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1635444444
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_32
timestamp 1635444444
transform 1 0 4048 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_40
timestamp 1635444444
transform 1 0 4784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1635444444
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1635444444
transform 1 0 5060 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1635444444
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_59
timestamp 1635444444
transform 1 0 6532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_71
timestamp 1635444444
transform 1 0 7636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1635444444
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1635444444
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1635444444
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_107
timestamp 1635444444
transform 1 0 10948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1955_
timestamp 1635444444
transform 1 0 9476 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1635444444
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _1264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 11868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _1372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 12236 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_2_134
timestamp 1635444444
transform 1 0 13432 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_151
timestamp 1635444444
transform 1 0 14996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1635444444
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1512_
timestamp 1635444444
transform 1 0 14076 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_2_157
timestamp 1635444444
transform 1 0 15548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1635444444
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1756_
timestamp 1635444444
transform 1 0 15640 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1758_
timestamp 1635444444
transform 1 0 16836 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1635444444
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1635444444
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1635444444
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1518_
timestamp 1635444444
transform -1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1635444444
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_208
timestamp 1635444444
transform 1 0 20240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_217
timestamp 1635444444
transform 1 0 21068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1013_
timestamp 1635444444
transform -1 0 21068 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 19412 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_226
timestamp 1635444444
transform 1 0 21896 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_233
timestamp 1635444444
transform 1 0 22540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_240
timestamp 1635444444
transform 1 0 23184 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1014_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 21896 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1635444444
transform 1 0 22264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1635444444
transform 1 0 22908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1635444444
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1635444444
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1635444444
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1635444444
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_289
timestamp 1635444444
transform 1 0 27692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1635444444
transform 1 0 28152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1635444444
transform 1 0 28520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1635444444
transform 1 0 28888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1635444444
transform 1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1635444444
transform 1 0 28612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_312
timestamp 1635444444
transform 1 0 29808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635444444
transform -1 0 30820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1635444444
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1635444444
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1635444444
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_21
timestamp 1635444444
transform 1 0 3036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1635444444
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635444444
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1635444444
transform 1 0 1748 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1635444444
transform 1 0 2668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_28
timestamp 1635444444
transform 1 0 3680 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_43
timestamp 1635444444
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _1172_
timestamp 1635444444
transform 1 0 4232 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1635444444
transform -1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1635444444
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1635444444
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1635444444
transform 1 0 6348 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_3_73
timestamp 1635444444
transform 1 0 7820 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_81
timestamp 1635444444
transform 1 0 8556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1076_
timestamp 1635444444
transform 1 0 8832 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_101
timestamp 1635444444
transform 1 0 10396 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1635444444
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 1635444444
transform 1 0 9660 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_97
timestamp 1635444444
transform 1 0 10028 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1376_
timestamp 1635444444
transform 1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp 1635444444
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_124
timestamp 1635444444
transform 1 0 12512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1635444444
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or3_1  _1016_
timestamp 1635444444
transform 1 0 12052 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 13248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1635444444
transform 1 0 13248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_136
timestamp 1635444444
transform 1 0 13616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1635444444
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1513_
timestamp 1635444444
transform -1 0 14628 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1754_
timestamp 1635444444
transform 1 0 14996 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1635444444
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1635444444
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1757_
timestamp 1635444444
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_178
timestamp 1635444444
transform 1 0 17480 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_186
timestamp 1635444444
transform 1 0 18216 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1635444444
transform 1 0 18400 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_204
timestamp 1635444444
transform 1 0 19872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1635444444
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1100_
timestamp 1635444444
transform 1 0 20240 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1635444444
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1635444444
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1635444444
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1635444444
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1635444444
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1635444444
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1635444444
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1635444444
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1635444444
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1635444444
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_293
timestamp 1635444444
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_297
timestamp 1635444444
transform 1 0 28428 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_301
timestamp 1635444444
transform 1 0 28796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1635444444
transform -1 0 29440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1635444444
transform -1 0 28796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_308
timestamp 1635444444
transform 1 0 29440 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_316
timestamp 1635444444
transform 1 0 30176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635444444
transform -1 0 30820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1635444444
transform 1 0 29808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1635444444
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1635444444
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635444444
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1635444444
transform 1 0 1380 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1635444444
transform -1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1635444444
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp 1635444444
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1635444444
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1635444444
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1174_
timestamp 1635444444
transform -1 0 5980 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1177_
timestamp 1635444444
transform 1 0 6348 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_66
timestamp 1635444444
transform 1 0 7176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_70
timestamp 1635444444
transform 1 0 7544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1635444444
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1635444444
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1077_
timestamp 1635444444
transform 1 0 8924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1078_
timestamp 1635444444
transform 1 0 7636 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1635444444
transform 1 0 10488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_107
timestamp 1635444444
transform 1 0 10948 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_94
timestamp 1635444444
transform 1 0 9752 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1635444444
transform 1 0 10672 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_116
timestamp 1635444444
transform 1 0 11776 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_124
timestamp 1635444444
transform 1 0 12512 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _1261_
timestamp 1635444444
transform -1 0 11776 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1501_
timestamp 1635444444
transform -1 0 13616 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1635444444
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_141
timestamp 1635444444
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1635444444
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1635444444
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14352 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1755_
timestamp 1635444444
transform 1 0 15088 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_161
timestamp 1635444444
transform 1 0 15916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_171
timestamp 1635444444
transform 1 0 16836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1517_
timestamp 1635444444
transform 1 0 16284 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_178
timestamp 1635444444
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_182
timestamp 1635444444
transform 1 0 17848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1635444444
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1635444444
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1102_
timestamp 1635444444
transform 1 0 17940 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1635444444
transform 1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1635444444
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_217
timestamp 1635444444
transform 1 0 21068 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1635444444
transform 1 0 19596 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_4_229
timestamp 1635444444
transform 1 0 22172 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1635444444
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1635444444
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1635444444
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1635444444
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1635444444
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1635444444
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1635444444
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1635444444
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1635444444
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp 1635444444
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_316
timestamp 1635444444
transform 1 0 30176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635444444
transform -1 0 30820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1635444444
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1635444444
transform 1 0 29900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1635444444
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635444444
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1166_
timestamp 1635444444
transform -1 0 3496 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1635444444
transform 1 0 1380 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_5_26
timestamp 1635444444
transform 1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_30
timestamp 1635444444
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_40
timestamp 1635444444
transform 1 0 4784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1169_
timestamp 1635444444
transform 1 0 3956 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1635444444
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1635444444
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp 1635444444
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1635444444
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1635444444
transform -1 0 8096 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1635444444
transform 1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_76
timestamp 1635444444
transform 1 0 8096 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1954_
timestamp 1635444444
transform 1 0 8464 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_104
timestamp 1635444444
transform 1 0 10672 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1635444444
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_96
timestamp 1635444444
transform 1 0 9936 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1635444444
transform -1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1635444444
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_120
timestamp 1635444444
transform 1 0 12144 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_128
timestamp 1635444444
transform 1 0 12880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1635444444
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1504_
timestamp 1635444444
transform 1 0 11592 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1751_
timestamp 1635444444
transform 1 0 12972 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_138
timestamp 1635444444
transform 1 0 13800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_146
timestamp 1635444444
transform 1 0 14536 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1109_
timestamp 1635444444
transform -1 0 15916 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1502_
timestamp 1635444444
transform -1 0 14536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1635444444
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1635444444
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1635444444
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1635444444
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1635444444
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1519_
timestamp 1635444444
transform 1 0 17112 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_180
timestamp 1635444444
transform 1 0 17664 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_190
timestamp 1635444444
transform 1 0 18584 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1521_
timestamp 1635444444
transform -1 0 18584 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_202
timestamp 1635444444
transform 1 0 19688 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1944_
timestamp 1635444444
transform -1 0 21344 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1635444444
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1635444444
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1635444444
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1635444444
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1635444444
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1635444444
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1635444444
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1635444444
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1635444444
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1635444444
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1635444444
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_305
timestamp 1635444444
transform 1 0 29164 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_311
timestamp 1635444444
transform 1 0 29716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_316
timestamp 1635444444
transform 1 0 30176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635444444
transform -1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1635444444
transform 1 0 29808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1635444444
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1635444444
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_21
timestamp 1635444444
transform 1 0 3036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1635444444
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635444444
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635444444
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1635444444
transform 1 0 1840 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1635444444
transform 1 0 1564 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1635444444
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1635444444
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_29
timestamp 1635444444
transform 1 0 3772 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1635444444
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1635444444
transform 1 0 4140 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1635444444
transform 1 0 3956 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_6_49
timestamp 1635444444
transform 1 0 5612 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_55
timestamp 1635444444
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1635444444
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1635444444
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1635444444
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_63
timestamp 1635444444
transform 1 0 6900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1635444444
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1176_
timestamp 1635444444
transform 1 0 6256 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_1  _1647_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 6900 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1635444444
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1635444444
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1635444444
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_73
timestamp 1635444444
transform 1 0 7820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_79
timestamp 1635444444
transform 1 0 8372 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_84
timestamp 1635444444
transform 1 0 8832 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1635444444
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_1  _1662_
timestamp 1635444444
transform -1 0 7820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_wb_clk_i
timestamp 1635444444
transform 1 0 8464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1635444444
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_101
timestamp 1635444444
transform 1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1635444444
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_90
timestamp 1635444444
transform 1 0 9384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1074_
timestamp 1635444444
transform -1 0 10396 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_2  _1828_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 11592 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _1746_
timestamp 1635444444
transform 1 0 11960 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1508_
timestamp 1635444444
transform 1 0 11868 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1635444444
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1635444444
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_114
timestamp 1635444444
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1503_
timestamp 1635444444
transform -1 0 13984 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_7_129
timestamp 1635444444
transform 1 0 12972 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_123
timestamp 1635444444
transform 1 0 12420 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_127
timestamp 1635444444
transform 1 0 12788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1254_
timestamp 1635444444
transform -1 0 13616 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1635444444
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_147
timestamp 1635444444
transform 1 0 14628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_140
timestamp 1635444444
transform 1 0 13984 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1635444444
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1510_
timestamp 1635444444
transform -1 0 14628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1635444444
transform 1 0 14352 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1635444444
transform 1 0 14996 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1635444444
transform 1 0 15272 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_174
timestamp 1635444444
transform 1 0 17112 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1635444444
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1635444444
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1937_
timestamp 1635444444
transform 1 0 15640 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1940_
timestamp 1635444444
transform -1 0 18124 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_6_187
timestamp 1635444444
transform 1 0 18308 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1635444444
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_185
timestamp 1635444444
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1635444444
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1104_
timestamp 1635444444
transform 1 0 17480 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1635444444
transform -1 0 19964 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_207
timestamp 1635444444
transform 1 0 20148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_214
timestamp 1635444444
transform 1 0 20792 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_205
timestamp 1635444444
transform 1 0 19964 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1635444444
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1096_
timestamp 1635444444
transform 1 0 20332 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1099_
timestamp 1635444444
transform 1 0 19228 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1690_
timestamp 1635444444
transform -1 0 20792 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_226
timestamp 1635444444
transform 1 0 21896 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_238
timestamp 1635444444
transform 1 0 23000 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1635444444
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1635444444
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1635444444
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1635444444
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1635444444
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1635444444
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1635444444
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1635444444
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1635444444
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1635444444
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1635444444
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1635444444
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1635444444
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1635444444
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1635444444
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1635444444
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1635444444
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1635444444
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1635444444
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp 1635444444
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_316
timestamp 1635444444
transform 1 0 30176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_317
timestamp 1635444444
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635444444
transform -1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635444444
transform -1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1635444444
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 29808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1635444444
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_19
timestamp 1635444444
transform 1 0 2852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1635444444
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635444444
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1159_
timestamp 1635444444
transform -1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1164_
timestamp 1635444444
transform 1 0 1656 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1635444444
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_38
timestamp 1635444444
transform 1 0 4600 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_42
timestamp 1635444444
transform 1 0 4968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1635444444
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1635444444
transform -1 0 5336 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1168_
timestamp 1635444444
transform 1 0 3772 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_46
timestamp 1635444444
transform 1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1635444444
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_2  _1673_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 5704 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1635444444
transform -1 0 8464 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1635444444
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1635444444
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1953_
timestamp 1635444444
transform 1 0 8924 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_101
timestamp 1635444444
transform 1 0 10396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_109
timestamp 1635444444
transform 1 0 11132 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1073_
timestamp 1635444444
transform -1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_117
timestamp 1635444444
transform 1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_129
timestamp 1635444444
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1750_
timestamp 1635444444
transform -1 0 12972 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1635444444
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1635444444
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_145
timestamp 1635444444
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1635444444
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1108_
timestamp 1635444444
transform 1 0 14536 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_8_156
timestamp 1635444444
transform 1 0 15456 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1635444444
transform 1 0 16100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_167
timestamp 1635444444
transform 1 0 16468 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1107_
timestamp 1635444444
transform 1 0 16560 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1635444444
transform 1 0 15824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_177
timestamp 1635444444
transform 1 0 17388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_181
timestamp 1635444444
transform 1 0 17756 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_186
timestamp 1635444444
transform 1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1635444444
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1635444444
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1085_
timestamp 1635444444
transform 1 0 17848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp 1635444444
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_207
timestamp 1635444444
transform 1 0 20148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1098_
timestamp 1635444444
transform 1 0 19320 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1946_
timestamp 1635444444
transform 1 0 20516 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1635444444
transform 1 0 21988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1635444444
transform 1 0 23092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1635444444
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1635444444
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1635444444
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1635444444
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1635444444
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1635444444
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1635444444
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1635444444
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 1635444444
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_316
timestamp 1635444444
transform 1 0 30176 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635444444
transform -1 0 30820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1635444444
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1729_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 29900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_13
timestamp 1635444444
transform 1 0 2300 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_19
timestamp 1635444444
transform 1 0 2852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1635444444
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635444444
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1162_
timestamp 1635444444
transform 1 0 1472 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1165_
timestamp 1635444444
transform -1 0 3864 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1635444444
transform 1 0 3864 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1167_
timestamp 1635444444
transform 1 0 4232 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_9_44
timestamp 1635444444
transform 1 0 5152 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1635444444
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1635444444
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1635444444
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1178_
timestamp 1635444444
transform 1 0 6716 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_wb_clk_i
timestamp 1635444444
transform -1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_70
timestamp 1635444444
transform 1 0 7544 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1635444444
transform 1 0 8280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1080_
timestamp 1635444444
transform 1 0 8464 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 1635444444
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_89
timestamp 1635444444
transform 1 0 9292 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _1298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 10672 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_116
timestamp 1635444444
transform 1 0 11776 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_126
timestamp 1635444444
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1635444444
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1507_
timestamp 1635444444
transform -1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1509_
timestamp 1635444444
transform -1 0 12696 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1752_
timestamp 1635444444
transform -1 0 13892 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_139
timestamp 1635444444
transform 1 0 13892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_146
timestamp 1635444444
transform 1 0 14536 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1505_
timestamp 1635444444
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1635444444
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1635444444
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1635444444
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_173
timestamp 1635444444
transform 1 0 17020 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1635444444
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1103_
timestamp 1635444444
transform -1 0 18032 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1111_
timestamp 1635444444
transform 1 0 15272 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1635444444
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_192
timestamp 1635444444
transform 1 0 18768 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1072_
timestamp 1635444444
transform -1 0 18768 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_198
timestamp 1635444444
transform 1 0 19320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1635444444
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1635444444
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1091_
timestamp 1635444444
transform 1 0 19412 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1095_
timestamp 1635444444
transform -1 0 21068 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1635444444
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1635444444
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1947_
timestamp 1635444444
transform 1 0 21804 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_241
timestamp 1635444444
transform 1 0 23276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_253
timestamp 1635444444
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_265
timestamp 1635444444
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1635444444
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1635444444
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1635444444
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1635444444
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_305
timestamp 1635444444
transform 1 0 29164 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_311
timestamp 1635444444
transform 1 0 29716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_316
timestamp 1635444444
transform 1 0 30176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635444444
transform -1 0 30820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1635444444
transform 1 0 29808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_6
timestamp 1635444444
transform 1 0 1656 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635444444
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1157_
timestamp 1635444444
transform 1 0 2392 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1635444444
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1635444444
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1635444444
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 1635444444
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1635444444
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1163_
timestamp 1635444444
transform 1 0 3956 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1635444444
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_60
timestamp 1635444444
transform 1 0 6624 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1071_
timestamp 1635444444
transform 1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1173_
timestamp 1635444444
transform 1 0 5704 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_10_68
timestamp 1635444444
transform 1 0 7360 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1635444444
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1635444444
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1635444444
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1079_
timestamp 1635444444
transform 1 0 8096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1262_
timestamp 1635444444
transform -1 0 9476 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_10_101
timestamp 1635444444
transform 1 0 10396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_91
timestamp 1635444444
transform 1 0 9476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1255_
timestamp 1635444444
transform -1 0 11224 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1285_
timestamp 1635444444
transform -1 0 10396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_110
timestamp 1635444444
transform 1 0 11224 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1635444444
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1511_
timestamp 1635444444
transform -1 0 13524 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1749_
timestamp 1635444444
transform -1 0 12604 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1635444444
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1635444444
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1635444444
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1635444444
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1635444444
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_157
timestamp 1635444444
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_167
timestamp 1635444444
transform 1 0 16468 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_171
timestamp 1635444444
transform 1 0 16836 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1097_
timestamp 1635444444
transform 1 0 16928 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1110_
timestamp 1635444444
transform 1 0 15640 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_176
timestamp 1635444444
transform 1 0 17296 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_190
timestamp 1635444444
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1635444444
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1088_
timestamp 1635444444
transform 1 0 17664 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 1635444444
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_201
timestamp 1635444444
transform 1 0 19596 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_218
timestamp 1635444444
transform 1 0 21160 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1945_
timestamp 1635444444
transform 1 0 19688 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_231
timestamp 1635444444
transform 1 0 22356 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _1094_
timestamp 1635444444
transform 1 0 21528 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1635444444
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1635444444
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1635444444
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1635444444
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1635444444
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1635444444
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1635444444
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1635444444
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1635444444
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_309
timestamp 1635444444
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_317
timestamp 1635444444
transform 1 0 30268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635444444
transform -1 0 30820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1635444444
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_19
timestamp 1635444444
transform 1 0 2852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635444444
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1635444444
transform 1 0 1380 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_31
timestamp 1635444444
transform 1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1155_
timestamp 1635444444
transform -1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1635444444
transform 1 0 4324 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1635444444
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1635444444
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1635444444
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1635444444
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1175_
timestamp 1635444444
transform 1 0 6440 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_67
timestamp 1635444444
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_75
timestamp 1635444444
transform 1 0 8004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1075_
timestamp 1635444444
transform 1 0 8372 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1635444444
transform -1 0 8004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1635444444
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_89
timestamp 1635444444
transform 1 0 9292 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1635444444
transform 1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1747_
timestamp 1635444444
transform 1 0 10212 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_122
timestamp 1635444444
transform 1 0 12328 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_130
timestamp 1635444444
transform 1 0 13064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1635444444
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1748_
timestamp 1635444444
transform 1 0 11500 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_142
timestamp 1635444444
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1116_
timestamp 1635444444
transform 1 0 13340 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1635444444
transform 1 0 14536 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1635444444
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1635444444
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1938_
timestamp 1635444444
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_185
timestamp 1635444444
transform 1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1951_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 18492 0 -1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1635444444
transform 1 0 20240 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1635444444
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_234
timestamp 1635444444
transform 1 0 22632 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1635444444
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1093_
timestamp 1635444444
transform 1 0 21804 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_246
timestamp 1635444444
transform 1 0 23736 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_258
timestamp 1635444444
transform 1 0 24840 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_270
timestamp 1635444444
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1635444444
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1635444444
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1635444444
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1635444444
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_305
timestamp 1635444444
transform 1 0 29164 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_311
timestamp 1635444444
transform 1 0 29716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_316
timestamp 1635444444
transform 1 0 30176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635444444
transform -1 0 30820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1635444444
transform 1 0 29808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_12
timestamp 1635444444
transform 1 0 2208 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_6
timestamp 1635444444
transform 1 0 1656 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635444444
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1161_
timestamp 1635444444
transform 1 0 2300 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1635444444
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1635444444
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1635444444
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1635444444
transform 1 0 3772 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_45
timestamp 1635444444
transform 1 0 5244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_53
timestamp 1635444444
transform 1 0 5980 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_61
timestamp 1635444444
transform 1 0 6716 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1171_
timestamp 1635444444
transform -1 0 5980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1635444444
transform -1 0 8280 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_12_78
timestamp 1635444444
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1635444444
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1084_
timestamp 1635444444
transform 1 0 8924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_101
timestamp 1635444444
transform 1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_108
timestamp 1635444444
transform 1 0 11040 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_94
timestamp 1635444444
transform 1 0 9752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1252_
timestamp 1635444444
transform 1 0 10120 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1253_
timestamp 1635444444
transform -1 0 11040 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_115
timestamp 1635444444
transform 1 0 11684 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_123
timestamp 1635444444
transform 1 0 12420 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1106_
timestamp 1635444444
transform 1 0 12696 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1506_
timestamp 1635444444
transform -1 0 11684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1635444444
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1635444444
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1635444444
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1635444444
transform 1 0 14260 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_159
timestamp 1635444444
transform 1 0 15732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1635444444
transform 1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_wb_clk_i
timestamp 1635444444
transform -1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_wb_clk_i
timestamp 1635444444
transform 1 0 16836 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_175
timestamp 1635444444
transform 1 0 17204 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_181
timestamp 1635444444
transform 1 0 17756 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1635444444
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1635444444
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1635444444
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1089_
timestamp 1635444444
transform 1 0 17848 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1635444444
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_203
timestamp 1635444444
transform 1 0 19780 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_210
timestamp 1635444444
transform 1 0 20424 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1092_
timestamp 1635444444
transform 1 0 21160 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1713_
timestamp 1635444444
transform 1 0 19504 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1723_
timestamp 1635444444
transform 1 0 20148 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1635444444
transform 1 0 21988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1635444444
transform 1 0 23092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1635444444
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1635444444
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1635444444
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1635444444
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1635444444
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1635444444
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1635444444
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1635444444
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_309
timestamp 1635444444
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_317
timestamp 1635444444
transform 1 0 30268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635444444
transform -1 0 30820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1635444444
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1635444444
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1158_
timestamp 1635444444
transform 1 0 1472 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635444444
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635444444
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1635444444
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_6
timestamp 1635444444
transform 1 0 1656 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1635444444
transform -1 0 2944 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1160_
timestamp 1635444444
transform 1 0 2576 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1635444444
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_14
timestamp 1635444444
transform 1 0 2392 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1635444444
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_25
timestamp 1635444444
transform 1 0 3404 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_31
timestamp 1635444444
transform 1 0 3956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_41
timestamp 1635444444
transform 1 0 4876 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1635444444
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1170_
timestamp 1635444444
transform 1 0 4048 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1635444444
transform 1 0 3772 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__a22oi_1  _1694_
timestamp 1635444444
transform 1 0 5980 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1112_
timestamp 1635444444
transform -1 0 5612 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_45
timestamp 1635444444
transform 1 0 5244 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp 1635444444
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _1686_
timestamp 1635444444
transform -1 0 6992 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1645_
timestamp 1635444444
transform -1 0 7268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1635444444
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_59
timestamp 1635444444
transform 1 0 6532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 1635444444
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1635444444
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_64
timestamp 1635444444
transform 1 0 6992 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_76
timestamp 1635444444
transform 1 0 8096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_67
timestamp 1635444444
transform 1 0 7268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1635444444
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1635444444
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1635444444
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1635444444
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1646_
timestamp 1635444444
transform -1 0 8004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1952_
timestamp 1635444444
transform 1 0 8280 0 -1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_13_103
timestamp 1635444444
transform 1 0 10580 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1635444444
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_97
timestamp 1635444444
transform 1 0 10028 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_94
timestamp 1635444444
transform 1 0 9752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_98
timestamp 1635444444
transform 1 0 10120 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1263_
timestamp 1635444444
transform -1 0 9752 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1635444444
transform 1 0 10212 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1635444444
transform -1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1635444444
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_124
timestamp 1635444444
transform 1 0 12512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_115
timestamp 1635444444
transform 1 0 11684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1635444444
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1115_
timestamp 1635444444
transform -1 0 12512 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1635444444
transform 1 0 12052 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1635444444
transform -1 0 14352 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_144
timestamp 1635444444
transform 1 0 14352 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1635444444
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1635444444
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_150
timestamp 1635444444
transform 1 0 14904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1635444444
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1114_
timestamp 1635444444
transform -1 0 15548 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1121_
timestamp 1635444444
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_157
timestamp 1635444444
transform 1 0 15548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1635444444
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1635444444
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_158
timestamp 1635444444
transform 1 0 15640 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_172
timestamp 1635444444
transform 1 0 16928 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1635444444
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1666_
timestamp 1635444444
transform 1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _1667_
timestamp 1635444444
transform 1 0 16376 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1635444444
transform 1 0 15272 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1665_
timestamp 1635444444
transform 1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1090_
timestamp 1635444444
transform 1 0 18124 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_184
timestamp 1635444444
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1635444444
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_176
timestamp 1635444444
transform 1 0 17296 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1635444444
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1635444444
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1635444444
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1635444444
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1950_
timestamp 1635444444
transform 1 0 17848 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_198
timestamp 1635444444
transform 1 0 19320 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1635444444
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1635444444
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_197
timestamp 1635444444
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_205
timestamp 1635444444
transform 1 0 19964 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_211
timestamp 1635444444
transform 1 0 20516 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1702_
timestamp 1635444444
transform 1 0 19688 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1703_
timestamp 1635444444
transform -1 0 20516 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1635444444
transform -1 0 22540 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1635444444
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1635444444
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1635444444
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1949_
timestamp 1635444444
transform 1 0 21804 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_13_241
timestamp 1635444444
transform 1 0 23276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_253
timestamp 1635444444
transform 1 0 24380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1635444444
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1635444444
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1635444444
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1635444444
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_265
timestamp 1635444444
transform 1 0 25484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1635444444
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1635444444
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1635444444
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1635444444
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1635444444
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1635444444
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1635444444
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1635444444
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1635444444
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_317
timestamp 1635444444
transform 1 0 30268 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1635444444
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_309
timestamp 1635444444
transform 1 0 29532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_316
timestamp 1635444444
transform 1 0 30176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635444444
transform -1 0 30820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635444444
transform -1 0 30820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1635444444
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1635444444
transform 1 0 29808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_20
timestamp 1635444444
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1635444444
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635444444
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1635444444
transform 1 0 1472 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_32
timestamp 1635444444
transform 1 0 4048 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_40
timestamp 1635444444
transform 1 0 4784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _1700_
timestamp 1635444444
transform 1 0 5060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1635444444
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1635444444
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1635444444
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_64
timestamp 1635444444
transform 1 0 6992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1635444444
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1720_
timestamp 1635444444
transform -1 0 6992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_72
timestamp 1635444444
transform 1 0 7728 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_78
timestamp 1635444444
transform 1 0 8280 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_83
timestamp 1635444444
transform 1 0 8740 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_87
timestamp 1635444444
transform 1 0 9108 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1635444444
transform -1 0 8740 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1635444444
transform -1 0 7728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1635444444
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_93
timestamp 1635444444
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_97
timestamp 1635444444
transform 1 0 10028 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1127_
timestamp 1635444444
transform 1 0 10120 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _1277_
timestamp 1635444444
transform 1 0 9200 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1635444444
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1635444444
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1635444444
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1635444444
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1113_
timestamp 1635444444
transform 1 0 12328 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1635444444
transform 1 0 11592 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_132
timestamp 1635444444
transform 1 0 13248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1635444444
transform 1 0 13984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_145
timestamp 1635444444
transform 1 0 14444 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1649_
timestamp 1635444444
transform -1 0 15272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1651_
timestamp 1635444444
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_154
timestamp 1635444444
transform 1 0 15272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1635444444
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1635444444
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1635444444
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1668_
timestamp 1635444444
transform 1 0 16744 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_1  _1678_
timestamp 1635444444
transform 1 0 15640 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1635444444
transform 1 0 17572 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_186
timestamp 1635444444
transform 1 0 18216 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1677_
timestamp 1635444444
transform 1 0 17940 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1705_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 18768 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1635444444
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_211
timestamp 1635444444
transform 1 0 20516 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1635444444
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1706_
timestamp 1635444444
transform 1 0 19688 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1714_
timestamp 1635444444
transform -1 0 21160 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1635444444
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1635444444
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1635444444
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1635444444
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1635444444
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1635444444
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1635444444
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1635444444
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1635444444
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1635444444
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1635444444
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_317
timestamp 1635444444
transform 1 0 30268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635444444
transform -1 0 30820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 1635444444
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_6
timestamp 1635444444
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635444444
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1635444444
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1635444444
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1635444444
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 1635444444
transform 1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1635444444
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_50
timestamp 1635444444
transform 1 0 5704 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_62
timestamp 1635444444
transform 1 0 6808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_1  _1711_
timestamp 1635444444
transform 1 0 5152 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1927_
timestamp 1635444444
transform -1 0 8372 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1635444444
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1635444444
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1635444444
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or4b_2  _1265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_101
timestamp 1635444444
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_105
timestamp 1635444444
transform 1 0 10764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1635444444
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1635444444
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1125_
timestamp 1635444444
transform 1 0 10856 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_115
timestamp 1635444444
transform 1 0 11684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_123
timestamp 1635444444
transform 1 0 12420 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1120_
timestamp 1635444444
transform 1 0 12788 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1635444444
transform 1 0 12052 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1635444444
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_150
timestamp 1635444444
transform 1 0 14904 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1635444444
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1119_
timestamp 1635444444
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_167
timestamp 1635444444
transform 1 0 16468 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _1655_
timestamp 1635444444
transform 1 0 16836 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1656_
timestamp 1635444444
transform 1 0 15640 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_177
timestamp 1635444444
transform 1 0 17388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_185
timestamp 1635444444
transform 1 0 18124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1635444444
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1635444444
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1370_
timestamp 1635444444
transform -1 0 18124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1675_
timestamp 1635444444
transform 1 0 18492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1635444444
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_212
timestamp 1635444444
transform 1 0 20608 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1716_
timestamp 1635444444
transform 1 0 19780 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1724_
timestamp 1635444444
transform -1 0 21252 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_219
timestamp 1635444444
transform 1 0 21252 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_231
timestamp 1635444444
transform 1 0 22356 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_243
timestamp 1635444444
transform 1 0 23460 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1635444444
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1635444444
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1635444444
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1635444444
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1635444444
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1635444444
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1635444444
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1635444444
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_309
timestamp 1635444444
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_317
timestamp 1635444444
transform 1 0 30268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635444444
transform -1 0 30820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1635444444
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_6
timestamp 1635444444
transform 1 0 1656 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635444444
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1156_
timestamp 1635444444
transform 1 0 2392 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1635444444
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_23
timestamp 1635444444
transform 1 0 3220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_43
timestamp 1635444444
transform 1 0 5060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1635444444
transform 1 0 3588 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_47
timestamp 1635444444
transform 1 0 5428 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1635444444
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_60
timestamp 1635444444
transform 1 0 6624 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1635444444
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1129_
timestamp 1635444444
transform 1 0 6992 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1638_
timestamp 1635444444
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_wb_clk_i
timestamp 1635444444
transform 1 0 5520 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_73
timestamp 1635444444
transform 1 0 7820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1635444444
transform 1 0 8188 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1635444444
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_93
timestamp 1635444444
transform 1 0 9660 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1128_
timestamp 1635444444
transform 1 0 10212 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1635444444
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_121
timestamp 1635444444
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1635444444
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1931_
timestamp 1635444444
transform 1 0 12420 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1635444444
transform 1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1635444444
transform 1 0 14260 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1635444444
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1635444444
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1635444444
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_173
timestamp 1635444444
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1635444444
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1679_
timestamp 1635444444
transform 1 0 17112 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_183
timestamp 1635444444
transform 1 0 17940 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_195
timestamp 1635444444
transform 1 0 19044 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1691_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 18308 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_212
timestamp 1635444444
transform 1 0 20608 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1682_
timestamp 1635444444
transform 1 0 20976 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1726_
timestamp 1635444444
transform 1 0 19780 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1635444444
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1635444444
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1635444444
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1635444444
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1635444444
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1635444444
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1635444444
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1635444444
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1635444444
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1635444444
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1635444444
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1731_
timestamp 1635444444
transform -1 0 29440 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_308
timestamp 1635444444
transform 1 0 29440 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_316
timestamp 1635444444
transform 1 0 30176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635444444
transform -1 0 30820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1635444444
transform 1 0 29808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1635444444
transform 1 0 2392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1635444444
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1635444444
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635444444
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1153_
timestamp 1635444444
transform -1 0 2392 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1635444444
transform -1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1635444444
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1635444444
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1635444444
transform 1 0 3772 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_45
timestamp 1635444444
transform 1 0 5244 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_51
timestamp 1635444444
transform 1 0 5796 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_61
timestamp 1635444444
transform 1 0 6716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1648_
timestamp 1635444444
transform 1 0 5888 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1722_
timestamp 1635444444
transform 1 0 7084 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_74
timestamp 1635444444
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1635444444
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1635444444
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1635444444
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_101
timestamp 1635444444
transform 1 0 10396 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1635444444
transform 1 0 9660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1356_
timestamp 1635444444
transform 1 0 9200 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1360_
timestamp 1635444444
transform -1 0 10396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1635444444
transform 1 0 10948 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_123
timestamp 1635444444
transform 1 0 12420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1123_
timestamp 1635444444
transform -1 0 13616 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1635444444
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1635444444
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1635444444
transform 1 0 14076 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1635444444
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_171
timestamp 1635444444
transform 1 0 16836 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1650_
timestamp 1635444444
transform 1 0 15916 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  FILLER_18_179
timestamp 1635444444
transform 1 0 17572 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1635444444
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1635444444
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _1683_
timestamp 1635444444
transform 1 0 17848 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1635444444
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_213
timestamp 1635444444
transform 1 0 20700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_4  _1044_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 20056 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1715_
timestamp 1635444444
transform 1 0 19228 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_18_225
timestamp 1635444444
transform 1 0 21804 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_237
timestamp 1635444444
transform 1 0 22908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1635444444
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1635444444
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1635444444
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1635444444
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1635444444
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1635444444
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1635444444
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1635444444
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_309
timestamp 1635444444
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_316
timestamp 1635444444
transform 1 0 30176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635444444
transform -1 0 30820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1635444444
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1658_
timestamp 1635444444
transform 1 0 29900 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_20
timestamp 1635444444
transform 1 0 2944 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1635444444
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_10
timestamp 1635444444
transform 1 0 2024 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1635444444
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635444444
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635444444
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1151_
timestamp 1635444444
transform 1 0 2392 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1685_
timestamp 1635444444
transform -1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1635444444
transform 1 0 1472 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__o221a_1  _1154_
timestamp 1635444444
transform 1 0 3312 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1635444444
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1635444444
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1635444444
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_wb_clk_i
timestamp 1635444444
transform -1 0 4876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1146_
timestamp 1635444444
transform -1 0 4508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1635444444
transform 1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_37
timestamp 1635444444
transform 1 0 4508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_41
timestamp 1635444444
transform 1 0 4876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_33
timestamp 1635444444
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _1721_
timestamp 1635444444
transform 1 0 5244 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1663_
timestamp 1635444444
transform 1 0 5796 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_50
timestamp 1635444444
transform 1 0 5704 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_44
timestamp 1635444444
transform 1 0 5152 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1635444444
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1642_
timestamp 1635444444
transform -1 0 7636 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1635444444
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_60
timestamp 1635444444
transform 1 0 6624 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1635444444
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1635444444
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_71
timestamp 1635444444
transform 1 0 7636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1635444444
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_68
timestamp 1635444444
transform 1 0 7360 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1635444444
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1635444444
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1635444444
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1358_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8740 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1652_
timestamp 1635444444
transform -1 0 8464 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1676_
timestamp 1635444444
transform 1 0 8004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_103
timestamp 1635444444
transform 1 0 10580 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1635444444
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_88
timestamp 1635444444
transform 1 0 9200 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1635444444
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_93
timestamp 1635444444
transform 1 0 9660 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1118_
timestamp 1635444444
transform 1 0 10672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1357_
timestamp 1635444444
transform 1 0 9292 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _1384_
timestamp 1635444444
transform 1 0 9568 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1635444444
transform 1 0 10212 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_19_116
timestamp 1635444444
transform 1 0 11776 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_124
timestamp 1635444444
transform 1 0 12512 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_128
timestamp 1635444444
transform 1 0 12880 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1635444444
transform 1 0 11684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_124
timestamp 1635444444
transform 1 0 12512 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1635444444
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1359_
timestamp 1635444444
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 12512 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1380_
timestamp 1635444444
transform -1 0 12880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1635444444
transform -1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1635444444
transform -1 0 13616 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1635444444
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_132
timestamp 1635444444
transform 1 0 13248 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_138
timestamp 1635444444
transform 1 0 13800 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_wb_clk_i
timestamp 1635444444
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1639_
timestamp 1635444444
transform -1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1635444444
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_147
timestamp 1635444444
transform 1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1635444444
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_146
timestamp 1635444444
transform 1 0 14536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1574_
timestamp 1635444444
transform -1 0 15456 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_19_151
timestamp 1635444444
transform 1 0 14996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1635444444
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1635444444
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_156
timestamp 1635444444
transform 1 0 15456 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_169
timestamp 1635444444
transform 1 0 16652 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1635444444
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1575_
timestamp 1635444444
transform 1 0 15364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1643_
timestamp 1635444444
transform 1 0 16192 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1657_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 17296 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1704_
timestamp 1635444444
transform 1 0 17664 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1688_
timestamp 1635444444
transform -1 0 18124 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_20_177
timestamp 1635444444
transform 1 0 17388 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_176
timestamp 1635444444
transform 1 0 17296 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1635444444
transform 1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_185
timestamp 1635444444
transform 1 0 18124 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_192
timestamp 1635444444
transform 1 0 18768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1635444444
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1725_
timestamp 1635444444
transform 1 0 19136 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1635444444
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1635444444
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_201
timestamp 1635444444
transform 1 0 19596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_212
timestamp 1635444444
transform 1 0 20608 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_201
timestamp 1635444444
transform 1 0 19596 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_207
timestamp 1635444444
transform 1 0 20148 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_216
timestamp 1635444444
transform 1 0 20976 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0914_
timestamp 1635444444
transform -1 0 19596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1669_
timestamp 1635444444
transform -1 0 20608 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1727_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 20976 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1635444444
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1635444444
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_228
timestamp 1635444444
transform 1 0 22080 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_240
timestamp 1635444444
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1635444444
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1635444444
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1635444444
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1635444444
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1635444444
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1635444444
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1635444444
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1635444444
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1635444444
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1635444444
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1635444444
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1635444444
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_305
timestamp 1635444444
transform 1 0 29164 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1635444444
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1635444444
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_316
timestamp 1635444444
transform 1 0 30176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1635444444
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1635444444
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_316
timestamp 1635444444
transform 1 0 30176 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635444444
transform -1 0 30820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635444444
transform -1 0 30820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1635444444
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1670_
timestamp 1635444444
transform 1 0 29900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1635444444
transform 1 0 29808 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_12
timestamp 1635444444
transform 1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635444444
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1149_
timestamp 1635444444
transform 1 0 2576 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1152_
timestamp 1635444444
transform -1 0 2208 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_26
timestamp 1635444444
transform 1 0 3496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1635444444
transform 1 0 4692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_43
timestamp 1635444444
transform 1 0 5060 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1150_
timestamp 1635444444
transform 1 0 3864 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1635444444
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1635444444
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1635444444
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_61
timestamp 1635444444
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1635444444
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1660_
timestamp 1635444444
transform 1 0 5152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1687_
timestamp 1635444444
transform 1 0 6808 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1635444444
transform 1 0 7636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_83
timestamp 1635444444
transform 1 0 8740 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1286_
timestamp 1635444444
transform -1 0 9568 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_103
timestamp 1635444444
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_92
timestamp 1635444444
transform 1 0 9568 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_98
timestamp 1635444444
transform 1 0 10120 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1126_
timestamp 1635444444
transform 1 0 10212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1635444444
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1635444444
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_121
timestamp 1635444444
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1635444444
transform 1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_131
timestamp 1635444444
transform 1 0 13156 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1635444444
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_wb_clk_i
timestamp 1635444444
transform -1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_138
timestamp 1635444444
transform 1 0 13800 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1635444444
transform 1 0 14812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1028_
timestamp 1635444444
transform 1 0 13248 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1641_
timestamp 1635444444
transform -1 0 14812 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1635444444
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1635444444
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _1528_
timestamp 1635444444
transform 1 0 15180 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_4  _1644_
timestamp 1635444444
transform -1 0 17848 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_21_182
timestamp 1635444444
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_186
timestamp 1635444444
transform 1 0 18216 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1982_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 19872 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_21_204
timestamp 1635444444
transform 1 0 19872 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1664_
timestamp 1635444444
transform 1 0 20424 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1635444444
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1635444444
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_229
timestamp 1635444444
transform 1 0 22172 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_240
timestamp 1635444444
transform 1 0 23184 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1635444444
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1375_
timestamp 1635444444
transform 1 0 22264 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_21_252
timestamp 1635444444
transform 1 0 24288 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_264
timestamp 1635444444
transform 1 0 25392 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1635444444
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1635444444
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1635444444
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1635444444
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_305
timestamp 1635444444
transform 1 0 29164 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_316
timestamp 1635444444
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635444444
transform -1 0 30820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1697_
timestamp 1635444444
transform 1 0 29900 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1635444444
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1635444444
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635444444
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1635444444
transform 1 0 1472 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1635444444
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1635444444
transform -1 0 5244 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_45
timestamp 1635444444
transform 1 0 5244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_49
timestamp 1635444444
transform 1 0 5612 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_59
timestamp 1635444444
transform 1 0 6532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1674_
timestamp 1635444444
transform 1 0 5704 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1695_
timestamp 1635444444
transform 1 0 6900 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_72
timestamp 1635444444
transform 1 0 7728 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1635444444
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1635444444
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1653_
timestamp 1635444444
transform 1 0 8096 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1858_
timestamp 1635444444
transform 1 0 8924 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_22_102
timestamp 1635444444
transform 1 0 10488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_114
timestamp 1635444444
transform 1 0 11592 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1635444444
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_127
timestamp 1635444444
transform 1 0 12788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1017_
timestamp 1635444444
transform 1 0 12420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1378_
timestamp 1635444444
transform -1 0 12052 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1379_
timestamp 1635444444
transform -1 0 13616 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1635444444
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1635444444
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1635444444
transform 1 0 14812 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1635444444
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1026_
timestamp 1635444444
transform -1 0 14812 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_156
timestamp 1635444444
transform 1 0 15456 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_166
timestamp 1635444444
transform 1 0 16376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1560_
timestamp 1635444444
transform -1 0 15456 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1573_
timestamp 1635444444
transform -1 0 16376 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_2  _1654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 17664 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_22_180
timestamp 1635444444
transform 1 0 17664 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1635444444
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1635444444
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1635444444
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1696_
timestamp 1635444444
transform -1 0 18676 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1635444444
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_201
timestamp 1635444444
transform 1 0 19596 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_209
timestamp 1635444444
transform 1 0 20332 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1659_
timestamp 1635444444
transform 1 0 20700 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1680_
timestamp 1635444444
transform -1 0 20332 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_22_223
timestamp 1635444444
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_234
timestamp 1635444444
transform 1 0 22632 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _1707_
timestamp 1635444444
transform -1 0 22632 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1635444444
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1635444444
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1635444444
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1635444444
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1635444444
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1635444444
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1635444444
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1732_
timestamp 1635444444
transform -1 0 29072 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_309
timestamp 1635444444
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_316
timestamp 1635444444
transform 1 0 30176 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635444444
transform -1 0 30820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1635444444
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1689_
timestamp 1635444444
transform 1 0 29900 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_13
timestamp 1635444444
transform 1 0 2300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_6
timestamp 1635444444
transform 1 0 1656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1635444444
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1147_
timestamp 1635444444
transform 1 0 2668 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1635444444
transform -1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1635444444
transform 1 0 2024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_26
timestamp 1635444444
transform 1 0 3496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1635444444
transform 1 0 3864 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_46
timestamp 1635444444
transform 1 0 5336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1635444444
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1635444444
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1701_
timestamp 1635444444
transform 1 0 6348 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_66
timestamp 1635444444
transform 1 0 7176 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1635444444
transform 1 0 8280 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_82
timestamp 1635444444
transform 1 0 8648 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_86
timestamp 1635444444
transform 1 0 9016 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1635444444
transform 1 0 8740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1635444444
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1635444444
transform -1 0 11040 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1635444444
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1635444444
transform 1 0 13156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1635444444
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _1739_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 13156 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_141
timestamp 1635444444
transform 1 0 14076 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1019_
timestamp 1635444444
transform -1 0 14076 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1981_
timestamp 1635444444
transform 1 0 14444 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1635444444
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_174
timestamp 1635444444
transform 1 0 17112 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1635444444
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1021_
timestamp 1635444444
transform 1 0 16652 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_23_187
timestamp 1635444444
transform 1 0 18308 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0896_
timestamp 1635444444
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1635444444
transform -1 0 18308 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_23_197
timestamp 1635444444
transform 1 0 19228 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_205
timestamp 1635444444
transform 1 0 19964 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_216
timestamp 1635444444
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _1717_
timestamp 1635444444
transform -1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_230
timestamp 1635444444
transform 1 0 22264 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1635444444
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1374_
timestamp 1635444444
transform 1 0 21804 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_23_242
timestamp 1635444444
transform 1 0 23368 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_254
timestamp 1635444444
transform 1 0 24472 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_266
timestamp 1635444444
transform 1 0 25576 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1635444444
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1635444444
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1635444444
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1635444444
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1708_
timestamp 1635444444
transform 1 0 29164 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_308
timestamp 1635444444
transform 1 0 29440 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_316
timestamp 1635444444
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1635444444
transform -1 0 30820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1635444444
transform 1 0 29808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_10
timestamp 1635444444
transform 1 0 2024 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1635444444
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_6
timestamp 1635444444
transform 1 0 1656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1635444444
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1145_
timestamp 1635444444
transform 1 0 2116 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1635444444
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_38
timestamp 1635444444
transform 1 0 4600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1635444444
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1144_
timestamp 1635444444
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1671_
timestamp 1635444444
transform 1 0 4968 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_45
timestamp 1635444444
transform 1 0 5244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_58
timestamp 1635444444
transform 1 0 6440 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1635444444
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1635444444
transform 1 0 6808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1712_
timestamp 1635444444
transform 1 0 5612 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_72
timestamp 1635444444
transform 1 0 7728 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1635444444
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1635444444
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1635444444
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1295_
timestamp 1635444444
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1698_
timestamp 1635444444
transform 1 0 7452 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1719_
timestamp 1635444444
transform 1 0 8096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1635444444
transform 1 0 9660 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1854_
timestamp 1635444444
transform 1 0 10028 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1635444444
transform 1 0 11592 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1635444444
transform 1 0 11960 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1635444444
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1635444444
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1635444444
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0903_
timestamp 1635444444
transform 1 0 14444 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_154
timestamp 1635444444
transform 1 0 15272 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_165
timestamp 1635444444
transform 1 0 16284 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_171
timestamp 1635444444
transform 1 0 16836 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1535_
timestamp 1635444444
transform 1 0 16928 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1539_
timestamp 1635444444
transform -1 0 16284 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_176
timestamp 1635444444
transform 1 0 17296 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_186
timestamp 1635444444
transform 1 0 18216 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1635444444
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1635444444
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or3_2  _1022_
timestamp 1635444444
transform 1 0 17664 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1635444444
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_204
timestamp 1635444444
transform 1 0 19872 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_212
timestamp 1635444444
transform 1 0 20608 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0897_
timestamp 1635444444
transform -1 0 20608 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1020_
timestamp 1635444444
transform -1 0 19872 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1046_
timestamp 1635444444
transform -1 0 21344 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_220
timestamp 1635444444
transform 1 0 21344 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_228
timestamp 1635444444
transform 1 0 22080 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_240
timestamp 1635444444
transform 1 0 23184 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1534_
timestamp 1635444444
transform -1 0 22080 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1635444444
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1635444444
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1635444444
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1635444444
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1635444444
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1635444444
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1635444444
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_309
timestamp 1635444444
transform 1 0 29532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_316
timestamp 1635444444
transform 1 0 30176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1635444444
transform -1 0 30820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1635444444
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1681_
timestamp 1635444444
transform 1 0 29900 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_12
timestamp 1635444444
transform 1 0 2208 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_6
timestamp 1635444444
transform 1 0 1656 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1635444444
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1635444444
transform 1 0 2300 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1635444444
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_29
timestamp 1635444444
transform 1 0 3772 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_43
timestamp 1635444444
transform 1 0 5060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1142_
timestamp 1635444444
transform 1 0 4140 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1635444444
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_57
timestamp 1635444444
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1635444444
transform 1 0 6808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1635444444
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1117_
timestamp 1635444444
transform 1 0 6440 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1640_
timestamp 1635444444
transform 1 0 5428 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_75
timestamp 1635444444
transform 1 0 8004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1288_
timestamp 1635444444
transform 1 0 8740 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1296_
timestamp 1635444444
transform -1 0 8004 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1635444444
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1635444444
transform 1 0 9660 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1297_
timestamp 1635444444
transform 1 0 10028 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1635444444
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1635444444
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_125
timestamp 1635444444
transform 1 0 12604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1635444444
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1369_
timestamp 1635444444
transform 1 0 12328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_133
timestamp 1635444444
transform 1 0 13340 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_141
timestamp 1635444444
transform 1 0 14076 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_150
timestamp 1635444444
transform 1 0 14904 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1024_
timestamp 1635444444
transform -1 0 14904 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 13432 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_25_162
timestamp 1635444444
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1635444444
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0899_
timestamp 1635444444
transform 1 0 16652 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_178
timestamp 1635444444
transform 1 0 17480 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_194
timestamp 1635444444
transform 1 0 18952 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0902_
timestamp 1635444444
transform 1 0 18216 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_202
timestamp 1635444444
transform 1 0 19688 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1984_
timestamp 1635444444
transform 1 0 19872 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1635444444
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1635444444
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1635444444
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1635444444
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1635444444
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1635444444
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1635444444
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1635444444
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1635444444
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1635444444
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1635444444
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1635444444
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_317
timestamp 1635444444
transform 1 0 30268 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1635444444
transform -1 0 30820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_10
timestamp 1635444444
transform 1 0 2024 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1635444444
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_6
timestamp 1635444444
transform 1 0 1656 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_19
timestamp 1635444444
transform 1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1635444444
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1635444444
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1134_
timestamp 1635444444
transform 1 0 2116 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1635444444
transform 1 0 1380 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1635444444
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1635444444
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_29
timestamp 1635444444
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_26
timestamp 1635444444
transform 1 0 3496 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1635444444
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1635444444
transform 1 0 4048 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1635444444
transform 1 0 4324 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1635444444
transform -1 0 3496 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_51
timestamp 1635444444
transform 1 0 5796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_58
timestamp 1635444444
transform 1 0 6440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1635444444
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1635444444
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_63
timestamp 1635444444
transform 1 0 6900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1635444444
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1270_
timestamp 1635444444
transform 1 0 6164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1271_
timestamp 1635444444
transform 1 0 6532 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1635444444
transform 1 0 6808 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_26_78
timestamp 1635444444
transform 1 0 8280 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_83
timestamp 1635444444
transform 1 0 8740 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1635444444
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1289_
timestamp 1635444444
transform 1 0 8924 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1293_
timestamp 1635444444
transform 1 0 9108 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1635444444
transform 1 0 7268 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_26_107
timestamp 1635444444
transform 1 0 10948 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_95
timestamp 1635444444
transform 1 0 9844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1635444444
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_96
timestamp 1635444444
transform 1 0 9936 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1635444444
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_123
timestamp 1635444444
transform 1 0 12420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1635444444
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1635444444
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1635444444
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _0884_
timestamp 1635444444
transform 1 0 11868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 13616 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1957_
timestamp 1635444444
transform 1 0 11960 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1635444444
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1635444444
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_134
timestamp 1635444444
transform 1 0 13432 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_141
timestamp 1635444444
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_145
timestamp 1635444444
transform 1 0 14444 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1635444444
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0905_
timestamp 1635444444
transform 1 0 14536 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1635444444
transform 1 0 13800 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1980_
timestamp 1635444444
transform 1 0 14812 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_26_168
timestamp 1635444444
transform 1 0 16560 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_155
timestamp 1635444444
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_162
timestamp 1635444444
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_172
timestamp 1635444444
transform 1 0 16928 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1635444444
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1635444444
transform -1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1541_
timestamp 1635444444
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1983_
timestamp 1635444444
transform 1 0 16928 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1635444444
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1635444444
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1635444444
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_196
timestamp 1635444444
transform 1 0 19136 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1635444444
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1635444444
transform -1 0 19136 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1561_
timestamp 1635444444
transform 1 0 17296 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_26_206
timestamp 1635444444
transform 1 0 20056 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_209
timestamp 1635444444
transform 1 0 20332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _0898_
timestamp 1635444444
transform -1 0 20056 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1730_
timestamp 1635444444
transform 1 0 19504 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1985_
timestamp 1635444444
transform 1 0 20608 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_26_228
timestamp 1635444444
transform 1 0 22080 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_240
timestamp 1635444444
transform 1 0 23184 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1635444444
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1635444444
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1635444444
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1635444444
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1635444444
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1635444444
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1635444444
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1635444444
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1635444444
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1635444444
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1635444444
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1635444444
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1635444444
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1635444444
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1635444444
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1635444444
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1635444444
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1635444444
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1635444444
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_309
timestamp 1635444444
transform 1 0 29532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_316
timestamp 1635444444
transform 1 0 30176 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_317
timestamp 1635444444
transform 1 0 30268 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1635444444
transform -1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1635444444
transform -1 0 30820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1635444444
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1635444444
transform 1 0 29808 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_14
timestamp 1635444444
transform 1 0 2392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1635444444
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1635444444
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1635444444
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1141_
timestamp 1635444444
transform -1 0 2392 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1635444444
transform -1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1635444444
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_39
timestamp 1635444444
transform 1 0 4692 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1635444444
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1140_
timestamp 1635444444
transform 1 0 3772 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_28_45
timestamp 1635444444
transform 1 0 5244 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_49
timestamp 1635444444
transform 1 0 5612 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1283_
timestamp 1635444444
transform 1 0 6348 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1661_
timestamp 1635444444
transform 1 0 5336 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_67
timestamp 1635444444
transform 1 0 7268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1635444444
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1635444444
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1635444444
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1290_
timestamp 1635444444
transform 1 0 7636 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1635444444
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1635444444
transform 1 0 9752 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_110
timestamp 1635444444
transform 1 0 11224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_130
timestamp 1635444444
transform 1 0 13064 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1635444444
transform 1 0 11592 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1635444444
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1635444444
transform 1 0 14812 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1635444444
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _1067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 14812 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1635444444
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1635444444
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1540_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 15180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1562_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 17848 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1809_
timestamp 1635444444
transform -1 0 16744 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_182
timestamp 1635444444
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1635444444
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1635444444
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1635444444
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1583_
timestamp 1635444444
transform 1 0 18216 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_200
timestamp 1635444444
transform 1 0 19504 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_210
timestamp 1635444444
transform 1 0 20424 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_217
timestamp 1635444444
transform 1 0 21068 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1584_
timestamp 1635444444
transform -1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1604_
timestamp 1635444444
transform -1 0 21068 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1624_
timestamp 1635444444
transform 1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_229
timestamp 1635444444
transform 1 0 22172 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_241
timestamp 1635444444
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1635444444
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1635444444
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1635444444
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1635444444
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1635444444
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1635444444
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1635444444
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1635444444
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1635444444
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_316
timestamp 1635444444
transform 1 0 30176 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1635444444
transform -1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1635444444
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1733_
timestamp 1635444444
transform 1 0 29900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_16
timestamp 1635444444
transform 1 0 2576 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1635444444
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1635444444
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1139_
timestamp 1635444444
transform 1 0 1748 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_24
timestamp 1635444444
transform 1 0 3312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_35
timestamp 1635444444
transform 1 0 4324 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_43
timestamp 1635444444
transform 1 0 5060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1130_
timestamp 1635444444
transform -1 0 5060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1143_
timestamp 1635444444
transform 1 0 3496 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1635444444
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1635444444
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_60
timestamp 1635444444
transform 1 0 6624 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1635444444
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1138_
timestamp 1635444444
transform -1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1709_
timestamp 1635444444
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1710_
timestamp 1635444444
transform 1 0 6992 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_67
timestamp 1635444444
transform 1 0 7268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_79
timestamp 1635444444
transform 1 0 8372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1292_
timestamp 1635444444
transform 1 0 8924 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_101
timestamp 1635444444
transform 1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1635444444
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_94
timestamp 1635444444
transform 1 0 9752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1430_
timestamp 1635444444
transform -1 0 10396 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_129
timestamp 1635444444
transform 1 0 12972 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1635444444
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1635444444
transform 1 0 11500 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_29_135
timestamp 1635444444
transform 1 0 13524 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_140
timestamp 1635444444
transform 1 0 13984 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_148
timestamp 1635444444
transform 1 0 14720 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1066_
timestamp 1635444444
transform 1 0 13616 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1773_
timestamp 1635444444
transform 1 0 14996 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_160
timestamp 1635444444
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1635444444
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1563_
timestamp 1635444444
transform -1 0 17572 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1635444444
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1635444444
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1585_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 19136 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_29_207
timestamp 1635444444
transform 1 0 20148 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_216
timestamp 1635444444
transform 1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1605_
timestamp 1635444444
transform 1 0 19504 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1625_
timestamp 1635444444
transform 1 0 20516 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_29_228
timestamp 1635444444
transform 1 0 22080 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_240
timestamp 1635444444
transform 1 0 23184 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1635444444
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1623_
timestamp 1635444444
transform -1 0 22080 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_252
timestamp 1635444444
transform 1 0 24288 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_264
timestamp 1635444444
transform 1 0 25392 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1635444444
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1635444444
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1635444444
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1635444444
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_305
timestamp 1635444444
transform 1 0 29164 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_311
timestamp 1635444444
transform 1 0 29716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_316
timestamp 1635444444
transform 1 0 30176 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1635444444
transform -1 0 30820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1635444444
transform 1 0 29808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1635444444
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1635444444
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1635444444
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1635444444
transform 1 0 1840 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1635444444
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp 1635444444
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_41
timestamp 1635444444
transform 1 0 4876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1635444444
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1131_
timestamp 1635444444
transform 1 0 4048 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_48
timestamp 1635444444
transform 1 0 5520 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1672_
timestamp 1635444444
transform 1 0 5244 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1635444444
transform -1 0 7360 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1635444444
transform 1 0 7360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1635444444
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1635444444
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1294_
timestamp 1635444444
transform 1 0 8924 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_106
timestamp 1635444444
transform 1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_94
timestamp 1635444444
transform 1 0 9752 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1105_
timestamp 1635444444
transform -1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_114
timestamp 1635444444
transform 1 0 11592 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_122
timestamp 1635444444
transform 1 0 12328 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_127
timestamp 1635444444
transform 1 0 12788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1068_
timestamp 1635444444
transform -1 0 12788 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1148_
timestamp 1635444444
transform 1 0 11224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1635444444
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_145
timestamp 1635444444
transform 1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1635444444
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1542_
timestamp 1635444444
transform -1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1772_
timestamp 1635444444
transform -1 0 15640 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_30_158
timestamp 1635444444
transform 1 0 15640 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  _1371_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 16192 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_180
timestamp 1635444444
transform 1 0 17664 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_188
timestamp 1635444444
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1635444444
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1586_
timestamp 1635444444
transform -1 0 18400 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_206
timestamp 1635444444
transform 1 0 20056 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1635444444
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1626_
timestamp 1635444444
transform -1 0 20700 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1781_
timestamp 1635444444
transform 1 0 21068 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1788_
timestamp 1635444444
transform 1 0 19228 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_226
timestamp 1635444444
transform 1 0 21896 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_238
timestamp 1635444444
transform 1 0 23000 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1635444444
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1635444444
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1635444444
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1635444444
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1635444444
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1635444444
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1635444444
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1635444444
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_309
timestamp 1635444444
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_317
timestamp 1635444444
transform 1 0 30268 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1635444444
transform -1 0 30820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1635444444
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_13
timestamp 1635444444
transform 1 0 2300 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_19
timestamp 1635444444
transform 1 0 2852 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 1635444444
transform 1 0 1380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1635444444
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1132_
timestamp 1635444444
transform -1 0 3864 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1137_
timestamp 1635444444
transform 1 0 1472 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_30
timestamp 1635444444
transform 1 0 3864 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1635444444
transform 1 0 4232 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_31_50
timestamp 1635444444
transform 1 0 5704 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1635444444
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_61
timestamp 1635444444
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1635444444
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1862_
timestamp 1635444444
transform 1 0 6808 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1635444444
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1442_
timestamp 1635444444
transform -1 0 9292 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_102
timestamp 1635444444
transform 1 0 10488 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_89
timestamp 1635444444
transform 1 0 9292 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1635444444
transform -1 0 10488 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1635444444
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1635444444
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1635444444
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 11868 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 1635444444
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1958_
timestamp 1635444444
transform -1 0 15548 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_157
timestamp 1635444444
transform 1 0 15548 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1635444444
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1635444444
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1635444444
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1524_
timestamp 1635444444
transform -1 0 17112 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_31_178
timestamp 1635444444
transform 1 0 17480 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_188
timestamp 1635444444
transform 1 0 18400 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1776_
timestamp 1635444444
transform 1 0 17572 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1815_
timestamp 1635444444
transform 1 0 18768 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_31_201
timestamp 1635444444
transform 1 0 19596 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_207
timestamp 1635444444
transform 1 0 20148 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1635444444
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1779_
timestamp 1635444444
transform 1 0 20240 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1635444444
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1635444444
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1635444444
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1635444444
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1635444444
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1635444444
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1635444444
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1635444444
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1635444444
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1635444444
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1635444444
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_305
timestamp 1635444444
transform 1 0 29164 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_311
timestamp 1635444444
transform 1 0 29716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_316
timestamp 1635444444
transform 1 0 30176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1635444444
transform -1 0 30820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1635444444
transform 1 0 29808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1635444444
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1635444444
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1635444444
transform 1 0 1748 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1635444444
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1635444444
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_38
timestamp 1635444444
transform 1 0 4600 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1635444444
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1133_
timestamp 1635444444
transform 1 0 3772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_46
timestamp 1635444444
transform 1 0 5336 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_51
timestamp 1635444444
transform 1 0 5796 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_64
timestamp 1635444444
transform 1 0 6992 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 1635444444
transform -1 0 5796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1284_
timestamp 1635444444
transform 1 0 6164 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_75
timestamp 1635444444
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1635444444
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1635444444
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1635444444
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1278_
timestamp 1635444444
transform -1 0 8004 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_32_109
timestamp 1635444444
transform 1 0 11132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1635444444
transform 1 0 9292 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1635444444
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1388_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 10396 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1390_
timestamp 1635444444
transform 1 0 9384 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_32_129
timestamp 1635444444
transform 1 0 12972 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1635444444
transform 1 0 11500 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1635444444
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_149
timestamp 1635444444
transform 1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1635444444
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1635444444
transform -1 0 13616 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_164
timestamp 1635444444
transform 1 0 16192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_172
timestamp 1635444444
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1526_
timestamp 1635444444
transform -1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 15548 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_32_185
timestamp 1635444444
transform 1 0 18124 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1635444444
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1635444444
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1777_
timestamp 1635444444
transform 1 0 17296 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_32_200
timestamp 1635444444
transform 1 0 19504 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_206
timestamp 1635444444
transform 1 0 20056 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_214
timestamp 1635444444
transform 1 0 20792 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1635444444
transform -1 0 19504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1627_
timestamp 1635444444
transform 1 0 21160 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1635_
timestamp 1635444444
transform 1 0 20148 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1635444444
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1635444444
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1635444444
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1635444444
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1635444444
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1635444444
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1635444444
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1635444444
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1635444444
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1635444444
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1635444444
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp 1635444444
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_317
timestamp 1635444444
transform 1 0 30268 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1635444444
transform -1 0 30820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1635444444
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1136_
timestamp 1635444444
transform 1 0 1656 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1135_
timestamp 1635444444
transform 1 0 1472 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1635444444
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1635444444
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1635444444
transform 1 0 1380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1635444444
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1635444444
transform 1 0 2852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_13
timestamp 1635444444
transform 1 0 2300 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1635444444
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1635444444
transform 1 0 3036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_22
timestamp 1635444444
transform 1 0 3128 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1635444444
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_32
timestamp 1635444444
transform 1 0 4048 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_39
timestamp 1635444444
transform 1 0 4692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1635444444
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1684_
timestamp 1635444444
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1635444444
transform 1 0 3680 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1635444444
transform 1 0 4416 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1699_
timestamp 1635444444
transform 1 0 5520 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1282_
timestamp 1635444444
transform 1 0 5980 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_51
timestamp 1635444444
transform 1 0 5796 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1635444444
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_44
timestamp 1635444444
transform 1 0 5152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1281_
timestamp 1635444444
transform 1 0 6440 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1635444444
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_62
timestamp 1635444444
transform 1 0 6808 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1635444444
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1635444444
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1400_
timestamp 1635444444
transform -1 0 7728 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_72
timestamp 1635444444
transform 1 0 7728 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_74
timestamp 1635444444
transform 1 0 7912 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_66
timestamp 1635444444
transform 1 0 7176 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1387_
timestamp 1635444444
transform -1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1635444444
transform -1 0 8556 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1635444444
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_81
timestamp 1635444444
transform 1 0 8556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1425_
timestamp 1635444444
transform -1 0 9476 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1300_
timestamp 1635444444
transform -1 0 9384 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1635444444
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1635444444
transform 1 0 9844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_90
timestamp 1635444444
transform 1 0 9384 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_91
timestamp 1635444444
transform 1 0 9476 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0979_
timestamp 1635444444
transform -1 0 10672 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0883_
timestamp 1635444444
transform 1 0 10488 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_98
timestamp 1635444444
transform 1 0 10120 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_104
timestamp 1635444444
transform 1 0 10672 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_98
timestamp 1635444444
transform 1 0 10120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1189_
timestamp 1635444444
transform -1 0 11408 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1635444444
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_122
timestamp 1635444444
transform 1 0 12328 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_112
timestamp 1635444444
transform 1 0 11408 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_124
timestamp 1635444444
transform 1 0 12512 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_130
timestamp 1635444444
transform 1 0 13064 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1635444444
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1179_
timestamp 1635444444
transform -1 0 13616 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1205_
timestamp 1635444444
transform 1 0 11500 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1635444444
transform 1 0 13432 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1635444444
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1635444444
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_137
timestamp 1635444444
transform 1 0 13708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1770_
timestamp 1635444444
transform -1 0 15640 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1529_
timestamp 1635444444
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 14628 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_148
timestamp 1635444444
transform 1 0 14720 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_144
timestamp 1635444444
transform 1 0 14352 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_147
timestamp 1635444444
transform 1 0 14628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1771_
timestamp 1635444444
transform 1 0 14996 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1635444444
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1635444444
transform 1 0 16928 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_158
timestamp 1635444444
transform 1 0 15640 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1635444444
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1525_
timestamp 1635444444
transform -1 0 16928 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1769_
timestamp 1635444444
transform -1 0 17204 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_184
timestamp 1635444444
transform 1 0 18032 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_188
timestamp 1635444444
transform 1 0 18400 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1635444444
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_175
timestamp 1635444444
transform 1 0 17204 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_188
timestamp 1635444444
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1635444444
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1606_
timestamp 1635444444
transform 1 0 18492 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1778_
timestamp 1635444444
transform 1 0 19136 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1790_
timestamp 1635444444
transform 1 0 17572 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1635444444
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1635444444
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_204
timestamp 1635444444
transform 1 0 19872 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_210
timestamp 1635444444
transform 1 0 20424 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1620_
timestamp 1635444444
transform 1 0 19228 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _1637_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 20332 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1787_
timestamp 1635444444
transform 1 0 20516 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_33_234
timestamp 1635444444
transform 1 0 22632 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_220
timestamp 1635444444
transform 1 0 21344 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_232
timestamp 1635444444
transform 1 0 22448 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1635444444
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1742_
timestamp 1635444444
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_33_246
timestamp 1635444444
transform 1 0 23736 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_258
timestamp 1635444444
transform 1 0 24840 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1635444444
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1635444444
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1635444444
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_270
timestamp 1635444444
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1635444444
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1635444444
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1635444444
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1635444444
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1635444444
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1635444444
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_305
timestamp 1635444444
transform 1 0 29164 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1635444444
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1635444444
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 1635444444
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1635444444
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_309
timestamp 1635444444
transform 1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_316
timestamp 1635444444
transform 1 0 30176 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1635444444
transform -1 0 30820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1635444444
transform -1 0 30820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1635444444
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1734_
timestamp 1635444444
transform 1 0 29900 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1635444444
transform 1 0 29808 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1635444444
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1635444444
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1635444444
transform 1 0 1656 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_22
timestamp 1635444444
transform 1 0 3128 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_29
timestamp 1635444444
transform 1 0 3772 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_37
timestamp 1635444444
transform 1 0 4508 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_43
timestamp 1635444444
transform 1 0 5060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1267_
timestamp 1635444444
transform -1 0 5060 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1635444444
transform 1 0 3496 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1635444444
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1635444444
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1272_
timestamp 1635444444
transform -1 0 7268 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1385_
timestamp 1635444444
transform -1 0 5888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_67
timestamp 1635444444
transform 1 0 7268 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_73
timestamp 1635444444
transform 1 0 7820 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_78
timestamp 1635444444
transform 1 0 8280 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1303_
timestamp 1635444444
transform 1 0 8648 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1397_
timestamp 1635444444
transform -1 0 8280 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_103
timestamp 1635444444
transform 1 0 10580 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1635444444
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_92
timestamp 1635444444
transform 1 0 9568 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_99
timestamp 1635444444
transform 1 0 10212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1204_
timestamp 1635444444
transform 1 0 10672 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1389_
timestamp 1635444444
transform -1 0 10212 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1635444444
transform 1 0 11500 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_130
timestamp 1635444444
transform 1 0 13064 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1635444444
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1635444444
transform 1 0 11592 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_35_142
timestamp 1635444444
transform 1 0 14168 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_150
timestamp 1635444444
transform 1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_162
timestamp 1635444444
transform 1 0 16008 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1635444444
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1537_
timestamp 1635444444
transform 1 0 16652 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1766_
timestamp 1635444444
transform -1 0 16008 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1635444444
transform 1 0 17480 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_191
timestamp 1635444444
transform 1 0 18676 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  _1622_
timestamp 1635444444
transform 1 0 19044 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1791_
timestamp 1635444444
transform 1 0 17848 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1635444444
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_211
timestamp 1635444444
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1636_
timestamp 1635444444
transform 1 0 20056 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1635444444
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1635444444
transform 1 0 22264 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1635444444
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _0913_
timestamp 1635444444
transform -1 0 22264 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_35_242
timestamp 1635444444
transform 1 0 23368 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_254
timestamp 1635444444
transform 1 0 24472 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_266
timestamp 1635444444
transform 1 0 25576 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1635444444
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1635444444
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1635444444
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1635444444
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1635444444
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_317
timestamp 1635444444
transform 1 0 30268 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1635444444
transform -1 0 30820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1635444444
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1635444444
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1635444444
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1635444444
transform 1 0 1840 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1635444444
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp 1635444444
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_37
timestamp 1635444444
transform 1 0 4508 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1635444444
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1268_
timestamp 1635444444
transform -1 0 5612 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_36_49
timestamp 1635444444
transform 1 0 5612 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1635444444
transform 1 0 6164 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_71
timestamp 1635444444
transform 1 0 7636 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_79
timestamp 1635444444
transform 1 0 8372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1635444444
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1635444444
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1302_
timestamp 1635444444
transform 1 0 8924 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_wb_clk_i
timestamp 1635444444
transform 1 0 8004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_108
timestamp 1635444444
transform 1 0 11040 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_95
timestamp 1635444444
transform 1 0 9844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1309_
timestamp 1635444444
transform 1 0 10212 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_36_123
timestamp 1635444444
transform 1 0 12420 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _1216_
timestamp 1635444444
transform 1 0 11592 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_135
timestamp 1635444444
transform 1 0 13524 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1635444444
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1635444444
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1635444444
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_153
timestamp 1635444444
transform 1 0 15180 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_161
timestamp 1635444444
transform 1 0 15916 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_1  _1536_
timestamp 1635444444
transform 1 0 15364 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_1  _1538_
timestamp 1635444444
transform 1 0 16652 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_36_176
timestamp 1635444444
transform 1 0 17296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1635444444
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1635444444
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1635444444
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1805_
timestamp 1635444444
transform 1 0 17664 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_36_202
timestamp 1635444444
transform 1 0 19688 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_210
timestamp 1635444444
transform 1 0 20424 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _1621_
timestamp 1635444444
transform -1 0 19688 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1801_
timestamp 1635444444
transform 1 0 20608 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_221
timestamp 1635444444
transform 1 0 21436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_234
timestamp 1635444444
transform 1 0 22632 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1800_
timestamp 1635444444
transform 1 0 21804 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_36_246
timestamp 1635444444
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1635444444
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1635444444
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1635444444
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1635444444
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1635444444
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1635444444
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1635444444
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_309
timestamp 1635444444
transform 1 0 29532 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_317
timestamp 1635444444
transform 1 0 30268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1635444444
transform -1 0 30820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1635444444
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_13
timestamp 1635444444
transform 1 0 2300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_20
timestamp 1635444444
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_6
timestamp 1635444444
transform 1 0 1656 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1635444444
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1635444444
transform -1 0 1656 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1635444444
transform -1 0 2300 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1635444444
transform -1 0 2944 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1635444444
transform 1 0 4048 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 1635444444
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1635444444
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1280_
timestamp 1635444444
transform -1 0 7176 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_37_66
timestamp 1635444444
transform 1 0 7176 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1635444444
transform 1 0 7728 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1635444444
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_88
timestamp 1635444444
transform 1 0 9200 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1635444444
transform -1 0 11040 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_37_122
timestamp 1635444444
transform 1 0 12328 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1635444444
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1218_
timestamp 1635444444
transform 1 0 11500 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1635444444
transform 1 0 12696 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_37_142
timestamp 1635444444
transform 1 0 14168 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1635444444
transform 1 0 14996 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1543_
timestamp 1635444444
transform 1 0 14720 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1635444444
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1635444444
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1635444444
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1820_
timestamp 1635444444
transform 1 0 16652 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_37_178
timestamp 1635444444
transform 1 0 17480 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_186
timestamp 1635444444
transform 1 0 18216 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _1765_
timestamp 1635444444
transform -1 0 19228 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_197
timestamp 1635444444
transform 1 0 19228 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_210
timestamp 1635444444
transform 1 0 20424 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1040_
timestamp 1635444444
transform -1 0 21252 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1783_
timestamp 1635444444
transform 1 0 19596 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 1635444444
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1635444444
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_225
timestamp 1635444444
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1635444444
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_8  _1738_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 24288 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_37_252
timestamp 1635444444
transform 1 0 24288 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_264
timestamp 1635444444
transform 1 0 25392 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1635444444
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1635444444
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1635444444
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1635444444
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_305
timestamp 1635444444
transform 1 0 29164 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_311
timestamp 1635444444
transform 1 0 29716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_316
timestamp 1635444444
transform 1 0 30176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1635444444
transform -1 0 30820 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1635444444
transform 1 0 29808 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_18
timestamp 1635444444
transform 1 0 2760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_6
timestamp 1635444444
transform 1 0 1656 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1635444444
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1635444444
transform -1 0 1656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1635444444
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1635444444
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1635444444
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1635444444
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1276_
timestamp 1635444444
transform -1 0 4968 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1635444444
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1635444444
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_38_75
timestamp 1635444444
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1635444444
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1635444444
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1301_
timestamp 1635444444
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1391_
timestamp 1635444444
transform -1 0 8004 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_38_88
timestamp 1635444444
transform 1 0 9200 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _1849_
timestamp 1635444444
transform 1 0 9752 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_38_111
timestamp 1635444444
transform 1 0 11316 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_119
timestamp 1635444444
transform 1 0 12052 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1635444444
transform 1 0 12144 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1635444444
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1635444444
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_147
timestamp 1635444444
transform 1 0 14628 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1635444444
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_1  _1609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 15272 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_154
timestamp 1635444444
transform 1 0 15272 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_161
timestamp 1635444444
transform 1 0 15916 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_165
timestamp 1635444444
transform 1 0 16284 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1629_
timestamp 1635444444
transform 1 0 15640 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1819_
timestamp 1635444444
transform -1 0 17204 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_175
timestamp 1635444444
transform 1 0 17204 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_179
timestamp 1635444444
transform 1 0 17572 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_183
timestamp 1635444444
transform 1 0 17940 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1635444444
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1635444444
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1530_
timestamp 1635444444
transform -1 0 18584 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1533_
timestamp 1635444444
transform -1 0 17940 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_203
timestamp 1635444444
transform 1 0 19780 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_214
timestamp 1635444444
transform 1 0 20792 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1041_
timestamp 1635444444
transform -1 0 19780 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1042_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 20148 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_38_231
timestamp 1635444444
transform 1 0 22356 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_240
timestamp 1635444444
transform 1 0 23184 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _1033_
timestamp 1635444444
transform -1 0 22356 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1035_
timestamp 1635444444
transform -1 0 23184 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1635444444
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1635444444
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1635444444
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1635444444
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1635444444
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1635444444
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1635444444
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 1635444444
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_317
timestamp 1635444444
transform 1 0 30268 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1635444444
transform -1 0 30820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1635444444
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_13
timestamp 1635444444
transform 1 0 2300 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_19
timestamp 1635444444
transform 1 0 2852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_7
timestamp 1635444444
transform 1 0 1748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1635444444
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1635444444
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1392_
timestamp 1635444444
transform -1 0 3312 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1635444444
transform 1 0 1380 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1635444444
transform -1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_25
timestamp 1635444444
transform 1 0 3404 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_40
timestamp 1635444444
transform 1 0 4784 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1635444444
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1635444444
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1273_
timestamp 1635444444
transform -1 0 4784 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1867_
timestamp 1635444444
transform 1 0 3772 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_wb_clk_i
timestamp 1635444444
transform -1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1275_
timestamp 1635444444
transform -1 0 6532 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_46
timestamp 1635444444
transform 1 0 5336 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1635444444
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1796_
timestamp 1635444444
transform 1 0 6900 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1386_
timestamp 1635444444
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1635444444
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_59
timestamp 1635444444
transform 1 0 6532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_60
timestamp 1635444444
transform 1 0 6624 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1635444444
transform -1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_64
timestamp 1635444444
transform 1 0 6992 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1308_
timestamp 1635444444
transform -1 0 8648 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_72
timestamp 1635444444
transform 1 0 7728 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_73
timestamp 1635444444
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1635444444
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1401_
timestamp 1635444444
transform -1 0 9568 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1396_
timestamp 1635444444
transform -1 0 8372 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1635444444
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1635444444
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_79
timestamp 1635444444
transform 1 0 8372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_82
timestamp 1635444444
transform 1 0 8648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1306_
timestamp 1635444444
transform 1 0 9016 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_39_103
timestamp 1635444444
transform 1 0 10580 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1635444444
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_95
timestamp 1635444444
transform 1 0 9844 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_103
timestamp 1635444444
transform 1 0 10580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_92
timestamp 1635444444
transform 1 0 9568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1414_
timestamp 1635444444
transform -1 0 11224 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1418_
timestamp 1635444444
transform 1 0 9936 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_wb_clk_i
timestamp 1635444444
transform 1 0 10672 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_122
timestamp 1635444444
transform 1 0 12328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_110
timestamp 1635444444
transform 1 0 11224 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_116
timestamp 1635444444
transform 1 0 11776 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_126
timestamp 1635444444
transform 1 0 12696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1635444444
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1190_
timestamp 1635444444
transform 1 0 11500 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1202_
timestamp 1635444444
transform 1 0 11868 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1416_
timestamp 1635444444
transform 1 0 13064 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1635444444
transform 1 0 12696 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1635444444
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1635444444
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 14444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1607_
timestamp 1635444444
transform 1 0 14536 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1635444444
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_145
timestamp 1635444444
transform 1 0 14444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_141
timestamp 1635444444
transform 1 0 14076 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_142
timestamp 1635444444
transform 1 0 14168 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1630_
timestamp 1635444444
transform 1 0 14812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_151
timestamp 1635444444
transform 1 0 14996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1635444444
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_157
timestamp 1635444444
transform 1 0 15548 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_161
timestamp 1635444444
transform 1 0 15916 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_171
timestamp 1635444444
transform 1 0 16836 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1635444444
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1557_
timestamp 1635444444
transform 1 0 16008 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o221ai_2  _1558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1789_
timestamp 1635444444
transform -1 0 16192 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_39_181
timestamp 1635444444
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_194
timestamp 1635444444
transform 1 0 18952 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_177
timestamp 1635444444
transform 1 0 17388 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_187
timestamp 1635444444
transform 1 0 18308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1635444444
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1635444444
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1775_
timestamp 1635444444
transform -1 0 18308 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1804_
timestamp 1635444444
transform 1 0 18124 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1635444444
transform -1 0 19780 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1037_
timestamp 1635444444
transform -1 0 20332 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1635444444
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_200
timestamp 1635444444
transform 1 0 19504 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_203
timestamp 1635444444
transform 1 0 19780 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1039_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 20148 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_4  _0894_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 21620 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1635444444
transform 1 0 20700 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1635444444
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1635444444
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0912_
timestamp 1635444444
transform 1 0 22172 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0911_
timestamp 1635444444
transform 1 0 21988 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1635444444
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_223
timestamp 1635444444
transform 1 0 21620 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1635444444
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1635444444
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0886_
timestamp 1635444444
transform -1 0 23184 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_240
timestamp 1635444444
transform 1 0 23184 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_232
timestamp 1635444444
transform 1 0 22448 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_239
timestamp 1635444444
transform 1 0 23092 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_246
timestamp 1635444444
transform 1 0 23736 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_258
timestamp 1635444444
transform 1 0 24840 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1635444444
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1635444444
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1635444444
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1635444444
transform 1 0 23460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0893_
timestamp 1635444444
transform -1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_270
timestamp 1635444444
transform 1 0 25944 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1635444444
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1635444444
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1635444444
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1635444444
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1635444444
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1635444444
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_305
timestamp 1635444444
transform 1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1635444444
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1635444444
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_316
timestamp 1635444444
transform 1 0 30176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1635444444
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_309
timestamp 1635444444
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_316
timestamp 1635444444
transform 1 0 30176 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1635444444
transform -1 0 30820 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1635444444
transform -1 0 30820 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1635444444
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1735_
timestamp 1635444444
transform 1 0 29900 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1635444444
transform 1 0 29808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_19
timestamp 1635444444
transform 1 0 2852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_7
timestamp 1635444444
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1635444444
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1635444444
transform -1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_25
timestamp 1635444444
transform 1 0 3404 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_33
timestamp 1635444444
transform 1 0 4140 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1403_
timestamp 1635444444
transform -1 0 3404 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1635444444
transform -1 0 5888 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1635444444
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_57
timestamp 1635444444
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1635444444
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1402_
timestamp 1635444444
transform -1 0 7728 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_41_72
timestamp 1635444444
transform 1 0 7728 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_79
timestamp 1635444444
transform 1 0 8372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_85
timestamp 1635444444
transform 1 0 8924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1307_
timestamp 1635444444
transform 1 0 9016 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1398_
timestamp 1635444444
transform 1 0 8096 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_107
timestamp 1635444444
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_94
timestamp 1635444444
transform 1 0 9752 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1212_
timestamp 1635444444
transform -1 0 10948 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1635444444
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_122
timestamp 1635444444
transform 1 0 12328 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1635444444
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1214_
timestamp 1635444444
transform 1 0 11500 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1635444444
transform -1 0 14352 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_144
timestamp 1635444444
transform 1 0 14352 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_151
timestamp 1635444444
transform 1 0 14996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1544_
timestamp 1635444444
transform 1 0 14720 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1635444444
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1635444444
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_172
timestamp 1635444444
transform 1 0 16928 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1635444444
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1590_
timestamp 1635444444
transform 1 0 15364 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1628_
timestamp 1635444444
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_185
timestamp 1635444444
transform 1 0 18124 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_194
timestamp 1635444444
transform 1 0 18952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1531_
timestamp 1635444444
transform 1 0 18676 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1774_
timestamp 1635444444
transform -1 0 18124 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_41_201
timestamp 1635444444
transform 1 0 19596 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_208
timestamp 1635444444
transform 1 0 20240 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1635444444
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1635444444
transform -1 0 21068 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1635444444
transform -1 0 19596 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1527_
timestamp 1635444444
transform 1 0 19964 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1635444444
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_234
timestamp 1635444444
transform 1 0 22632 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1635444444
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0892_
timestamp 1635444444
transform 1 0 23000 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1802_
timestamp 1635444444
transform 1 0 21804 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_41_243
timestamp 1635444444
transform 1 0 23460 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_255
timestamp 1635444444
transform 1 0 24564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_267
timestamp 1635444444
transform 1 0 25668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1635444444
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1635444444
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1635444444
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1635444444
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1635444444
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_317
timestamp 1635444444
transform 1 0 30268 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1635444444
transform -1 0 30820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1635444444
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1635444444
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1635444444
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1635444444
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1635444444
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_41
timestamp 1635444444
transform 1 0 4876 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1635444444
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_47
timestamp 1635444444
transform 1 0 5428 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_52
timestamp 1635444444
transform 1 0 5888 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_59
timestamp 1635444444
transform 1 0 6532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1415_
timestamp 1635444444
transform 1 0 6256 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1795_
timestamp 1635444444
transform 1 0 6900 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_wb_clk_i
timestamp 1635444444
transform -1 0 5888 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_72
timestamp 1635444444
transform 1 0 7728 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_79
timestamp 1635444444
transform 1 0 8372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1635444444
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1635444444
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1399_
timestamp 1635444444
transform 1 0 8096 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1419_
timestamp 1635444444
transform -1 0 9752 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_42_102
timestamp 1635444444
transform 1 0 10488 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_94
timestamp 1635444444
transform 1 0 9752 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_98
timestamp 1635444444
transform 1 0 10120 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1208_
timestamp 1635444444
transform -1 0 10488 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_126
timestamp 1635444444
transform 1 0 12696 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1635444444
transform 1 0 11224 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1635444444
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_144
timestamp 1635444444
transform 1 0 14352 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_152
timestamp 1635444444
transform 1 0 15088 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1635444444
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1587_
timestamp 1635444444
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_wb_clk_i
timestamp 1635444444
transform 1 0 14720 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_158
timestamp 1635444444
transform 1 0 15640 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_164
timestamp 1635444444
transform 1 0 16192 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_168
timestamp 1635444444
transform 1 0 16560 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1556_
timestamp 1635444444
transform -1 0 16192 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1786_
timestamp 1635444444
transform -1 0 17480 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_42_178
timestamp 1635444444
transform 1 0 17480 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_186
timestamp 1635444444
transform 1 0 18216 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1635444444
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1635444444
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1532_
timestamp 1635444444
transform -1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_197
timestamp 1635444444
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_204
timestamp 1635444444
transform 1 0 19872 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_216
timestamp 1635444444
transform 1 0 20976 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1050_
timestamp 1635444444
transform 1 0 19504 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1051_
timestamp 1635444444
transform 1 0 20240 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_222
timestamp 1635444444
transform 1 0 21528 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_226
timestamp 1635444444
transform 1 0 21896 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_238
timestamp 1635444444
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1635444444
transform 1 0 21620 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1635444444
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1635444444
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1635444444
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1635444444
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1635444444
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1635444444
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1635444444
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1635444444
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_309
timestamp 1635444444
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_317
timestamp 1635444444
transform 1 0 30268 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1635444444
transform -1 0 30820 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1635444444
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_19
timestamp 1635444444
transform 1 0 2852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_7
timestamp 1635444444
transform 1 0 1748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1635444444
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1635444444
transform -1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_25
timestamp 1635444444
transform 1 0 3404 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _1269_
timestamp 1635444444
transform -1 0 5244 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1420_
timestamp 1635444444
transform -1 0 3404 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_45
timestamp 1635444444
transform 1 0 5244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1635444444
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_64
timestamp 1635444444
transform 1 0 6992 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1635444444
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__o31a_1  _1196_
timestamp 1635444444
transform -1 0 6992 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1408_
timestamp 1635444444
transform -1 0 5888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_74
timestamp 1635444444
transform 1 0 7912 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_87
timestamp 1635444444
transform 1 0 9108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1793_
timestamp 1635444444
transform 1 0 8280 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1635444444
transform -1 0 7912 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1635444444
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1848_
timestamp 1635444444
transform 1 0 9476 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1635444444
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_117
timestamp 1635444444
transform 1 0 11868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_127
timestamp 1635444444
transform 1 0 12788 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1635444444
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1200_
timestamp 1635444444
transform 1 0 11960 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1635444444
transform -1 0 13524 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_135
timestamp 1635444444
transform 1 0 13524 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_147
timestamp 1635444444
transform 1 0 14628 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_151
timestamp 1635444444
transform 1 0 14996 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1588_
timestamp 1635444444
transform 1 0 14720 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1635444444
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1635444444
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1635444444
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1565_
timestamp 1635444444
transform 1 0 16928 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1780_
timestamp 1635444444
transform -1 0 16192 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_43_175
timestamp 1635444444
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_188
timestamp 1635444444
transform 1 0 18400 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_196
timestamp 1635444444
transform 1 0 19136 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1816_
timestamp 1635444444
transform 1 0 17572 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_43_207
timestamp 1635444444
transform 1 0 20148 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1056_
timestamp 1635444444
transform 1 0 19412 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1058_
timestamp 1635444444
transform 1 0 20516 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1635444444
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_228
timestamp 1635444444
transform 1 0 22080 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_240
timestamp 1635444444
transform 1 0 23184 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1635444444
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1635444444
transform -1 0 22080 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_252
timestamp 1635444444
transform 1 0 24288 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_264
timestamp 1635444444
transform 1 0 25392 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1635444444
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1635444444
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1635444444
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1635444444
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_305
timestamp 1635444444
transform 1 0 29164 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_311
timestamp 1635444444
transform 1 0 29716 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_316
timestamp 1635444444
transform 1 0 30176 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1635444444
transform -1 0 30820 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1635444444
transform 1 0 29808 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_19
timestamp 1635444444
transform 1 0 2852 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_7
timestamp 1635444444
transform 1 0 1748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1635444444
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1411_
timestamp 1635444444
transform -1 0 3312 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1635444444
transform -1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1635444444
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1635444444
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1635444444
transform -1 0 5244 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_44_45
timestamp 1635444444
transform 1 0 5244 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_57
timestamp 1635444444
transform 1 0 6348 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_63
timestamp 1635444444
transform 1 0 6900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1274_
timestamp 1635444444
transform -1 0 6348 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1794_
timestamp 1635444444
transform 1 0 6992 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_73
timestamp 1635444444
transform 1 0 7820 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1635444444
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_85
timestamp 1635444444
transform 1 0 8924 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1635444444
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1305_
timestamp 1635444444
transform 1 0 9016 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1406_
timestamp 1635444444
transform -1 0 8464 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_101
timestamp 1635444444
transform 1 0 10396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_94
timestamp 1635444444
transform 1 0 9752 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1417_
timestamp 1635444444
transform -1 0 10396 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_113
timestamp 1635444444
transform 1 0 11500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_126
timestamp 1635444444
transform 1 0 12696 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _1197_
timestamp 1635444444
transform 1 0 11868 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1635444444
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_141
timestamp 1635444444
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_147
timestamp 1635444444
transform 1 0 14628 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1635444444
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1545_
timestamp 1635444444
transform 1 0 14996 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1589_
timestamp 1635444444
transform 1 0 14168 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_44_154
timestamp 1635444444
transform 1 0 15272 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_161
timestamp 1635444444
transform 1 0 15916 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_168
timestamp 1635444444
transform 1 0 16560 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1546_
timestamp 1635444444
transform 1 0 15640 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1570_
timestamp 1635444444
transform -1 0 16560 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_176
timestamp 1635444444
transform 1 0 17296 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_182
timestamp 1635444444
transform 1 0 17848 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1635444444
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1635444444
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1635444444
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1600_
timestamp 1635444444
transform 1 0 17388 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1603_
timestamp 1635444444
transform 1 0 18216 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1635444444
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_206
timestamp 1635444444
transform 1 0 20056 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_210
timestamp 1635444444
transform 1 0 20424 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1052_
timestamp 1635444444
transform 1 0 20516 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o211ai_1  _1057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 19504 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_220
timestamp 1635444444
transform 1 0 21344 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_240
timestamp 1635444444
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1960_
timestamp 1635444444
transform 1 0 21712 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1635444444
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1635444444
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1635444444
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1635444444
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1635444444
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1635444444
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1635444444
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_309
timestamp 1635444444
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_317
timestamp 1635444444
transform 1 0 30268 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1635444444
transform -1 0 30820 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1635444444
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_19
timestamp 1635444444
transform 1 0 2852 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_7
timestamp 1635444444
transform 1 0 1748 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1635444444
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1635444444
transform -1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_31
timestamp 1635444444
transform 1 0 3956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1868_
timestamp 1635444444
transform -1 0 5888 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1635444444
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_61
timestamp 1635444444
transform 1 0 6716 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1635444444
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1410_
timestamp 1635444444
transform 1 0 7084 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1635444444
transform -1 0 6716 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_74
timestamp 1635444444
transform 1 0 7912 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_78
timestamp 1635444444
transform 1 0 8280 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_83
timestamp 1635444444
transform 1 0 8740 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1304_
timestamp 1635444444
transform 1 0 9108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1635444444
transform -1 0 8740 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1635444444
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_95
timestamp 1635444444
transform 1 0 9844 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1199_
timestamp 1635444444
transform 1 0 10212 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1635444444
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_121
timestamp 1635444444
transform 1 0 12236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1635444444
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1635444444
transform 1 0 12604 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1635444444
transform 1 0 11868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_141
timestamp 1635444444
transform 1 0 14076 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1568_
timestamp 1635444444
transform -1 0 15272 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_154
timestamp 1635444444
transform 1 0 15272 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1635444444
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1635444444
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1635444444
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1635444444
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1569_
timestamp 1635444444
transform 1 0 15640 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1803_
timestamp 1635444444
transform 1 0 16836 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_180
timestamp 1635444444
transform 1 0 17664 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_184
timestamp 1635444444
transform 1 0 18032 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_194
timestamp 1635444444
transform 1 0 18952 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1813_
timestamp 1635444444
transform 1 0 18124 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1635444444
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_215
timestamp 1635444444
transform 1 0 20884 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0888_
timestamp 1635444444
transform -1 0 19964 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1054_
timestamp 1635444444
transform -1 0 20884 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1635444444
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1635444444
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1959_
timestamp 1635444444
transform 1 0 21804 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_45_241
timestamp 1635444444
transform 1 0 23276 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_253
timestamp 1635444444
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_265
timestamp 1635444444
transform 1 0 25484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1635444444
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1635444444
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1635444444
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1635444444
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_305
timestamp 1635444444
transform 1 0 29164 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_316
timestamp 1635444444
transform 1 0 30176 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1635444444
transform -1 0 30820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1736_
timestamp 1635444444
transform 1 0 29900 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1635444444
transform -1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1635444444
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1635444444
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_7
timestamp 1635444444
transform 1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1456_
timestamp 1635444444
transform 1 0 2116 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1427_
timestamp 1635444444
transform -1 0 3312 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1083_
timestamp 1635444444
transform 1 0 2852 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_18
timestamp 1635444444
transform 1 0 2760 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_14
timestamp 1635444444
transform 1 0 2392 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_15
timestamp 1635444444
transform 1 0 2484 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1635444444
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1433_
timestamp 1635444444
transform -1 0 3864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1635444444
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_23
timestamp 1635444444
transform 1 0 3220 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1635444444
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1635444444
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1082_
timestamp 1635444444
transform -1 0 4600 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_38
timestamp 1635444444
transform 1 0 4600 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_33
timestamp 1635444444
transform 1 0 4140 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_42
timestamp 1635444444
transform 1 0 4968 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_30
timestamp 1635444444
transform 1 0 3864 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__o31a_1  _1198_
timestamp 1635444444
transform -1 0 6164 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_46_46
timestamp 1635444444
transform 1 0 5336 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _1438_
timestamp 1635444444
transform -1 0 6808 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1191_
timestamp 1635444444
transform 1 0 6532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1635444444
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1635444444
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1635444444
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_55
timestamp 1635444444
transform 1 0 6164 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_62
timestamp 1635444444
transform 1 0 6808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_62
timestamp 1635444444
transform 1 0 6808 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1437_
timestamp 1635444444
transform -1 0 7728 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1409_
timestamp 1635444444
transform 1 0 7176 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_47_72
timestamp 1635444444
transform 1 0 7728 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_73
timestamp 1635444444
transform 1 0 7820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1432_
timestamp 1635444444
transform 1 0 8464 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1426_
timestamp 1635444444
transform 1 0 8924 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1407_
timestamp 1635444444
transform -1 0 8464 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1635444444
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1635444444
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_87
timestamp 1635444444
transform 1 0 9108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_102
timestamp 1635444444
transform 1 0 10488 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_107
timestamp 1635444444
transform 1 0 10948 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_94
timestamp 1635444444
transform 1 0 9752 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1635444444
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_91
timestamp 1635444444
transform 1 0 9476 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1192_
timestamp 1635444444
transform -1 0 10948 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1635444444
transform 1 0 9568 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_46_127
timestamp 1635444444
transform 1 0 12788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_116
timestamp 1635444444
transform 1 0 11776 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_124
timestamp 1635444444
transform 1 0 12512 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1635444444
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1195_
timestamp 1635444444
transform -1 0 12512 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1424_
timestamp 1635444444
transform -1 0 11776 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1635444444
transform 1 0 11316 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1635444444
transform 1 0 12880 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1635444444
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_141
timestamp 1635444444
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_150
timestamp 1635444444
transform 1 0 14904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_144
timestamp 1635444444
transform 1 0 14352 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_152
timestamp 1635444444
transform 1 0 15088 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1635444444
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0916_
timestamp 1635444444
transform -1 0 15088 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1591_
timestamp 1635444444
transform -1 0 14904 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1592_
timestamp 1635444444
transform 1 0 15272 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1567_
timestamp 1635444444
transform 1 0 15456 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1635444444
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_158
timestamp 1635444444
transform 1 0 15640 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1810_
timestamp 1635444444
transform -1 0 17020 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1580_
timestamp 1635444444
transform 1 0 16652 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1635444444
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1635444444
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_174
timestamp 1635444444
transform 1 0 17112 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_173
timestamp 1635444444
transform 1 0 17020 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_181
timestamp 1635444444
transform 1 0 17756 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1635444444
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_191
timestamp 1635444444
transform 1 0 18676 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1635444444
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1601_
timestamp 1635444444
transform 1 0 17848 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1814_
timestamp 1635444444
transform 1 0 17940 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1818_
timestamp 1635444444
transform 1 0 19044 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_46_201
timestamp 1635444444
transform 1 0 19596 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_211
timestamp 1635444444
transform 1 0 20516 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_204
timestamp 1635444444
transform 1 0 19872 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_216
timestamp 1635444444
transform 1 0 20976 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1045_
timestamp 1635444444
transform -1 0 20516 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1047_
timestamp 1635444444
transform -1 0 20976 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1055_
timestamp 1635444444
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_219
timestamp 1635444444
transform 1 0 21252 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_230
timestamp 1635444444
transform 1 0 22264 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_228
timestamp 1635444444
transform 1 0 22080 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_240
timestamp 1635444444
transform 1 0 23184 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1635444444
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0889_
timestamp 1635444444
transform 1 0 21344 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1635444444
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_242
timestamp 1635444444
transform 1 0 23368 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1635444444
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1635444444
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_252
timestamp 1635444444
transform 1 0 24288 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1635444444
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1635444444
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1635444444
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_264
timestamp 1635444444
transform 1 0 25392 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1635444444
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1635444444
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1635444444
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1635444444
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1635444444
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1635444444
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_305
timestamp 1635444444
transform 1 0 29164 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1635444444
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1635444444
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_316
timestamp 1635444444
transform 1 0 30176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_316
timestamp 1635444444
transform 1 0 30176 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1635444444
transform -1 0 30820 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1635444444
transform -1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1635444444
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1718_
timestamp 1635444444
transform 1 0 29900 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1635444444
transform 1 0 29808 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_13
timestamp 1635444444
transform 1 0 2300 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_17
timestamp 1635444444
transform 1 0 2668 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_7
timestamp 1635444444
transform 1 0 1748 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1635444444
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1439_
timestamp 1635444444
transform -1 0 3312 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1444_
timestamp 1635444444
transform 1 0 2392 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1635444444
transform -1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1635444444
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_32
timestamp 1635444444
transform 1 0 4048 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1635444444
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1635444444
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 4048 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1338_
timestamp 1635444444
transform 1 0 4600 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_56
timestamp 1635444444
transform 1 0 6256 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1635444444
transform -1 0 6256 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1798_
timestamp 1635444444
transform 1 0 6624 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_48_69
timestamp 1635444444
transform 1 0 7452 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1635444444
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1635444444
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1431_
timestamp 1635444444
transform -1 0 8464 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1797_
timestamp 1635444444
transform 1 0 8924 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_48_101
timestamp 1635444444
transform 1 0 10396 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_94
timestamp 1635444444
transform 1 0 9752 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1203_
timestamp 1635444444
transform 1 0 10948 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1423_
timestamp 1635444444
transform -1 0 10396 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_111
timestamp 1635444444
transform 1 0 11316 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_119
timestamp 1635444444
transform 1 0 12052 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1188_
timestamp 1635444444
transform 1 0 11684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1194_
timestamp 1635444444
transform -1 0 13340 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1635444444
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1635444444
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_144
timestamp 1635444444
transform 1 0 14352 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_152
timestamp 1635444444
transform 1 0 15088 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1635444444
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0900_
timestamp 1635444444
transform 1 0 14720 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1579_
timestamp 1635444444
transform -1 0 14352 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_160
timestamp 1635444444
transform 1 0 15824 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_168
timestamp 1635444444
transform 1 0 16560 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_173
timestamp 1635444444
transform 1 0 17020 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1564_
timestamp 1635444444
transform -1 0 17020 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_wb_clk_i
timestamp 1635444444
transform 1 0 15456 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_181
timestamp 1635444444
transform 1 0 17756 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_190
timestamp 1635444444
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1635444444
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__o311a_1  _1602_
timestamp 1635444444
transform 1 0 17848 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1635444444
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_205
timestamp 1635444444
transform 1 0 19964 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_214
timestamp 1635444444
transform 1 0 20792 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_1  _1048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 20148 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_48_222
timestamp 1635444444
transform 1 0 21528 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1635444444
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_1  _1367_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 21804 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1635444444
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1635444444
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1635444444
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1635444444
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1635444444
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1635444444
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1635444444
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1635444444
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1635444444
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_309
timestamp 1635444444
transform 1 0 29532 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_316
timestamp 1635444444
transform 1 0 30176 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1635444444
transform -1 0 30820 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1635444444
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1635444444
transform 1 0 29808 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_14
timestamp 1635444444
transform 1 0 2392 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_21
timestamp 1635444444
transform 1 0 3036 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_7
timestamp 1635444444
transform 1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1635444444
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1449_
timestamp 1635444444
transform -1 0 2392 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1453_
timestamp 1635444444
transform 1 0 2760 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1635444444
transform -1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1635444444
transform 1 0 3772 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_49_45
timestamp 1635444444
transform 1 0 5244 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_52
timestamp 1635444444
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_57
timestamp 1635444444
transform 1 0 6348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1635444444
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1339_
timestamp 1635444444
transform 1 0 5612 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1792_
timestamp 1635444444
transform 1 0 6900 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_72
timestamp 1635444444
transform 1 0 7728 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_79
timestamp 1635444444
transform 1 0 8372 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1635444444
transform 1 0 8096 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1799_
timestamp 1635444444
transform 1 0 9108 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_49_104
timestamp 1635444444
transform 1 0 10672 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1635444444
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_96
timestamp 1635444444
transform 1 0 9936 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1635444444
transform -1 0 11040 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1635444444
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_121
timestamp 1635444444
transform 1 0 12236 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_127
timestamp 1635444444
transform 1 0 12788 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1635444444
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1187_
timestamp 1635444444
transform -1 0 12788 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_141
timestamp 1635444444
transform 1 0 14076 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_149
timestamp 1635444444
transform 1 0 14812 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__a221o_1  _1215_
timestamp 1635444444
transform 1 0 13340 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1635444444
transform 1 0 14996 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_49_156
timestamp 1635444444
transform 1 0 15456 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1635444444
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1635444444
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1365_
timestamp 1635444444
transform 1 0 15824 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1806_
timestamp 1635444444
transform 1 0 16652 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_49_178
timestamp 1635444444
transform 1 0 17480 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_193
timestamp 1635444444
transform 1 0 18860 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1599_
timestamp 1635444444
transform 1 0 18216 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_49_203
timestamp 1635444444
transform 1 0 19780 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_211
timestamp 1635444444
transform 1 0 20516 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_218
timestamp 1635444444
transform 1 0 21160 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0920_
timestamp 1635444444
transform 1 0 20792 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1032_
timestamp 1635444444
transform 1 0 19412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1635444444
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1961_
timestamp 1635444444
transform 1 0 21804 0 -1 29376
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_49_244
timestamp 1635444444
transform 1 0 23552 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_256
timestamp 1635444444
transform 1 0 24656 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_268
timestamp 1635444444
transform 1 0 25760 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1635444444
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1635444444
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1635444444
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1635444444
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_317
timestamp 1635444444
transform 1 0 30268 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1635444444
transform -1 0 30820 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_14
timestamp 1635444444
transform 1 0 2392 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_7
timestamp 1635444444
transform 1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1635444444
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1330_
timestamp 1635444444
transform -1 0 3220 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1447_
timestamp 1635444444
transform 1 0 2116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1635444444
transform -1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1635444444
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1635444444
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_32
timestamp 1635444444
transform 1 0 4048 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_39
timestamp 1635444444
transform 1 0 4692 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1635444444
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1329_
timestamp 1635444444
transform -1 0 4048 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1332_
timestamp 1635444444
transform -1 0 4692 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1635444444
transform -1 0 6532 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_59
timestamp 1635444444
transform 1 0 6532 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_wb_clk_i
timestamp 1635444444
transform 1 0 6900 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_67
timestamp 1635444444
transform 1 0 7268 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_74
timestamp 1635444444
transform 1 0 7912 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1635444444
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1635444444
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1635444444
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1436_
timestamp 1635444444
transform 1 0 7636 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_109
timestamp 1635444444
transform 1 0 11132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1635444444
transform 1 0 9660 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_50_117
timestamp 1635444444
transform 1 0 11868 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_131
timestamp 1635444444
transform 1 0 13156 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1181_
timestamp 1635444444
transform 1 0 11500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1185_
timestamp 1635444444
transform 1 0 12236 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1635444444
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_141
timestamp 1635444444
transform 1 0 14076 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1635444444
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1635444444
transform 1 0 14168 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_50_158
timestamp 1635444444
transform 1 0 15640 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1581_
timestamp 1635444444
transform -1 0 17204 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_50_175
timestamp 1635444444
transform 1 0 17204 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1635444444
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1635444444
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1764_
timestamp 1635444444
transform -1 0 18768 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_203
timestamp 1635444444
transform 1 0 19780 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_207
timestamp 1635444444
transform 1 0 20148 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_215
timestamp 1635444444
transform 1 0 20884 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1366_
timestamp 1635444444
transform -1 0 20884 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1582_
timestamp 1635444444
transform -1 0 19780 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_221
timestamp 1635444444
transform 1 0 21436 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_227
timestamp 1635444444
transform 1 0 21988 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1031_
timestamp 1635444444
transform 1 0 21528 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1832_
timestamp 1635444444
transform 1 0 22356 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1635444444
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1635444444
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1635444444
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1635444444
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1635444444
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1635444444
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1635444444
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1635444444
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_309
timestamp 1635444444
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_317
timestamp 1635444444
transform 1 0 30268 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1635444444
transform -1 0 30820 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1635444444
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_15
timestamp 1635444444
transform 1 0 2484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1635444444
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_7
timestamp 1635444444
transform 1 0 1748 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1635444444
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1446_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1840 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1635444444
transform 1 0 2852 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_51_35
timestamp 1635444444
transform 1 0 4324 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_42
timestamp 1635444444
transform 1 0 4968 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1335_
timestamp 1635444444
transform -1 0 4968 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_49
timestamp 1635444444
transform 1 0 5612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1635444444
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1635444444
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1315_
timestamp 1635444444
transform 1 0 5336 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1340_
timestamp 1635444444
transform -1 0 7176 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_51_66
timestamp 1635444444
transform 1 0 7176 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_75
timestamp 1635444444
transform 1 0 8004 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_82
timestamp 1635444444
transform 1 0 8648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_86
timestamp 1635444444
transform 1 0 9016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1395_
timestamp 1635444444
transform 1 0 7728 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1405_
timestamp 1635444444
transform 1 0 8372 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1429_
timestamp 1635444444
transform -1 0 9384 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 1635444444
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_90
timestamp 1635444444
transform 1 0 9384 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1209_
timestamp 1635444444
transform -1 0 11040 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_122
timestamp 1635444444
transform 1 0 12328 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_126
timestamp 1635444444
transform 1 0 12696 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1635444444
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1193_
timestamp 1635444444
transform 1 0 12788 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1213_
timestamp 1635444444
transform 1 0 11500 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_137
timestamp 1635444444
transform 1 0 13708 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_149
timestamp 1635444444
transform 1 0 14812 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1201_
timestamp 1635444444
transform 1 0 14076 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_157
timestamp 1635444444
transform 1 0 15548 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1635444444
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1635444444
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1566_
timestamp 1635444444
transform 1 0 15916 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1807_
timestamp 1635444444
transform 1 0 16652 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1635444444
transform 1 0 15180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_178
timestamp 1635444444
transform 1 0 17480 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_186
timestamp 1635444444
transform 1 0 18216 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0901_
timestamp 1635444444
transform 1 0 17848 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_2  _1373_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 18584 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_51_197
timestamp 1635444444
transform 1 0 19228 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_208
timestamp 1635444444
transform 1 0 20240 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_214
timestamp 1635444444
transform 1 0 20792 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_218
timestamp 1635444444
transform 1 0 21160 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1635444444
transform 1 0 20884 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1030_
timestamp 1635444444
transform -1 0 20240 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_51_225
timestamp 1635444444
transform 1 0 21804 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_233
timestamp 1635444444
transform 1 0 22540 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_238
timestamp 1635444444
transform 1 0 23000 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1635444444
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1368_
timestamp 1635444444
transform 1 0 22724 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_250
timestamp 1635444444
transform 1 0 24104 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_262
timestamp 1635444444
transform 1 0 25208 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_274
timestamp 1635444444
transform 1 0 26312 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1635444444
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1635444444
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1635444444
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1737_
timestamp 1635444444
transform -1 0 29440 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_308
timestamp 1635444444
transform 1 0 29440 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_316
timestamp 1635444444
transform 1 0 30176 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1635444444
transform -1 0 30820 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1635444444
transform 1 0 29808 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_16
timestamp 1635444444
transform 1 0 2576 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_3
timestamp 1635444444
transform 1 0 1380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_16
timestamp 1635444444
transform 1 0 2576 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1635444444
transform 1 0 1380 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1635444444
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1635444444
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1448_
timestamp 1635444444
transform 1 0 1932 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1450_
timestamp 1635444444
transform 1 0 1932 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1635444444
transform 1 0 2944 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1635444444
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_32
timestamp 1635444444
transform 1 0 4048 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_24
timestamp 1635444444
transform 1 0 3312 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_34
timestamp 1635444444
transform 1 0 4232 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1635444444
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1316_
timestamp 1635444444
transform 1 0 4784 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1331_
timestamp 1635444444
transform -1 0 4232 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1334_
timestamp 1635444444
transform -1 0 5244 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1336_
timestamp 1635444444
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_45
timestamp 1635444444
transform 1 0 5244 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_65
timestamp 1635444444
transform 1 0 7084 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_50
timestamp 1635444444
transform 1 0 5704 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1635444444
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1337_
timestamp 1635444444
transform -1 0 7176 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1635444444
transform 1 0 5612 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _1383_
timestamp 1635444444
transform 1 0 7544 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_66
timestamp 1635444444
transform 1 0 7176 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  net99_2
timestamp 1635444444
transform -1 0 8464 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1394_
timestamp 1635444444
transform -1 0 8464 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_73
timestamp 1635444444
transform 1 0 7820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_73
timestamp 1635444444
transform 1 0 7820 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _1404_
timestamp 1635444444
transform -1 0 9476 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1393_
timestamp 1635444444
transform 1 0 8832 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1635444444
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_80
timestamp 1635444444
transform 1 0 8464 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1635444444
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_87
timestamp 1635444444
transform 1 0 9108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1413_
timestamp 1635444444
transform 1 0 9844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1412_
timestamp 1635444444
transform 1 0 9476 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_97
timestamp 1635444444
transform 1 0 10028 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_91
timestamp 1635444444
transform 1 0 9476 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1422_
timestamp 1635444444
transform 1 0 10488 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1421_
timestamp 1635444444
transform 1 0 10396 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1635444444
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_98
timestamp 1635444444
transform 1 0 10120 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_105
timestamp 1635444444
transform 1 0 10764 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1206_
timestamp 1635444444
transform 1 0 11132 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_52_118
timestamp 1635444444
transform 1 0 11960 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1635444444
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_113
timestamp 1635444444
transform 1 0 11500 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_124
timestamp 1635444444
transform 1 0 12512 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1635444444
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1182_
timestamp 1635444444
transform -1 0 13248 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1186_
timestamp 1635444444
transform 1 0 12880 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1207_
timestamp 1635444444
transform -1 0 12512 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1635444444
transform 1 0 13248 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1635444444
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_136
timestamp 1635444444
transform 1 0 13616 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_148
timestamp 1635444444
transform 1 0 14720 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1635444444
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1635444444
transform 1 0 14260 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_52_159
timestamp 1635444444
transform 1 0 15732 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_167
timestamp 1635444444
transform 1 0 16468 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_154
timestamp 1635444444
transform 1 0 15272 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1635444444
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_169
timestamp 1635444444
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1635444444
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1744_
timestamp 1635444444
transform 1 0 15364 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1808_
timestamp 1635444444
transform -1 0 17480 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1812_
timestamp 1635444444
transform -1 0 17756 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_52_178
timestamp 1635444444
transform 1 0 17480 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1635444444
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1635444444
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_181
timestamp 1635444444
transform 1 0 17756 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_196
timestamp 1635444444
transform 1 0 19136 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1635444444
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1578_
timestamp 1635444444
transform -1 0 18492 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1743_
timestamp 1635444444
transform -1 0 19136 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0972_
timestamp 1635444444
transform -1 0 20608 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0922_
timestamp 1635444444
transform 1 0 19964 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_204
timestamp 1635444444
transform 1 0 19872 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_201
timestamp 1635444444
transform 1 0 19596 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1635444444
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1635444444
transform -1 0 20976 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0890_
timestamp 1635444444
transform -1 0 21436 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1635444444
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_209
timestamp 1635444444
transform 1 0 20332 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_212
timestamp 1635444444
transform 1 0 20608 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1635444444
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1635444444
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_228
timestamp 1635444444
transform 1 0 22080 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_240
timestamp 1635444444
transform 1 0 23184 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1635444444
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1635444444
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1635444444
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1635444444
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1635444444
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_252
timestamp 1635444444
transform 1 0 24288 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1635444444
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1635444444
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1635444444
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_264
timestamp 1635444444
transform 1 0 25392 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1635444444
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1635444444
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1635444444
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1635444444
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1635444444
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1635444444
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1635444444
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1635444444
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_309
timestamp 1635444444
transform 1 0 29532 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_316
timestamp 1635444444
transform 1 0 30176 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_317
timestamp 1635444444
transform 1 0 30268 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1635444444
transform -1 0 30820 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1635444444
transform -1 0 30820 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1635444444
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1728_
timestamp 1635444444
transform 1 0 29900 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_16
timestamp 1635444444
transform 1 0 2576 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_3
timestamp 1635444444
transform 1 0 1380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1635444444
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1451_
timestamp 1635444444
transform 1 0 2944 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1452_
timestamp 1635444444
transform 1 0 1932 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_54_23
timestamp 1635444444
transform 1 0 3220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1635444444
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_29
timestamp 1635444444
transform 1 0 3772 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_36
timestamp 1635444444
transform 1 0 4416 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1635444444
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1314_
timestamp 1635444444
transform -1 0 4416 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1320_
timestamp 1635444444
transform -1 0 5704 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_54_50
timestamp 1635444444
transform 1 0 5704 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_54
timestamp 1635444444
transform 1 0 6072 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_58
timestamp 1635444444
transform 1 0 6440 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_65
timestamp 1635444444
transform 1 0 7084 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0957_
timestamp 1635444444
transform 1 0 6808 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0961_
timestamp 1635444444
transform 1 0 6164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_72
timestamp 1635444444
transform 1 0 7728 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_79
timestamp 1635444444
transform 1 0 8372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1635444444
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_85
timestamp 1635444444
transform 1 0 8924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1635444444
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0960_
timestamp 1635444444
transform -1 0 7728 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1635444444
transform 1 0 8096 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_105
timestamp 1635444444
transform 1 0 10764 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_109
timestamp 1635444444
transform 1 0 11132 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_97
timestamp 1635444444
transform 1 0 10028 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1217_
timestamp 1635444444
transform 1 0 10396 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1428_
timestamp 1635444444
transform -1 0 10028 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_126
timestamp 1635444444
transform 1 0 12696 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1635444444
transform 1 0 11224 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_wb_clk_i
timestamp 1635444444
transform -1 0 13432 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_134
timestamp 1635444444
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1635444444
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1635444444
transform 1 0 14076 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_54_157
timestamp 1635444444
transform 1 0 15548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_169
timestamp 1635444444
transform 1 0 16652 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_181
timestamp 1635444444
transform 1 0 17756 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_187
timestamp 1635444444
transform 1 0 18308 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1635444444
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1635444444
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1343_
timestamp 1635444444
transform -1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_197
timestamp 1635444444
transform 1 0 19228 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_205
timestamp 1635444444
transform 1 0 19964 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_209
timestamp 1635444444
transform 1 0 20332 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0923_
timestamp 1635444444
transform -1 0 19964 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _1313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 21252 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_54_219
timestamp 1635444444
transform 1 0 21252 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_231
timestamp 1635444444
transform 1 0 22356 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_243
timestamp 1635444444
transform 1 0 23460 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1635444444
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1635444444
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1635444444
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1635444444
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1635444444
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1635444444
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1635444444
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1635444444
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_309
timestamp 1635444444
transform 1 0 29532 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_316
timestamp 1635444444
transform 1 0 30176 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1635444444
transform -1 0 30820 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1635444444
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1635444444
transform 1 0 29808 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_15
timestamp 1635444444
transform 1 0 2484 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_21
timestamp 1635444444
transform 1 0 3036 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_7
timestamp 1635444444
transform 1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1635444444
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1635444444
transform -1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1635444444
transform -1 0 2484 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_25
timestamp 1635444444
transform 1 0 3404 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_38
timestamp 1635444444
transform 1 0 4600 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1326_
timestamp 1635444444
transform 1 0 3128 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1327_
timestamp 1635444444
transform -1 0 4600 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1635444444
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1635444444
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_61
timestamp 1635444444
transform 1 0 6716 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1635444444
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  _0980_
timestamp 1635444444
transform 1 0 5336 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1971_
timestamp 1635444444
transform 1 0 6808 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_78
timestamp 1635444444
transform 1 0 8280 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1972_
timestamp 1635444444
transform 1 0 8648 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1635444444
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_98
timestamp 1635444444
transform 1 0 10120 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1062_
timestamp 1635444444
transform -1 0 11040 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_130
timestamp 1635444444
transform 1 0 13064 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1635444444
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1881_
timestamp 1635444444
transform 1 0 11500 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_55_150
timestamp 1635444444
transform 1 0 14904 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1635444444
transform 1 0 13432 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_55_154
timestamp 1635444444
transform 1 0 15272 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_158
timestamp 1635444444
transform 1 0 15640 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1635444444
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_169
timestamp 1635444444
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_173
timestamp 1635444444
transform 1 0 17020 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1635444444
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1635444444
transform 1 0 15364 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0924_
timestamp 1635444444
transform 1 0 17112 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_55_183
timestamp 1635444444
transform 1 0 17940 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1355_
timestamp 1635444444
transform 1 0 18492 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_55_198
timestamp 1635444444
transform 1 0 19320 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_4  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 21344 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1635444444
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_230
timestamp 1635444444
transform 1 0 22264 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1635444444
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1312_
timestamp 1635444444
transform -1 0 22264 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_55_242
timestamp 1635444444
transform 1 0 23368 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_254
timestamp 1635444444
transform 1 0 24472 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_266
timestamp 1635444444
transform 1 0 25576 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1635444444
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1635444444
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1635444444
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1635444444
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1635444444
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_317
timestamp 1635444444
transform 1 0 30268 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1635444444
transform -1 0 30820 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_15
timestamp 1635444444
transform 1 0 2484 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1635444444
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_7
timestamp 1635444444
transform 1 0 1748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1635444444
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1325_
timestamp 1635444444
transform 1 0 2852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1455_
timestamp 1635444444
transform 1 0 1840 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_56_22
timestamp 1635444444
transform 1 0 3128 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1635444444
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1635444444
transform 1 0 3772 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_45
timestamp 1635444444
transform 1 0 5244 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_53
timestamp 1635444444
transform 1 0 5980 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_61
timestamp 1635444444
transform 1 0 6716 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_65
timestamp 1635444444
transform 1 0 7084 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0956_
timestamp 1635444444
transform -1 0 7084 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1240_
timestamp 1635444444
transform -1 0 5980 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1635444444
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_85
timestamp 1635444444
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1635444444
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0959_
timestamp 1635444444
transform 1 0 7636 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_56_105
timestamp 1635444444
transform 1 0 10764 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1973_
timestamp 1635444444
transform 1 0 9292 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_56_120
timestamp 1635444444
transform 1 0 12144 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__o221ai_1  _1211_
timestamp 1635444444
transform -1 0 12144 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_56_132
timestamp 1635444444
transform 1 0 13248 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_56_141
timestamp 1635444444
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_149
timestamp 1635444444
transform 1 0 14812 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1635444444
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _1979_
timestamp 1635444444
transform 1 0 14996 0 1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_56_168
timestamp 1635444444
transform 1 0 16560 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1978_
timestamp 1635444444
transform 1 0 16928 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_56_188
timestamp 1635444444
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1635444444
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_206
timestamp 1635444444
transform 1 0 20056 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _1345_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 19228 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1767_
timestamp 1635444444
transform -1 0 21620 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_56_223
timestamp 1635444444
transform 1 0 21620 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_232
timestamp 1635444444
transform 1 0 22448 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_1  _0973_
timestamp 1635444444
transform -1 0 22448 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_56_244
timestamp 1635444444
transform 1 0 23552 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1635444444
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1635444444
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1635444444
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1635444444
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1635444444
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1635444444
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1635444444
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_309
timestamp 1635444444
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_317
timestamp 1635444444
transform 1 0 30268 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1635444444
transform -1 0 30820 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1635444444
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_14
timestamp 1635444444
transform 1 0 2392 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_7
timestamp 1635444444
transform 1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1635444444
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1322_
timestamp 1635444444
transform -1 0 3220 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1635444444
transform 1 0 2116 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1635444444
transform -1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_23
timestamp 1635444444
transform 1 0 3220 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_36
timestamp 1635444444
transform 1 0 4416 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1324_
timestamp 1635444444
transform -1 0 4416 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_57_44
timestamp 1635444444
transform 1 0 5152 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1635444444
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1635444444
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_60
timestamp 1635444444
transform 1 0 6624 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1635444444
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0944_
timestamp 1635444444
transform -1 0 6624 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1248_
timestamp 1635444444
transform -1 0 5612 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_68
timestamp 1635444444
transform 1 0 7360 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_79
timestamp 1635444444
transform 1 0 8372 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_86
timestamp 1635444444
transform 1 0 9016 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0952_
timestamp 1635444444
transform 1 0 8740 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0963_
timestamp 1635444444
transform -1 0 8372 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_107
timestamp 1635444444
transform 1 0 10948 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_93
timestamp 1635444444
transform 1 0 9660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0933_
timestamp 1635444444
transform 1 0 10028 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _0953_
timestamp 1635444444
transform -1 0 9660 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1635444444
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_123
timestamp 1635444444
transform 1 0 12420 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_127
timestamp 1635444444
transform 1 0 12788 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1635444444
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0950_
timestamp 1635444444
transform 1 0 11500 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_2  _1895_
timestamp 1635444444
transform 1 0 12880 0 -1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_57_145
timestamp 1635444444
transform 1 0 14444 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0917_
timestamp 1635444444
transform 1 0 14996 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_159
timestamp 1635444444
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1635444444
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1635444444
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_173
timestamp 1635444444
transform 1 0 17020 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1635444444
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1635444444
transform -1 0 17572 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_57_179
timestamp 1635444444
transform 1 0 17572 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_57_194
timestamp 1635444444
transform 1 0 18952 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _1745_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 18952 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_57_200
timestamp 1635444444
transform 1 0 19504 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_206
timestamp 1635444444
transform 1 0 20056 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1635444444
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0928_
timestamp 1635444444
transform 1 0 19596 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0930_
timestamp 1635444444
transform 1 0 20424 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1635444444
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_228
timestamp 1635444444
transform 1 0 22080 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_235
timestamp 1635444444
transform 1 0 22724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1635444444
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1635444444
transform 1 0 21804 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1362_
timestamp 1635444444
transform -1 0 22724 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_247
timestamp 1635444444
transform 1 0 23828 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_259
timestamp 1635444444
transform 1 0 24932 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_271
timestamp 1635444444
transform 1 0 26036 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1635444444
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1635444444
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1635444444
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1635444444
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_305
timestamp 1635444444
transform 1 0 29164 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_311
timestamp 1635444444
transform 1 0 29716 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_316
timestamp 1635444444
transform 1 0 30176 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1635444444
transform -1 0 30820 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1635444444
transform 1 0 29808 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_15
timestamp 1635444444
transform 1 0 2484 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1635444444
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_7
timestamp 1635444444
transform 1 0 1748 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1635444444
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1458_
timestamp 1635444444
transform 1 0 1840 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1635444444
transform -1 0 3220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_23
timestamp 1635444444
transform 1 0 3220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1635444444
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1635444444
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1635444444
transform 1 0 3772 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_58_45
timestamp 1635444444
transform 1 0 5244 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_53
timestamp 1635444444
transform 1 0 5980 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_57
timestamp 1635444444
transform 1 0 6348 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_64
timestamp 1635444444
transform 1 0 6992 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0906__1
timestamp 1635444444
transform -1 0 6992 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0907_
timestamp 1635444444
transform -1 0 6348 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_71
timestamp 1635444444
transform 1 0 7636 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_80
timestamp 1635444444
transform 1 0 8464 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1635444444
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1635444444
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1635444444
transform 1 0 8188 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0945_
timestamp 1635444444
transform 1 0 7360 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_89
timestamp 1635444444
transform 1 0 9292 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_99
timestamp 1635444444
transform 1 0 10212 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0955_
timestamp 1635444444
transform -1 0 10212 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1975_
timestamp 1635444444
transform 1 0 10580 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_119
timestamp 1635444444
transform 1 0 12052 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_131
timestamp 1635444444
transform 1 0 13156 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1183_
timestamp 1635444444
transform 1 0 12420 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1635444444
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_149
timestamp 1635444444
transform 1 0 14812 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1635444444
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1184_
timestamp 1635444444
transform -1 0 14812 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_155
timestamp 1635444444
transform 1 0 15364 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_159
timestamp 1635444444
transform 1 0 15732 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_166
timestamp 1635444444
transform 1 0 16376 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0918_
timestamp 1635444444
transform 1 0 15456 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0919_
timestamp 1635444444
transform 1 0 16100 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_178
timestamp 1635444444
transform 1 0 17480 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_185
timestamp 1635444444
transform 1 0 18124 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1635444444
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1635444444
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1344_
timestamp 1635444444
transform 1 0 18492 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1354_
timestamp 1635444444
transform 1 0 17848 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_197
timestamp 1635444444
transform 1 0 19228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_206
timestamp 1635444444
transform 1 0 20056 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_217
timestamp 1635444444
transform 1 0 21068 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1635444444
transform -1 0 20056 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1223_
timestamp 1635444444
transform 1 0 20424 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_58_223
timestamp 1635444444
transform 1 0 21620 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_227
timestamp 1635444444
transform 1 0 21988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_239
timestamp 1635444444
transform 1 0 23092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1361_
timestamp 1635444444
transform 1 0 21712 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1635444444
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1635444444
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1635444444
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1635444444
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1635444444
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1635444444
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1635444444
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1635444444
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_309
timestamp 1635444444
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_317
timestamp 1635444444
transform 1 0 30268 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1635444444
transform -1 0 30820 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1635444444
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1635444444
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1635444444
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_7
timestamp 1635444444
transform 1 0 1748 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_3
timestamp 1635444444
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_7
timestamp 1635444444
transform 1 0 1748 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1635444444
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1462_
timestamp 1635444444
transform -1 0 2484 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1460_
timestamp 1635444444
transform 1 0 1840 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_60_15
timestamp 1635444444
transform 1 0 2484 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_15
timestamp 1635444444
transform 1 0 2484 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1635444444
transform -1 0 3220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1323_
timestamp 1635444444
transform 1 0 2852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1321_
timestamp 1635444444
transform -1 0 4324 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1635444444
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_29
timestamp 1635444444
transform 1 0 3772 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1635444444
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_23
timestamp 1635444444
transform 1 0 3220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_22
timestamp 1635444444
transform 1 0 3128 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1317_
timestamp 1635444444
transform -1 0 5520 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1310_
timestamp 1635444444
transform 1 0 4232 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_37
timestamp 1635444444
transform 1 0 4508 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_33
timestamp 1635444444
transform 1 0 4140 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_35
timestamp 1635444444
transform 1 0 4324 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1635444444
transform 1 0 4876 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_59_48
timestamp 1635444444
transform 1 0 5520 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_63
timestamp 1635444444
transform 1 0 6900 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_57
timestamp 1635444444
transform 1 0 6348 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_63
timestamp 1635444444
transform 1 0 6900 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1635444444
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _1382_
timestamp 1635444444
transform 1 0 6348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1970_
timestamp 1635444444
transform -1 0 8464 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_59_69
timestamp 1635444444
transform 1 0 7452 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_79
timestamp 1635444444
transform 1 0 8372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1635444444
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1635444444
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0932_
timestamp 1635444444
transform 1 0 8924 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _0967_
timestamp 1635444444
transform -1 0 8372 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1974_
timestamp 1635444444
transform 1 0 8924 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1635444444
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_95
timestamp 1635444444
transform 1 0 9844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_101
timestamp 1635444444
transform 1 0 10396 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_108
timestamp 1635444444
transform 1 0 11040 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0940_
timestamp 1635444444
transform -1 0 11040 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0943_
timestamp 1635444444
transform 1 0 10212 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_59_117
timestamp 1635444444
transform 1 0 11868 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_121
timestamp 1635444444
transform 1 0 12236 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_114
timestamp 1635444444
transform 1 0 11592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1635444444
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0904_
timestamp 1635444444
transform -1 0 11868 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1882_
timestamp 1635444444
transform 1 0 11684 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1894_
timestamp 1635444444
transform 1 0 12328 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_59_139
timestamp 1635444444
transform 1 0 13892 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_132
timestamp 1635444444
transform 1 0 13248 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1635444444
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_145
timestamp 1635444444
transform 1 0 14444 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1635444444
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1829_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 14536 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1830_
timestamp 1635444444
transform 1 0 14260 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1635444444
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_169
timestamp 1635444444
transform 1 0 16652 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_167
timestamp 1635444444
transform 1 0 16468 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1635444444
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1811_
timestamp 1635444444
transform 1 0 16928 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_59_181
timestamp 1635444444
transform 1 0 17756 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_188
timestamp 1635444444
transform 1 0 18400 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_192
timestamp 1635444444
transform 1 0 18768 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_175
timestamp 1635444444
transform 1 0 17204 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1635444444
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1635444444
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _1346_
timestamp 1635444444
transform 1 0 18860 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1347_
timestamp 1635444444
transform -1 0 18400 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1635444444
transform 1 0 17296 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_59_201
timestamp 1635444444
transform 1 0 19596 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_210
timestamp 1635444444
transform 1 0 20424 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp 1635444444
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_201
timestamp 1635444444
transform 1 0 19596 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_211
timestamp 1635444444
transform 1 0 20516 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1635444444
transform 1 0 20148 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1523_
timestamp 1635444444
transform -1 0 21436 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1762_
timestamp 1635444444
transform 1 0 19688 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1635444444
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1635444444
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1635444444
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1635444444
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1635444444
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1635444444
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1635444444
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1635444444
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1635444444
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1635444444
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1635444444
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1635444444
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1635444444
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1635444444
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1635444444
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1635444444
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1635444444
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1635444444
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1635444444
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_305
timestamp 1635444444
transform 1 0 29164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1635444444
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1635444444
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_316
timestamp 1635444444
transform 1 0 30176 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1635444444
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_309
timestamp 1635444444
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_317
timestamp 1635444444
transform 1 0 30268 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1635444444
transform -1 0 30820 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1635444444
transform -1 0 30820 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1635444444
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1635444444
transform -1 0 30176 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_61_15
timestamp 1635444444
transform 1 0 2484 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_21
timestamp 1635444444
transform 1 0 3036 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1635444444
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_7
timestamp 1635444444
transform 1 0 1748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1635444444
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1464_
timestamp 1635444444
transform 1 0 1840 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_61_38
timestamp 1635444444
transform 1 0 4600 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1311_
timestamp 1635444444
transform -1 0 5244 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1635444444
transform 1 0 3128 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_61_45
timestamp 1635444444
transform 1 0 5244 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_52
timestamp 1635444444
transform 1 0 5888 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_57
timestamp 1635444444
transform 1 0 6348 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_61
timestamp 1635444444
transform 1 0 6716 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_65
timestamp 1635444444
transform 1 0 7084 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1635444444
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0964_
timestamp 1635444444
transform 1 0 6808 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1328_
timestamp 1635444444
transform -1 0 5888 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_73
timestamp 1635444444
transform 1 0 7820 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_78
timestamp 1635444444
transform 1 0 8280 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_86
timestamp 1635444444
transform 1 0 9016 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0946_
timestamp 1635444444
transform 1 0 8004 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_106
timestamp 1635444444
transform 1 0 10856 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_97
timestamp 1635444444
transform 1 0 10028 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0941_
timestamp 1635444444
transform -1 0 10856 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0951_
timestamp 1635444444
transform -1 0 10028 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_61_116
timestamp 1635444444
transform 1 0 11776 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_128
timestamp 1635444444
transform 1 0 12880 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1635444444
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1342_
timestamp 1635444444
transform 1 0 11500 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_140
timestamp 1635444444
transform 1 0 13984 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_152
timestamp 1635444444
transform 1 0 15088 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1635444444
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1635444444
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1817_
timestamp 1635444444
transform -1 0 17480 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_61_178
timestamp 1635444444
transform 1 0 17480 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_187
timestamp 1635444444
transform 1 0 18308 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_193
timestamp 1635444444
transform 1 0 18860 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _1350_
timestamp 1635444444
transform 1 0 18952 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1576_
timestamp 1635444444
transform 1 0 17848 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_61_202
timestamp 1635444444
transform 1 0 19688 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_209
timestamp 1635444444
transform 1 0 20332 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0921_
timestamp 1635444444
transform 1 0 20700 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1222_
timestamp 1635444444
transform -1 0 20332 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_219
timestamp 1635444444
transform 1 0 21252 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1635444444
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1635444444
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1635444444
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1635444444
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1635444444
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1635444444
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1635444444
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1635444444
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1635444444
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1635444444
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1635444444
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1635444444
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_317
timestamp 1635444444
transform 1 0 30268 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1635444444
transform -1 0 30820 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_14
timestamp 1635444444
transform 1 0 2392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1635444444
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_7
timestamp 1635444444
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1635444444
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1319_
timestamp 1635444444
transform 1 0 2760 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1454_
timestamp 1635444444
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1635444444
transform -1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1635444444
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_32
timestamp 1635444444
transform 1 0 4048 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_36
timestamp 1635444444
transform 1 0 4416 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_40
timestamp 1635444444
transform 1 0 4784 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1635444444
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1318_
timestamp 1635444444
transform -1 0 4048 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1341_
timestamp 1635444444
transform 1 0 4508 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_47
timestamp 1635444444
transform 1 0 5428 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_61
timestamp 1635444444
transform 1 0 6716 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1249_
timestamp 1635444444
transform -1 0 5428 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1381_
timestamp 1635444444
transform -1 0 6716 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _1435_
timestamp 1635444444
transform 1 0 7084 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_71
timestamp 1635444444
transform 1 0 7636 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_78
timestamp 1635444444
transform 1 0 8280 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1635444444
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0947_
timestamp 1635444444
transform -1 0 9200 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0965_
timestamp 1635444444
transform 1 0 8004 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_109
timestamp 1635444444
transform 1 0 11132 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_88
timestamp 1635444444
transform 1 0 9200 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_95
timestamp 1635444444
transform 1 0 9844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_99
timestamp 1635444444
transform 1 0 10212 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0939_
timestamp 1635444444
transform 1 0 10304 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1004_
timestamp 1635444444
transform 1 0 9568 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_116
timestamp 1635444444
transform 1 0 11776 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_128
timestamp 1635444444
transform 1 0 12880 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1465_
timestamp 1635444444
transform 1 0 11500 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_144
timestamp 1635444444
transform 1 0 14352 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1635444444
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1595_
timestamp 1635444444
transform 1 0 14076 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1824_
timestamp 1635444444
transform 1 0 14904 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_62_171
timestamp 1635444444
transform 1 0 16836 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_175
timestamp 1635444444
transform 1 0 17204 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_179
timestamp 1635444444
transform 1 0 17572 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_187
timestamp 1635444444
transform 1 0 18308 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_191
timestamp 1635444444
transform 1 0 18676 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1635444444
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1635444444
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1351_
timestamp 1635444444
transform -1 0 18676 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1577_
timestamp 1635444444
transform 1 0 17296 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_197
timestamp 1635444444
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_205
timestamp 1635444444
transform 1 0 19964 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_212
timestamp 1635444444
transform 1 0 20608 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_216
timestamp 1635444444
transform 1 0 20976 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0948_
timestamp 1635444444
transform 1 0 21068 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1522_
timestamp 1635444444
transform -1 0 20608 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_227
timestamp 1635444444
transform 1 0 21988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_239
timestamp 1635444444
transform 1 0 23092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1635444444
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1635444444
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1635444444
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1635444444
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1635444444
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1635444444
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1635444444
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1635444444
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_309
timestamp 1635444444
transform 1 0 29532 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_317
timestamp 1635444444
transform 1 0 30268 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1635444444
transform -1 0 30820 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1635444444
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_15
timestamp 1635444444
transform 1 0 2484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_7
timestamp 1635444444
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1635444444
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0992_
timestamp 1635444444
transform 1 0 2852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1635444444
transform -1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1635444444
transform 1 0 2116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_22
timestamp 1635444444
transform 1 0 3128 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_29
timestamp 1635444444
transform 1 0 3772 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_36
timestamp 1635444444
transform 1 0 4416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_43
timestamp 1635444444
transform 1 0 5060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0993_
timestamp 1635444444
transform 1 0 3496 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1250_
timestamp 1635444444
transform 1 0 4784 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1635444444
transform 1 0 4140 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_50
timestamp 1635444444
transform 1 0 5704 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1635444444
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1635444444
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0968_
timestamp 1635444444
transform -1 0 5704 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1434_
timestamp 1635444444
transform 1 0 6532 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_63_69
timestamp 1635444444
transform 1 0 7452 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_86
timestamp 1635444444
transform 1 0 9016 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1005_
timestamp 1635444444
transform 1 0 8188 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_63_108
timestamp 1635444444
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_95
timestamp 1635444444
transform 1 0 9844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0908_
timestamp 1635444444
transform 1 0 9568 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0935_
timestamp 1635444444
transform 1 0 10212 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_63_129
timestamp 1635444444
transform 1 0 12972 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1635444444
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1977_
timestamp 1635444444
transform 1 0 11500 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_63_136
timestamp 1635444444
transform 1 0 13616 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_149
timestamp 1635444444
transform 1 0 14812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1210_
timestamp 1635444444
transform 1 0 13340 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 14812 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_63_160
timestamp 1635444444
transform 1 0 15824 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_169
timestamp 1635444444
transform 1 0 16652 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1635444444
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1594_
timestamp 1635444444
transform -1 0 15824 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1768_
timestamp 1635444444
transform -1 0 17572 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_63_179
timestamp 1635444444
transform 1 0 17572 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1635444444
transform 1 0 18308 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_63_203
timestamp 1635444444
transform 1 0 19780 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_216
timestamp 1635444444
transform 1 0 20976 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1761_
timestamp 1635444444
transform 1 0 20148 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_63_231
timestamp 1635444444
transform 1 0 22356 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1635444444
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0966_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 22356 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_243
timestamp 1635444444
transform 1 0 23460 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_255
timestamp 1635444444
transform 1 0 24564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_267
timestamp 1635444444
transform 1 0 25668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1635444444
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1635444444
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1635444444
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1635444444
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_305
timestamp 1635444444
transform 1 0 29164 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_316
timestamp 1635444444
transform 1 0 30176 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1635444444
transform -1 0 30820 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1635444444
transform 1 0 29900 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1635444444
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1635444444
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1635444444
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1635444444
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1467_
timestamp 1635444444
transform 1 0 1840 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1635444444
transform 1 0 2852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1635444444
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1635444444
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_32
timestamp 1635444444
transform 1 0 4048 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_39
timestamp 1635444444
transform 1 0 4692 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1635444444
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0989_
timestamp 1635444444
transform -1 0 4048 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1459_
timestamp 1635444444
transform 1 0 4416 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_47
timestamp 1635444444
transform 1 0 5428 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_64
timestamp 1635444444
transform 1 0 6992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1635444444
transform 1 0 5520 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_64_74
timestamp 1635444444
transform 1 0 7912 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1635444444
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1635444444
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _1440_
timestamp 1635444444
transform 1 0 7360 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1962_
timestamp 1635444444
transform -1 0 10396 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_101
timestamp 1635444444
transform 1 0 10396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_105
timestamp 1635444444
transform 1 0 10764 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1976_
timestamp 1635444444
transform 1 0 10856 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_64_122
timestamp 1635444444
transform 1 0 12328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_130
timestamp 1635444444
transform 1 0 13064 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1612_
timestamp 1635444444
transform 1 0 12696 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1635444444
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_144
timestamp 1635444444
transform 1 0 14352 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1635444444
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1571_
timestamp 1635444444
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1823_
timestamp 1635444444
transform 1 0 14904 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_64_171
timestamp 1635444444
transform 1 0 16836 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1635444444
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1635444444
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1763_
timestamp 1635444444
transform -1 0 18400 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_64_200
timestamp 1635444444
transform 1 0 19504 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_211
timestamp 1635444444
transform 1 0 20516 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1221_
timestamp 1635444444
transform -1 0 20516 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1349_
timestamp 1635444444
transform -1 0 19504 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_223
timestamp 1635444444
transform 1 0 21620 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_235
timestamp 1635444444
transform 1 0 22724 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1635444444
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1635444444
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1635444444
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1635444444
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1635444444
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1635444444
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1635444444
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1635444444
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1635444444
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 1635444444
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_317
timestamp 1635444444
transform 1 0 30268 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1635444444
transform -1 0 30820 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1635444444
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_16
timestamp 1635444444
transform 1 0 2576 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_20
timestamp 1635444444
transform 1 0 2944 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_3
timestamp 1635444444
transform 1 0 1380 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1635444444
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1472_
timestamp 1635444444
transform -1 0 2576 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1965_
timestamp 1635444444
transform -1 0 4508 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_37
timestamp 1635444444
transform 1 0 4508 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_41
timestamp 1635444444
transform 1 0 4876 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0978_
timestamp 1635444444
transform -1 0 5888 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_65_52
timestamp 1635444444
transform 1 0 5888 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1635444444
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0981_
timestamp 1635444444
transform 1 0 6348 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_65_67
timestamp 1635444444
transform 1 0 7268 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_78
timestamp 1635444444
transform 1 0 8280 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1002_
timestamp 1635444444
transform 1 0 8648 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1003_
timestamp 1635444444
transform 1 0 8004 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_106
timestamp 1635444444
transform 1 0 10856 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_91
timestamp 1635444444
transform 1 0 9476 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_95
timestamp 1635444444
transform 1 0 9844 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_99
timestamp 1635444444
transform 1 0 10212 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0925_
timestamp 1635444444
transform 1 0 10580 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0937_
timestamp 1635444444
transform 1 0 9936 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_116
timestamp 1635444444
transform 1 0 11776 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_124
timestamp 1635444444
transform 1 0 12512 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_131
timestamp 1635444444
transform 1 0 13156 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1635444444
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0926_
timestamp 1635444444
transform -1 0 11776 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1610_
timestamp 1635444444
transform -1 0 13156 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_65_137
timestamp 1635444444
transform 1 0 13708 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_144
timestamp 1635444444
transform 1 0 14352 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_151
timestamp 1635444444
transform 1 0 14996 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1593_
timestamp 1635444444
transform -1 0 14996 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1596_
timestamp 1635444444
transform 1 0 13800 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_163
timestamp 1635444444
transform 1 0 16100 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1635444444
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1635444444
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_174
timestamp 1635444444
transform 1 0 17112 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1635444444
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1598_
timestamp 1635444444
transform -1 0 17112 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_183
timestamp 1635444444
transform 1 0 17940 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_190
timestamp 1635444444
transform 1 0 18584 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1348_
timestamp 1635444444
transform 1 0 18308 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1597_
timestamp 1635444444
transform -1 0 17940 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _1835_
timestamp 1635444444
transform 1 0 18952 0 -1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_65_211
timestamp 1635444444
transform 1 0 20516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1635444444
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_231
timestamp 1635444444
transform 1 0 22356 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1635444444
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0962_
timestamp 1635444444
transform -1 0 22356 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_243
timestamp 1635444444
transform 1 0 23460 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_255
timestamp 1635444444
transform 1 0 24564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_267
timestamp 1635444444
transform 1 0 25668 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1635444444
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1635444444
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1635444444
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1635444444
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1635444444
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_317
timestamp 1635444444
transform 1 0 30268 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1635444444
transform -1 0 30820 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1474_
timestamp 1635444444
transform 1 0 1840 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1470_
timestamp 1635444444
transform 1 0 1472 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1635444444
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1635444444
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_67_7
timestamp 1635444444
transform 1 0 1748 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_3
timestamp 1635444444
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_3
timestamp 1635444444
transform 1 0 1380 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1635444444
transform 1 0 2852 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0994_
timestamp 1635444444
transform -1 0 3312 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_67_15
timestamp 1635444444
transform 1 0 2484 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_11
timestamp 1635444444
transform 1 0 2116 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1635444444
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_29
timestamp 1635444444
transform 1 0 3772 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_23
timestamp 1635444444
transform 1 0 3220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_29
timestamp 1635444444
transform 1 0 3772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_39
timestamp 1635444444
transform 1 0 4692 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1635444444
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0991_
timestamp 1635444444
transform -1 0 4692 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1966_
timestamp 1635444444
transform 1 0 3956 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1635444444
transform -1 0 5888 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0976_
timestamp 1635444444
transform 1 0 5796 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_67_52
timestamp 1635444444
transform 1 0 5888 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_47
timestamp 1635444444
transform 1 0 5428 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_47
timestamp 1635444444
transform 1 0 5428 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1251_
timestamp 1635444444
transform -1 0 7912 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1635444444
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_61
timestamp 1635444444
transform 1 0 6716 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_57
timestamp 1635444444
transform 1 0 6348 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_61
timestamp 1635444444
transform 1 0 6716 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1635444444
transform 1 0 6808 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_66_74
timestamp 1635444444
transform 1 0 7912 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1635444444
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_78
timestamp 1635444444
transform 1 0 8280 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_86
timestamp 1635444444
transform 1 0 9016 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1635444444
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0999_
timestamp 1635444444
transform 1 0 8924 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_66_102
timestamp 1635444444
transform 1 0 10488 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_107
timestamp 1635444444
transform 1 0 10948 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_94
timestamp 1635444444
transform 1 0 9752 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_104
timestamp 1635444444
transform 1 0 10672 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0936_
timestamp 1635444444
transform -1 0 10948 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1963_
timestamp 1635444444
transform 1 0 9200 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_66_119
timestamp 1635444444
transform 1 0 12052 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_125
timestamp 1635444444
transform 1 0 12604 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1635444444
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_125
timestamp 1635444444
transform 1 0 12604 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_129
timestamp 1635444444
transform 1 0 12972 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1635444444
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1611_
timestamp 1635444444
transform -1 0 12604 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1613_
timestamp 1635444444
transform 1 0 12972 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_2  _1617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 13892 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_66_134
timestamp 1635444444
transform 1 0 13432 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_144
timestamp 1635444444
transform 1 0 14352 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_139
timestamp 1635444444
transform 1 0 13892 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1635444444
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1614_
timestamp 1635444444
transform -1 0 14352 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1827_
timestamp 1635444444
transform 1 0 14260 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_12  FILLER_66_156
timestamp 1635444444
transform 1 0 15456 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_168
timestamp 1635444444
transform 1 0 16560 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_164
timestamp 1635444444
transform 1 0 16192 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1635444444
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1635444444
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_180
timestamp 1635444444
transform 1 0 17664 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_191
timestamp 1635444444
transform 1 0 18676 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1635444444
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_181
timestamp 1635444444
transform 1 0 17756 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_189
timestamp 1635444444
transform 1 0 18492 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1635444444
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0998_
timestamp 1635444444
transform -1 0 17664 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1352_
timestamp 1635444444
transform 1 0 18400 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1782_
timestamp 1635444444
transform -1 0 19596 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_200
timestamp 1635444444
transform 1 0 19504 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_212
timestamp 1635444444
transform 1 0 20608 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_201
timestamp 1635444444
transform 1 0 19596 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_205
timestamp 1635444444
transform 1 0 19964 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_209
timestamp 1635444444
transform 1 0 20332 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1353_
timestamp 1635444444
transform -1 0 19504 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1635444444
transform -1 0 20332 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_224
timestamp 1635444444
transform 1 0 21712 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_236
timestamp 1635444444
transform 1 0 22816 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_221
timestamp 1635444444
transform 1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1635444444
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1635444444
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1635444444
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_248
timestamp 1635444444
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1635444444
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1635444444
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1635444444
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1635444444
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1635444444
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1635444444
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1635444444
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1635444444
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1635444444
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1635444444
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1635444444
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1635444444
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1635444444
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1635444444
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1635444444
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_309
timestamp 1635444444
transform 1 0 29532 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_316
timestamp 1635444444
transform 1 0 30176 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_317
timestamp 1635444444
transform 1 0 30268 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1635444444
transform -1 0 30820 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1635444444
transform -1 0 30820 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1635444444
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1635444444
transform 1 0 29900 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_15
timestamp 1635444444
transform 1 0 2484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_7
timestamp 1635444444
transform 1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1635444444
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0987_
timestamp 1635444444
transform -1 0 3128 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1635444444
transform -1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1635444444
transform -1 0 2484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_22
timestamp 1635444444
transform 1 0 3128 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_32
timestamp 1635444444
transform 1 0 4048 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_36
timestamp 1635444444
transform 1 0 4416 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_40
timestamp 1635444444
transform 1 0 4784 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1635444444
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0990_
timestamp 1635444444
transform 1 0 3772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1246_
timestamp 1635444444
transform 1 0 4508 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_47
timestamp 1635444444
transform 1 0 5428 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_54
timestamp 1635444444
transform 1 0 6072 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1231_
timestamp 1635444444
transform -1 0 6072 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1245_
timestamp 1635444444
transform -1 0 5428 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1247_
timestamp 1635444444
transform 1 0 6440 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_68_67
timestamp 1635444444
transform 1 0 7268 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_75
timestamp 1635444444
transform 1 0 8004 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_80
timestamp 1635444444
transform 1 0 8464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_85
timestamp 1635444444
transform 1 0 8924 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1635444444
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0995_
timestamp 1635444444
transform -1 0 8464 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_106
timestamp 1635444444
transform 1 0 10856 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_89
timestamp 1635444444
transform 1 0 9292 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1964_
timestamp 1635444444
transform 1 0 9384 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_68_118
timestamp 1635444444
transform 1 0 11960 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_124
timestamp 1635444444
transform 1 0 12512 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_130
timestamp 1635444444
transform 1 0 13064 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1615_
timestamp 1635444444
transform 1 0 12604 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_68_138
timestamp 1635444444
transform 1 0 13800 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_141
timestamp 1635444444
transform 1 0 14076 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1635444444
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1826_
timestamp 1635444444
transform 1 0 14628 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_68_168
timestamp 1635444444
transform 1 0 16560 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1784_
timestamp 1635444444
transform -1 0 17756 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_68_181
timestamp 1635444444
transform 1 0 17756 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_190
timestamp 1635444444
transform 1 0 18584 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1635444444
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1554_
timestamp 1635444444
transform 1 0 18124 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_68_200
timestamp 1635444444
transform 1 0 19504 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_213
timestamp 1635444444
transform 1 0 20700 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1619_
timestamp 1635444444
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1741_
timestamp 1635444444
transform -1 0 20700 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_68_227
timestamp 1635444444
transform 1 0 21988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_239
timestamp 1635444444
transform 1 0 23092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _0958_
timestamp 1635444444
transform -1 0 21988 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1635444444
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1635444444
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1635444444
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1635444444
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1635444444
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1635444444
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1635444444
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1635444444
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_309
timestamp 1635444444
transform 1 0 29532 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_316
timestamp 1635444444
transform 1 0 30176 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1635444444
transform -1 0 30820 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1635444444
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1635444444
transform 1 0 29900 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_15
timestamp 1635444444
transform 1 0 2484 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_3
timestamp 1635444444
transform 1 0 1380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_7
timestamp 1635444444
transform 1 0 1748 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1635444444
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1476_
timestamp 1635444444
transform 1 0 1840 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1967_
timestamp 1635444444
transform 1 0 2852 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_69_35
timestamp 1635444444
transform 1 0 4324 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_43
timestamp 1635444444
transform 1 0 5060 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_52
timestamp 1635444444
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_57
timestamp 1635444444
transform 1 0 6348 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_61
timestamp 1635444444
transform 1 0 6716 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_65
timestamp 1635444444
transform 1 0 7084 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1635444444
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1635444444
transform 1 0 6808 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1484_
timestamp 1635444444
transform -1 0 5888 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_69_72
timestamp 1635444444
transform 1 0 7728 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_78
timestamp 1635444444
transform 1 0 8280 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_82
timestamp 1635444444
transform 1 0 8648 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0996_
timestamp 1635444444
transform 1 0 9016 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1000_
timestamp 1635444444
transform 1 0 8372 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1243_
timestamp 1635444444
transform 1 0 7452 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_108
timestamp 1635444444
transform 1 0 11040 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_89
timestamp 1635444444
transform 1 0 9292 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_96
timestamp 1635444444
transform 1 0 9936 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0997_
timestamp 1635444444
transform -1 0 9936 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1635444444
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_125
timestamp 1635444444
transform 1 0 12604 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1635444444
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1821_
timestamp 1635444444
transform 1 0 12788 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_69_148
timestamp 1635444444
transform 1 0 14720 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_156
timestamp 1635444444
transform 1 0 15456 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_162
timestamp 1635444444
transform 1 0 16008 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_172
timestamp 1635444444
transform 1 0 16928 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1635444444
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1548_
timestamp 1635444444
transform 1 0 15548 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1552_
timestamp 1635444444
transform -1 0 16928 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_187
timestamp 1635444444
transform 1 0 18308 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_196
timestamp 1635444444
transform 1 0 19136 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1618_
timestamp 1635444444
transform 1 0 18676 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1785_
timestamp 1635444444
transform 1 0 17480 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_69_202
timestamp 1635444444
transform 1 0 19688 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_208
timestamp 1635444444
transform 1 0 20240 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1633_
timestamp 1635444444
transform 1 0 19780 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1635444444
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1635444444
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1635444444
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1635444444
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1635444444
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1635444444
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1635444444
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1635444444
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1635444444
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1635444444
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1635444444
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1635444444
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_317
timestamp 1635444444
transform 1 0 30268 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1635444444
transform -1 0 30820 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_15
timestamp 1635444444
transform 1 0 2484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 1635444444
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_70_7
timestamp 1635444444
transform 1 0 1748 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1635444444
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0986_
timestamp 1635444444
transform 1 0 2576 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1635444444
transform -1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1635444444
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_38
timestamp 1635444444
transform 1 0 4600 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1635444444
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0988_
timestamp 1635444444
transform -1 0 4600 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1466_
timestamp 1635444444
transform 1 0 4968 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_70_45
timestamp 1635444444
transform 1 0 5244 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_51
timestamp 1635444444
transform 1 0 5796 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_61
timestamp 1635444444
transform 1 0 6716 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1225_
timestamp 1635444444
transform 1 0 7084 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1244_
timestamp 1635444444
transform 1 0 5888 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_70_75
timestamp 1635444444
transform 1 0 8004 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1635444444
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1635444444
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1001_
timestamp 1635444444
transform 1 0 8924 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_107
timestamp 1635444444
transform 1 0 10948 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_88
timestamp 1635444444
transform 1 0 9200 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_95
timestamp 1635444444
transform 1 0 9844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1481_
timestamp 1635444444
transform 1 0 9568 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_119
timestamp 1635444444
transform 1 0 12052 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_125
timestamp 1635444444
transform 1 0 12604 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1616_
timestamp 1635444444
transform -1 0 13248 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1631_
timestamp 1635444444
transform -1 0 12604 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_132
timestamp 1635444444
transform 1 0 13248 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_141
timestamp 1635444444
transform 1 0 14076 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1635444444
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _1740_
timestamp 1635444444
transform -1 0 15272 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_70_154
timestamp 1635444444
transform 1 0 15272 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_162
timestamp 1635444444
transform 1 0 16008 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1825_
timestamp 1635444444
transform 1 0 16100 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_70_184
timestamp 1635444444
transform 1 0 18032 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_191
timestamp 1635444444
transform 1 0 18676 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1635444444
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1635444444
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1635444444
transform 1 0 18400 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1635444444
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1635444444
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1635444444
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1635444444
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1635444444
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1635444444
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1635444444
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1635444444
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1635444444
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1635444444
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1635444444
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1635444444
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1635444444
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_309
timestamp 1635444444
transform 1 0 29532 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_317
timestamp 1635444444
transform 1 0 30268 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1635444444
transform -1 0 30820 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1635444444
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_13
timestamp 1635444444
transform 1 0 2300 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_21
timestamp 1635444444
transform 1 0 3036 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_7
timestamp 1635444444
transform 1 0 1748 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1635444444
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1479_
timestamp 1635444444
transform -1 0 3036 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1635444444
transform -1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_34
timestamp 1635444444
transform 1 0 4232 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_41
timestamp 1635444444
transform 1 0 4876 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0985_
timestamp 1635444444
transform -1 0 4232 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1242_
timestamp 1635444444
transform 1 0 4600 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_52
timestamp 1635444444
transform 1 0 5888 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_57
timestamp 1635444444
transform 1 0 6348 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1635444444
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _1486_
timestamp 1635444444
transform -1 0 5888 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1635444444
transform -1 0 8004 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_75
timestamp 1635444444
transform 1 0 8004 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1226_
timestamp 1635444444
transform 1 0 8372 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_71_101
timestamp 1635444444
transform 1 0 10396 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_109
timestamp 1635444444
transform 1 0 11132 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_89
timestamp 1635444444
transform 1 0 9292 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1635444444
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1635444444
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__mux4_1  _1822_
timestamp 1635444444
transform 1 0 12604 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_71_146
timestamp 1635444444
transform 1 0 14536 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_150
timestamp 1635444444
transform 1 0 14904 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1547_
timestamp 1635444444
transform 1 0 14996 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_154
timestamp 1635444444
transform 1 0 15272 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_163
timestamp 1635444444
transform 1 0 16100 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1635444444
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_173
timestamp 1635444444
transform 1 0 17020 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1635444444
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _1550_
timestamp 1635444444
transform 1 0 16652 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1551_
timestamp 1635444444
transform 1 0 15640 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1635444444
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1635444444
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _1553_
timestamp 1635444444
transform 1 0 17388 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1635444444
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1635444444
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1635444444
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_231
timestamp 1635444444
transform 1 0 22356 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1635444444
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0954_
timestamp 1635444444
transform -1 0 22356 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_243
timestamp 1635444444
transform 1 0 23460 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_255
timestamp 1635444444
transform 1 0 24564 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_267
timestamp 1635444444
transform 1 0 25668 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1635444444
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1635444444
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1635444444
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1635444444
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_305
timestamp 1635444444
transform 1 0 29164 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_316
timestamp 1635444444
transform 1 0 30176 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1635444444
transform -1 0 30820 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1635444444
transform 1 0 29900 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1635444444
transform -1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1635444444
transform 1 0 1656 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1635444444
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1635444444
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_7
timestamp 1635444444
transform 1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_9
timestamp 1635444444
transform 1 0 1932 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_3
timestamp 1635444444
transform 1 0 1380 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1468_
timestamp 1635444444
transform 1 0 2116 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0983_
timestamp 1635444444
transform -1 0 3128 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_14
timestamp 1635444444
transform 1 0 2392 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_17
timestamp 1635444444
transform 1 0 2668 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1968_
timestamp 1635444444
transform 1 0 2760 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_72_22
timestamp 1635444444
transform 1 0 3128 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_32
timestamp 1635444444
transform 1 0 4048 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_34
timestamp 1635444444
transform 1 0 4232 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_41
timestamp 1635444444
transform 1 0 4876 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1635444444
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0982_
timestamp 1635444444
transform -1 0 5244 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1469_
timestamp 1635444444
transform 1 0 3772 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1477_
timestamp 1635444444
transform 1 0 4600 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1488_
timestamp 1635444444
transform -1 0 5888 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1482_
timestamp 1635444444
transform -1 0 6256 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_73_52
timestamp 1635444444
transform 1 0 5888 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_45
timestamp 1635444444
transform 1 0 5244 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1238_
timestamp 1635444444
transform 1 0 6716 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1236_
timestamp 1635444444
transform -1 0 6992 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1635444444
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_57
timestamp 1635444444
transform 1 0 6348 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_60
timestamp 1635444444
transform 1 0 6624 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_56
timestamp 1635444444
transform 1 0 6256 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_64
timestamp 1635444444
transform 1 0 6992 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_64
timestamp 1635444444
transform 1 0 6992 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1635444444
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1635444444
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_72
timestamp 1635444444
transform 1 0 7728 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1635444444
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1239_
timestamp 1635444444
transform 1 0 8924 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1241_
timestamp 1635444444
transform 1 0 7360 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1635444444
transform -1 0 9384 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_100
timestamp 1635444444
transform 1 0 10304 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_88
timestamp 1635444444
transform 1 0 9200 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_102
timestamp 1635444444
transform 1 0 10488 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_90
timestamp 1635444444
transform 1 0 9384 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_112
timestamp 1635444444
transform 1 0 11408 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_124
timestamp 1635444444
transform 1 0 12512 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_130
timestamp 1635444444
transform 1 0 13064 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1635444444
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1635444444
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1635444444
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1635444444
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1632_
timestamp 1635444444
transform 1 0 12788 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_138
timestamp 1635444444
transform 1 0 13800 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1635444444
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1635444444
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1635444444
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1635444444
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_153
timestamp 1635444444
transform 1 0 15180 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_164
timestamp 1635444444
transform 1 0 16192 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1635444444
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1635444444
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1635444444
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1635444444
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1549_
timestamp 1635444444
transform -1 0 16192 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_176
timestamp 1635444444
transform 1 0 17296 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_188
timestamp 1635444444
transform 1 0 18400 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1635444444
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1635444444
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1635444444
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1635444444
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_209
timestamp 1635444444
transform 1 0 20332 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_217
timestamp 1635444444
transform 1 0 21068 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1635444444
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1635444444
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_227
timestamp 1635444444
transform 1 0 21988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_239
timestamp 1635444444
transform 1 0 23092 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1635444444
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1635444444
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1635444444
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1635444444
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0949_
timestamp 1635444444
transform -1 0 21988 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1635444444
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1635444444
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1635444444
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1635444444
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1635444444
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1635444444
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1635444444
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1635444444
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1635444444
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1635444444
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1635444444
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1635444444
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1635444444
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1635444444
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1635444444
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1635444444
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_309
timestamp 1635444444
transform 1 0 29532 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_317
timestamp 1635444444
transform 1 0 30268 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_73_317
timestamp 1635444444
transform 1 0 30268 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1635444444
transform -1 0 30820 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1635444444
transform -1 0 30820 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1635444444
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_14
timestamp 1635444444
transform 1 0 2392 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_20
timestamp 1635444444
transform 1 0 2944 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_7
timestamp 1635444444
transform 1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1635444444
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0970_
timestamp 1635444444
transform 1 0 3036 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1471_
timestamp 1635444444
transform -1 0 2392 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1635444444
transform -1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_24
timestamp 1635444444
transform 1 0 3312 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_29
timestamp 1635444444
transform 1 0 3772 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1635444444
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1635444444
transform 1 0 4140 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_74_49
timestamp 1635444444
transform 1 0 5612 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_60
timestamp 1635444444
transform 1 0 6624 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1237_
timestamp 1635444444
transform -1 0 7820 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1491_
timestamp 1635444444
transform -1 0 6624 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_74_73
timestamp 1635444444
transform 1 0 7820 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_80
timestamp 1635444444
transform 1 0 8464 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1635444444
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1219_
timestamp 1635444444
transform 1 0 8924 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1228_
timestamp 1635444444
transform 1 0 8188 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_100
timestamp 1635444444
transform 1 0 10304 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_88
timestamp 1635444444
transform 1 0 9200 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_112
timestamp 1635444444
transform 1 0 11408 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_124
timestamp 1635444444
transform 1 0 12512 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_136
timestamp 1635444444
transform 1 0 13616 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1635444444
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1635444444
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1635444444
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1635444444
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1635444444
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1635444444
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1635444444
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1635444444
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1635444444
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1635444444
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1635444444
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1635444444
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1635444444
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1635444444
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1635444444
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1635444444
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1635444444
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1635444444
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1635444444
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1635444444
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1635444444
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_309
timestamp 1635444444
transform 1 0 29532 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_316
timestamp 1635444444
transform 1 0 30176 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1635444444
transform -1 0 30820 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1635444444
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1635444444
transform 1 0 29900 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_18
timestamp 1635444444
transform 1 0 2760 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_7
timestamp 1635444444
transform 1 0 1748 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1635444444
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0984_
timestamp 1635444444
transform 1 0 2484 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1635444444
transform -1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_26
timestamp 1635444444
transform 1 0 3496 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_31
timestamp 1635444444
transform 1 0 3956 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_38
timestamp 1635444444
transform 1 0 4600 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1635444444
transform -1 0 3956 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1485_
timestamp 1635444444
transform 1 0 4324 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1490_
timestamp 1635444444
transform -1 0 5244 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_45
timestamp 1635444444
transform 1 0 5244 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_52
timestamp 1635444444
transform 1 0 5888 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_57
timestamp 1635444444
transform 1 0 6348 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1635444444
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1235_
timestamp 1635444444
transform 1 0 5612 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1635444444
transform 1 0 6716 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_75_77
timestamp 1635444444
transform 1 0 8188 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_83
timestamp 1635444444
transform 1 0 8740 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1635444444
transform -1 0 10304 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_75_100
timestamp 1635444444
transform 1 0 10304 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1635444444
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1635444444
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1635444444
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1635444444
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1635444444
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1635444444
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1635444444
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1635444444
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1635444444
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_181
timestamp 1635444444
transform 1 0 17756 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_190
timestamp 1635444444
transform 1 0 18584 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _0942_
timestamp 1635444444
transform -1 0 18584 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_202
timestamp 1635444444
transform 1 0 19688 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_214
timestamp 1635444444
transform 1 0 20792 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_222
timestamp 1635444444
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1635444444
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1635444444
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1635444444
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1635444444
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1635444444
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1635444444
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1635444444
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1635444444
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1635444444
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1635444444
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1635444444
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_317
timestamp 1635444444
transform 1 0 30268 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1635444444
transform -1 0 30820 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_16
timestamp 1635444444
transform 1 0 2576 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_3
timestamp 1635444444
transform 1 0 1380 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_9
timestamp 1635444444
transform 1 0 1932 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1635444444
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1473_
timestamp 1635444444
transform 1 0 1656 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1475_
timestamp 1635444444
transform -1 0 2576 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1483_
timestamp 1635444444
transform 1 0 2944 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_23
timestamp 1635444444
transform 1 0 3220 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1635444444
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_32
timestamp 1635444444
transform 1 0 4048 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1635444444
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1478_
timestamp 1635444444
transform -1 0 4048 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_76_44
timestamp 1635444444
transform 1 0 5152 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_52
timestamp 1635444444
transform 1 0 5888 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_58
timestamp 1635444444
transform 1 0 6440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_62
timestamp 1635444444
transform 1 0 6808 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1232_
timestamp 1635444444
transform -1 0 6808 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1493_
timestamp 1635444444
transform -1 0 5888 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_76_70
timestamp 1635444444
transform 1 0 7544 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_80
timestamp 1635444444
transform 1 0 8464 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1635444444
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1230_
timestamp 1635444444
transform 1 0 7636 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1635444444
transform 1 0 8924 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_101
timestamp 1635444444
transform 1 0 10396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_113
timestamp 1635444444
transform 1 0 11500 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_125
timestamp 1635444444
transform 1 0 12604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_137
timestamp 1635444444
transform 1 0 13708 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1635444444
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1635444444
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1635444444
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1635444444
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_177
timestamp 1635444444
transform 1 0 17388 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_183
timestamp 1635444444
transform 1 0 17940 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_190
timestamp 1635444444
transform 1 0 18584 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1635444444
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__and2_2  _0934_
timestamp 1635444444
transform -1 0 18584 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1635444444
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1635444444
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1635444444
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1635444444
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1635444444
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1635444444
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1635444444
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1635444444
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1635444444
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1635444444
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1635444444
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1635444444
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1635444444
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_309
timestamp 1635444444
transform 1 0 29532 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_317
timestamp 1635444444
transform 1 0 30268 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1635444444
transform -1 0 30820 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1635444444
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_14
timestamp 1635444444
transform 1 0 2392 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_21
timestamp 1635444444
transform 1 0 3036 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_7
timestamp 1635444444
transform 1 0 1748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1635444444
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1480_
timestamp 1635444444
transform 1 0 2116 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1487_
timestamp 1635444444
transform 1 0 2760 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1635444444
transform -1 0 1748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_28
timestamp 1635444444
transform 1 0 3680 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_41
timestamp 1635444444
transform 1 0 4876 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1489_
timestamp 1635444444
transform 1 0 3404 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1499_
timestamp 1635444444
transform 1 0 4232 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_77_52
timestamp 1635444444
transform 1 0 5888 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_60
timestamp 1635444444
transform 1 0 6624 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1635444444
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1233_
timestamp 1635444444
transform 1 0 6348 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1234_
timestamp 1635444444
transform -1 0 7820 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1495_
timestamp 1635444444
transform -1 0 5888 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_77_73
timestamp 1635444444
transform 1 0 7820 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_86
timestamp 1635444444
transform 1 0 9016 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1227_
timestamp 1635444444
transform 1 0 8188 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1635444444
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1635444444
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1220_
timestamp 1635444444
transform 1 0 9384 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1635444444
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1635444444
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1635444444
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1635444444
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1635444444
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1635444444
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1635444444
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1635444444
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1635444444
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1635444444
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_181
timestamp 1635444444
transform 1 0 17756 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_190
timestamp 1635444444
transform 1 0 18584 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _0938_
timestamp 1635444444
transform -1 0 18584 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_202
timestamp 1635444444
transform 1 0 19688 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_214
timestamp 1635444444
transform 1 0 20792 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_222
timestamp 1635444444
transform 1 0 21528 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1635444444
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1635444444
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1635444444
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1635444444
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1635444444
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1635444444
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1635444444
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1635444444
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1635444444
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1635444444
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_305
timestamp 1635444444
transform 1 0 29164 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_316
timestamp 1635444444
transform 1 0 30176 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1635444444
transform -1 0 30820 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1635444444
transform 1 0 29900 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_15
timestamp 1635444444
transform 1 0 2484 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_7
timestamp 1635444444
transform 1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1635444444
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1635444444
transform 1 0 2852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1635444444
transform -1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1635444444
transform -1 0 2484 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_22
timestamp 1635444444
transform 1 0 3128 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_32
timestamp 1635444444
transform 1 0 4048 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_39
timestamp 1635444444
transform 1 0 4692 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1635444444
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1494_
timestamp 1635444444
transform 1 0 3772 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 1635444444
transform 1 0 4416 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_78_52
timestamp 1635444444
transform 1 0 5888 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1497_
timestamp 1635444444
transform -1 0 5888 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1635444444
transform 1 0 6624 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_78_76
timestamp 1635444444
transform 1 0 8096 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1635444444
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1229_
timestamp 1635444444
transform -1 0 9200 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_100
timestamp 1635444444
transform 1 0 10304 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_88
timestamp 1635444444
transform 1 0 9200 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_112
timestamp 1635444444
transform 1 0 11408 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_124
timestamp 1635444444
transform 1 0 12512 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_136
timestamp 1635444444
transform 1 0 13616 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1635444444
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1635444444
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1635444444
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1635444444
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1635444444
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1635444444
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1635444444
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1635444444
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1635444444
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1635444444
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1635444444
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1635444444
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1635444444
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1635444444
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1635444444
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1635444444
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1635444444
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1635444444
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1635444444
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1635444444
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1635444444
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_309
timestamp 1635444444
transform 1 0 29532 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_316
timestamp 1635444444
transform 1 0 30176 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1635444444
transform -1 0 30820 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1635444444
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1635444444
transform 1 0 29900 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_15
timestamp 1635444444
transform 1 0 2484 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_7
timestamp 1635444444
transform 1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1635444444
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1635444444
transform -1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1635444444
transform -1 0 2484 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1635444444
transform -1 0 3220 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_23
timestamp 1635444444
transform 1 0 3220 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_27
timestamp 1635444444
transform 1 0 3588 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_32
timestamp 1635444444
transform 1 0 4048 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1635444444
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1635444444
transform 1 0 3680 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1635444444
transform 1 0 3772 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1635444444
transform 1 0 4416 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1635444444
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1635444444
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1635444444
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1635444444
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1635444444
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_81
timestamp 1635444444
transform 1 0 8556 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_85
timestamp 1635444444
transform 1 0 8924 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1635444444
transform 1 0 8832 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_109
timestamp 1635444444
transform 1 0 11132 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_97
timestamp 1635444444
transform 1 0 10028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1635444444
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1635444444
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1635444444
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_137
timestamp 1635444444
transform 1 0 13708 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_141
timestamp 1635444444
transform 1 0 14076 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1635444444
transform 1 0 13984 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_153
timestamp 1635444444
transform 1 0 15180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_165
timestamp 1635444444
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1635444444
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1635444444
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1635444444
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_193
timestamp 1635444444
transform 1 0 18860 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1635444444
transform 1 0 19136 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_197
timestamp 1635444444
transform 1 0 19228 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_209
timestamp 1635444444
transform 1 0 20332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_221
timestamp 1635444444
transform 1 0 21436 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1635444444
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1635444444
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1635444444
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_249
timestamp 1635444444
transform 1 0 24012 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_253
timestamp 1635444444
transform 1 0 24380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1635444444
transform 1 0 24288 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_265
timestamp 1635444444
transform 1 0 25484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_277
timestamp 1635444444
transform 1 0 26588 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1635444444
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1635444444
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1635444444
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_305
timestamp 1635444444
transform 1 0 29164 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_309
timestamp 1635444444
transform 1 0 29532 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_316
timestamp 1635444444
transform 1 0 30176 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1635444444
transform -1 0 30820 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1635444444
transform 1 0 29440 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1635444444
transform 1 0 29900 0 -1 45696
box -38 -48 314 592
<< labels >>
rlabel metal3 s 31200 3680 32000 3800 6 hb_clk_o
port 0 nsew signal tristate
rlabel metal3 s 31200 5312 32000 5432 6 hb_clkn_o
port 1 nsew signal tristate
rlabel metal3 s 31200 2184 32000 2304 6 hb_csn_o
port 2 nsew signal tristate
rlabel metal3 s 31200 36184 32000 36304 6 hb_dq_i[0]
port 3 nsew signal input
rlabel metal3 s 31200 37816 32000 37936 6 hb_dq_i[1]
port 4 nsew signal input
rlabel metal3 s 31200 39312 32000 39432 6 hb_dq_i[2]
port 5 nsew signal input
rlabel metal3 s 31200 40944 32000 41064 6 hb_dq_i[3]
port 6 nsew signal input
rlabel metal3 s 31200 42440 32000 42560 6 hb_dq_i[4]
port 7 nsew signal input
rlabel metal3 s 31200 43936 32000 44056 6 hb_dq_i[5]
port 8 nsew signal input
rlabel metal3 s 31200 45568 32000 45688 6 hb_dq_i[6]
port 9 nsew signal input
rlabel metal3 s 31200 47064 32000 47184 6 hb_dq_i[7]
port 10 nsew signal input
rlabel metal3 s 31200 9936 32000 10056 6 hb_dq_o[0]
port 11 nsew signal tristate
rlabel metal3 s 31200 13064 32000 13184 6 hb_dq_o[1]
port 12 nsew signal tristate
rlabel metal3 s 31200 16056 32000 16176 6 hb_dq_o[2]
port 13 nsew signal tristate
rlabel metal3 s 31200 19184 32000 19304 6 hb_dq_o[3]
port 14 nsew signal tristate
rlabel metal3 s 31200 22312 32000 22432 6 hb_dq_o[4]
port 15 nsew signal tristate
rlabel metal3 s 31200 25440 32000 25560 6 hb_dq_o[5]
port 16 nsew signal tristate
rlabel metal3 s 31200 28432 32000 28552 6 hb_dq_o[6]
port 17 nsew signal tristate
rlabel metal3 s 31200 31560 32000 31680 6 hb_dq_o[7]
port 18 nsew signal tristate
rlabel metal3 s 31200 11432 32000 11552 6 hb_dq_oen[0]
port 19 nsew signal tristate
rlabel metal3 s 31200 14560 32000 14680 6 hb_dq_oen[1]
port 20 nsew signal tristate
rlabel metal3 s 31200 17688 32000 17808 6 hb_dq_oen[2]
port 21 nsew signal tristate
rlabel metal3 s 31200 20816 32000 20936 6 hb_dq_oen[3]
port 22 nsew signal tristate
rlabel metal3 s 31200 23808 32000 23928 6 hb_dq_oen[4]
port 23 nsew signal tristate
rlabel metal3 s 31200 26936 32000 27056 6 hb_dq_oen[5]
port 24 nsew signal tristate
rlabel metal3 s 31200 30064 32000 30184 6 hb_dq_oen[6]
port 25 nsew signal tristate
rlabel metal3 s 31200 33192 32000 33312 6 hb_dq_oen[7]
port 26 nsew signal tristate
rlabel metal3 s 31200 688 32000 808 6 hb_rstn_o
port 27 nsew signal tristate
rlabel metal3 s 31200 34688 32000 34808 6 hb_rwds_i
port 28 nsew signal input
rlabel metal3 s 31200 6808 32000 6928 6 hb_rwds_o
port 29 nsew signal tristate
rlabel metal3 s 31200 8304 32000 8424 6 hb_rwds_oen
port 30 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 rst_i
port 31 nsew signal input
rlabel metal4 s 5909 2128 6229 45744 6 vccd1
port 32 nsew power input
rlabel metal4 s 15839 2128 16159 45744 6 vccd1
port 32 nsew power input
rlabel metal4 s 25770 2128 26090 45744 6 vccd1
port 32 nsew power input
rlabel metal4 s 10874 2128 11194 45744 6 vssd1
port 33 nsew ground input
rlabel metal4 s 20805 2128 21125 45744 6 vssd1
port 33 nsew ground input
rlabel metal2 s 1122 0 1178 800 6 wb_clk_i
port 34 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wb_rst_i
port 35 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 wbs_ack_o
port 36 nsew signal tristate
rlabel metal2 s 7930 0 7986 800 6 wbs_adr_i[0]
port 37 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[10]
port 38 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[11]
port 39 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_adr_i[12]
port 40 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[13]
port 41 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[14]
port 42 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[15]
port 43 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[16]
port 44 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[17]
port 45 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_adr_i[18]
port 46 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[19]
port 47 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[1]
port 48 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_adr_i[20]
port 49 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[21]
port 50 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[22]
port 51 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[23]
port 52 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[24]
port 53 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_adr_i[25]
port 54 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_adr_i[26]
port 55 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[27]
port 56 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[28]
port 57 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[29]
port 58 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_adr_i[2]
port 59 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[30]
port 60 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_adr_i[31]
port 61 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[3]
port 62 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_adr_i[4]
port 63 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_adr_i[5]
port 64 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[6]
port 65 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[7]
port 66 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_adr_i[8]
port 67 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[9]
port 68 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_cyc_i
port 69 nsew signal input
rlabel metal3 s 0 280 800 400 6 wbs_dat_i[0]
port 70 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 wbs_dat_i[10]
port 71 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 wbs_dat_i[11]
port 72 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 wbs_dat_i[12]
port 73 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 wbs_dat_i[13]
port 74 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 wbs_dat_i[14]
port 75 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 wbs_dat_i[15]
port 76 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 wbs_dat_i[16]
port 77 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 wbs_dat_i[17]
port 78 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 wbs_dat_i[18]
port 79 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 wbs_dat_i[19]
port 80 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wbs_dat_i[1]
port 81 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 wbs_dat_i[20]
port 82 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 wbs_dat_i[21]
port 83 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 wbs_dat_i[22]
port 84 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 wbs_dat_i[23]
port 85 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 wbs_dat_i[24]
port 86 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 wbs_dat_i[25]
port 87 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wbs_dat_i[26]
port 88 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 wbs_dat_i[27]
port 89 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 wbs_dat_i[28]
port 90 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 wbs_dat_i[29]
port 91 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 wbs_dat_i[2]
port 92 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 wbs_dat_i[30]
port 93 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wbs_dat_i[31]
port 94 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 wbs_dat_i[3]
port 95 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 wbs_dat_i[4]
port 96 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 wbs_dat_i[5]
port 97 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 wbs_dat_i[6]
port 98 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 wbs_dat_i[7]
port 99 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wbs_dat_i[8]
port 100 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wbs_dat_i[9]
port 101 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 wbs_dat_o[0]
port 102 nsew signal tristate
rlabel metal3 s 0 31288 800 31408 6 wbs_dat_o[10]
port 103 nsew signal tristate
rlabel metal3 s 0 31968 800 32088 6 wbs_dat_o[11]
port 104 nsew signal tristate
rlabel metal3 s 0 32648 800 32768 6 wbs_dat_o[12]
port 105 nsew signal tristate
rlabel metal3 s 0 33464 800 33584 6 wbs_dat_o[13]
port 106 nsew signal tristate
rlabel metal3 s 0 34144 800 34264 6 wbs_dat_o[14]
port 107 nsew signal tristate
rlabel metal3 s 0 34960 800 35080 6 wbs_dat_o[15]
port 108 nsew signal tristate
rlabel metal3 s 0 35640 800 35760 6 wbs_dat_o[16]
port 109 nsew signal tristate
rlabel metal3 s 0 36456 800 36576 6 wbs_dat_o[17]
port 110 nsew signal tristate
rlabel metal3 s 0 37136 800 37256 6 wbs_dat_o[18]
port 111 nsew signal tristate
rlabel metal3 s 0 37816 800 37936 6 wbs_dat_o[19]
port 112 nsew signal tristate
rlabel metal3 s 0 24624 800 24744 6 wbs_dat_o[1]
port 113 nsew signal tristate
rlabel metal3 s 0 38632 800 38752 6 wbs_dat_o[20]
port 114 nsew signal tristate
rlabel metal3 s 0 39312 800 39432 6 wbs_dat_o[21]
port 115 nsew signal tristate
rlabel metal3 s 0 40128 800 40248 6 wbs_dat_o[22]
port 116 nsew signal tristate
rlabel metal3 s 0 40808 800 40928 6 wbs_dat_o[23]
port 117 nsew signal tristate
rlabel metal3 s 0 41624 800 41744 6 wbs_dat_o[24]
port 118 nsew signal tristate
rlabel metal3 s 0 42304 800 42424 6 wbs_dat_o[25]
port 119 nsew signal tristate
rlabel metal3 s 0 42984 800 43104 6 wbs_dat_o[26]
port 120 nsew signal tristate
rlabel metal3 s 0 43800 800 43920 6 wbs_dat_o[27]
port 121 nsew signal tristate
rlabel metal3 s 0 44480 800 44600 6 wbs_dat_o[28]
port 122 nsew signal tristate
rlabel metal3 s 0 45296 800 45416 6 wbs_dat_o[29]
port 123 nsew signal tristate
rlabel metal3 s 0 25304 800 25424 6 wbs_dat_o[2]
port 124 nsew signal tristate
rlabel metal3 s 0 45976 800 46096 6 wbs_dat_o[30]
port 125 nsew signal tristate
rlabel metal3 s 0 46792 800 46912 6 wbs_dat_o[31]
port 126 nsew signal tristate
rlabel metal3 s 0 26120 800 26240 6 wbs_dat_o[3]
port 127 nsew signal tristate
rlabel metal3 s 0 26800 800 26920 6 wbs_dat_o[4]
port 128 nsew signal tristate
rlabel metal3 s 0 27480 800 27600 6 wbs_dat_o[5]
port 129 nsew signal tristate
rlabel metal3 s 0 28296 800 28416 6 wbs_dat_o[6]
port 130 nsew signal tristate
rlabel metal3 s 0 28976 800 29096 6 wbs_dat_o[7]
port 131 nsew signal tristate
rlabel metal3 s 0 29792 800 29912 6 wbs_dat_o[8]
port 132 nsew signal tristate
rlabel metal3 s 0 30472 800 30592 6 wbs_dat_o[9]
port 133 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 wbs_sel_i[0]
port 134 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_sel_i[1]
port 135 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_sel_i[2]
port 136 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_sel_i[3]
port 137 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_stb_i
port 138 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_we_i
port 139 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32000 48000
<< end >>
